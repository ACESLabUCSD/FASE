
module MAC_TG_N32 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047;
  wire   [31:0] o_reg;

  DFF \o_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[0])
         );
  DFF \o_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[1])
         );
  DFF \o_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[2])
         );
  DFF \o_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[3])
         );
  DFF \o_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[4])
         );
  DFF \o_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[5])
         );
  DFF \o_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[6])
         );
  DFF \o_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[7])
         );
  DFF \o_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[8])
         );
  DFF \o_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[9])
         );
  DFF \o_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[10]) );
  DFF \o_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[11]) );
  DFF \o_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[12]) );
  DFF \o_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[13]) );
  DFF \o_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[14]) );
  DFF \o_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[15]) );
  DFF \o_reg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[16]) );
  DFF \o_reg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[17]) );
  DFF \o_reg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[18]) );
  DFF \o_reg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[19]) );
  DFF \o_reg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[20]) );
  DFF \o_reg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[21]) );
  DFF \o_reg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[22]) );
  DFF \o_reg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[23]) );
  DFF \o_reg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[24]) );
  DFF \o_reg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[25]) );
  DFF \o_reg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[26]) );
  DFF \o_reg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[27]) );
  DFF \o_reg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[28]) );
  DFF \o_reg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[29]) );
  DFF \o_reg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[30]) );
  DFF \o_reg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[31]) );
  MUX U35 ( .IN0(n4344), .IN1(n33), .SEL(n3981), .F(n4332) );
  IV U36 ( .A(n3980), .Z(n33) );
  MUX U37 ( .IN0(n3953), .IN1(n34), .SEL(n3954), .F(n3935) );
  IV U38 ( .A(n3955), .Z(n34) );
  MUX U39 ( .IN0(n3519), .IN1(n35), .SEL(n3520), .F(n3479) );
  IV U40 ( .A(n3521), .Z(n35) );
  MUX U41 ( .IN0(n761), .IN1(n36), .SEL(n762), .F(n725) );
  IV U42 ( .A(n763), .Z(n36) );
  MUX U43 ( .IN0(n1088), .IN1(n37), .SEL(n1089), .F(n1021) );
  IV U44 ( .A(n1090), .Z(n37) );
  MUX U45 ( .IN0(n1146), .IN1(n38), .SEL(n1147), .F(n1079) );
  IV U46 ( .A(n1148), .Z(n38) );
  MUX U47 ( .IN0(n1175), .IN1(n39), .SEL(n1176), .F(n1108) );
  IV U48 ( .A(n1177), .Z(n39) );
  MUX U49 ( .IN0(n663), .IN1(n40), .SEL(n664), .F(n640) );
  IV U50 ( .A(n665), .Z(n40) );
  MUX U51 ( .IN0(n795), .IN1(n41), .SEL(n796), .F(n756) );
  IV U52 ( .A(n797), .Z(n41) );
  MUX U53 ( .IN0(n861), .IN1(n42), .SEL(n862), .F(n804) );
  IV U54 ( .A(n863), .Z(n42) );
  MUX U55 ( .IN0(n1045), .IN1(n43), .SEL(n1046), .F(n987) );
  IV U56 ( .A(n1047), .Z(n43) );
  MUX U57 ( .IN0(n1375), .IN1(n44), .SEL(n1376), .F(n1301) );
  IV U58 ( .A(n1377), .Z(n44) );
  MUX U59 ( .IN0(n1415), .IN1(n45), .SEL(n1416), .F(n1322) );
  IV U60 ( .A(n1417), .Z(n45) );
  MUX U61 ( .IN0(n1737), .IN1(n46), .SEL(n1738), .F(n1644) );
  IV U62 ( .A(n1739), .Z(n46) );
  MUX U63 ( .IN0(n2503), .IN1(n47), .SEL(n2504), .F(n2471) );
  IV U64 ( .A(n2505), .Z(n47) );
  MUX U65 ( .IN0(n2591), .IN1(n48), .SEL(n2592), .F(n2543) );
  IV U66 ( .A(n2593), .Z(n48) );
  MUX U67 ( .IN0(n2164), .IN1(n49), .SEL(n2165), .F(n2089) );
  IV U68 ( .A(n2166), .Z(n49) );
  MUX U69 ( .IN0(n2728), .IN1(n50), .SEL(n2729), .F(n2679) );
  IV U70 ( .A(n2730), .Z(n50) );
  MUX U71 ( .IN0(n938), .IN1(n51), .SEL(n939), .F(n884) );
  IV U72 ( .A(n940), .Z(n51) );
  MUX U73 ( .IN0(n1655), .IN1(n52), .SEL(n1656), .F(n1566) );
  IV U74 ( .A(n1657), .Z(n52) );
  MUX U75 ( .IN0(n3559), .IN1(n53), .SEL(n3560), .F(n3519) );
  IV U76 ( .A(n3561), .Z(n53) );
  MUX U77 ( .IN0(n4332), .IN1(n54), .SEL(n3963), .F(n4320) );
  IV U78 ( .A(n3962), .Z(n54) );
  XNOR U79 ( .A(n3947), .B(n3932), .Z(n3936) );
  XNOR U80 ( .A(n3576), .B(n3539), .Z(n3543) );
  MUX U81 ( .IN0(n3399), .IN1(n55), .SEL(n3400), .F(n3359) );
  IV U82 ( .A(n3401), .Z(n55) );
  XNOR U83 ( .A(n3893), .B(n3878), .Z(n3882) );
  MUX U84 ( .IN0(n4424), .IN1(n56), .SEL(n4425), .F(n4412) );
  IV U85 ( .A(n4426), .Z(n56) );
  XNOR U86 ( .A(n4838), .B(n4829), .Z(n4703) );
  MUX U87 ( .IN0(n4111), .IN1(n4113), .SEL(n4112), .F(n4089) );
  MUX U88 ( .IN0(n3199), .IN1(n57), .SEL(n3200), .F(n3159) );
  IV U89 ( .A(n3201), .Z(n57) );
  MUX U90 ( .IN0(n4672), .IN1(n4674), .SEL(n4673), .F(n4650) );
  MUX U91 ( .IN0(n3115), .IN1(n58), .SEL(n3116), .F(n3075) );
  IV U92 ( .A(n3117), .Z(n58) );
  XNOR U93 ( .A(n3785), .B(n3770), .Z(n3774) );
  MUX U94 ( .IN0(n4404), .IN1(n4074), .SEL(n4076), .F(n4392) );
  MUX U95 ( .IN0(n4041), .IN1(n59), .SEL(n4042), .F(n4019) );
  IV U96 ( .A(n4043), .Z(n59) );
  MUX U97 ( .IN0(n4796), .IN1(n4635), .SEL(n4637), .F(n4784) );
  MUX U98 ( .IN0(n2947), .IN1(n60), .SEL(n2948), .F(n2875) );
  IV U99 ( .A(n2949), .Z(n60) );
  MUX U100 ( .IN0(n3701), .IN1(n61), .SEL(n3702), .F(n2977) );
  IV U101 ( .A(n3703), .Z(n61) );
  MUX U102 ( .IN0(n692), .IN1(n62), .SEL(n693), .F(n659) );
  IV U103 ( .A(n694), .Z(n62) );
  MUX U104 ( .IN0(n1288), .IN1(n63), .SEL(n1289), .F(n1216) );
  IV U105 ( .A(n1290), .Z(n63) );
  MUX U106 ( .IN0(n2620), .IN1(n64), .SEL(n2621), .F(n2587) );
  IV U107 ( .A(n2622), .Z(n64) );
  MUX U108 ( .IN0(n2960), .IN1(n65), .SEL(n2961), .F(n2888) );
  IV U109 ( .A(n2962), .Z(n65) );
  MUX U110 ( .IN0(n804), .IN1(n66), .SEL(n805), .F(n765) );
  IV U111 ( .A(n806), .Z(n66) );
  MUX U112 ( .IN0(n902), .IN1(n67), .SEL(n903), .F(n852) );
  IV U113 ( .A(n904), .Z(n67) );
  MUX U114 ( .IN0(n1025), .IN1(n68), .SEL(n1026), .F(n967) );
  IV U115 ( .A(n1027), .Z(n68) );
  MUX U116 ( .IN0(n1179), .IN1(n69), .SEL(n1180), .F(n1112) );
  IV U117 ( .A(n1181), .Z(n69) );
  MUX U118 ( .IN0(n1202), .IN1(n70), .SEL(n1203), .F(n1131) );
  IV U119 ( .A(n1204), .Z(n70) );
  MUX U120 ( .IN0(n1301), .IN1(n71), .SEL(n1302), .F(n1229) );
  IV U121 ( .A(n1303), .Z(n71) );
  MUX U122 ( .IN0(n1644), .IN1(n72), .SEL(n1645), .F(n1554) );
  IV U123 ( .A(n1646), .Z(n72) );
  MUX U124 ( .IN0(n1617), .IN1(n73), .SEL(n1618), .F(n1527) );
  IV U125 ( .A(n1619), .Z(n73) );
  MUX U126 ( .IN0(n1591), .IN1(n74), .SEL(n1592), .F(n1501) );
  IV U127 ( .A(n1593), .Z(n74) );
  MUX U128 ( .IN0(n1663), .IN1(n75), .SEL(n1664), .F(n1570) );
  IV U129 ( .A(n1665), .Z(n75) );
  MUX U130 ( .IN0(n1728), .IN1(n76), .SEL(n1729), .F(n1635) );
  IV U131 ( .A(n1730), .Z(n76) );
  MUX U132 ( .IN0(n1967), .IN1(n77), .SEL(n1968), .F(n1895) );
  IV U133 ( .A(n1969), .Z(n77) );
  MUX U134 ( .IN0(n2543), .IN1(n78), .SEL(n2544), .F(n2512) );
  IV U135 ( .A(n2545), .Z(n78) );
  MUX U136 ( .IN0(n2534), .IN1(n79), .SEL(n2535), .F(n2503) );
  IV U137 ( .A(n2536), .Z(n79) );
  MUX U138 ( .IN0(n2089), .IN1(n80), .SEL(n2090), .F(n2020) );
  IV U139 ( .A(n2091), .Z(n80) );
  MUX U140 ( .IN0(n2062), .IN1(n81), .SEL(n2063), .F(n1993) );
  IV U141 ( .A(n2064), .Z(n81) );
  MUX U142 ( .IN0(n2255), .IN1(n82), .SEL(n2256), .F(n2183) );
  IV U143 ( .A(n2257), .Z(n82) );
  MUX U144 ( .IN0(n2705), .IN1(n83), .SEL(n2706), .F(n2658) );
  IV U145 ( .A(n2707), .Z(n83) );
  MUX U146 ( .IN0(n2714), .IN1(n84), .SEL(n2715), .F(n2667) );
  IV U147 ( .A(n2716), .Z(n84) );
  MUX U148 ( .IN0(n2377), .IN1(n85), .SEL(n2378), .F(n2308) );
  IV U149 ( .A(n2379), .Z(n85) );
  MUX U150 ( .IN0(n2747), .IN1(n86), .SEL(n2748), .F(n2728) );
  IV U151 ( .A(n2749), .Z(n86) );
  MUX U152 ( .IN0(n687), .IN1(n87), .SEL(n688), .F(n655) );
  IV U153 ( .A(n689), .Z(n87) );
  MUX U154 ( .IN0(n1141), .IN1(n88), .SEL(n1142), .F(n1074) );
  IV U155 ( .A(n1143), .Z(n88) );
  MUX U156 ( .IN0(n1450), .IN1(n89), .SEL(n1451), .F(n1357) );
  IV U157 ( .A(n1452), .Z(n89) );
  MUX U158 ( .IN0(n1855), .IN1(n90), .SEL(n1856), .F(n1719) );
  IV U159 ( .A(n1857), .Z(n90) );
  MUX U160 ( .IN0(n2218), .IN1(n91), .SEL(n2219), .F(n2146) );
  IV U161 ( .A(n2220), .Z(n91) );
  MUX U162 ( .IN0(n995), .IN1(n92), .SEL(n996), .F(n938) );
  IV U163 ( .A(n997), .Z(n92) );
  MUX U164 ( .IN0(n2599), .IN1(n93), .SEL(n2103), .F(n2551) );
  IV U165 ( .A(n2102), .Z(n93) );
  ANDN U166 ( .A(n1581), .B(n1582), .Z(n1491) );
  MUX U167 ( .IN0(n1812), .IN1(n94), .SEL(n1748), .F(n1671) );
  IV U168 ( .A(n1747), .Z(n94) );
  MUX U169 ( .IN0(n3555), .IN1(n95), .SEL(n3556), .F(n3515) );
  IV U170 ( .A(n3557), .Z(n95) );
  MUX U171 ( .IN0(n3949), .IN1(n96), .SEL(n3950), .F(n3931) );
  IV U172 ( .A(n3951), .Z(n96) );
  MUX U173 ( .IN0(n3935), .IN1(n97), .SEL(n3936), .F(n3917) );
  IV U174 ( .A(n3937), .Z(n97) );
  XNOR U175 ( .A(n3536), .B(n3499), .Z(n3503) );
  XNOR U176 ( .A(n4314), .B(n4305), .Z(n3927) );
  XNOR U177 ( .A(n3473), .B(n3436), .Z(n3440) );
  MUX U178 ( .IN0(n3338), .IN1(n98), .SEL(n3339), .F(n3298) );
  IV U179 ( .A(n3340), .Z(n98) );
  MUX U180 ( .IN0(n3319), .IN1(n99), .SEL(n3320), .F(n3279) );
  IV U181 ( .A(n3321), .Z(n99) );
  XNOR U182 ( .A(n4266), .B(n4257), .Z(n3855) );
  MUX U183 ( .IN0(n3845), .IN1(n100), .SEL(n3846), .F(n3827) );
  IV U184 ( .A(n3847), .Z(n100) );
  XNOR U185 ( .A(n4434), .B(n4425), .Z(n4120) );
  MUX U186 ( .IN0(n4133), .IN1(n101), .SEL(n4134), .F(n4111) );
  IV U187 ( .A(n4135), .Z(n101) );
  MUX U188 ( .IN0(n4844), .IN1(n4721), .SEL(n4722), .F(n4832) );
  MUX U189 ( .IN0(n4716), .IN1(n102), .SEL(n4717), .F(n4694) );
  IV U190 ( .A(n4718), .Z(n102) );
  MUX U191 ( .IN0(n4816), .IN1(n103), .SEL(n4817), .F(n4804) );
  IV U192 ( .A(n4818), .Z(n103) );
  XNOR U193 ( .A(n3256), .B(n3219), .Z(n3223) );
  MUX U194 ( .IN0(n4646), .IN1(n104), .SEL(n4647), .F(n4624) );
  IV U195 ( .A(n4648), .Z(n104) );
  MUX U196 ( .IN0(n3159), .IN1(n105), .SEL(n3160), .F(n3119) );
  IV U197 ( .A(n3161), .Z(n105) );
  XNOR U198 ( .A(n4218), .B(n4209), .Z(n3783) );
  MUX U199 ( .IN0(n3773), .IN1(n106), .SEL(n3774), .F(n3755) );
  IV U200 ( .A(n3775), .Z(n106) );
  MUX U201 ( .IN0(n3075), .IN1(n107), .SEL(n3076), .F(n3035) );
  IV U202 ( .A(n3077), .Z(n107) );
  MUX U203 ( .IN0(n4392), .IN1(n4052), .SEL(n4054), .F(n4380) );
  MUX U204 ( .IN0(n4045), .IN1(n4047), .SEL(n4046), .F(n4023) );
  MUX U205 ( .IN0(n3102), .IN1(n108), .SEL(n3103), .F(n3062) );
  IV U206 ( .A(n3104), .Z(n108) );
  MUX U207 ( .IN0(n4606), .IN1(n4608), .SEL(n4607), .F(n4584) );
  MUX U208 ( .IN0(n4772), .IN1(n4591), .SEL(n4593), .F(n4760) );
  MUX U209 ( .IN0(n907), .IN1(n109), .SEL(n908), .F(n857) );
  IV U210 ( .A(n909), .Z(n109) );
  MUX U211 ( .IN0(n954), .IN1(n110), .SEL(n955), .F(n898) );
  IV U212 ( .A(n956), .Z(n110) );
  MUX U213 ( .IN0(n1041), .IN1(n111), .SEL(n1042), .F(n983) );
  IV U214 ( .A(n1043), .Z(n111) );
  MUX U215 ( .IN0(n1437), .IN1(n112), .SEL(n1438), .F(n1344) );
  IV U216 ( .A(n1439), .Z(n112) );
  MUX U217 ( .IN0(n1541), .IN1(n113), .SEL(n1542), .F(n1455) );
  IV U218 ( .A(n1543), .Z(n113) );
  MUX U219 ( .IN0(n1587), .IN1(n114), .SEL(n1588), .F(n1497) );
  IV U220 ( .A(n1589), .Z(n114) );
  MUX U221 ( .IN0(n2477), .IN1(n115), .SEL(n2478), .F(n1800) );
  IV U222 ( .A(n2479), .Z(n115) );
  MUX U223 ( .IN0(n1963), .IN1(n116), .SEL(n1964), .F(n1891) );
  IV U224 ( .A(n1965), .Z(n116) );
  MUX U225 ( .IN0(n2085), .IN1(n117), .SEL(n2086), .F(n2016) );
  IV U226 ( .A(n2087), .Z(n117) );
  MUX U227 ( .IN0(n2076), .IN1(n118), .SEL(n2077), .F(n2007) );
  IV U228 ( .A(n2078), .Z(n118) );
  MUX U229 ( .IN0(n2251), .IN1(n119), .SEL(n2252), .F(n2179) );
  IV U230 ( .A(n2253), .Z(n119) );
  MUX U231 ( .IN0(n2364), .IN1(n120), .SEL(n2365), .F(n2295) );
  IV U232 ( .A(n2366), .Z(n120) );
  MUX U233 ( .IN0(n2448), .IN1(n121), .SEL(n2449), .F(n2373) );
  IV U234 ( .A(n2450), .Z(n121) );
  MUX U235 ( .IN0(n2421), .IN1(n122), .SEL(n2422), .F(n2346) );
  IV U236 ( .A(n2423), .Z(n122) );
  MUX U237 ( .IN0(n2811), .IN1(n123), .SEL(n2812), .F(n2778) );
  IV U238 ( .A(n2813), .Z(n123) );
  MUX U239 ( .IN0(n2835), .IN1(n124), .SEL(n2836), .F(n2743) );
  IV U240 ( .A(n2837), .Z(n124) );
  MUX U241 ( .IN0(n2977), .IN1(n125), .SEL(n2978), .F(n2906) );
  IV U242 ( .A(n2979), .Z(n125) );
  MUX U243 ( .IN0(n729), .IN1(n126), .SEL(n730), .F(n696) );
  IV U244 ( .A(n731), .Z(n126) );
  MUX U245 ( .IN0(n1083), .IN1(n127), .SEL(n1084), .F(n1016) );
  IV U246 ( .A(n1085), .Z(n127) );
  MUX U247 ( .IN0(n1159), .IN1(n128), .SEL(n1160), .F(n1092) );
  IV U248 ( .A(n1161), .Z(n128) );
  MUX U249 ( .IN0(n1249), .IN1(n129), .SEL(n1250), .F(n1179) );
  IV U250 ( .A(n1251), .Z(n129) );
  MUX U251 ( .IN0(n1274), .IN1(n130), .SEL(n1275), .F(n1202) );
  IV U252 ( .A(n1276), .Z(n130) );
  MUX U253 ( .IN0(n1366), .IN1(n131), .SEL(n1367), .F(n1292) );
  IV U254 ( .A(n1368), .Z(n131) );
  MUX U255 ( .IN0(n1468), .IN1(n132), .SEL(n1469), .F(n1375) );
  IV U256 ( .A(n1470), .Z(n132) );
  MUX U257 ( .IN0(n1873), .IN1(n133), .SEL(n1874), .F(n1737) );
  IV U258 ( .A(n1875), .Z(n133) );
  MUX U259 ( .IN0(n1846), .IN1(n134), .SEL(n1847), .F(n1710) );
  IV U260 ( .A(n1848), .Z(n134) );
  MUX U261 ( .IN0(n1820), .IN1(n135), .SEL(n1821), .F(n1684) );
  IV U262 ( .A(n1822), .Z(n135) );
  MUX U263 ( .IN0(n1939), .IN1(n136), .SEL(n1940), .F(n1864) );
  IV U264 ( .A(n1941), .Z(n136) );
  MUX U265 ( .IN0(n2111), .IN1(n137), .SEL(n2112), .F(n2036) );
  IV U266 ( .A(n2113), .Z(n137) );
  MUX U267 ( .IN0(n2615), .IN1(n138), .SEL(n2616), .F(n2582) );
  IV U268 ( .A(n2617), .Z(n138) );
  MUX U269 ( .IN0(n2624), .IN1(n139), .SEL(n2625), .F(n2591) );
  IV U270 ( .A(n2626), .Z(n139) );
  MUX U271 ( .IN0(n2227), .IN1(n140), .SEL(n2228), .F(n2155) );
  IV U272 ( .A(n2229), .Z(n140) );
  MUX U273 ( .IN0(n2308), .IN1(n141), .SEL(n2309), .F(n2236) );
  IV U274 ( .A(n2310), .Z(n141) );
  MUX U275 ( .IN0(n2281), .IN1(n142), .SEL(n2282), .F(n2209) );
  IV U276 ( .A(n2283), .Z(n142) );
  MUX U277 ( .IN0(n2399), .IN1(n143), .SEL(n2400), .F(n2324) );
  IV U278 ( .A(n2401), .Z(n143) );
  MUX U279 ( .IN0(n2824), .IN1(n144), .SEL(n2825), .F(n2791) );
  IV U280 ( .A(n2826), .Z(n144) );
  MUX U281 ( .IN0(n787), .IN1(n145), .SEL(n788), .F(n750) );
  IV U282 ( .A(n789), .Z(n145) );
  MUX U283 ( .IN0(n146), .IN1(n1065), .SEL(n1066), .F(n998) );
  IV U284 ( .A(n1067), .Z(n146) );
  MUX U285 ( .IN0(n1283), .IN1(n147), .SEL(n1284), .F(n1211) );
  IV U286 ( .A(n1285), .Z(n147) );
  MUX U287 ( .IN0(n1570), .IN1(n148), .SEL(n1571), .F(n1481) );
  IV U288 ( .A(n1572), .Z(n148) );
  MUX U289 ( .IN0(n1432), .IN1(n149), .SEL(n1433), .F(n1339) );
  IV U290 ( .A(n1434), .Z(n149) );
  MUX U291 ( .IN0(n1626), .IN1(n150), .SEL(n1627), .F(n1536) );
  IV U292 ( .A(n1628), .Z(n150) );
  MUX U293 ( .IN0(n2002), .IN1(n151), .SEL(n2003), .F(n1930) );
  IV U294 ( .A(n2004), .Z(n151) );
  MUX U295 ( .IN0(n1984), .IN1(n152), .SEL(n1985), .F(n1912) );
  IV U296 ( .A(n1986), .Z(n152) );
  MUX U297 ( .IN0(n2679), .IN1(n153), .SEL(n2680), .F(n2633) );
  IV U298 ( .A(n2681), .Z(n153) );
  MUX U299 ( .IN0(n2696), .IN1(n154), .SEL(n2697), .F(n2649) );
  IV U300 ( .A(n2698), .Z(n154) );
  MUX U301 ( .IN0(n2434), .IN1(n155), .SEL(n2435), .F(n2359) );
  IV U302 ( .A(n2436), .Z(n155) );
  MUX U303 ( .IN0(n875), .IN1(n156), .SEL(n876), .F(n820) );
  IV U304 ( .A(n877), .Z(n156) );
  MUX U305 ( .IN0(n884), .IN1(n157), .SEL(n885), .F(n830) );
  IV U306 ( .A(n886), .Z(n157) );
  MUX U307 ( .IN0(n1120), .IN1(n158), .SEL(n1121), .F(n1053) );
  IV U308 ( .A(n1122), .Z(n158) );
  MUX U309 ( .IN0(n1828), .IN1(n159), .SEL(n1829), .F(n1692) );
  IV U310 ( .A(n1830), .Z(n159) );
  MUX U311 ( .IN0(n2119), .IN1(n160), .SEL(n2120), .F(n2044) );
  IV U312 ( .A(n2121), .Z(n160) );
  MUX U313 ( .IN0(n2642), .IN1(n161), .SEL(n2175), .F(n2599) );
  IV U314 ( .A(n2174), .Z(n161) );
  MUX U315 ( .IN0(n1578), .IN1(n162), .SEL(n1579), .F(n1488) );
  IV U316 ( .A(n1580), .Z(n162) );
  ANDN U317 ( .A(n1887), .B(n1886), .Z(n1883) );
  MUX U318 ( .IN0(n3569), .IN1(n3587), .SEL(n3570), .F(n3529) );
  MUX U319 ( .IN0(n3578), .IN1(n163), .SEL(n3579), .F(n3538) );
  IV U320 ( .A(n3580), .Z(n163) );
  XNOR U321 ( .A(n4338), .B(n4329), .Z(n3963) );
  MUX U322 ( .IN0(n3921), .IN1(n3938), .SEL(n3922), .F(n3903) );
  XNOR U323 ( .A(n3513), .B(n3476), .Z(n3480) );
  MUX U324 ( .IN0(n3585), .IN1(n164), .SEL(n2969), .F(n3545) );
  IV U325 ( .A(n2968), .Z(n164) );
  XNOR U326 ( .A(n3929), .B(n3914), .Z(n3918) );
  XNOR U327 ( .A(n3496), .B(n3459), .Z(n3463) );
  XNOR U328 ( .A(n4302), .B(n4293), .Z(n3909) );
  MUX U329 ( .IN0(n3359), .IN1(n165), .SEL(n3360), .F(n3319) );
  IV U330 ( .A(n3361), .Z(n165) );
  XNOR U331 ( .A(n3875), .B(n3860), .Z(n3864) );
  MUX U332 ( .IN0(n3275), .IN1(n166), .SEL(n3276), .F(n3235) );
  IV U333 ( .A(n3277), .Z(n166) );
  XNOR U334 ( .A(n3376), .B(n3339), .Z(n3343) );
  MUX U335 ( .IN0(n4440), .IN1(n167), .SEL(n4139), .F(n4428) );
  IV U336 ( .A(n4138), .Z(n167) );
  MUX U337 ( .IN0(n4418), .IN1(n4429), .SEL(n4419), .F(n4406) );
  XNOR U338 ( .A(n3821), .B(n3806), .Z(n3810) );
  XNOR U339 ( .A(n4242), .B(n4233), .Z(n3819) );
  MUX U340 ( .IN0(n4412), .IN1(n168), .SEL(n4413), .F(n4400) );
  IV U341 ( .A(n4414), .Z(n168) );
  XNOR U342 ( .A(n4710), .B(n4691), .Z(n4695) );
  XNOR U343 ( .A(n4105), .B(n4086), .Z(n4090) );
  MUX U344 ( .IN0(n4820), .IN1(n4679), .SEL(n4681), .F(n4808) );
  MUX U345 ( .IN0(n3119), .IN1(n169), .SEL(n3120), .F(n3079) );
  IV U346 ( .A(n3121), .Z(n169) );
  XNOR U347 ( .A(n3176), .B(n3139), .Z(n3143) );
  XNOR U348 ( .A(n4206), .B(n4197), .Z(n3765) );
  MUX U349 ( .IN0(n3755), .IN1(n170), .SEL(n3756), .F(n3737) );
  IV U350 ( .A(n3757), .Z(n170) );
  MUX U351 ( .IN0(n4628), .IN1(n4630), .SEL(n4629), .F(n4606) );
  MUX U352 ( .IN0(n3035), .IN1(n171), .SEL(n3036), .F(n2995) );
  IV U353 ( .A(n3037), .Z(n171) );
  MUX U354 ( .IN0(n3715), .IN1(n172), .SEL(n3716), .F(n3697) );
  IV U355 ( .A(n3717), .Z(n172) );
  MUX U356 ( .IN0(n4380), .IN1(n4030), .SEL(n4032), .F(n4368) );
  MUX U357 ( .IN0(n4023), .IN1(n4025), .SEL(n4024), .F(n4001) );
  XNOR U358 ( .A(n4778), .B(n4769), .Z(n4593) );
  MUX U359 ( .IN0(n4580), .IN1(n173), .SEL(n4581), .F(n4550) );
  IV U360 ( .A(n4582), .Z(n173) );
  XNOR U361 ( .A(n4170), .B(n4161), .Z(n3711) );
  MUX U362 ( .IN0(n3022), .IN1(n174), .SEL(n3023), .F(n2951) );
  IV U363 ( .A(n3024), .Z(n174) );
  MUX U364 ( .IN0(n1155), .IN1(n175), .SEL(n1156), .F(n1088) );
  IV U365 ( .A(n1157), .Z(n175) );
  MUX U366 ( .IN0(n1116), .IN1(n1182), .SEL(n1117), .F(n1049) );
  MUX U367 ( .IN0(n1245), .IN1(n176), .SEL(n1246), .F(n1175) );
  IV U368 ( .A(n1247), .Z(n176) );
  MUX U369 ( .IN0(n1362), .IN1(n177), .SEL(n1363), .F(n1288) );
  IV U370 ( .A(n1364), .Z(n177) );
  MUX U371 ( .IN0(n1733), .IN1(n178), .SEL(n1734), .F(n1640) );
  IV U372 ( .A(n1735), .Z(n178) );
  MUX U373 ( .IN0(n1724), .IN1(n179), .SEL(n1725), .F(n1631) );
  IV U374 ( .A(n1726), .Z(n179) );
  MUX U375 ( .IN0(n1800), .IN1(n180), .SEL(n1801), .F(n1659) );
  IV U376 ( .A(n1802), .Z(n180) );
  MUX U377 ( .IN0(n1842), .IN1(n181), .SEL(n1843), .F(n1706) );
  IV U378 ( .A(n1844), .Z(n181) );
  MUX U379 ( .IN0(n2487), .IN1(n2515), .SEL(n2488), .F(n1808) );
  MUX U380 ( .IN0(n2032), .IN1(n182), .SEL(n2033), .F(n1963) );
  IV U381 ( .A(n2034), .Z(n182) );
  MUX U382 ( .IN0(n2160), .IN1(n183), .SEL(n2161), .F(n2085) );
  IV U383 ( .A(n2162), .Z(n183) );
  MUX U384 ( .IN0(n2205), .IN1(n184), .SEL(n2206), .F(n2133) );
  IV U385 ( .A(n2207), .Z(n184) );
  MUX U386 ( .IN0(n2654), .IN1(n185), .SEL(n2655), .F(n2611) );
  IV U387 ( .A(n2656), .Z(n185) );
  MUX U388 ( .IN0(n2787), .IN1(n186), .SEL(n2788), .F(n2710) );
  IV U389 ( .A(n2789), .Z(n186) );
  MUX U390 ( .IN0(n2743), .IN1(n187), .SEL(n2744), .F(n2724) );
  IV U391 ( .A(n2745), .Z(n187) );
  XNOR U392 ( .A(n4752), .B(n4753), .Z(n4569) );
  MUX U393 ( .IN0(n659), .IN1(n188), .SEL(n660), .F(n638) );
  IV U394 ( .A(n661), .Z(n188) );
  MUX U395 ( .IN0(n696), .IN1(n189), .SEL(n697), .F(n663) );
  IV U396 ( .A(n698), .Z(n189) );
  MUX U397 ( .IN0(n756), .IN1(n190), .SEL(n757), .F(n719) );
  IV U398 ( .A(n758), .Z(n190) );
  MUX U399 ( .IN0(n911), .IN1(n191), .SEL(n912), .F(n861) );
  IV U400 ( .A(n913), .Z(n191) );
  MUX U401 ( .IN0(n958), .IN1(n192), .SEL(n959), .F(n902) );
  IV U402 ( .A(n960), .Z(n192) );
  MUX U403 ( .IN0(n987), .IN1(n193), .SEL(n988), .F(n928) );
  IV U404 ( .A(n989), .Z(n193) );
  MUX U405 ( .IN0(n1220), .IN1(n194), .SEL(n1221), .F(n1150) );
  IV U406 ( .A(n1222), .Z(n194) );
  MUX U407 ( .IN0(n1441), .IN1(n195), .SEL(n1442), .F(n1348) );
  IV U408 ( .A(n1443), .Z(n195) );
  MUX U409 ( .IN0(n1545), .IN1(n196), .SEL(n1546), .F(n1459) );
  IV U410 ( .A(n1547), .Z(n196) );
  MUX U411 ( .IN0(n1501), .IN1(n197), .SEL(n1502), .F(n1415) );
  IV U412 ( .A(n1503), .Z(n197) );
  MUX U413 ( .IN0(n1895), .IN1(n198), .SEL(n1896), .F(n1820) );
  IV U414 ( .A(n1897), .Z(n198) );
  MUX U415 ( .IN0(n2512), .IN1(n199), .SEL(n2513), .F(n2481) );
  IV U416 ( .A(n2514), .Z(n199) );
  MUX U417 ( .IN0(n2020), .IN1(n200), .SEL(n2021), .F(n1948) );
  IV U418 ( .A(n2022), .Z(n200) );
  MUX U419 ( .IN0(n2011), .IN1(n201), .SEL(n2012), .F(n1939) );
  IV U420 ( .A(n2013), .Z(n201) );
  MUX U421 ( .IN0(n1993), .IN1(n202), .SEL(n1994), .F(n1921) );
  IV U422 ( .A(n1995), .Z(n202) );
  MUX U423 ( .IN0(n2183), .IN1(n203), .SEL(n2184), .F(n2111) );
  IV U424 ( .A(n2185), .Z(n203) );
  MUX U425 ( .IN0(n2667), .IN1(n204), .SEL(n2668), .F(n2624) );
  IV U426 ( .A(n2669), .Z(n204) );
  MUX U427 ( .IN0(n2299), .IN1(n205), .SEL(n2300), .F(n2227) );
  IV U428 ( .A(n2301), .Z(n205) );
  MUX U429 ( .IN0(n2350), .IN1(n206), .SEL(n2351), .F(n2281) );
  IV U430 ( .A(n2352), .Z(n206) );
  MUX U431 ( .IN0(n2782), .IN1(n207), .SEL(n2783), .F(n2705) );
  IV U432 ( .A(n2784), .Z(n207) );
  MUX U433 ( .IN0(n2839), .IN1(n208), .SEL(n2840), .F(n2747) );
  IV U434 ( .A(n2841), .Z(n208) );
  MUX U435 ( .IN0(n5026), .IN1(n209), .SEL(n4933), .F(n2452) );
  IV U436 ( .A(n4932), .Z(n209) );
  MUX U437 ( .IN0(n4525), .IN1(n210), .SEL(n4526), .F(n2399) );
  IV U438 ( .A(n4527), .Z(n210) );
  MUX U439 ( .IN0(n2888), .IN1(n211), .SEL(n2889), .F(n2824) );
  IV U440 ( .A(n2890), .Z(n211) );
  MUX U441 ( .IN0(n2942), .IN1(n212), .SEL(n2943), .F(n2870) );
  IV U442 ( .A(n2944), .Z(n212) );
  MUX U443 ( .IN0(n716), .IN1(n213), .SEL(n717), .F(n687) );
  IV U444 ( .A(n718), .Z(n213) );
  MUX U445 ( .IN0(n1074), .IN1(n214), .SEL(n1075), .F(n1007) );
  IV U446 ( .A(n1076), .Z(n214) );
  MUX U447 ( .IN0(n1128), .IN1(n215), .SEL(n1129), .F(n1065) );
  IV U448 ( .A(n1130), .Z(n215) );
  XNOR U449 ( .A(n1462), .B(n1372), .Z(n1376) );
  MUX U450 ( .IN0(n1608), .IN1(n216), .SEL(n1609), .F(n1518) );
  IV U451 ( .A(n1610), .Z(n216) );
  MUX U452 ( .IN0(n2526), .IN1(n217), .SEL(n2527), .F(n2497) );
  IV U453 ( .A(n2528), .Z(n217) );
  MUX U454 ( .IN0(n2071), .IN1(n218), .SEL(n2072), .F(n2002) );
  IV U455 ( .A(n2073), .Z(n218) );
  MUX U456 ( .IN0(n2053), .IN1(n219), .SEL(n2054), .F(n1984) );
  IV U457 ( .A(n2055), .Z(n219) );
  MUX U458 ( .IN0(n2359), .IN1(n220), .SEL(n2360), .F(n2290) );
  IV U459 ( .A(n2361), .Z(n220) );
  MUX U460 ( .IN0(n1187), .IN1(n221), .SEL(n1188), .F(n1120) );
  IV U461 ( .A(n1189), .Z(n221) );
  MUX U462 ( .IN0(n1481), .IN1(n222), .SEL(n1482), .F(n1396) );
  IV U463 ( .A(n1483), .Z(n222) );
  MUX U464 ( .IN0(n1509), .IN1(n223), .SEL(n1510), .F(n1423) );
  IV U465 ( .A(n1511), .Z(n223) );
  XNOR U466 ( .A(n1655), .B(n1791), .Z(n1784) );
  MUX U467 ( .IN0(n2633), .IN1(n224), .SEL(n2634), .F(n2555) );
  IV U468 ( .A(n2635), .Z(n224) );
  MUX U469 ( .IN0(n2191), .IN1(n225), .SEL(n2192), .F(n2119) );
  IV U470 ( .A(n2193), .Z(n225) );
  MUX U471 ( .IN0(n2689), .IN1(n226), .SEL(n2247), .F(n2642) );
  IV U472 ( .A(n2246), .Z(n226) );
  MUX U473 ( .IN0(n4533), .IN1(n227), .SEL(n2934), .F(n2407) );
  IV U474 ( .A(n2933), .Z(n227) );
  MUX U475 ( .IN0(n778), .IN1(n228), .SEL(n779), .F(n743) );
  IV U476 ( .A(n780), .Z(n228) );
  MUX U477 ( .IN0(n1404), .IN1(n229), .SEL(n1405), .F(n1311) );
  IV U478 ( .A(n1406), .Z(n229) );
  ANDN U479 ( .A(n1883), .B(n1882), .Z(n1674) );
  MUX U480 ( .IN0(n230), .IN1(n1956), .SEL(n1756), .F(n1884) );
  IV U481 ( .A(n1755), .Z(n230) );
  MUX U482 ( .IN0(n231), .IN1(n2388), .SEL(n1780), .F(n2316) );
  IV U483 ( .A(n1779), .Z(n231) );
  MUX U484 ( .IN0(n3957), .IN1(n3974), .SEL(n3958), .F(n3939) );
  MUX U485 ( .IN0(n4334), .IN1(n4345), .SEL(n4335), .F(n4322) );
  MUX U486 ( .IN0(n3515), .IN1(n232), .SEL(n3516), .F(n3475) );
  IV U487 ( .A(n3517), .Z(n232) );
  MUX U488 ( .IN0(n3582), .IN1(n233), .SEL(n3583), .F(n3542) );
  IV U489 ( .A(n3584), .Z(n233) );
  MUX U490 ( .IN0(n3538), .IN1(n234), .SEL(n3539), .F(n3498) );
  IV U491 ( .A(n3540), .Z(n234) );
  MUX U492 ( .IN0(n3964), .IN1(n235), .SEL(n3685), .F(n3946) );
  IV U493 ( .A(n3684), .Z(n235) );
  XNOR U494 ( .A(n4326), .B(n4317), .Z(n3945) );
  MUX U495 ( .IN0(n3913), .IN1(n236), .SEL(n3914), .F(n3895) );
  IV U496 ( .A(n3915), .Z(n236) );
  MUX U497 ( .IN0(n3917), .IN1(n237), .SEL(n3918), .F(n3899) );
  IV U498 ( .A(n3919), .Z(n237) );
  MUX U499 ( .IN0(n3533), .IN1(n238), .SEL(n3534), .F(n3493) );
  IV U500 ( .A(n3535), .Z(n238) );
  XNOR U501 ( .A(n3433), .B(n3396), .Z(n3400) );
  XNOR U502 ( .A(n4290), .B(n4281), .Z(n3891) );
  XNOR U503 ( .A(n3416), .B(n3379), .Z(n3383) );
  MUX U504 ( .IN0(n3849), .IN1(n3866), .SEL(n3850), .F(n3831) );
  XNOR U505 ( .A(n3857), .B(n3842), .Z(n3846) );
  MUX U506 ( .IN0(n4129), .IN1(n239), .SEL(n4130), .F(n4107) );
  IV U507 ( .A(n4131), .Z(n239) );
  MUX U508 ( .IN0(n3279), .IN1(n240), .SEL(n3280), .F(n3239) );
  IV U509 ( .A(n3281), .Z(n240) );
  MUX U510 ( .IN0(n3235), .IN1(n241), .SEL(n3236), .F(n3195) );
  IV U511 ( .A(n3237), .Z(n241) );
  XNOR U512 ( .A(n4254), .B(n4245), .Z(n3837) );
  MUX U513 ( .IN0(n4690), .IN1(n242), .SEL(n4691), .F(n4668) );
  IV U514 ( .A(n4692), .Z(n242) );
  XNOR U515 ( .A(n3296), .B(n3259), .Z(n3263) );
  MUX U516 ( .IN0(n4428), .IN1(n4118), .SEL(n4120), .F(n4416) );
  MUX U517 ( .IN0(n4406), .IN1(n4417), .SEL(n4407), .F(n4394) );
  MUX U518 ( .IN0(n4832), .IN1(n4701), .SEL(n4703), .F(n4820) );
  XNOR U519 ( .A(n3803), .B(n3788), .Z(n3792) );
  MUX U520 ( .IN0(n3178), .IN1(n243), .SEL(n3179), .F(n3138) );
  IV U521 ( .A(n3180), .Z(n243) );
  MUX U522 ( .IN0(n4400), .IN1(n244), .SEL(n4401), .F(n4388) );
  IV U523 ( .A(n4402), .Z(n244) );
  MUX U524 ( .IN0(n4089), .IN1(n4091), .SEL(n4090), .F(n4067) );
  MUX U525 ( .IN0(n4491), .IN1(n245), .SEL(n4492), .F(n4475) );
  IV U526 ( .A(n4493), .Z(n245) );
  MUX U527 ( .IN0(n4900), .IN1(n4905), .SEL(n4901), .F(n4885) );
  MUX U528 ( .IN0(n4895), .IN1(n246), .SEL(n4896), .F(n4879) );
  IV U529 ( .A(n4897), .Z(n246) );
  MUX U530 ( .IN0(n4804), .IN1(n247), .SEL(n4805), .F(n4792) );
  IV U531 ( .A(n4806), .Z(n247) );
  MUX U532 ( .IN0(n4798), .IN1(n4809), .SEL(n4799), .F(n4786) );
  MUX U533 ( .IN0(n3639), .IN1(n248), .SEL(n3640), .F(n3623) );
  IV U534 ( .A(n3641), .Z(n248) );
  XNOR U535 ( .A(n4037), .B(n4038), .Z(n4047) );
  MUX U536 ( .IN0(n4993), .IN1(n249), .SEL(n4994), .F(n4977) );
  IV U537 ( .A(n4995), .Z(n249) );
  MUX U538 ( .IN0(n4650), .IN1(n4652), .SEL(n4651), .F(n4628) );
  MUX U539 ( .IN0(n4212), .IN1(n250), .SEL(n3783), .F(n4200) );
  IV U540 ( .A(n3782), .Z(n250) );
  XNOR U541 ( .A(n4015), .B(n4016), .Z(n4025) );
  XNOR U542 ( .A(n4598), .B(n4599), .Z(n4608) );
  MUX U543 ( .IN0(n3079), .IN1(n251), .SEL(n3080), .F(n3039) );
  IV U544 ( .A(n3081), .Z(n251) );
  MUX U545 ( .IN0(n4196), .IN1(n252), .SEL(n4197), .F(n4184) );
  IV U546 ( .A(n4198), .Z(n252) );
  MUX U547 ( .IN0(n3737), .IN1(n253), .SEL(n3738), .F(n3719) );
  IV U548 ( .A(n3739), .Z(n253) );
  XNOR U549 ( .A(n4374), .B(n4365), .Z(n4010) );
  XNOR U550 ( .A(n3993), .B(n3994), .Z(n4003) );
  MUX U551 ( .IN0(n3997), .IN1(n254), .SEL(n3998), .F(n3967) );
  IV U552 ( .A(n3999), .Z(n254) );
  MUX U553 ( .IN0(n4784), .IN1(n4613), .SEL(n4615), .F(n4772) );
  MUX U554 ( .IN0(n3003), .IN1(n3042), .SEL(n3004), .F(n2964) );
  XNOR U555 ( .A(n3096), .B(n3059), .Z(n3063) );
  MUX U556 ( .IN0(n3697), .IN1(n255), .SEL(n3698), .F(n2973) );
  IV U557 ( .A(n3699), .Z(n255) );
  MUX U558 ( .IN0(n4750), .IN1(n4761), .SEL(n4751), .F(n4543) );
  MUX U559 ( .IN0(n4756), .IN1(n256), .SEL(n4757), .F(n4744) );
  IV U560 ( .A(n4758), .Z(n256) );
  MUX U561 ( .IN0(n4558), .IN1(n4573), .SEL(n4559), .F(n4529) );
  MUX U562 ( .IN0(n2956), .IN1(n257), .SEL(n2957), .F(n2884) );
  IV U563 ( .A(n2958), .Z(n257) );
  MUX U564 ( .IN0(n733), .IN1(n768), .SEL(n734), .F(n700) );
  MUX U565 ( .IN0(n889), .IN1(n942), .SEL(n890), .F(n837) );
  MUX U566 ( .IN0(n898), .IN1(n258), .SEL(n899), .F(n846) );
  IV U567 ( .A(n900), .Z(n258) );
  MUX U568 ( .IN0(n1096), .IN1(n1162), .SEL(n1097), .F(n1029) );
  MUX U569 ( .IN0(n1216), .IN1(n259), .SEL(n1217), .F(n1146) );
  IV U570 ( .A(n1218), .Z(n259) );
  MUX U571 ( .IN0(n1262), .IN1(n1334), .SEL(n1263), .F(n1192) );
  MUX U572 ( .IN0(n1371), .IN1(n260), .SEL(n1372), .F(n1297) );
  IV U573 ( .A(n1373), .Z(n260) );
  MUX U574 ( .IN0(n1523), .IN1(n261), .SEL(n1524), .F(n1437) );
  IV U575 ( .A(n1525), .Z(n261) );
  MUX U576 ( .IN0(n1648), .IN1(n1740), .SEL(n1649), .F(n1558) );
  MUX U577 ( .IN0(n1680), .IN1(n262), .SEL(n1681), .F(n1587) );
  IV U578 ( .A(n1682), .Z(n262) );
  MUX U579 ( .IN0(n1860), .IN1(n263), .SEL(n1861), .F(n1724) );
  IV U580 ( .A(n1862), .Z(n263) );
  MUX U581 ( .IN0(n1989), .IN1(n264), .SEL(n1990), .F(n1917) );
  IV U582 ( .A(n1991), .Z(n264) );
  MUX U583 ( .IN0(n2547), .IN1(n2594), .SEL(n2548), .F(n2516) );
  MUX U584 ( .IN0(n2611), .IN1(n265), .SEL(n2612), .F(n2576) );
  IV U585 ( .A(n2613), .Z(n265) );
  MUX U586 ( .IN0(n2223), .IN1(n266), .SEL(n2224), .F(n2151) );
  IV U587 ( .A(n2225), .Z(n266) );
  MUX U588 ( .IN0(n2277), .IN1(n267), .SEL(n2278), .F(n2205) );
  IV U589 ( .A(n2279), .Z(n267) );
  MUX U590 ( .IN0(n2373), .IN1(n268), .SEL(n2374), .F(n2304) );
  IV U591 ( .A(n2375), .Z(n268) );
  MUX U592 ( .IN0(n2320), .IN1(n269), .SEL(n2321), .F(n2251) );
  IV U593 ( .A(n2322), .Z(n269) );
  MUX U594 ( .IN0(n2751), .IN1(n2842), .SEL(n2752), .F(n2732) );
  MUX U595 ( .IN0(n4938), .IN1(n270), .SEL(n4939), .F(n2439) );
  IV U596 ( .A(n4940), .Z(n270) );
  MUX U597 ( .IN0(n4164), .IN1(n271), .SEL(n3711), .F(n2929) );
  IV U598 ( .A(n3710), .Z(n271) );
  MUX U599 ( .IN0(n765), .IN1(n272), .SEL(n766), .F(n729) );
  IV U600 ( .A(n767), .Z(n272) );
  MUX U601 ( .IN0(n1016), .IN1(n273), .SEL(n1017), .F(n958) );
  IV U602 ( .A(n1018), .Z(n273) );
  MUX U603 ( .IN0(n983), .IN1(n274), .SEL(n984), .F(n926) );
  IV U604 ( .A(n985), .Z(n274) );
  MUX U605 ( .IN0(n1112), .IN1(n275), .SEL(n1113), .F(n1045) );
  IV U606 ( .A(n1114), .Z(n275) );
  MUX U607 ( .IN0(n1292), .IN1(n276), .SEL(n1293), .F(n1220) );
  IV U608 ( .A(n1294), .Z(n276) );
  MUX U609 ( .IN0(n1348), .IN1(n277), .SEL(n1349), .F(n1274) );
  IV U610 ( .A(n1350), .Z(n277) );
  MUX U611 ( .IN0(n1635), .IN1(n278), .SEL(n1636), .F(n1545) );
  IV U612 ( .A(n1637), .Z(n278) );
  MUX U613 ( .IN0(n1710), .IN1(n279), .SEL(n1711), .F(n1617) );
  IV U614 ( .A(n1712), .Z(n279) );
  MUX U615 ( .IN0(n1804), .IN1(n280), .SEL(n1805), .F(n1663) );
  IV U616 ( .A(n1806), .Z(n280) );
  MUX U617 ( .IN0(n2080), .IN1(n281), .SEL(n2081), .F(n2011) );
  IV U618 ( .A(n2082), .Z(n281) );
  MUX U619 ( .IN0(n2137), .IN1(n282), .SEL(n2138), .F(n2062) );
  IV U620 ( .A(n2139), .Z(n282) );
  MUX U621 ( .IN0(n2658), .IN1(n283), .SEL(n2659), .F(n2615) );
  IV U622 ( .A(n2660), .Z(n283) );
  MUX U623 ( .IN0(n2368), .IN1(n284), .SEL(n2369), .F(n2299) );
  IV U624 ( .A(n2370), .Z(n284) );
  MUX U625 ( .IN0(n2791), .IN1(n285), .SEL(n2792), .F(n2714) );
  IV U626 ( .A(n2793), .Z(n285) );
  MUX U627 ( .IN0(n2452), .IN1(n286), .SEL(n2453), .F(n2377) );
  IV U628 ( .A(n2454), .Z(n286) );
  MUX U629 ( .IN0(n2425), .IN1(n287), .SEL(n2426), .F(n2350) );
  IV U630 ( .A(n2427), .Z(n287) );
  MUX U631 ( .IN0(n2879), .IN1(n288), .SEL(n2880), .F(n2815) );
  IV U632 ( .A(n2881), .Z(n288) );
  MUX U633 ( .IN0(n2906), .IN1(n289), .SEL(n2907), .F(n2839) );
  IV U634 ( .A(n2908), .Z(n289) );
  XNOR U635 ( .A(n4548), .B(n4522), .Z(n4526) );
  MUX U636 ( .IN0(n640), .IN1(n290), .SEL(n641), .F(n621) );
  IV U637 ( .A(n642), .Z(n290) );
  MUX U638 ( .IN0(n719), .IN1(n753), .SEL(n721), .F(n681) );
  MUX U639 ( .IN0(n841), .IN1(n291), .SEL(n842), .F(n787) );
  IV U640 ( .A(n843), .Z(n291) );
  XNOR U641 ( .A(n961), .B(n908), .Z(n912) );
  XNOR U642 ( .A(n1223), .B(n1156), .Z(n1160) );
  MUX U643 ( .IN0(n1266), .IN1(n292), .SEL(n1267), .F(n1196) );
  IV U644 ( .A(n1268), .Z(n292) );
  MUX U645 ( .IN0(n1357), .IN1(n293), .SEL(n1358), .F(n1283) );
  IV U646 ( .A(n1359), .Z(n293) );
  XNOR U647 ( .A(n1409), .B(n1319), .Z(n1323) );
  XNOR U648 ( .A(n1638), .B(n1551), .Z(n1555) );
  MUX U649 ( .IN0(n1719), .IN1(n294), .SEL(n1720), .F(n1626) );
  IV U650 ( .A(n1721), .Z(n294) );
  MUX U651 ( .IN0(n1837), .IN1(n295), .SEL(n1838), .F(n1701) );
  IV U652 ( .A(n1839), .Z(n295) );
  MUX U653 ( .IN0(n2471), .IN1(n2500), .SEL(n2473), .F(n1787) );
  XNOR U654 ( .A(n1942), .B(n1870), .Z(n1874) );
  XNOR U655 ( .A(n2585), .B(n2540), .Z(n2544) );
  MUX U656 ( .IN0(n2571), .IN1(n296), .SEL(n2572), .F(n2526) );
  IV U657 ( .A(n2573), .Z(n296) );
  XNOR U658 ( .A(n2158), .B(n2086), .Z(n2090) );
  MUX U659 ( .IN0(n2146), .IN1(n297), .SEL(n2147), .F(n2071) );
  IV U660 ( .A(n2148), .Z(n297) );
  XNOR U661 ( .A(n2105), .B(n2033), .Z(n2037) );
  MUX U662 ( .IN0(n2200), .IN1(n298), .SEL(n2201), .F(n2128) );
  IV U663 ( .A(n2202), .Z(n298) );
  XNOR U664 ( .A(n2723), .B(n2677), .Z(n2680) );
  MUX U665 ( .IN0(n299), .IN1(n2764), .SEL(n2765), .F(n2736) );
  IV U666 ( .A(n2766), .Z(n299) );
  MUX U667 ( .IN0(n2806), .IN1(n300), .SEL(n2807), .F(n2773) );
  IV U668 ( .A(n2808), .Z(n300) );
  MUX U669 ( .IN0(n4928), .IN1(n301), .SEL(n4538), .F(n2434) );
  IV U670 ( .A(n4537), .Z(n301) );
  ANDN U671 ( .A(n617), .B(n618), .Z(n610) );
  MUX U672 ( .IN0(n302), .IN1(n998), .SEL(n999), .F(n937) );
  IV U673 ( .A(n1000), .Z(n302) );
  MUX U674 ( .IN0(n1053), .IN1(n303), .SEL(n1054), .F(n995) );
  IV U675 ( .A(n1055), .Z(n303) );
  MUX U676 ( .IN0(n1423), .IN1(n304), .SEL(n1424), .F(n1330) );
  IV U677 ( .A(n1425), .Z(n304) );
  MUX U678 ( .IN0(n1903), .IN1(n305), .SEL(n1904), .F(n1828) );
  IV U679 ( .A(n1905), .Z(n305) );
  MUX U680 ( .IN0(n2263), .IN1(n306), .SEL(n2264), .F(n2191) );
  IV U681 ( .A(n2265), .Z(n306) );
  MUX U682 ( .IN0(n307), .IN1(n2739), .SEL(n2387), .F(n2689) );
  IV U683 ( .A(n2386), .Z(n307) );
  XNOR U684 ( .A(n778), .B(n828), .Z(n817) );
  AND U685 ( .A(n1399), .B(n1400), .Z(n1398) );
  MUX U686 ( .IN0(n308), .IN1(n1671), .SEL(n1672), .F(n1578) );
  IV U687 ( .A(n1673), .Z(n308) );
  ANDN U688 ( .A(n1959), .B(n1958), .Z(n1887) );
  MUX U689 ( .IN0(n309), .IN1(n2100), .SEL(n1764), .F(n2028) );
  IV U690 ( .A(n1763), .Z(n309) );
  MUX U691 ( .IN0(n310), .IN1(n2460), .SEL(n2461), .F(n2388) );
  IV U692 ( .A(n2462), .Z(n310) );
  MUX U693 ( .IN0(n628), .IN1(o_reg[29]), .SEL(n629), .F(n595) );
  AND U694 ( .A(n739), .B(n740), .Z(n706) );
  MUX U695 ( .IN0(n919), .IN1(o_reg[21]), .SEL(n920), .F(n869) );
  ANDN U696 ( .A(n1169), .B(n1170), .Z(n1102) );
  MUX U697 ( .IN0(o_reg[15]), .IN1(n1309), .SEL(n1310), .F(n1237) );
  MUX U698 ( .IN0(n1745), .IN1(o_reg[10]), .SEL(n579), .F(n1652) );
  MUX U699 ( .IN0(o_reg[4]), .IN1(n1769), .SEL(n585), .F(n1765) );
  MUX U700 ( .IN0(n4340), .IN1(n311), .SEL(n4341), .F(n4328) );
  IV U701 ( .A(n4342), .Z(n311) );
  MUX U702 ( .IN0(n3931), .IN1(n312), .SEL(n3932), .F(n3913) );
  IV U703 ( .A(n3933), .Z(n312) );
  XNOR U704 ( .A(n3553), .B(n3516), .Z(n3520) );
  MUX U705 ( .IN0(n4322), .IN1(n4333), .SEL(n4323), .F(n4310) );
  MUX U706 ( .IN0(n3483), .IN1(n3522), .SEL(n3484), .F(n3443) );
  MUX U707 ( .IN0(n3489), .IN1(n3528), .SEL(n3490), .F(n3449) );
  MUX U708 ( .IN0(n3542), .IN1(n313), .SEL(n3543), .F(n3502) );
  IV U709 ( .A(n3544), .Z(n313) );
  MUX U710 ( .IN0(n3498), .IN1(n314), .SEL(n3499), .F(n3458) );
  IV U711 ( .A(n3500), .Z(n314) );
  MUX U712 ( .IN0(n3946), .IN1(n315), .SEL(n3551), .F(n3928) );
  IV U713 ( .A(n3549), .Z(n315) );
  MUX U714 ( .IN0(n4308), .IN1(n316), .SEL(n3927), .F(n4296) );
  IV U715 ( .A(n3926), .Z(n316) );
  MUX U716 ( .IN0(n3899), .IN1(n317), .SEL(n3900), .F(n3881) );
  IV U717 ( .A(n3901), .Z(n317) );
  MUX U718 ( .IN0(n3493), .IN1(n318), .SEL(n3494), .F(n3453) );
  IV U719 ( .A(n3495), .Z(n318) );
  MUX U720 ( .IN0(n4292), .IN1(n319), .SEL(n4293), .F(n4280) );
  IV U721 ( .A(n4294), .Z(n319) );
  MUX U722 ( .IN0(n3859), .IN1(n320), .SEL(n3860), .F(n3841) );
  IV U723 ( .A(n3861), .Z(n320) );
  XNOR U724 ( .A(n3393), .B(n3356), .Z(n3360) );
  MUX U725 ( .IN0(n3323), .IN1(n3362), .SEL(n3324), .F(n3283) );
  MUX U726 ( .IN0(n3329), .IN1(n3368), .SEL(n3330), .F(n3289) );
  MUX U727 ( .IN0(n3382), .IN1(n321), .SEL(n3383), .F(n3342) );
  IV U728 ( .A(n3384), .Z(n321) );
  MUX U729 ( .IN0(n3874), .IN1(n322), .SEL(n3391), .F(n3856) );
  IV U730 ( .A(n3389), .Z(n322) );
  MUX U731 ( .IN0(n3298), .IN1(n323), .SEL(n3299), .F(n3258) );
  IV U732 ( .A(n3300), .Z(n323) );
  MUX U733 ( .IN0(n4834), .IN1(n4845), .SEL(n4835), .F(n4822) );
  MUX U734 ( .IN0(n4260), .IN1(n324), .SEL(n3855), .F(n4248) );
  IV U735 ( .A(n3854), .Z(n324) );
  MUX U736 ( .IN0(n3827), .IN1(n325), .SEL(n3828), .F(n3809) );
  IV U737 ( .A(n3829), .Z(n325) );
  MUX U738 ( .IN0(n3333), .IN1(n326), .SEL(n3334), .F(n3293) );
  IV U739 ( .A(n3335), .Z(n326) );
  MUX U740 ( .IN0(n4828), .IN1(n327), .SEL(n4829), .F(n4816) );
  IV U741 ( .A(n4830), .Z(n327) );
  MUX U742 ( .IN0(n3239), .IN1(n328), .SEL(n3240), .F(n3199) );
  IV U743 ( .A(n3241), .Z(n328) );
  MUX U744 ( .IN0(n3195), .IN1(n329), .SEL(n3196), .F(n3155) );
  IV U745 ( .A(n3197), .Z(n329) );
  MUX U746 ( .IN0(n4244), .IN1(n330), .SEL(n4245), .F(n4232) );
  IV U747 ( .A(n4246), .Z(n330) );
  MUX U748 ( .IN0(n3787), .IN1(n331), .SEL(n3788), .F(n3769) );
  IV U749 ( .A(n3789), .Z(n331) );
  XNOR U750 ( .A(n4127), .B(n4108), .Z(n4112) );
  XNOR U751 ( .A(n4081), .B(n4082), .Z(n4091) );
  MUX U752 ( .IN0(n4694), .IN1(n4696), .SEL(n4695), .F(n4672) );
  MUX U753 ( .IN0(n4668), .IN1(n332), .SEL(n4669), .F(n4646) );
  IV U754 ( .A(n4670), .Z(n332) );
  MUX U755 ( .IN0(n3163), .IN1(n3202), .SEL(n3164), .F(n3123) );
  MUX U756 ( .IN0(n3777), .IN1(n3794), .SEL(n3778), .F(n3759) );
  MUX U757 ( .IN0(n3169), .IN1(n3208), .SEL(n3170), .F(n3129) );
  MUX U758 ( .IN0(n3222), .IN1(n333), .SEL(n3223), .F(n3182) );
  IV U759 ( .A(n3224), .Z(n333) );
  XNOR U760 ( .A(n4410), .B(n4401), .Z(n4076) );
  XNOR U761 ( .A(n4059), .B(n4060), .Z(n4069) );
  MUX U762 ( .IN0(n4063), .IN1(n334), .SEL(n4064), .F(n4041) );
  IV U763 ( .A(n4065), .Z(n334) );
  MUX U764 ( .IN0(n4640), .IN1(n4661), .SEL(n4641), .F(n4618) );
  MUX U765 ( .IN0(n3802), .IN1(n335), .SEL(n3231), .F(n3784) );
  IV U766 ( .A(n3229), .Z(n335) );
  MUX U767 ( .IN0(n3138), .IN1(n336), .SEL(n3139), .F(n3098) );
  IV U768 ( .A(n3140), .Z(n336) );
  MUX U769 ( .IN0(n4382), .IN1(n4393), .SEL(n4383), .F(n4370) );
  MUX U770 ( .IN0(n4500), .IN1(n4157), .SEL(n4158), .F(n4485) );
  MUX U771 ( .IN0(n4475), .IN1(n4490), .SEL(n4477), .F(n4459) );
  MUX U772 ( .IN0(n4904), .IN1(n4740), .SEL(n4741), .F(n4889) );
  MUX U773 ( .IN0(n4879), .IN1(n4894), .SEL(n4881), .F(n4863) );
  MUX U774 ( .IN0(n4808), .IN1(n4657), .SEL(n4659), .F(n4796) );
  MUX U775 ( .IN0(n4786), .IN1(n4797), .SEL(n4787), .F(n4774) );
  MUX U776 ( .IN0(n3173), .IN1(n337), .SEL(n3174), .F(n3133) );
  IV U777 ( .A(n3175), .Z(n337) );
  MUX U778 ( .IN0(n3648), .IN1(n3592), .SEL(n3593), .F(n3633) );
  MUX U779 ( .IN0(n3623), .IN1(n3638), .SEL(n3625), .F(n3607) );
  MUX U780 ( .IN0(n5002), .IN1(n4934), .SEL(n4935), .F(n4987) );
  MUX U781 ( .IN0(n4780), .IN1(n338), .SEL(n4781), .F(n4768) );
  IV U782 ( .A(n4782), .Z(n338) );
  MUX U783 ( .IN0(n4200), .IN1(n339), .SEL(n3765), .F(n4188) );
  IV U784 ( .A(n3764), .Z(n339) );
  XNOR U785 ( .A(n3749), .B(n3734), .Z(n3738) );
  XOR U786 ( .A(n3081), .B(n3080), .Z(n3095) );
  MUX U787 ( .IN0(n4178), .IN1(n4189), .SEL(n4179), .F(n4166) );
  XNOR U788 ( .A(n4622), .B(n4603), .Z(n4607) );
  XNOR U789 ( .A(n4576), .B(n4577), .Z(n4586) );
  MUX U790 ( .IN0(n4184), .IN1(n340), .SEL(n4185), .F(n4172) );
  IV U791 ( .A(n4186), .Z(n340) );
  MUX U792 ( .IN0(n3705), .IN1(n3722), .SEL(n3706), .F(n2981) );
  MUX U793 ( .IN0(n3009), .IN1(n3048), .SEL(n3010), .F(n2938) );
  MUX U794 ( .IN0(n4368), .IN1(n4008), .SEL(n4010), .F(n4356) );
  XNOR U795 ( .A(n4017), .B(n3998), .Z(n4002) );
  XNOR U796 ( .A(n3977), .B(n3978), .Z(n3973) );
  MUX U797 ( .IN0(n5029), .IN1(n5032), .SEL(n5030), .F(n5022) );
  MUX U798 ( .IN0(n4944), .IN1(n4966), .SEL(n4946), .F(n4924) );
  XNOR U799 ( .A(n4560), .B(n4561), .Z(n4556) );
  MUX U800 ( .IN0(n4550), .IN1(n341), .SEL(n4551), .F(n4521) );
  IV U801 ( .A(n4552), .Z(n341) );
  MUX U802 ( .IN0(n2964), .IN1(n3002), .SEL(n2965), .F(n2892) );
  MUX U803 ( .IN0(n2999), .IN1(n342), .SEL(n3000), .F(n2960) );
  IV U804 ( .A(n3001), .Z(n342) );
  MUX U805 ( .IN0(n3730), .IN1(n343), .SEL(n3071), .F(n3712) );
  IV U806 ( .A(n3069), .Z(n343) );
  XNOR U807 ( .A(n3056), .B(n3019), .Z(n3023) );
  MUX U808 ( .IN0(n783), .IN1(n836), .SEL(n784), .F(n746) );
  MUX U809 ( .IN0(n915), .IN1(n970), .SEL(n916), .F(n865) );
  MUX U810 ( .IN0(n963), .IN1(n344), .SEL(n964), .F(n907) );
  IV U811 ( .A(n965), .Z(n344) );
  MUX U812 ( .IN0(n1079), .IN1(n345), .SEL(n1080), .F(n1012) );
  IV U813 ( .A(n1081), .Z(n345) );
  MUX U814 ( .IN0(n1225), .IN1(n346), .SEL(n1226), .F(n1155) );
  IV U815 ( .A(n1227), .Z(n346) );
  MUX U816 ( .IN0(n1183), .IN1(n1252), .SEL(n1184), .F(n1116) );
  MUX U817 ( .IN0(n1379), .IN1(n1471), .SEL(n1380), .F(n1305) );
  MUX U818 ( .IN0(n1318), .IN1(n347), .SEL(n1319), .F(n1245) );
  IV U819 ( .A(n1320), .Z(n347) );
  MUX U820 ( .IN0(n1335), .IN1(n1427), .SEL(n1336), .F(n1262) );
  MUX U821 ( .IN0(n1344), .IN1(n348), .SEL(n1345), .F(n1270) );
  IV U822 ( .A(n1346), .Z(n348) );
  MUX U823 ( .IN0(n1505), .IN1(n1594), .SEL(n1506), .F(n1419) );
  MUX U824 ( .IN0(n1741), .IN1(n1876), .SEL(n1742), .F(n1648) );
  MUX U825 ( .IN0(n1706), .IN1(n349), .SEL(n1707), .F(n1613) );
  IV U826 ( .A(n1708), .Z(n349) );
  MUX U827 ( .IN0(n1899), .IN1(n1970), .SEL(n1900), .F(n1824) );
  MUX U828 ( .IN0(n2007), .IN1(n350), .SEL(n2008), .F(n1935) );
  IV U829 ( .A(n2009), .Z(n350) );
  MUX U830 ( .IN0(n2058), .IN1(n351), .SEL(n2059), .F(n1989) );
  IV U831 ( .A(n2060), .Z(n351) );
  MUX U832 ( .IN0(n2587), .IN1(n352), .SEL(n2588), .F(n2539) );
  IV U833 ( .A(n2589), .Z(n352) );
  MUX U834 ( .IN0(n2187), .IN1(n2258), .SEL(n2188), .F(n2115) );
  MUX U835 ( .IN0(n2295), .IN1(n353), .SEL(n2296), .F(n2223) );
  IV U836 ( .A(n2297), .Z(n353) );
  MUX U837 ( .IN0(n2718), .IN1(n2794), .SEL(n2719), .F(n2671) );
  MUX U838 ( .IN0(n2381), .IN1(n2455), .SEL(n2382), .F(n2312) );
  MUX U839 ( .IN0(n2778), .IN1(n354), .SEL(n2779), .F(n2701) );
  IV U840 ( .A(n2780), .Z(n354) );
  MUX U841 ( .IN0(n2820), .IN1(n355), .SEL(n2821), .F(n2787) );
  IV U842 ( .A(n2822), .Z(n355) );
  XNOR U843 ( .A(n3695), .B(n2974), .Z(n2978) );
  MUX U844 ( .IN0(n852), .IN1(n356), .SEL(n853), .F(n795) );
  IV U845 ( .A(n854), .Z(n356) );
  MUX U846 ( .IN0(n1092), .IN1(n357), .SEL(n1093), .F(n1025) );
  IV U847 ( .A(n1094), .Z(n357) );
  MUX U848 ( .IN0(n1150), .IN1(n358), .SEL(n1151), .F(n1083) );
  IV U849 ( .A(n1152), .Z(n358) );
  MUX U850 ( .IN0(n1808), .IN1(n2486), .SEL(n1809), .F(n1667) );
  MUX U851 ( .IN0(n1527), .IN1(n359), .SEL(n1528), .F(n1441) );
  IV U852 ( .A(n1529), .Z(n359) );
  MUX U853 ( .IN0(n1864), .IN1(n360), .SEL(n1865), .F(n1728) );
  IV U854 ( .A(n1866), .Z(n360) );
  MUX U855 ( .IN0(n1921), .IN1(n361), .SEL(n1922), .F(n1846) );
  IV U856 ( .A(n1923), .Z(n361) );
  MUX U857 ( .IN0(n2732), .IN1(n2750), .SEL(n2733), .F(n2683) );
  MUX U858 ( .IN0(n2582), .IN1(n362), .SEL(n2583), .F(n2534) );
  IV U859 ( .A(n2584), .Z(n362) );
  MUX U860 ( .IN0(n2155), .IN1(n363), .SEL(n2156), .F(n2080) );
  IV U861 ( .A(n2157), .Z(n363) );
  MUX U862 ( .IN0(n2209), .IN1(n364), .SEL(n2210), .F(n2137) );
  IV U863 ( .A(n2211), .Z(n364) );
  MUX U864 ( .IN0(n2443), .IN1(n365), .SEL(n2444), .F(n2368) );
  IV U865 ( .A(n2445), .Z(n365) );
  MUX U866 ( .IN0(n2815), .IN1(n366), .SEL(n2816), .F(n2782) );
  IV U867 ( .A(n2817), .Z(n366) );
  MUX U868 ( .IN0(n4748), .IN1(n367), .SEL(n4564), .F(n2425) );
  IV U869 ( .A(n4563), .Z(n367) );
  MUX U870 ( .IN0(n2929), .IN1(n368), .SEL(n2930), .F(n2855) );
  IV U871 ( .A(n2931), .Z(n368) );
  XNOR U872 ( .A(n658), .B(n638), .Z(n641) );
  XNOR U873 ( .A(n798), .B(n762), .Z(n766) );
  MUX U874 ( .IN0(n893), .IN1(n369), .SEL(n894), .F(n841) );
  IV U875 ( .A(n895), .Z(n369) );
  MUX U876 ( .IN0(n1211), .IN1(n370), .SEL(n1212), .F(n1141) );
  IV U877 ( .A(n1213), .Z(n370) );
  XNOR U878 ( .A(n1173), .B(n1109), .Z(n1113) );
  MUX U879 ( .IN0(n1196), .IN1(n371), .SEL(n1197), .F(n1128) );
  IV U880 ( .A(n1198), .Z(n371) );
  XNOR U881 ( .A(n1453), .B(n1363), .Z(n1367) );
  XNOR U882 ( .A(n1548), .B(n1465), .Z(n1469) );
  XNOR U883 ( .A(n1585), .B(n1498), .Z(n1502) );
  MUX U884 ( .IN0(n1701), .IN1(n372), .SEL(n1702), .F(n1608) );
  IV U885 ( .A(n1703), .Z(n372) );
  XNOR U886 ( .A(n1867), .B(n1734), .Z(n1738) );
  XNOR U887 ( .A(n2475), .B(n1801), .Z(n1805) );
  MUX U888 ( .IN0(n2468), .IN1(n373), .SEL(n2469), .F(n1793) );
  IV U889 ( .A(n2470), .Z(n373) );
  MUX U890 ( .IN0(n1930), .IN1(n374), .SEL(n1931), .F(n1855) );
  IV U891 ( .A(n1932), .Z(n374) );
  XNOR U892 ( .A(n1889), .B(n1817), .Z(n1821) );
  MUX U893 ( .IN0(n2606), .IN1(n375), .SEL(n2607), .F(n2571) );
  IV U894 ( .A(n2608), .Z(n375) );
  XNOR U895 ( .A(n2230), .B(n2161), .Z(n2165) );
  XNOR U896 ( .A(n2177), .B(n2108), .Z(n2112) );
  MUX U897 ( .IN0(n2290), .IN1(n376), .SEL(n2291), .F(n2218) );
  IV U898 ( .A(n2292), .Z(n376) );
  MUX U899 ( .IN0(n2272), .IN1(n377), .SEL(n2273), .F(n2200) );
  IV U900 ( .A(n2274), .Z(n377) );
  XNOR U901 ( .A(n2708), .B(n2664), .Z(n2668) );
  XNOR U902 ( .A(n2741), .B(n2725), .Z(n2729) );
  XNOR U903 ( .A(n2446), .B(n2374), .Z(n2378) );
  XNOR U904 ( .A(n2393), .B(n2321), .Z(n2325) );
  MUX U905 ( .IN0(n2852), .IN1(n378), .SEL(n2853), .F(n2764) );
  IV U906 ( .A(n2854), .Z(n378) );
  MUX U907 ( .IN0(n2870), .IN1(n379), .SEL(n2871), .F(n2806) );
  IV U908 ( .A(n2872), .Z(n379) );
  MUX U909 ( .IN0(n644), .IN1(n666), .SEL(n645), .F(n624) );
  MUX U910 ( .IN0(n380), .IN1(n655), .SEL(n656), .F(n636) );
  IV U911 ( .A(n657), .Z(n380) );
  XOR U912 ( .A(n930), .B(n929), .Z(n936) );
  MUX U913 ( .IN0(n1257), .IN1(n381), .SEL(n1258), .F(n1187) );
  IV U914 ( .A(n1259), .Z(n381) );
  XNOR U915 ( .A(n1395), .B(n1396), .Z(n1401) );
  MUX U916 ( .IN0(n1599), .IN1(n382), .SEL(n1600), .F(n1509) );
  IV U917 ( .A(n1601), .Z(n382) );
  XOR U918 ( .A(n1572), .B(n1571), .Z(n1565) );
  MUX U919 ( .IN0(n1975), .IN1(n383), .SEL(n1976), .F(n1903) );
  IV U920 ( .A(n1977), .Z(n383) );
  MUX U921 ( .IN0(n2799), .IN1(n384), .SEL(n2391), .F(n2739) );
  IV U922 ( .A(n2390), .Z(n384) );
  MUX U923 ( .IN0(n2407), .IN1(n385), .SEL(n2408), .F(n2332) );
  IV U924 ( .A(n2409), .Z(n385) );
  XOR U925 ( .A(n951), .B(n950), .Z(n940) );
  MUX U926 ( .IN0(n1488), .IN1(n386), .SEL(n1489), .F(n1404) );
  IV U927 ( .A(n1490), .Z(n386) );
  AND U928 ( .A(n1674), .B(n1675), .Z(n1581) );
  MUX U929 ( .IN0(n387), .IN1(n1884), .SEL(n1752), .F(n1812) );
  IV U930 ( .A(n1751), .Z(n387) );
  MUX U931 ( .IN0(n388), .IN1(n2551), .SEL(n2099), .F(n1959) );
  IV U932 ( .A(n2098), .Z(n388) );
  MUX U933 ( .IN0(n389), .IN1(n2172), .SEL(n1768), .F(n2100) );
  IV U934 ( .A(n1767), .Z(n389) );
  MUX U935 ( .IN0(n390), .IN1(n2896), .SEL(n2897), .F(n2460) );
  IV U936 ( .A(n2898), .Z(n390) );
  MUX U937 ( .IN0(o_reg[27]), .IN1(n671), .SEL(n672), .F(n648) );
  AND U938 ( .A(n814), .B(n815), .Z(n775) );
  AND U939 ( .A(n1035), .B(n1036), .Z(n977) );
  MUX U940 ( .IN0(n1167), .IN1(o_reg[17]), .SEL(n1168), .F(n1100) );
  MUX U941 ( .IN0(n1562), .IN1(o_reg[12]), .SEL(n1563), .F(n1476) );
  MUX U942 ( .IN0(o_reg[8]), .IN1(n1753), .SEL(n581), .F(n1749) );
  MUX U943 ( .IN0(n1773), .IN1(o_reg[3]), .SEL(n615), .F(n1769) );
  MUX U944 ( .IN0(n3563), .IN1(n3680), .SEL(n3564), .F(n3523) );
  MUX U945 ( .IN0(n3939), .IN1(n3956), .SEL(n3940), .F(n3921) );
  MUX U946 ( .IN0(n3529), .IN1(n3568), .SEL(n3530), .F(n3489) );
  MUX U947 ( .IN0(n4328), .IN1(n391), .SEL(n4329), .F(n4316) );
  IV U948 ( .A(n4330), .Z(n391) );
  MUX U949 ( .IN0(n3573), .IN1(n392), .SEL(n3574), .F(n3533) );
  IV U950 ( .A(n3575), .Z(n392) );
  MUX U951 ( .IN0(n3479), .IN1(n393), .SEL(n3480), .F(n3439) );
  IV U952 ( .A(n3481), .Z(n393) );
  MUX U953 ( .IN0(n3458), .IN1(n394), .SEL(n3459), .F(n3418) );
  IV U954 ( .A(n3460), .Z(n394) );
  MUX U955 ( .IN0(n3403), .IN1(n3442), .SEL(n3404), .F(n3363) );
  MUX U956 ( .IN0(n3395), .IN1(n395), .SEL(n3396), .F(n3355) );
  IV U957 ( .A(n3397), .Z(n395) );
  MUX U958 ( .IN0(n3928), .IN1(n396), .SEL(n3511), .F(n3910) );
  IV U959 ( .A(n3509), .Z(n396) );
  MUX U960 ( .IN0(n3462), .IN1(n397), .SEL(n3463), .F(n3422) );
  IV U961 ( .A(n3464), .Z(n397) );
  MUX U962 ( .IN0(n4296), .IN1(n398), .SEL(n3909), .F(n4284) );
  IV U963 ( .A(n3908), .Z(n398) );
  MUX U964 ( .IN0(n3867), .IN1(n3884), .SEL(n3868), .F(n3849) );
  MUX U965 ( .IN0(n3881), .IN1(n399), .SEL(n3882), .F(n3863) );
  IV U966 ( .A(n3883), .Z(n399) );
  MUX U967 ( .IN0(n4274), .IN1(n4285), .SEL(n4275), .F(n4262) );
  MUX U968 ( .IN0(n4280), .IN1(n400), .SEL(n4281), .F(n4268) );
  IV U969 ( .A(n4282), .Z(n400) );
  MUX U970 ( .IN0(n3841), .IN1(n401), .SEL(n3842), .F(n3823) );
  IV U971 ( .A(n3843), .Z(n401) );
  MUX U972 ( .IN0(n3413), .IN1(n402), .SEL(n3414), .F(n3373) );
  IV U973 ( .A(n3415), .Z(n402) );
  XNOR U974 ( .A(n3313), .B(n3276), .Z(n3280) );
  MUX U975 ( .IN0(n4123), .IN1(n4154), .SEL(n4124), .F(n4101) );
  MUX U976 ( .IN0(n4436), .IN1(n403), .SEL(n4437), .F(n4424) );
  IV U977 ( .A(n4438), .Z(n403) );
  MUX U978 ( .IN0(n4430), .IN1(n4441), .SEL(n4431), .F(n4418) );
  MUX U979 ( .IN0(n4840), .IN1(n404), .SEL(n4841), .F(n4828) );
  IV U980 ( .A(n4842), .Z(n404) );
  MUX U981 ( .IN0(n4706), .IN1(n4737), .SEL(n4707), .F(n4684) );
  MUX U982 ( .IN0(n3243), .IN1(n3282), .SEL(n3244), .F(n3203) );
  MUX U983 ( .IN0(n3856), .IN1(n405), .SEL(n3351), .F(n3838) );
  IV U984 ( .A(n3349), .Z(n405) );
  MUX U985 ( .IN0(n3302), .IN1(n406), .SEL(n3303), .F(n3262) );
  IV U986 ( .A(n3304), .Z(n406) );
  MUX U987 ( .IN0(n4822), .IN1(n4833), .SEL(n4823), .F(n4810) );
  MUX U988 ( .IN0(n4248), .IN1(n407), .SEL(n3837), .F(n4236) );
  IV U989 ( .A(n3836), .Z(n407) );
  MUX U990 ( .IN0(n3795), .IN1(n3812), .SEL(n3796), .F(n3777) );
  MUX U991 ( .IN0(n3809), .IN1(n408), .SEL(n3810), .F(n3791) );
  IV U992 ( .A(n3811), .Z(n408) );
  MUX U993 ( .IN0(n409), .IN1(n4136), .SEL(n3687), .F(n4114) );
  IV U994 ( .A(n3686), .Z(n409) );
  MUX U995 ( .IN0(n4226), .IN1(n4237), .SEL(n4227), .F(n4214) );
  MUX U996 ( .IN0(n410), .IN1(n4719), .SEL(n4540), .F(n4697) );
  IV U997 ( .A(n4539), .Z(n410) );
  MUX U998 ( .IN0(n4232), .IN1(n411), .SEL(n4233), .F(n4220) );
  IV U999 ( .A(n4234), .Z(n411) );
  MUX U1000 ( .IN0(n3769), .IN1(n412), .SEL(n3770), .F(n3751) );
  IV U1001 ( .A(n3771), .Z(n412) );
  MUX U1002 ( .IN0(n3253), .IN1(n413), .SEL(n3254), .F(n3213) );
  IV U1003 ( .A(n3255), .Z(n413) );
  XNOR U1004 ( .A(n3193), .B(n3156), .Z(n3160) );
  MUX U1005 ( .IN0(n4416), .IN1(n4096), .SEL(n4098), .F(n4404) );
  MUX U1006 ( .IN0(n4496), .IN1(n4501), .SEL(n4497), .F(n4481) );
  XNOR U1007 ( .A(n4688), .B(n4669), .Z(n4673) );
  XNOR U1008 ( .A(n4814), .B(n4805), .Z(n4659) );
  XNOR U1009 ( .A(n4642), .B(n4643), .Z(n4652) );
  MUX U1010 ( .IN0(n3644), .IN1(n3649), .SEL(n3645), .F(n3629) );
  MUX U1011 ( .IN0(n4035), .IN1(n4056), .SEL(n4036), .F(n4013) );
  MUX U1012 ( .IN0(n4388), .IN1(n414), .SEL(n4389), .F(n4376) );
  IV U1013 ( .A(n4390), .Z(n414) );
  XNOR U1014 ( .A(n4083), .B(n4064), .Z(n4068) );
  MUX U1015 ( .IN0(n4510), .IN1(n4515), .SEL(n4511), .F(n4506) );
  MUX U1016 ( .IN0(n4885), .IN1(n4899), .SEL(n4887), .F(n4869) );
  MUX U1017 ( .IN0(n4914), .IN1(n4919), .SEL(n4915), .F(n4910) );
  XNOR U1018 ( .A(n4620), .B(n4621), .Z(n4630) );
  MUX U1019 ( .IN0(n3083), .IN1(n3122), .SEL(n3084), .F(n3043) );
  MUX U1020 ( .IN0(n3784), .IN1(n415), .SEL(n3191), .F(n3766) );
  IV U1021 ( .A(n3189), .Z(n415) );
  MUX U1022 ( .IN0(n3142), .IN1(n416), .SEL(n3143), .F(n3102) );
  IV U1023 ( .A(n3144), .Z(n416) );
  MUX U1024 ( .IN0(n3658), .IN1(n3663), .SEL(n3659), .F(n3654) );
  XNOR U1025 ( .A(n4384), .B(n4385), .Z(n4052) );
  MUX U1026 ( .IN0(n4146), .IN1(n4151), .SEL(n4147), .F(n4142) );
  MUX U1027 ( .IN0(n4983), .IN1(n4997), .SEL(n4985), .F(n4967) );
  MUX U1028 ( .IN0(n5012), .IN1(n5017), .SEL(n5013), .F(n5008) );
  MUX U1029 ( .IN0(n4729), .IN1(n4734), .SEL(n4730), .F(n4725) );
  XNOR U1030 ( .A(n4788), .B(n4789), .Z(n4635) );
  MUX U1031 ( .IN0(n4602), .IN1(n417), .SEL(n4603), .F(n4580) );
  IV U1032 ( .A(n4604), .Z(n417) );
  XNOR U1033 ( .A(n4194), .B(n4185), .Z(n3747) );
  MUX U1034 ( .IN0(n3723), .IN1(n3740), .SEL(n3724), .F(n3705) );
  MUX U1035 ( .IN0(n3058), .IN1(n418), .SEL(n3059), .F(n3018) );
  IV U1036 ( .A(n3060), .Z(n418) );
  XNOR U1037 ( .A(n3073), .B(n3036), .Z(n3040) );
  MUX U1038 ( .IN0(n3672), .IN1(n3677), .SEL(n3673), .F(n3668) );
  MUX U1039 ( .IN0(n4358), .IN1(n4369), .SEL(n4359), .F(n4346) );
  XNOR U1040 ( .A(n3731), .B(n3716), .Z(n3720) );
  MUX U1041 ( .IN0(n3093), .IN1(n419), .SEL(n3094), .F(n3053) );
  IV U1042 ( .A(n3095), .Z(n419) );
  MUX U1043 ( .IN0(n3967), .IN1(n420), .SEL(n3968), .F(n3949) );
  IV U1044 ( .A(n3969), .Z(n420) );
  XNOR U1045 ( .A(n4362), .B(n4353), .Z(n3988) );
  MUX U1046 ( .IN0(n4001), .IN1(n4003), .SEL(n4002), .F(n3971) );
  MUX U1047 ( .IN0(n2938), .IN1(n3008), .SEL(n2939), .F(n2866) );
  MUX U1048 ( .IN0(n857), .IN1(n421), .SEL(n858), .F(n800) );
  IV U1049 ( .A(n859), .Z(n421) );
  MUX U1050 ( .IN0(n971), .IN1(n1028), .SEL(n972), .F(n915) );
  MUX U1051 ( .IN0(n1003), .IN1(n1069), .SEL(n1004), .F(n943) );
  MUX U1052 ( .IN0(n1012), .IN1(n422), .SEL(n1013), .F(n954) );
  IV U1053 ( .A(n1014), .Z(n422) );
  MUX U1054 ( .IN0(n1049), .IN1(n1115), .SEL(n1050), .F(n991) );
  MUX U1055 ( .IN0(n1233), .IN1(n1304), .SEL(n1234), .F(n1163) );
  MUX U1056 ( .IN0(n1279), .IN1(n1352), .SEL(n1280), .F(n1207) );
  MUX U1057 ( .IN0(n1326), .IN1(n1418), .SEL(n1327), .F(n1253) );
  MUX U1058 ( .IN0(n1464), .IN1(n423), .SEL(n1465), .F(n1371) );
  IV U1059 ( .A(n1466), .Z(n423) );
  MUX U1060 ( .IN0(n1622), .IN1(n1714), .SEL(n1623), .F(n1532) );
  MUX U1061 ( .IN0(n1631), .IN1(n424), .SEL(n1632), .F(n1541) );
  IV U1062 ( .A(n1633), .Z(n424) );
  MUX U1063 ( .IN0(n1604), .IN1(n1696), .SEL(n1605), .F(n1514) );
  MUX U1064 ( .IN0(n1613), .IN1(n425), .SEL(n1614), .F(n1523) );
  IV U1065 ( .A(n1615), .Z(n425) );
  MUX U1066 ( .IN0(n1688), .IN1(n1823), .SEL(n1689), .F(n1595) );
  MUX U1067 ( .IN0(n1952), .IN1(n2023), .SEL(n1953), .F(n1877) );
  MUX U1068 ( .IN0(n1998), .IN1(n2066), .SEL(n1999), .F(n1926) );
  MUX U1069 ( .IN0(n1980), .IN1(n2048), .SEL(n1981), .F(n1908) );
  MUX U1070 ( .IN0(n2522), .IN1(n2566), .SEL(n2523), .F(n2493) );
  MUX U1071 ( .IN0(n2040), .IN1(n2114), .SEL(n2041), .F(n1971) );
  MUX U1072 ( .IN0(n2133), .IN1(n426), .SEL(n2134), .F(n2058) );
  IV U1073 ( .A(n2135), .Z(n426) );
  MUX U1074 ( .IN0(n2628), .IN1(n2670), .SEL(n2629), .F(n2595) );
  MUX U1075 ( .IN0(n2240), .IN1(n2311), .SEL(n2241), .F(n2168) );
  MUX U1076 ( .IN0(n2286), .IN1(n2354), .SEL(n2287), .F(n2214) );
  MUX U1077 ( .IN0(n2268), .IN1(n2336), .SEL(n2269), .F(n2196) );
  MUX U1078 ( .IN0(n2692), .IN1(n2768), .SEL(n2693), .F(n2645) );
  MUX U1079 ( .IN0(n2328), .IN1(n2402), .SEL(n2329), .F(n2259) );
  MUX U1080 ( .IN0(n2439), .IN1(n427), .SEL(n2440), .F(n2364) );
  IV U1081 ( .A(n2441), .Z(n427) );
  MUX U1082 ( .IN0(n2828), .IN1(n2891), .SEL(n2829), .F(n2795) );
  MUX U1083 ( .IN0(n2843), .IN1(n2909), .SEL(n2844), .F(n2751) );
  MUX U1084 ( .IN0(n4744), .IN1(n428), .SEL(n4745), .F(n2421) );
  IV U1085 ( .A(n4746), .Z(n428) );
  XNOR U1086 ( .A(n5035), .B(n5036), .Z(n5026) );
  MUX U1087 ( .IN0(n4760), .IN1(n4569), .SEL(n4571), .F(n4748) );
  MUX U1088 ( .IN0(n4554), .IN1(n4556), .SEL(n4555), .F(n4525) );
  MUX U1089 ( .IN0(n3712), .IN1(n429), .SEL(n3031), .F(n3694) );
  IV U1090 ( .A(n3029), .Z(n429) );
  MUX U1091 ( .IN0(n700), .IN1(n732), .SEL(n701), .F(n667) );
  MUX U1092 ( .IN0(n1459), .IN1(n430), .SEL(n1460), .F(n1366) );
  IV U1093 ( .A(n1461), .Z(n430) );
  MUX U1094 ( .IN0(n2724), .IN1(n431), .SEL(n2725), .F(n2677) );
  IV U1095 ( .A(n2726), .Z(n431) );
  MUX U1096 ( .IN0(n2919), .IN1(n3689), .SEL(n2920), .F(n2848) );
  MUX U1097 ( .IN0(n4942), .IN1(n432), .SEL(n4931), .F(n2443) );
  IV U1098 ( .A(n4930), .Z(n432) );
  XNOR U1099 ( .A(n2954), .B(n2885), .Z(n2889) );
  XNOR U1100 ( .A(n2945), .B(n2876), .Z(n2880) );
  XNOR U1101 ( .A(n2971), .B(n2903), .Z(n2907) );
  XNOR U1102 ( .A(n4159), .B(n2927), .Z(n2930) );
  XNOR U1103 ( .A(n759), .B(n726), .Z(n730) );
  XNOR U1104 ( .A(n896), .B(n849), .Z(n853) );
  MUX U1105 ( .IN0(n1007), .IN1(n433), .SEL(n1008), .F(n947) );
  IV U1106 ( .A(n1009), .Z(n433) );
  XNOR U1107 ( .A(n1019), .B(n964), .Z(n968) );
  XNOR U1108 ( .A(n982), .B(n926), .Z(n929) );
  XNOR U1109 ( .A(n1214), .B(n1147), .Z(n1151) );
  XNOR U1110 ( .A(n1295), .B(n1226), .Z(n1230) );
  MUX U1111 ( .IN0(n1667), .IN1(n1807), .SEL(n1668), .F(n1574) );
  XNOR U1112 ( .A(n1316), .B(n1246), .Z(n1250) );
  XNOR U1113 ( .A(n1342), .B(n1271), .Z(n1275) );
  MUX U1114 ( .IN0(n1536), .IN1(n434), .SEL(n1537), .F(n1450) );
  IV U1115 ( .A(n1538), .Z(n434) );
  MUX U1116 ( .IN0(n1518), .IN1(n435), .SEL(n1519), .F(n1432) );
  IV U1117 ( .A(n1520), .Z(n435) );
  XNOR U1118 ( .A(n1731), .B(n1641), .Z(n1645) );
  XNOR U1119 ( .A(n1678), .B(n1588), .Z(n1592) );
  XNOR U1120 ( .A(n1933), .B(n1861), .Z(n1865) );
  XNOR U1121 ( .A(n1915), .B(n1843), .Z(n1847) );
  XNOR U1122 ( .A(n2506), .B(n2478), .Z(n2484) );
  MUX U1123 ( .IN0(n2497), .IN1(n436), .SEL(n2498), .F(n2468) );
  IV U1124 ( .A(n2499), .Z(n436) );
  XNOR U1125 ( .A(n2014), .B(n1945), .Z(n1949) );
  XNOR U1126 ( .A(n1961), .B(n1892), .Z(n1896) );
  XNOR U1127 ( .A(n2574), .B(n2531), .Z(n2535) );
  MUX U1128 ( .IN0(n2128), .IN1(n437), .SEL(n2129), .F(n2053) );
  IV U1129 ( .A(n2130), .Z(n437) );
  XNOR U1130 ( .A(n2618), .B(n2588), .Z(n2592) );
  XNOR U1131 ( .A(n2221), .B(n2152), .Z(n2156) );
  XNOR U1132 ( .A(n2302), .B(n2233), .Z(n2237) );
  XNOR U1133 ( .A(n2699), .B(n2655), .Z(n2659) );
  XNOR U1134 ( .A(n2318), .B(n2252), .Z(n2256) );
  XNOR U1135 ( .A(n2344), .B(n2278), .Z(n2282) );
  XNOR U1136 ( .A(n2785), .B(n2711), .Z(n2715) );
  MUX U1137 ( .IN0(n2773), .IN1(n438), .SEL(n2774), .F(n2696) );
  IV U1138 ( .A(n2775), .Z(n438) );
  MUX U1139 ( .IN0(n2416), .IN1(n439), .SEL(n2417), .F(n2341) );
  IV U1140 ( .A(n2418), .Z(n439) );
  XOR U1141 ( .A(n642), .B(n641), .Z(n635) );
  XNOR U1142 ( .A(n655), .B(n685), .Z(n678) );
  XNOR U1143 ( .A(n998), .B(n1063), .Z(n1056) );
  XOR U1144 ( .A(n1303), .B(n1302), .Z(n1285) );
  MUX U1145 ( .IN0(n1330), .IN1(n440), .SEL(n1331), .F(n1257) );
  IV U1146 ( .A(n1332), .Z(n440) );
  XOR U1147 ( .A(n1483), .B(n1482), .Z(n1479) );
  MUX U1148 ( .IN0(n1692), .IN1(n441), .SEL(n1693), .F(n1599) );
  IV U1149 ( .A(n1694), .Z(n441) );
  XOR U1150 ( .A(n2022), .B(n2021), .Z(n2004) );
  MUX U1151 ( .IN0(n2044), .IN1(n442), .SEL(n2045), .F(n1975) );
  IV U1152 ( .A(n2046), .Z(n442) );
  MUX U1153 ( .IN0(n443), .IN1(n2736), .SEL(n2737), .F(n2688) );
  IV U1154 ( .A(n2738), .Z(n443) );
  XOR U1155 ( .A(n2310), .B(n2309), .Z(n2292) );
  MUX U1156 ( .IN0(n2332), .IN1(n444), .SEL(n2333), .F(n2263) );
  IV U1157 ( .A(n2334), .Z(n444) );
  MUX U1158 ( .IN0(n2859), .IN1(n445), .SEL(n2860), .F(n2799) );
  IV U1159 ( .A(n2861), .Z(n445) );
  XOR U1160 ( .A(n2454), .B(n2453), .Z(n2436) );
  XOR U1161 ( .A(n752), .B(n751), .Z(n742) );
  XOR U1162 ( .A(n830), .B(n823), .Z(n874) );
  XOR U1163 ( .A(n1076), .B(n1075), .Z(n1055) );
  XNOR U1164 ( .A(n2551), .B(n2563), .Z(n2552) );
  MUX U1165 ( .IN0(n446), .IN1(n2244), .SEL(n1772), .F(n2172) );
  IV U1166 ( .A(n1771), .Z(n446) );
  XOR U1167 ( .A(n2933), .B(n2934), .Z(n2898) );
  NANDN U1168 ( .B(n631), .A(n630), .Z(n613) );
  MUX U1169 ( .IN0(n737), .IN1(o_reg[25]), .SEL(n738), .F(n704) );
  ANDN U1170 ( .A(n921), .B(n922), .Z(n871) );
  MUX U1171 ( .IN0(o_reg[19]), .IN1(n1033), .SEL(n1034), .F(n975) );
  ANDN U1172 ( .A(n1239), .B(n1240), .Z(n1169) );
  MUX U1173 ( .IN0(n1383), .IN1(o_reg[14]), .SEL(n1384), .F(n1309) );
  XNOR U1174 ( .A(n1581), .B(n1578), .Z(n1654) );
  MUX U1175 ( .IN0(n1757), .IN1(o_reg[7]), .SEL(n582), .F(n1753) );
  MUX U1176 ( .IN0(o_reg[2]), .IN1(n492), .SEL(n979), .F(n1773) );
  MUX U1177 ( .IN0(n4310), .IN1(n4321), .SEL(n4311), .F(n4298) );
  MUX U1178 ( .IN0(n3443), .IN1(n3482), .SEL(n3444), .F(n3403) );
  MUX U1179 ( .IN0(n3435), .IN1(n447), .SEL(n3436), .F(n3395) );
  IV U1180 ( .A(n3437), .Z(n447) );
  MUX U1181 ( .IN0(n3903), .IN1(n3920), .SEL(n3904), .F(n3885) );
  MUX U1182 ( .IN0(n3895), .IN1(n448), .SEL(n3896), .F(n3877) );
  IV U1183 ( .A(n3897), .Z(n448) );
  MUX U1184 ( .IN0(n3502), .IN1(n449), .SEL(n3503), .F(n3462) );
  IV U1185 ( .A(n3504), .Z(n449) );
  MUX U1186 ( .IN0(n3409), .IN1(n3448), .SEL(n3410), .F(n3369) );
  MUX U1187 ( .IN0(n3418), .IN1(n450), .SEL(n3419), .F(n3378) );
  IV U1188 ( .A(n3420), .Z(n450) );
  MUX U1189 ( .IN0(n3910), .IN1(n451), .SEL(n3471), .F(n3892) );
  IV U1190 ( .A(n3469), .Z(n451) );
  MUX U1191 ( .IN0(n3453), .IN1(n452), .SEL(n3454), .F(n3413) );
  IV U1192 ( .A(n3455), .Z(n452) );
  XNOR U1193 ( .A(n4278), .B(n4269), .Z(n3873) );
  MUX U1194 ( .IN0(n3863), .IN1(n453), .SEL(n3864), .F(n3845) );
  IV U1195 ( .A(n3865), .Z(n453) );
  XNOR U1196 ( .A(n3353), .B(n3316), .Z(n3320) );
  MUX U1197 ( .IN0(n4262), .IN1(n4273), .SEL(n4263), .F(n4250) );
  MUX U1198 ( .IN0(n3283), .IN1(n3322), .SEL(n3284), .F(n3243) );
  MUX U1199 ( .IN0(n3831), .IN1(n3848), .SEL(n3832), .F(n3813) );
  MUX U1200 ( .IN0(n3823), .IN1(n454), .SEL(n3824), .F(n3805) );
  IV U1201 ( .A(n3825), .Z(n454) );
  MUX U1202 ( .IN0(n3342), .IN1(n455), .SEL(n3343), .F(n3302) );
  IV U1203 ( .A(n3344), .Z(n455) );
  MUX U1204 ( .IN0(n4712), .IN1(n456), .SEL(n4713), .F(n4690) );
  IV U1205 ( .A(n4714), .Z(n456) );
  MUX U1206 ( .IN0(n3249), .IN1(n3288), .SEL(n3250), .F(n3209) );
  MUX U1207 ( .IN0(n3258), .IN1(n457), .SEL(n3259), .F(n3218) );
  IV U1208 ( .A(n3260), .Z(n457) );
  MUX U1209 ( .IN0(n4101), .IN1(n4122), .SEL(n4102), .F(n4079) );
  MUX U1210 ( .IN0(n4107), .IN1(n458), .SEL(n4108), .F(n4085) );
  IV U1211 ( .A(n4109), .Z(n458) );
  MUX U1212 ( .IN0(n4684), .IN1(n4705), .SEL(n4685), .F(n4662) );
  MUX U1213 ( .IN0(n3838), .IN1(n459), .SEL(n3311), .F(n3820) );
  IV U1214 ( .A(n3309), .Z(n459) );
  MUX U1215 ( .IN0(n3293), .IN1(n460), .SEL(n3294), .F(n3253) );
  IV U1216 ( .A(n3295), .Z(n460) );
  XNOR U1217 ( .A(n3233), .B(n3196), .Z(n3200) );
  XNOR U1218 ( .A(n4420), .B(n4421), .Z(n4118) );
  XNOR U1219 ( .A(n4826), .B(n4817), .Z(n4681) );
  MUX U1220 ( .IN0(n4810), .IN1(n4821), .SEL(n4811), .F(n4798) );
  XNOR U1221 ( .A(n4230), .B(n4221), .Z(n3801) );
  MUX U1222 ( .IN0(n3791), .IN1(n461), .SEL(n3792), .F(n3773) );
  IV U1223 ( .A(n3793), .Z(n461) );
  MUX U1224 ( .IN0(n4214), .IN1(n4225), .SEL(n4215), .F(n4202) );
  MUX U1225 ( .IN0(n3123), .IN1(n3162), .SEL(n3124), .F(n3083) );
  MUX U1226 ( .IN0(n3759), .IN1(n3776), .SEL(n3760), .F(n3741) );
  MUX U1227 ( .IN0(n3751), .IN1(n462), .SEL(n3752), .F(n3733) );
  IV U1228 ( .A(n3753), .Z(n462) );
  MUX U1229 ( .IN0(n3182), .IN1(n463), .SEL(n3183), .F(n3142) );
  IV U1230 ( .A(n3184), .Z(n463) );
  XNOR U1231 ( .A(n4398), .B(n4389), .Z(n4054) );
  MUX U1232 ( .IN0(n4067), .IN1(n4069), .SEL(n4068), .F(n4045) );
  MUX U1233 ( .IN0(n4481), .IN1(n4495), .SEL(n4483), .F(n4465) );
  XNOR U1234 ( .A(n4666), .B(n4647), .Z(n4651) );
  MUX U1235 ( .IN0(n3089), .IN1(n3128), .SEL(n3090), .F(n3049) );
  MUX U1236 ( .IN0(n3098), .IN1(n464), .SEL(n3099), .F(n3058) );
  IV U1237 ( .A(n3100), .Z(n464) );
  XNOR U1238 ( .A(n3113), .B(n3076), .Z(n3080) );
  MUX U1239 ( .IN0(n3629), .IN1(n3643), .SEL(n3631), .F(n3613) );
  MUX U1240 ( .IN0(n4013), .IN1(n4034), .SEL(n4014), .F(n3991) );
  MUX U1241 ( .IN0(n4370), .IN1(n4381), .SEL(n4371), .F(n4358) );
  MUX U1242 ( .IN0(n4019), .IN1(n465), .SEL(n4020), .F(n3997) );
  IV U1243 ( .A(n4021), .Z(n465) );
  MUX U1244 ( .IN0(n4459), .IN1(n4474), .SEL(n4461), .F(n4448) );
  MUX U1245 ( .IN0(n4977), .IN1(n4992), .SEL(n4979), .F(n4961) );
  MUX U1246 ( .IN0(n4869), .IN1(n4884), .SEL(n4871), .F(n4846) );
  MUX U1247 ( .IN0(n4863), .IN1(n4878), .SEL(n4865), .F(n4852) );
  XNOR U1248 ( .A(n4790), .B(n4781), .Z(n4615) );
  MUX U1249 ( .IN0(n4596), .IN1(n4617), .SEL(n4597), .F(n4574) );
  MUX U1250 ( .IN0(n3766), .IN1(n466), .SEL(n3151), .F(n3748) );
  IV U1251 ( .A(n3149), .Z(n466) );
  MUX U1252 ( .IN0(n3133), .IN1(n467), .SEL(n3134), .F(n3093) );
  IV U1253 ( .A(n3135), .Z(n467) );
  MUX U1254 ( .IN0(n3607), .IN1(n3622), .SEL(n3609), .F(n3596) );
  MUX U1255 ( .IN0(n4364), .IN1(n468), .SEL(n4365), .F(n4352) );
  IV U1256 ( .A(n4366), .Z(n468) );
  XNOR U1257 ( .A(n4512), .B(n4513), .Z(n4500) );
  MUX U1258 ( .IN0(n4967), .IN1(n4982), .SEL(n4969), .F(n4944) );
  XNOR U1259 ( .A(n4916), .B(n4917), .Z(n4904) );
  MUX U1260 ( .IN0(n4762), .IN1(n4773), .SEL(n4763), .F(n4750) );
  XNOR U1261 ( .A(n4182), .B(n4173), .Z(n3729) );
  MUX U1262 ( .IN0(n3719), .IN1(n469), .SEL(n3720), .F(n3701) );
  IV U1263 ( .A(n3721), .Z(n469) );
  XOR U1264 ( .A(n3041), .B(n3040), .Z(n3055) );
  XNOR U1265 ( .A(n3660), .B(n3661), .Z(n3648) );
  XNOR U1266 ( .A(n4148), .B(n4149), .Z(n4133) );
  MUX U1267 ( .IN0(n4166), .IN1(n4177), .SEL(n4167), .F(n3690) );
  XNOR U1268 ( .A(n5014), .B(n5015), .Z(n5002) );
  XNOR U1269 ( .A(n4731), .B(n4732), .Z(n4716) );
  XNOR U1270 ( .A(n4600), .B(n4581), .Z(n4585) );
  MUX U1271 ( .IN0(n2981), .IN1(n3704), .SEL(n2982), .F(n2910) );
  MUX U1272 ( .IN0(n2973), .IN1(n470), .SEL(n2974), .F(n2902) );
  IV U1273 ( .A(n2975), .Z(n470) );
  XNOR U1274 ( .A(n2993), .B(n2957), .Z(n2961) );
  XOR U1275 ( .A(n3001), .B(n3000), .Z(n3015) );
  MUX U1276 ( .IN0(n3971), .IN1(n3973), .SEL(n3972), .F(n3953) );
  MUX U1277 ( .IN0(n4356), .IN1(n3986), .SEL(n3988), .F(n4344) );
  MUX U1278 ( .IN0(n725), .IN1(n471), .SEL(n726), .F(n692) );
  IV U1279 ( .A(n727), .Z(n471) );
  MUX U1280 ( .IN0(n808), .IN1(n864), .SEL(n809), .F(n769) );
  MUX U1281 ( .IN0(n837), .IN1(n888), .SEL(n838), .F(n783) );
  MUX U1282 ( .IN0(n1029), .IN1(n1095), .SEL(n1030), .F(n971) );
  MUX U1283 ( .IN0(n1070), .IN1(n1136), .SEL(n1071), .F(n1003) );
  MUX U1284 ( .IN0(n1305), .IN1(n1378), .SEL(n1306), .F(n1233) );
  MUX U1285 ( .IN0(n1353), .IN1(n1445), .SEL(n1354), .F(n1279) );
  MUX U1286 ( .IN0(n1419), .IN1(n1504), .SEL(n1420), .F(n1326) );
  MUX U1287 ( .IN0(n1715), .IN1(n1850), .SEL(n1716), .F(n1622) );
  MUX U1288 ( .IN0(n1697), .IN1(n1832), .SEL(n1698), .F(n1604) );
  MUX U1289 ( .IN0(n1869), .IN1(n472), .SEL(n1870), .F(n1733) );
  IV U1290 ( .A(n1871), .Z(n472) );
  MUX U1291 ( .IN0(n1824), .IN1(n1898), .SEL(n1825), .F(n1688) );
  MUX U1292 ( .IN0(n1917), .IN1(n473), .SEL(n1918), .F(n1842) );
  IV U1293 ( .A(n1919), .Z(n473) );
  MUX U1294 ( .IN0(n2093), .IN1(n2167), .SEL(n2094), .F(n2024) );
  MUX U1295 ( .IN0(n2067), .IN1(n2141), .SEL(n2068), .F(n1998) );
  MUX U1296 ( .IN0(n2049), .IN1(n2123), .SEL(n2050), .F(n1980) );
  MUX U1297 ( .IN0(n2595), .IN1(n2627), .SEL(n2596), .F(n2547) );
  MUX U1298 ( .IN0(n2567), .IN1(n2601), .SEL(n2568), .F(n2522) );
  MUX U1299 ( .IN0(n2151), .IN1(n474), .SEL(n2152), .F(n2076) );
  IV U1300 ( .A(n2153), .Z(n474) );
  MUX U1301 ( .IN0(n2115), .IN1(n2186), .SEL(n2116), .F(n2040) );
  MUX U1302 ( .IN0(n2355), .IN1(n2429), .SEL(n2356), .F(n2286) );
  MUX U1303 ( .IN0(n2337), .IN1(n2411), .SEL(n2338), .F(n2268) );
  MUX U1304 ( .IN0(n2346), .IN1(n475), .SEL(n2347), .F(n2277) );
  IV U1305 ( .A(n2348), .Z(n475) );
  MUX U1306 ( .IN0(n2795), .IN1(n2827), .SEL(n2796), .F(n2718) );
  MUX U1307 ( .IN0(n2769), .IN1(n2801), .SEL(n2770), .F(n2692) );
  MUX U1308 ( .IN0(n2456), .IN1(n5043), .SEL(n2457), .F(n2381) );
  MUX U1309 ( .IN0(n2403), .IN1(n4528), .SEL(n2404), .F(n2328) );
  MUX U1310 ( .IN0(n2875), .IN1(n476), .SEL(n2876), .F(n2811) );
  IV U1311 ( .A(n2877), .Z(n476) );
  MUX U1312 ( .IN0(n2951), .IN1(n477), .SEL(n2952), .F(n2879) );
  IV U1313 ( .A(n2953), .Z(n477) );
  XNOR U1314 ( .A(n3666), .B(n3556), .Z(n3560) );
  MUX U1315 ( .IN0(n791), .IN1(n478), .SEL(n792), .F(n754) );
  IV U1316 ( .A(n793), .Z(n478) );
  MUX U1317 ( .IN0(n991), .IN1(n1048), .SEL(n992), .F(n932) );
  MUX U1318 ( .IN0(n1192), .IN1(n1261), .SEL(n1193), .F(n1124) );
  MUX U1319 ( .IN0(n1270), .IN1(n479), .SEL(n1271), .F(n1200) );
  IV U1320 ( .A(n1272), .Z(n479) );
  MUX U1321 ( .IN0(n1659), .IN1(n480), .SEL(n1660), .F(n1568) );
  IV U1322 ( .A(n1661), .Z(n480) );
  XNOR U1323 ( .A(n5027), .B(n5023), .Z(n4933) );
  XNOR U1324 ( .A(n4948), .B(n4939), .Z(n4931) );
  XNOR U1325 ( .A(n4754), .B(n4745), .Z(n4564) );
  MUX U1326 ( .IN0(n3694), .IN1(n481), .SEL(n2991), .F(n2923) );
  IV U1327 ( .A(n2989), .Z(n481) );
  MUX U1328 ( .IN0(n750), .IN1(n482), .SEL(n751), .F(n716) );
  IV U1329 ( .A(n752), .Z(n482) );
  XNOR U1330 ( .A(n855), .B(n801), .Z(n805) );
  XNOR U1331 ( .A(n1086), .B(n1022), .Z(n1026) );
  XNOR U1332 ( .A(n1077), .B(n1013), .Z(n1017) );
  XNOR U1333 ( .A(n1039), .B(n984), .Z(n988) );
  XNOR U1334 ( .A(n1243), .B(n1176), .Z(n1180) );
  XNOR U1335 ( .A(n1369), .B(n1298), .Z(n1302) );
  XNOR U1336 ( .A(n1360), .B(n1289), .Z(n1293) );
  MUX U1337 ( .IN0(n1339), .IN1(n483), .SEL(n1340), .F(n1266) );
  IV U1338 ( .A(n1341), .Z(n483) );
  XNOR U1339 ( .A(n1495), .B(n1412), .Z(n1416) );
  XNOR U1340 ( .A(n1629), .B(n1542), .Z(n1546) );
  XNOR U1341 ( .A(n1611), .B(n1524), .Z(n1528) );
  XNOR U1342 ( .A(n1814), .B(n1681), .Z(n1685) );
  MUX U1343 ( .IN0(n1912), .IN1(n484), .SEL(n1913), .F(n1837) );
  IV U1344 ( .A(n1914), .Z(n484) );
  XNOR U1345 ( .A(n2005), .B(n1936), .Z(n1940) );
  XNOR U1346 ( .A(n2537), .B(n2509), .Z(n2513) );
  XNOR U1347 ( .A(n2083), .B(n2017), .Z(n2021) );
  XNOR U1348 ( .A(n2030), .B(n1964), .Z(n1968) );
  MUX U1349 ( .IN0(n2683), .IN1(n2731), .SEL(n2684), .F(n2636) );
  XNOR U1350 ( .A(n2131), .B(n2059), .Z(n2063) );
  XNOR U1351 ( .A(n2609), .B(n2579), .Z(n2583) );
  XNOR U1352 ( .A(n2661), .B(n2621), .Z(n2625) );
  MUX U1353 ( .IN0(n2649), .IN1(n485), .SEL(n2650), .F(n2606) );
  IV U1354 ( .A(n2651), .Z(n485) );
  XNOR U1355 ( .A(n2249), .B(n2180), .Z(n2184) );
  XNOR U1356 ( .A(n2371), .B(n2305), .Z(n2309) );
  XNOR U1357 ( .A(n2362), .B(n2296), .Z(n2300) );
  MUX U1358 ( .IN0(n2341), .IN1(n486), .SEL(n2342), .F(n2272) );
  IV U1359 ( .A(n2343), .Z(n486) );
  XNOR U1360 ( .A(n2776), .B(n2702), .Z(n2706) );
  XNOR U1361 ( .A(n2818), .B(n2788), .Z(n2792) );
  XNOR U1362 ( .A(n2833), .B(n2744), .Z(n2748) );
  XNOR U1363 ( .A(n4519), .B(n2396), .Z(n2400) );
  MUX U1364 ( .IN0(n621), .IN1(n487), .SEL(n622), .F(n607) );
  IV U1365 ( .A(n623), .Z(n487) );
  XOR U1366 ( .A(n665), .B(n664), .Z(n657) );
  XOR U1367 ( .A(n877), .B(n876), .Z(n883) );
  XOR U1368 ( .A(n1094), .B(n1093), .Z(n1076) );
  XOR U1369 ( .A(n1047), .B(n1046), .Z(n1067) );
  XOR U1370 ( .A(n1161), .B(n1160), .Z(n1143) );
  MUX U1371 ( .IN0(n1574), .IN1(n1666), .SEL(n1575), .F(n1484) );
  XOR U1372 ( .A(n1377), .B(n1376), .Z(n1359) );
  XOR U1373 ( .A(n1470), .B(n1469), .Z(n1452) );
  XOR U1374 ( .A(n1556), .B(n1555), .Z(n1538) );
  XOR U1375 ( .A(n1739), .B(n1738), .Z(n1721) );
  XOR U1376 ( .A(n1806), .B(n1805), .Z(n1797) );
  XOR U1377 ( .A(n1875), .B(n1874), .Z(n1857) );
  XOR U1378 ( .A(n1950), .B(n1949), .Z(n1932) );
  XOR U1379 ( .A(n2166), .B(n2165), .Z(n2148) );
  XOR U1380 ( .A(n2238), .B(n2237), .Z(n2220) );
  XNOR U1381 ( .A(n2736), .B(n2762), .Z(n2755) );
  XOR U1382 ( .A(n2826), .B(n2825), .Z(n2808) );
  MUX U1383 ( .IN0(n2914), .IN1(n488), .SEL(n2915), .F(n2859) );
  IV U1384 ( .A(n2916), .Z(n488) );
  AND U1385 ( .A(n610), .B(n611), .Z(n609) );
  XOR U1386 ( .A(n689), .B(n688), .Z(n676) );
  XOR U1387 ( .A(n843), .B(n842), .Z(n834) );
  XOR U1388 ( .A(n895), .B(n894), .Z(n886) );
  XOR U1389 ( .A(n1213), .B(n1212), .Z(n1189) );
  ANDN U1390 ( .A(n1491), .B(n1492), .Z(n1399) );
  XOR U1391 ( .A(n1628), .B(n1627), .Z(n1601) );
  MUX U1392 ( .IN0(n2028), .IN1(n489), .SEL(n1760), .F(n1956) );
  IV U1393 ( .A(n1759), .Z(n489) );
  XOR U1394 ( .A(n2073), .B(n2072), .Z(n2046) );
  XOR U1395 ( .A(n2599), .B(n2558), .Z(n2632) );
  MUX U1396 ( .IN0(n2316), .IN1(n490), .SEL(n1776), .F(n2244) );
  IV U1397 ( .A(n1775), .Z(n490) );
  XOR U1398 ( .A(n2361), .B(n2360), .Z(n2334) );
  XOR U1399 ( .A(n2436), .B(n2435), .Z(n2409) );
  ANDN U1400 ( .A(n650), .B(n651), .Z(n630) );
  ANDN U1401 ( .A(n775), .B(n776), .Z(n739) );
  MUX U1402 ( .IN0(o_reg[23]), .IN1(n812), .SEL(n813), .F(n773) );
  ANDN U1403 ( .A(n977), .B(n978), .Z(n921) );
  MUX U1404 ( .IN0(n1100), .IN1(o_reg[18]), .SEL(n1101), .F(n1033) );
  MUX U1405 ( .IN0(n491), .IN1(n1311), .SEL(n1312), .F(n1239) );
  IV U1406 ( .A(n1313), .Z(n491) );
  MUX U1407 ( .IN0(n1476), .IN1(o_reg[13]), .SEL(n1477), .F(n1383) );
  XNOR U1408 ( .A(n1674), .B(n1671), .Z(n1783) );
  MUX U1409 ( .IN0(o_reg[9]), .IN1(n1749), .SEL(n580), .F(n1745) );
  MUX U1410 ( .IN0(o_reg[5]), .IN1(n1765), .SEL(n584), .F(n1761) );
  MUX U1411 ( .IN0(o_reg[1]), .IN1(n1781), .SEL(n1782), .F(n492) );
  IV U1412 ( .A(n492), .Z(n1777) );
  MUX U1413 ( .IN0(n595), .IN1(o_reg[30]), .SEL(n596), .F(n586) );
  MUX U1414 ( .IN0(n3523), .IN1(n3562), .SEL(n3524), .F(n3483) );
  MUX U1415 ( .IN0(n4320), .IN1(n493), .SEL(n3945), .F(n4308) );
  IV U1416 ( .A(n3944), .Z(n493) );
  MUX U1417 ( .IN0(n3439), .IN1(n494), .SEL(n3440), .F(n3399) );
  IV U1418 ( .A(n3441), .Z(n494) );
  MUX U1419 ( .IN0(n4304), .IN1(n495), .SEL(n4305), .F(n4292) );
  IV U1420 ( .A(n4306), .Z(n495) );
  XNOR U1421 ( .A(n3911), .B(n3896), .Z(n3900) );
  MUX U1422 ( .IN0(n3885), .IN1(n3902), .SEL(n3886), .F(n3867) );
  MUX U1423 ( .IN0(n4286), .IN1(n4297), .SEL(n4287), .F(n4274) );
  MUX U1424 ( .IN0(n3363), .IN1(n3402), .SEL(n3364), .F(n3323) );
  MUX U1425 ( .IN0(n3355), .IN1(n496), .SEL(n3356), .F(n3315) );
  IV U1426 ( .A(n3357), .Z(n496) );
  MUX U1427 ( .IN0(n3369), .IN1(n3408), .SEL(n3370), .F(n3329) );
  MUX U1428 ( .IN0(n3422), .IN1(n497), .SEL(n3423), .F(n3382) );
  IV U1429 ( .A(n3424), .Z(n497) );
  MUX U1430 ( .IN0(n3378), .IN1(n498), .SEL(n3379), .F(n3338) );
  IV U1431 ( .A(n3380), .Z(n498) );
  MUX U1432 ( .IN0(n3892), .IN1(n499), .SEL(n3431), .F(n3874) );
  IV U1433 ( .A(n3429), .Z(n499) );
  MUX U1434 ( .IN0(n4272), .IN1(n500), .SEL(n3873), .F(n4260) );
  IV U1435 ( .A(n3872), .Z(n500) );
  MUX U1436 ( .IN0(n3373), .IN1(n501), .SEL(n3374), .F(n3333) );
  IV U1437 ( .A(n3375), .Z(n501) );
  MUX U1438 ( .IN0(n4256), .IN1(n502), .SEL(n4257), .F(n4244) );
  IV U1439 ( .A(n4258), .Z(n502) );
  XNOR U1440 ( .A(n3839), .B(n3824), .Z(n3828) );
  MUX U1441 ( .IN0(n3813), .IN1(n3830), .SEL(n3814), .F(n3795) );
  XNOR U1442 ( .A(n3273), .B(n3236), .Z(n3240) );
  XNOR U1443 ( .A(n4103), .B(n4104), .Z(n4113) );
  MUX U1444 ( .IN0(n4238), .IN1(n4249), .SEL(n4239), .F(n4226) );
  XNOR U1445 ( .A(n4686), .B(n4687), .Z(n4696) );
  MUX U1446 ( .IN0(n3203), .IN1(n3242), .SEL(n3204), .F(n3163) );
  MUX U1447 ( .IN0(n3209), .IN1(n3248), .SEL(n3210), .F(n3169) );
  MUX U1448 ( .IN0(n3262), .IN1(n503), .SEL(n3263), .F(n3222) );
  IV U1449 ( .A(n3264), .Z(n503) );
  MUX U1450 ( .IN0(n3218), .IN1(n504), .SEL(n3219), .F(n3178) );
  IV U1451 ( .A(n3220), .Z(n504) );
  XNOR U1452 ( .A(n4422), .B(n4413), .Z(n4098) );
  MUX U1453 ( .IN0(n4085), .IN1(n505), .SEL(n4086), .F(n4063) );
  IV U1454 ( .A(n4087), .Z(n505) );
  XNOR U1455 ( .A(n4824), .B(n4825), .Z(n4701) );
  XNOR U1456 ( .A(n4664), .B(n4665), .Z(n4674) );
  MUX U1457 ( .IN0(n3820), .IN1(n506), .SEL(n3271), .F(n3802) );
  IV U1458 ( .A(n3269), .Z(n506) );
  MUX U1459 ( .IN0(n4057), .IN1(n4078), .SEL(n4058), .F(n4035) );
  MUX U1460 ( .IN0(n4394), .IN1(n4405), .SEL(n4395), .F(n4382) );
  XNOR U1461 ( .A(n4812), .B(n4813), .Z(n4679) );
  MUX U1462 ( .IN0(n4224), .IN1(n507), .SEL(n3801), .F(n4212) );
  IV U1463 ( .A(n3800), .Z(n507) );
  MUX U1464 ( .IN0(n3213), .IN1(n508), .SEL(n3214), .F(n3173) );
  IV U1465 ( .A(n3215), .Z(n508) );
  XNOR U1466 ( .A(n3153), .B(n3116), .Z(n3120) );
  MUX U1467 ( .IN0(n4792), .IN1(n509), .SEL(n4793), .F(n4780) );
  IV U1468 ( .A(n4794), .Z(n509) );
  XNOR U1469 ( .A(n4800), .B(n4801), .Z(n4657) );
  MUX U1470 ( .IN0(n4618), .IN1(n4639), .SEL(n4619), .F(n4596) );
  MUX U1471 ( .IN0(n4624), .IN1(n510), .SEL(n4625), .F(n4602) );
  IV U1472 ( .A(n4626), .Z(n510) );
  MUX U1473 ( .IN0(n4208), .IN1(n511), .SEL(n4209), .F(n4196) );
  IV U1474 ( .A(n4210), .Z(n511) );
  XNOR U1475 ( .A(n3767), .B(n3752), .Z(n3756) );
  MUX U1476 ( .IN0(n3741), .IN1(n3758), .SEL(n3742), .F(n3723) );
  XNOR U1477 ( .A(n4386), .B(n4377), .Z(n4032) );
  MUX U1478 ( .IN0(n4465), .IN1(n4480), .SEL(n4467), .F(n4442) );
  MUX U1479 ( .IN0(n4506), .IN1(n4509), .SEL(n4507), .F(n4491) );
  MUX U1480 ( .IN0(n4190), .IN1(n4201), .SEL(n4191), .F(n4178) );
  MUX U1481 ( .IN0(n4910), .IN1(n4913), .SEL(n4911), .F(n4895) );
  MUX U1482 ( .IN0(n4774), .IN1(n4785), .SEL(n4775), .F(n4762) );
  MUX U1483 ( .IN0(n3043), .IN1(n3082), .SEL(n3044), .F(n3003) );
  XNOR U1484 ( .A(n3136), .B(n3099), .Z(n3103) );
  MUX U1485 ( .IN0(n3049), .IN1(n3088), .SEL(n3050), .F(n3009) );
  MUX U1486 ( .IN0(n3613), .IN1(n3628), .SEL(n3615), .F(n3588) );
  MUX U1487 ( .IN0(n3654), .IN1(n3657), .SEL(n3655), .F(n3639) );
  XNOR U1488 ( .A(n4039), .B(n4020), .Z(n4024) );
  MUX U1489 ( .IN0(n4448), .IN1(n4458), .SEL(n4450), .F(n4436) );
  MUX U1490 ( .IN0(n5008), .IN1(n5011), .SEL(n5009), .F(n4993) );
  MUX U1491 ( .IN0(n4852), .IN1(n4862), .SEL(n4854), .F(n4840) );
  MUX U1492 ( .IN0(n3748), .IN1(n512), .SEL(n3111), .F(n3730) );
  IV U1493 ( .A(n3109), .Z(n512) );
  XNOR U1494 ( .A(n3033), .B(n2996), .Z(n3000) );
  MUX U1495 ( .IN0(n3668), .IN1(n3671), .SEL(n3669), .F(n3555) );
  MUX U1496 ( .IN0(n3975), .IN1(n3990), .SEL(n3976), .F(n3957) );
  MUX U1497 ( .IN0(n4352), .IN1(n513), .SEL(n4353), .F(n4340) );
  IV U1498 ( .A(n4354), .Z(n513) );
  XNOR U1499 ( .A(n4360), .B(n4361), .Z(n4008) );
  XNOR U1500 ( .A(n4498), .B(n4499), .Z(n4157) );
  MUX U1501 ( .IN0(n4950), .IN1(n4960), .SEL(n4952), .F(n4938) );
  XNOR U1502 ( .A(n4902), .B(n4903), .Z(n4740) );
  XNOR U1503 ( .A(n4766), .B(n4757), .Z(n4571) );
  MUX U1504 ( .IN0(n4584), .IN1(n4586), .SEL(n4585), .F(n4554) );
  MUX U1505 ( .IN0(n4176), .IN1(n514), .SEL(n3729), .F(n4164) );
  IV U1506 ( .A(n3728), .Z(n514) );
  XNOR U1507 ( .A(n3713), .B(n3698), .Z(n3702) );
  MUX U1508 ( .IN0(n3053), .IN1(n515), .SEL(n3054), .F(n3013) );
  IV U1509 ( .A(n3055), .Z(n515) );
  XNOR U1510 ( .A(n3646), .B(n3647), .Z(n3592) );
  XNOR U1511 ( .A(n4348), .B(n4349), .Z(n3986) );
  XNOR U1512 ( .A(n4140), .B(n4130), .Z(n4134) );
  MUX U1513 ( .IN0(n865), .IN1(n914), .SEL(n866), .F(n808) );
  MUX U1514 ( .IN0(n1137), .IN1(n1206), .SEL(n1138), .F(n1070) );
  MUX U1515 ( .IN0(n1446), .IN1(n1531), .SEL(n1447), .F(n1353) );
  MUX U1516 ( .IN0(n1455), .IN1(n516), .SEL(n1456), .F(n1362) );
  IV U1517 ( .A(n1457), .Z(n516) );
  MUX U1518 ( .IN0(n1428), .IN1(n1513), .SEL(n1429), .F(n1335) );
  MUX U1519 ( .IN0(n1558), .IN1(n1647), .SEL(n1559), .F(n1472) );
  MUX U1520 ( .IN0(n1550), .IN1(n517), .SEL(n1551), .F(n1464) );
  IV U1521 ( .A(n1552), .Z(n517) );
  MUX U1522 ( .IN0(n1497), .IN1(n518), .SEL(n1498), .F(n1411) );
  IV U1523 ( .A(n1499), .Z(n518) );
  MUX U1524 ( .IN0(n1851), .IN1(n1925), .SEL(n1852), .F(n1715) );
  MUX U1525 ( .IN0(n1833), .IN1(n1907), .SEL(n1834), .F(n1697) );
  MUX U1526 ( .IN0(n1944), .IN1(n519), .SEL(n1945), .F(n1869) );
  IV U1527 ( .A(n1946), .Z(n519) );
  MUX U1528 ( .IN0(n1935), .IN1(n520), .SEL(n1936), .F(n1860) );
  IV U1529 ( .A(n1937), .Z(n520) );
  MUX U1530 ( .IN0(n1891), .IN1(n521), .SEL(n1892), .F(n1816) );
  IV U1531 ( .A(n1893), .Z(n521) );
  MUX U1532 ( .IN0(n2508), .IN1(n522), .SEL(n2509), .F(n2477) );
  IV U1533 ( .A(n2510), .Z(n522) );
  MUX U1534 ( .IN0(n2024), .IN1(n2092), .SEL(n2025), .F(n1952) );
  MUX U1535 ( .IN0(n2142), .IN1(n2213), .SEL(n2143), .F(n2067) );
  MUX U1536 ( .IN0(n2124), .IN1(n2195), .SEL(n2125), .F(n2049) );
  MUX U1537 ( .IN0(n2602), .IN1(n2644), .SEL(n2603), .F(n2567) );
  MUX U1538 ( .IN0(n2232), .IN1(n523), .SEL(n2233), .F(n2160) );
  IV U1539 ( .A(n2234), .Z(n523) );
  MUX U1540 ( .IN0(n2179), .IN1(n524), .SEL(n2180), .F(n2107) );
  IV U1541 ( .A(n2181), .Z(n524) );
  MUX U1542 ( .IN0(n2663), .IN1(n525), .SEL(n2664), .F(n2620) );
  IV U1543 ( .A(n2665), .Z(n525) );
  MUX U1544 ( .IN0(n2312), .IN1(n2380), .SEL(n2313), .F(n2240) );
  MUX U1545 ( .IN0(n2430), .IN1(n4923), .SEL(n2431), .F(n2355) );
  MUX U1546 ( .IN0(n2412), .IN1(n4542), .SEL(n2413), .F(n2337) );
  MUX U1547 ( .IN0(n2802), .IN1(n2865), .SEL(n2803), .F(n2769) );
  MUX U1548 ( .IN0(n5022), .IN1(n526), .SEL(n5023), .F(n2448) );
  IV U1549 ( .A(n5024), .Z(n526) );
  MUX U1550 ( .IN0(n4529), .IN1(n4557), .SEL(n4530), .F(n2403) );
  MUX U1551 ( .IN0(n4521), .IN1(n527), .SEL(n4522), .F(n2395) );
  IV U1552 ( .A(n4523), .Z(n527) );
  MUX U1553 ( .IN0(n2884), .IN1(n528), .SEL(n2885), .F(n2820) );
  IV U1554 ( .A(n2886), .Z(n528) );
  MUX U1555 ( .IN0(n2910), .IN1(n2980), .SEL(n2911), .F(n2843) );
  XNOR U1556 ( .A(n5000), .B(n5001), .Z(n4934) );
  XNOR U1557 ( .A(n4723), .B(n4713), .Z(n4717) );
  XNOR U1558 ( .A(n4836), .B(n4837), .Z(n4721) );
  MUX U1559 ( .IN0(n4160), .IN1(n529), .SEL(n4161), .F(n2927) );
  IV U1560 ( .A(n4162), .Z(n529) );
  XOR U1561 ( .A(n2962), .B(n2961), .Z(n2944) );
  XNOR U1562 ( .A(n3016), .B(n2948), .Z(n2952) );
  XNOR U1563 ( .A(n3594), .B(n3579), .Z(n3583) );
  XNOR U1564 ( .A(n3965), .B(n3950), .Z(n3954) );
  MUX U1565 ( .IN0(n746), .IN1(n782), .SEL(n747), .F(n712) );
  XOR U1566 ( .A(n3561), .B(n3560), .Z(n3575) );
  MUX U1567 ( .IN0(n667), .IN1(n699), .SEL(n668), .F(n644) );
  XNOR U1568 ( .A(n723), .B(n693), .Z(n697) );
  XNOR U1569 ( .A(n790), .B(n754), .Z(n757) );
  MUX U1570 ( .IN0(n932), .IN1(n990), .SEL(n933), .F(n878) );
  XNOR U1571 ( .A(n905), .B(n858), .Z(n862) );
  XNOR U1572 ( .A(n952), .B(n899), .Z(n903) );
  XNOR U1573 ( .A(n1153), .B(n1089), .Z(n1093) );
  XNOR U1574 ( .A(n1144), .B(n1080), .Z(n1084) );
  XNOR U1575 ( .A(n1106), .B(n1042), .Z(n1046) );
  MUX U1576 ( .IN0(n1131), .IN1(n1199), .SEL(n1133), .F(n1059) );
  XNOR U1577 ( .A(n1435), .B(n1345), .Z(n1349) );
  XNOR U1578 ( .A(n1658), .B(n1568), .Z(n1571) );
  XNOR U1579 ( .A(n1722), .B(n1632), .Z(n1636) );
  XNOR U1580 ( .A(n1704), .B(n1614), .Z(n1618) );
  MUX U1581 ( .IN0(n2464), .IN1(n2492), .SEL(n2465), .F(n1791) );
  XNOR U1582 ( .A(n1987), .B(n1918), .Z(n1922) );
  XNOR U1583 ( .A(n2529), .B(n2501), .Z(n2504) );
  XNOR U1584 ( .A(n2149), .B(n2077), .Z(n2081) );
  XNOR U1585 ( .A(n2203), .B(n2134), .Z(n2138) );
  XNOR U1586 ( .A(n2652), .B(n2612), .Z(n2616) );
  MUX U1587 ( .IN0(n2848), .IN1(n2918), .SEL(n2849), .F(n2762) );
  XNOR U1588 ( .A(n2437), .B(n2365), .Z(n2369) );
  XNOR U1589 ( .A(n2419), .B(n2347), .Z(n2351) );
  XNOR U1590 ( .A(n2809), .B(n2779), .Z(n2783) );
  MUX U1591 ( .IN0(n4547), .IN1(n530), .SEL(n4536), .F(n2416) );
  IV U1592 ( .A(n4535), .Z(n530) );
  XNOR U1593 ( .A(n2900), .B(n2836), .Z(n2840) );
  MUX U1594 ( .IN0(n2923), .IN1(n531), .SEL(n2924), .F(n2852) );
  IV U1595 ( .A(n2925), .Z(n531) );
  XOR U1596 ( .A(n4932), .B(n4933), .Z(n4537) );
  XOR U1597 ( .A(n2890), .B(n2889), .Z(n2872) );
  XOR U1598 ( .A(n623), .B(n622), .Z(n619) );
  XOR U1599 ( .A(n731), .B(n730), .Z(n718) );
  XOR U1600 ( .A(n767), .B(n766), .Z(n752) );
  XOR U1601 ( .A(n913), .B(n912), .Z(n895) );
  XOR U1602 ( .A(n969), .B(n968), .Z(n951) );
  XOR U1603 ( .A(n1027), .B(n1026), .Z(n1009) );
  XOR U1604 ( .A(n1114), .B(n1113), .Z(n1130) );
  XOR U1605 ( .A(n1231), .B(n1230), .Z(n1213) );
  XOR U1606 ( .A(n1181), .B(n1180), .Z(n1198) );
  XOR U1607 ( .A(n1251), .B(n1250), .Z(n1268) );
  XOR U1608 ( .A(n1324), .B(n1323), .Z(n1341) );
  XOR U1609 ( .A(n1417), .B(n1416), .Z(n1434) );
  XOR U1610 ( .A(n1503), .B(n1502), .Z(n1520) );
  XOR U1611 ( .A(n1646), .B(n1645), .Z(n1628) );
  XOR U1612 ( .A(n1593), .B(n1592), .Z(n1610) );
  XOR U1613 ( .A(n1665), .B(n1664), .Z(n1657) );
  XOR U1614 ( .A(n1686), .B(n1685), .Z(n1703) );
  XOR U1615 ( .A(n1822), .B(n1821), .Z(n1839) );
  XOR U1616 ( .A(n2485), .B(n2484), .Z(n2470) );
  XOR U1617 ( .A(n1897), .B(n1896), .Z(n1914) );
  XOR U1618 ( .A(n2514), .B(n2513), .Z(n2499) );
  XOR U1619 ( .A(n1969), .B(n1968), .Z(n1986) );
  MUX U1620 ( .IN0(n2636), .IN1(n2682), .SEL(n2637), .F(n2563) );
  XOR U1621 ( .A(n2545), .B(n2544), .Z(n2528) );
  XOR U1622 ( .A(n2091), .B(n2090), .Z(n2073) );
  XOR U1623 ( .A(n2038), .B(n2037), .Z(n2055) );
  XOR U1624 ( .A(n2593), .B(n2592), .Z(n2573) );
  XOR U1625 ( .A(n2113), .B(n2112), .Z(n2130) );
  XOR U1626 ( .A(n2626), .B(n2625), .Z(n2608) );
  XOR U1627 ( .A(n2185), .B(n2184), .Z(n2202) );
  XOR U1628 ( .A(n2669), .B(n2668), .Z(n2651) );
  XOR U1629 ( .A(n2257), .B(n2256), .Z(n2274) );
  XOR U1630 ( .A(n2716), .B(n2715), .Z(n2698) );
  XOR U1631 ( .A(n2379), .B(n2378), .Z(n2361) );
  XOR U1632 ( .A(n2326), .B(n2325), .Z(n2343) );
  XOR U1633 ( .A(n2793), .B(n2792), .Z(n2775) );
  ANDN U1634 ( .A(n634), .B(n633), .Z(n617) );
  XOR U1635 ( .A(n789), .B(n788), .Z(n780) );
  XOR U1636 ( .A(n884), .B(n882), .Z(n924) );
  XOR U1637 ( .A(n1143), .B(n1142), .Z(n1122) );
  XOR U1638 ( .A(n1285), .B(n1284), .Z(n1259) );
  XOR U1639 ( .A(n1359), .B(n1358), .Z(n1332) );
  XOR U1640 ( .A(n1452), .B(n1451), .Z(n1425) );
  XOR U1641 ( .A(n1538), .B(n1537), .Z(n1511) );
  XOR U1642 ( .A(n1721), .B(n1720), .Z(n1694) );
  XOR U1643 ( .A(n1857), .B(n1856), .Z(n1830) );
  XOR U1644 ( .A(n1932), .B(n1931), .Z(n1905) );
  XOR U1645 ( .A(n2004), .B(n2003), .Z(n1977) );
  XOR U1646 ( .A(n2148), .B(n2147), .Z(n2121) );
  XOR U1647 ( .A(n2642), .B(n2640), .Z(n2675) );
  XOR U1648 ( .A(n2220), .B(n2219), .Z(n2193) );
  XOR U1649 ( .A(n2292), .B(n2291), .Z(n2265) );
  XOR U1650 ( .A(n2808), .B(n2807), .Z(n2861) );
  MUX U1651 ( .IN0(o_reg[28]), .IN1(n648), .SEL(n649), .F(n628) );
  AND U1652 ( .A(n706), .B(n707), .Z(n673) );
  MUX U1653 ( .IN0(n773), .IN1(o_reg[24]), .SEL(n774), .F(n737) );
  AND U1654 ( .A(n871), .B(n872), .Z(n814) );
  MUX U1655 ( .IN0(n975), .IN1(o_reg[20]), .SEL(n976), .F(n919) );
  ANDN U1656 ( .A(n1102), .B(n1103), .Z(n1035) );
  MUX U1657 ( .IN0(n1237), .IN1(o_reg[16]), .SEL(n1238), .F(n1167) );
  XNOR U1658 ( .A(n1311), .B(n1394), .Z(n1402) );
  XNOR U1659 ( .A(n1491), .B(n1488), .Z(n1564) );
  MUX U1660 ( .IN0(o_reg[11]), .IN1(n1652), .SEL(n1653), .F(n1562) );
  XNOR U1661 ( .A(n1883), .B(n1812), .Z(n1881) );
  MUX U1662 ( .IN0(o_reg[6]), .IN1(n1761), .SEL(n583), .F(n1757) );
  XOR U1663 ( .A(n2409), .B(n2408), .Z(n2462) );
  OR U1664 ( .A(n613), .B(n614), .Z(n588) );
  MUX U1665 ( .IN0(n3475), .IN1(n532), .SEL(n3476), .F(n3435) );
  IV U1666 ( .A(n3477), .Z(n532) );
  XOR U1667 ( .A(n3521), .B(n3520), .Z(n3535) );
  XOR U1668 ( .A(n3937), .B(n3936), .Z(n3549) );
  MUX U1669 ( .IN0(n3449), .IN1(n3488), .SEL(n3450), .F(n3409) );
  XOR U1670 ( .A(n3481), .B(n3480), .Z(n3495) );
  MUX U1671 ( .IN0(n4298), .IN1(n4309), .SEL(n4299), .F(n4286) );
  MUX U1672 ( .IN0(n4316), .IN1(n533), .SEL(n4317), .F(n4304) );
  IV U1673 ( .A(n4318), .Z(n533) );
  XOR U1674 ( .A(n3919), .B(n3918), .Z(n3509) );
  MUX U1675 ( .IN0(n3877), .IN1(n534), .SEL(n3878), .F(n3859) );
  IV U1676 ( .A(n3879), .Z(n534) );
  XOR U1677 ( .A(n3441), .B(n3440), .Z(n3455) );
  XOR U1678 ( .A(n3901), .B(n3900), .Z(n3469) );
  XNOR U1679 ( .A(n3456), .B(n3419), .Z(n3423) );
  XOR U1680 ( .A(n3401), .B(n3400), .Z(n3415) );
  MUX U1681 ( .IN0(n3315), .IN1(n535), .SEL(n3316), .F(n3275) );
  IV U1682 ( .A(n3317), .Z(n535) );
  MUX U1683 ( .IN0(n4284), .IN1(n536), .SEL(n3891), .F(n4272) );
  IV U1684 ( .A(n3890), .Z(n536) );
  XOR U1685 ( .A(n3883), .B(n3882), .Z(n3429) );
  XOR U1686 ( .A(n3361), .B(n3360), .Z(n3375) );
  XOR U1687 ( .A(n3865), .B(n3864), .Z(n3389) );
  MUX U1688 ( .IN0(n3289), .IN1(n3328), .SEL(n3290), .F(n3249) );
  XOR U1689 ( .A(n3321), .B(n3320), .Z(n3335) );
  MUX U1690 ( .IN0(n4250), .IN1(n4261), .SEL(n4251), .F(n4238) );
  MUX U1691 ( .IN0(n4268), .IN1(n537), .SEL(n4269), .F(n4256) );
  IV U1692 ( .A(n4270), .Z(n537) );
  XOR U1693 ( .A(n3847), .B(n3846), .Z(n3349) );
  XNOR U1694 ( .A(n3336), .B(n3299), .Z(n3303) );
  MUX U1695 ( .IN0(n3805), .IN1(n538), .SEL(n3806), .F(n3787) );
  IV U1696 ( .A(n3807), .Z(n538) );
  XOR U1697 ( .A(n3281), .B(n3280), .Z(n3295) );
  XOR U1698 ( .A(n3829), .B(n3828), .Z(n3309) );
  XOR U1699 ( .A(n3241), .B(n3240), .Z(n3255) );
  MUX U1700 ( .IN0(n4079), .IN1(n4100), .SEL(n4080), .F(n4057) );
  MUX U1701 ( .IN0(n4662), .IN1(n4683), .SEL(n4663), .F(n4640) );
  MUX U1702 ( .IN0(n3155), .IN1(n539), .SEL(n3156), .F(n3115) );
  IV U1703 ( .A(n3157), .Z(n539) );
  MUX U1704 ( .IN0(n4236), .IN1(n540), .SEL(n3819), .F(n4224) );
  IV U1705 ( .A(n3818), .Z(n540) );
  XOR U1706 ( .A(n3811), .B(n3810), .Z(n3269) );
  XOR U1707 ( .A(n3201), .B(n3200), .Z(n3215) );
  XNOR U1708 ( .A(n4408), .B(n4409), .Z(n4096) );
  XOR U1709 ( .A(n3793), .B(n3792), .Z(n3229) );
  XNOR U1710 ( .A(n3216), .B(n3179), .Z(n3183) );
  MUX U1711 ( .IN0(n3129), .IN1(n3168), .SEL(n3130), .F(n3089) );
  XOR U1712 ( .A(n3161), .B(n3160), .Z(n3175) );
  XNOR U1713 ( .A(n4396), .B(n4397), .Z(n4074) );
  MUX U1714 ( .IN0(n4202), .IN1(n4213), .SEL(n4203), .F(n4190) );
  MUX U1715 ( .IN0(n4220), .IN1(n541), .SEL(n4221), .F(n4208) );
  IV U1716 ( .A(n4222), .Z(n541) );
  MUX U1717 ( .IN0(n4998), .IN1(n5003), .SEL(n4999), .F(n4983) );
  XNOR U1718 ( .A(n4802), .B(n4793), .Z(n4637) );
  XOR U1719 ( .A(n3775), .B(n3774), .Z(n3189) );
  MUX U1720 ( .IN0(n3733), .IN1(n542), .SEL(n3734), .F(n3715) );
  IV U1721 ( .A(n3735), .Z(n542) );
  XOR U1722 ( .A(n3121), .B(n3120), .Z(n3135) );
  MUX U1723 ( .IN0(n4376), .IN1(n543), .SEL(n4377), .F(n4364) );
  IV U1724 ( .A(n4378), .Z(n543) );
  XNOR U1725 ( .A(n4061), .B(n4042), .Z(n4046) );
  XNOR U1726 ( .A(n4644), .B(n4625), .Z(n4629) );
  XOR U1727 ( .A(n3757), .B(n3756), .Z(n3149) );
  MUX U1728 ( .IN0(n3991), .IN1(n4012), .SEL(n3992), .F(n3975) );
  XNOR U1729 ( .A(n4372), .B(n4373), .Z(n4030) );
  MUX U1730 ( .IN0(n4142), .IN1(n4145), .SEL(n4143), .F(n4129) );
  MUX U1731 ( .IN0(n4442), .IN1(n4464), .SEL(n4444), .F(n4430) );
  MUX U1732 ( .IN0(n5033), .IN1(n5040), .SEL(n5034), .F(n5029) );
  MUX U1733 ( .IN0(n4961), .IN1(n4976), .SEL(n4963), .F(n4950) );
  MUX U1734 ( .IN0(n4725), .IN1(n4728), .SEL(n4726), .F(n4712) );
  MUX U1735 ( .IN0(n4846), .IN1(n4868), .SEL(n4848), .F(n4834) );
  MUX U1736 ( .IN0(n4768), .IN1(n544), .SEL(n4769), .F(n4756) );
  IV U1737 ( .A(n4770), .Z(n544) );
  XNOR U1738 ( .A(n4776), .B(n4777), .Z(n4613) );
  MUX U1739 ( .IN0(n4574), .IN1(n4595), .SEL(n4575), .F(n4558) );
  MUX U1740 ( .IN0(n3039), .IN1(n545), .SEL(n3040), .F(n2999) );
  IV U1741 ( .A(n3041), .Z(n545) );
  MUX U1742 ( .IN0(n2995), .IN1(n546), .SEL(n2996), .F(n2956) );
  IV U1743 ( .A(n2997), .Z(n546) );
  MUX U1744 ( .IN0(n4188), .IN1(n547), .SEL(n3747), .F(n4176) );
  IV U1745 ( .A(n3746), .Z(n547) );
  XOR U1746 ( .A(n3739), .B(n3738), .Z(n3109) );
  MUX U1747 ( .IN0(n3062), .IN1(n548), .SEL(n3063), .F(n3022) );
  IV U1748 ( .A(n3064), .Z(n548) );
  MUX U1749 ( .IN0(n3018), .IN1(n549), .SEL(n3019), .F(n2947) );
  IV U1750 ( .A(n3020), .Z(n549) );
  MUX U1751 ( .IN0(n3588), .IN1(n3612), .SEL(n3590), .F(n3569) );
  MUX U1752 ( .IN0(n3596), .IN1(n3606), .SEL(n3598), .F(n3578) );
  MUX U1753 ( .IN0(n4346), .IN1(n4357), .SEL(n4347), .F(n4334) );
  XNOR U1754 ( .A(n4504), .B(n4492), .Z(n4158) );
  XNOR U1755 ( .A(n4908), .B(n4896), .Z(n4741) );
  XNOR U1756 ( .A(n4764), .B(n4765), .Z(n4591) );
  XOR U1757 ( .A(n3721), .B(n3720), .Z(n3069) );
  XNOR U1758 ( .A(n3652), .B(n3640), .Z(n3593) );
  XNOR U1759 ( .A(n3674), .B(n3675), .Z(n3559) );
  XNOR U1760 ( .A(n3995), .B(n3968), .Z(n3972) );
  XNOR U1761 ( .A(n4446), .B(n4437), .Z(n4139) );
  MUX U1762 ( .IN0(n769), .IN1(n807), .SEL(n770), .F(n733) );
  MUX U1763 ( .IN0(n800), .IN1(n550), .SEL(n801), .F(n761) );
  IV U1764 ( .A(n802), .Z(n550) );
  MUX U1765 ( .IN0(n943), .IN1(n1002), .SEL(n944), .F(n889) );
  MUX U1766 ( .IN0(n1021), .IN1(n551), .SEL(n1022), .F(n963) );
  IV U1767 ( .A(n1023), .Z(n551) );
  MUX U1768 ( .IN0(n1163), .IN1(n1232), .SEL(n1164), .F(n1096) );
  MUX U1769 ( .IN0(n1108), .IN1(n552), .SEL(n1109), .F(n1041) );
  IV U1770 ( .A(n1110), .Z(n552) );
  MUX U1771 ( .IN0(n1207), .IN1(n1278), .SEL(n1208), .F(n1137) );
  MUX U1772 ( .IN0(n1297), .IN1(n553), .SEL(n1298), .F(n1225) );
  IV U1773 ( .A(n1299), .Z(n553) );
  MUX U1774 ( .IN0(n1253), .IN1(n1325), .SEL(n1254), .F(n1183) );
  MUX U1775 ( .IN0(n1472), .IN1(n1557), .SEL(n1473), .F(n1379) );
  MUX U1776 ( .IN0(n1411), .IN1(n554), .SEL(n1412), .F(n1318) );
  IV U1777 ( .A(n1413), .Z(n554) );
  MUX U1778 ( .IN0(n1532), .IN1(n1621), .SEL(n1533), .F(n1446) );
  MUX U1779 ( .IN0(n1514), .IN1(n1603), .SEL(n1515), .F(n1428) );
  MUX U1780 ( .IN0(n1640), .IN1(n555), .SEL(n1641), .F(n1550) );
  IV U1781 ( .A(n1642), .Z(n555) );
  MUX U1782 ( .IN0(n1595), .IN1(n1687), .SEL(n1596), .F(n1505) );
  MUX U1783 ( .IN0(n1877), .IN1(n1951), .SEL(n1878), .F(n1741) );
  MUX U1784 ( .IN0(n1816), .IN1(n556), .SEL(n1817), .F(n1680) );
  IV U1785 ( .A(n1818), .Z(n556) );
  MUX U1786 ( .IN0(n1926), .IN1(n1997), .SEL(n1927), .F(n1851) );
  MUX U1787 ( .IN0(n1908), .IN1(n1979), .SEL(n1909), .F(n1833) );
  MUX U1788 ( .IN0(n2516), .IN1(n2546), .SEL(n2517), .F(n2487) );
  MUX U1789 ( .IN0(n2016), .IN1(n557), .SEL(n2017), .F(n1944) );
  IV U1790 ( .A(n2018), .Z(n557) );
  MUX U1791 ( .IN0(n1971), .IN1(n2039), .SEL(n1972), .F(n1899) );
  MUX U1792 ( .IN0(n2539), .IN1(n558), .SEL(n2540), .F(n2508) );
  IV U1793 ( .A(n2541), .Z(n558) );
  MUX U1794 ( .IN0(n2168), .IN1(n2239), .SEL(n2169), .F(n2093) );
  MUX U1795 ( .IN0(n2107), .IN1(n559), .SEL(n2108), .F(n2032) );
  IV U1796 ( .A(n2109), .Z(n559) );
  MUX U1797 ( .IN0(n2214), .IN1(n2285), .SEL(n2215), .F(n2142) );
  MUX U1798 ( .IN0(n2196), .IN1(n2267), .SEL(n2197), .F(n2124) );
  MUX U1799 ( .IN0(n2671), .IN1(n2717), .SEL(n2672), .F(n2628) );
  MUX U1800 ( .IN0(n2645), .IN1(n2691), .SEL(n2646), .F(n2602) );
  MUX U1801 ( .IN0(n2304), .IN1(n560), .SEL(n2305), .F(n2232) );
  IV U1802 ( .A(n2306), .Z(n560) );
  MUX U1803 ( .IN0(n2259), .IN1(n2327), .SEL(n2260), .F(n2187) );
  MUX U1804 ( .IN0(n2701), .IN1(n561), .SEL(n2702), .F(n2654) );
  IV U1805 ( .A(n2703), .Z(n561) );
  MUX U1806 ( .IN0(n2710), .IN1(n562), .SEL(n2711), .F(n2663) );
  IV U1807 ( .A(n2712), .Z(n562) );
  MUX U1808 ( .IN0(n3690), .IN1(n4165), .SEL(n3691), .F(n2919) );
  MUX U1809 ( .IN0(n2395), .IN1(n563), .SEL(n2396), .F(n2320) );
  IV U1810 ( .A(n2397), .Z(n563) );
  MUX U1811 ( .IN0(n564), .IN1(n5044), .SEL(n5038), .F(n2456) );
  IV U1812 ( .A(n5039), .Z(n564) );
  MUX U1813 ( .IN0(n4924), .IN1(n4943), .SEL(n4925), .F(n2430) );
  MUX U1814 ( .IN0(n4543), .IN1(n4749), .SEL(n4544), .F(n2412) );
  MUX U1815 ( .IN0(n2892), .IN1(n2963), .SEL(n2893), .F(n2828) );
  MUX U1816 ( .IN0(n2866), .IN1(n2937), .SEL(n2867), .F(n2802) );
  MUX U1817 ( .IN0(n2902), .IN1(n565), .SEL(n2903), .F(n2835) );
  IV U1818 ( .A(n2904), .Z(n565) );
  MUX U1819 ( .IN0(n4172), .IN1(n566), .SEL(n4173), .F(n4160) );
  IV U1820 ( .A(n4174), .Z(n566) );
  XNOR U1821 ( .A(n5006), .B(n4994), .Z(n4935) );
  XNOR U1822 ( .A(n4850), .B(n4841), .Z(n4722) );
  XNOR U1823 ( .A(n4578), .B(n4551), .Z(n4555) );
  XOR U1824 ( .A(n3703), .B(n3702), .Z(n3029) );
  MUX U1825 ( .IN0(n3013), .IN1(n567), .SEL(n3014), .F(n2942) );
  IV U1826 ( .A(n3015), .Z(n567) );
  XNOR U1827 ( .A(n4350), .B(n4341), .Z(n3981) );
  XOR U1828 ( .A(n4135), .B(n4134), .Z(n3686) );
  MUX U1829 ( .IN0(n967), .IN1(n568), .SEL(n968), .F(n911) );
  IV U1830 ( .A(n969), .Z(n568) );
  MUX U1831 ( .IN0(n1229), .IN1(n569), .SEL(n1230), .F(n1159) );
  IV U1832 ( .A(n1231), .Z(n569) );
  MUX U1833 ( .IN0(n1322), .IN1(n570), .SEL(n1323), .F(n1249) );
  IV U1834 ( .A(n1324), .Z(n570) );
  MUX U1835 ( .IN0(n1554), .IN1(n571), .SEL(n1555), .F(n1468) );
  IV U1836 ( .A(n1556), .Z(n571) );
  MUX U1837 ( .IN0(n1684), .IN1(n572), .SEL(n1685), .F(n1591) );
  IV U1838 ( .A(n1686), .Z(n572) );
  MUX U1839 ( .IN0(n2493), .IN1(n2521), .SEL(n2494), .F(n2464) );
  MUX U1840 ( .IN0(n1948), .IN1(n573), .SEL(n1949), .F(n1873) );
  IV U1841 ( .A(n1950), .Z(n573) );
  MUX U1842 ( .IN0(n2530), .IN1(n574), .SEL(n2531), .F(n2501) );
  IV U1843 ( .A(n2532), .Z(n574) );
  MUX U1844 ( .IN0(n2036), .IN1(n575), .SEL(n2037), .F(n1967) );
  IV U1845 ( .A(n2038), .Z(n575) );
  MUX U1846 ( .IN0(n2236), .IN1(n576), .SEL(n2237), .F(n2164) );
  IV U1847 ( .A(n2238), .Z(n576) );
  MUX U1848 ( .IN0(n2324), .IN1(n577), .SEL(n2325), .F(n2255) );
  IV U1849 ( .A(n2326), .Z(n577) );
  XOR U1850 ( .A(n4718), .B(n4717), .Z(n4539) );
  XOR U1851 ( .A(n2979), .B(n2978), .Z(n2989) );
  XOR U1852 ( .A(n3955), .B(n3954), .Z(n3684) );
  MUX U1853 ( .IN0(n712), .IN1(n745), .SEL(n713), .F(n685) );
  XNOR U1854 ( .A(n690), .B(n660), .Z(n664) );
  XNOR U1855 ( .A(n844), .B(n792), .Z(n796) );
  MUX U1856 ( .IN0(n928), .IN1(n578), .SEL(n929), .F(n875) );
  IV U1857 ( .A(n930), .Z(n578) );
  XNOR U1858 ( .A(n1010), .B(n955), .Z(n959) );
  MUX U1859 ( .IN0(n1124), .IN1(n1191), .SEL(n1125), .F(n1063) );
  XNOR U1860 ( .A(n1286), .B(n1217), .Z(n1221) );
  XNOR U1861 ( .A(n1269), .B(n1200), .Z(n1203) );
  XNOR U1862 ( .A(n1539), .B(n1456), .Z(n1460) );
  XNOR U1863 ( .A(n1521), .B(n1438), .Z(n1442) );
  XNOR U1864 ( .A(n1798), .B(n1660), .Z(n1664) );
  XNOR U1865 ( .A(n1858), .B(n1725), .Z(n1729) );
  XNOR U1866 ( .A(n1840), .B(n1707), .Z(n1711) );
  XNOR U1867 ( .A(n2074), .B(n2008), .Z(n2012) );
  XNOR U1868 ( .A(n2056), .B(n1990), .Z(n1994) );
  XNOR U1869 ( .A(n2293), .B(n2224), .Z(n2228) );
  XNOR U1870 ( .A(n2275), .B(n2206), .Z(n2210) );
  MUX U1871 ( .IN0(n2855), .IN1(n2926), .SEL(n2857), .F(n2758) );
  XNOR U1872 ( .A(n5020), .B(n2449), .Z(n2453) );
  XNOR U1873 ( .A(n4936), .B(n2440), .Z(n2444) );
  XNOR U1874 ( .A(n4742), .B(n2422), .Z(n2426) );
  XNOR U1875 ( .A(n2882), .B(n2821), .Z(n2825) );
  XNOR U1876 ( .A(n2873), .B(n2812), .Z(n2816) );
  XOR U1877 ( .A(n4527), .B(n4526), .Z(n4535) );
  XOR U1878 ( .A(n2908), .B(n2907), .Z(n2925) );
  XOR U1879 ( .A(n3575), .B(n3574), .Z(n2968) );
  XOR U1880 ( .A(n698), .B(n697), .Z(n689) );
  XOR U1881 ( .A(n806), .B(n805), .Z(n789) );
  MUX U1882 ( .IN0(n878), .IN1(n931), .SEL(n879), .F(n828) );
  XOR U1883 ( .A(n863), .B(n862), .Z(n843) );
  XOR U1884 ( .A(n989), .B(n988), .Z(n1000) );
  XOR U1885 ( .A(n2635), .B(n2634), .Z(n2641) );
  XOR U1886 ( .A(n2681), .B(n2680), .Z(n2687) );
  XOR U1887 ( .A(n2730), .B(n2729), .Z(n2738) );
  XOR U1888 ( .A(n2749), .B(n2748), .Z(n2766) );
  XOR U1889 ( .A(n2401), .B(n2400), .Z(n2418) );
  XOR U1890 ( .A(n2841), .B(n2840), .Z(n2854) );
  XOR U1891 ( .A(n4537), .B(n4538), .Z(n2933) );
  XOR U1892 ( .A(n2872), .B(n2871), .Z(n2916) );
  MUX U1893 ( .IN0(n624), .IN1(n643), .SEL(n625), .F(n594) );
  XOR U1894 ( .A(n718), .B(n717), .Z(n709) );
  XOR U1895 ( .A(n1009), .B(n1008), .Z(n997) );
  MUX U1896 ( .IN0(n1484), .IN1(n1573), .SEL(n1485), .F(n1394) );
  XOR U1897 ( .A(n1565), .B(n1566), .Z(n1582) );
  XOR U1898 ( .A(n1797), .B(n1796), .Z(n1882) );
  XOR U1899 ( .A(n2470), .B(n2469), .Z(n1886) );
  XOR U1900 ( .A(n2499), .B(n2498), .Z(n1958) );
  XOR U1901 ( .A(n2528), .B(n2527), .Z(n2098) );
  XOR U1902 ( .A(n2573), .B(n2572), .Z(n2102) );
  XOR U1903 ( .A(n2608), .B(n2607), .Z(n2174) );
  XOR U1904 ( .A(n2651), .B(n2650), .Z(n2246) );
  XOR U1905 ( .A(n2698), .B(n2697), .Z(n2386) );
  XOR U1906 ( .A(n2775), .B(n2774), .Z(n2390) );
  XOR U1907 ( .A(n618), .B(n617), .Z(n631) );
  ANDN U1908 ( .A(n673), .B(n674), .Z(n650) );
  MUX U1909 ( .IN0(n704), .IN1(o_reg[26]), .SEL(n705), .F(n671) );
  XOR U1910 ( .A(n742), .B(n743), .Z(n776) );
  MUX U1911 ( .IN0(n869), .IN1(o_reg[22]), .SEL(n870), .F(n812) );
  XOR U1912 ( .A(n886), .B(n885), .Z(n922) );
  XOR U1913 ( .A(n940), .B(n939), .Z(n978) );
  XOR U1914 ( .A(n1055), .B(n1054), .Z(n1103) );
  XOR U1915 ( .A(n1122), .B(n1121), .Z(n1170) );
  XOR U1916 ( .A(n1189), .B(n1188), .Z(n1240) );
  XOR U1917 ( .A(n1259), .B(n1258), .Z(n1313) );
  XOR U1918 ( .A(n1332), .B(n1331), .Z(n1406) );
  XOR U1919 ( .A(n1425), .B(n1424), .Z(n1490) );
  XOR U1920 ( .A(n1511), .B(n1510), .Z(n1580) );
  XOR U1921 ( .A(n1601), .B(n1600), .Z(n1673) );
  XOR U1922 ( .A(n1694), .B(n1693), .Z(n1747) );
  XOR U1923 ( .A(n1830), .B(n1829), .Z(n1751) );
  XOR U1924 ( .A(n1905), .B(n1904), .Z(n1755) );
  XOR U1925 ( .A(n1977), .B(n1976), .Z(n1759) );
  XOR U1926 ( .A(n2046), .B(n2045), .Z(n1763) );
  XOR U1927 ( .A(n2121), .B(n2120), .Z(n1767) );
  XOR U1928 ( .A(n2193), .B(n2192), .Z(n1771) );
  XOR U1929 ( .A(n2265), .B(n2264), .Z(n1775) );
  XOR U1930 ( .A(n2334), .B(n2333), .Z(n1779) );
  XOR U1931 ( .A(n2462), .B(n1781), .Z(n2862) );
  MUX U1932 ( .IN0(o_reg[31]), .IN1(n586), .SEL(n587), .F(o[31]) );
  XOR U1933 ( .A(o_reg[10]), .B(n579), .Z(o[9]) );
  XNOR U1934 ( .A(o_reg[9]), .B(n580), .Z(o[8]) );
  XNOR U1935 ( .A(o_reg[8]), .B(n581), .Z(o[7]) );
  XOR U1936 ( .A(n582), .B(o_reg[7]), .Z(o[6]) );
  XNOR U1937 ( .A(o_reg[6]), .B(n583), .Z(o[5]) );
  XNOR U1938 ( .A(o_reg[5]), .B(n584), .Z(o[4]) );
  XNOR U1939 ( .A(o_reg[4]), .B(n585), .Z(o[3]) );
  XNOR U1940 ( .A(n587), .B(o_reg[31]), .Z(o[30]) );
  XNOR U1941 ( .A(n588), .B(n589), .Z(n587) );
  XOR U1942 ( .A(n590), .B(n591), .Z(n589) );
  XOR U1943 ( .A(n592), .B(n593), .Z(n591) );
  XOR U1944 ( .A(n594), .B(n586), .Z(n593) );
  XOR U1945 ( .A(n597), .B(n598), .Z(n592) );
  XOR U1946 ( .A(n599), .B(n600), .Z(n590) );
  XNOR U1947 ( .A(n601), .B(n602), .Z(n600) );
  AND U1948 ( .A(n603), .B(n604), .Z(n602) );
  NAND U1949 ( .A(n605), .B(n594), .Z(n604) );
  NANDN U1950 ( .B(n606), .A(n607), .Z(n603) );
  XOR U1951 ( .A(n608), .B(n609), .Z(n599) );
  NOR U1952 ( .A(n612), .B(n601), .Z(n608) );
  XOR U1953 ( .A(n615), .B(o_reg[3]), .Z(o[2]) );
  XOR U1954 ( .A(o_reg[30]), .B(n596), .Z(o[29]) );
  XOR U1955 ( .A(n616), .B(n614), .Z(n596) );
  XNOR U1956 ( .A(n611), .B(n597), .Z(n614) );
  IV U1957 ( .A(n610), .Z(n597) );
  XOR U1958 ( .A(n612), .B(n601), .Z(n611) );
  OR U1959 ( .A(n619), .B(n620), .Z(n601) );
  XNOR U1960 ( .A(n606), .B(n598), .Z(n612) );
  IV U1961 ( .A(n607), .Z(n598) );
  XNOR U1962 ( .A(n594), .B(n605), .Z(n606) );
  NAND U1963 ( .A(g_input[31]), .B(e_input[31]), .Z(n605) );
  XNOR U1964 ( .A(n627), .B(n624), .Z(n625) );
  XOR U1965 ( .A(n613), .B(n595), .Z(n616) );
  XOR U1966 ( .A(o_reg[29]), .B(n629), .Z(o[28]) );
  XOR U1967 ( .A(n632), .B(n631), .Z(n629) );
  XNOR U1968 ( .A(n619), .B(n620), .Z(n618) );
  NANDN U1969 ( .B(n635), .A(n636), .Z(n620) );
  XOR U1970 ( .A(n621), .B(n637), .Z(n622) );
  ANDN U1971 ( .A(n638), .B(n639), .Z(n637) );
  XNOR U1972 ( .A(n626), .B(n627), .Z(n623) );
  NAND U1973 ( .A(e_input[31]), .B(g_input[30]), .Z(n627) );
  XNOR U1974 ( .A(n624), .B(n643), .Z(n626) );
  AND U1975 ( .A(g_input[31]), .B(e_input[30]), .Z(n643) );
  XNOR U1976 ( .A(n647), .B(n644), .Z(n645) );
  XNOR U1977 ( .A(n630), .B(n628), .Z(n632) );
  XNOR U1978 ( .A(o_reg[28]), .B(n649), .Z(o[27]) );
  XNOR U1979 ( .A(n652), .B(n651), .Z(n649) );
  XOR U1980 ( .A(n634), .B(n633), .Z(n651) );
  OR U1981 ( .A(n653), .B(n654), .Z(n633) );
  XNOR U1982 ( .A(n635), .B(n636), .Z(n634) );
  XNOR U1983 ( .A(n662), .B(n639), .Z(n658) );
  NAND U1984 ( .A(e_input[29]), .B(g_input[31]), .Z(n639) );
  IV U1985 ( .A(n640), .Z(n662) );
  XNOR U1986 ( .A(n646), .B(n647), .Z(n642) );
  NAND U1987 ( .A(e_input[31]), .B(g_input[29]), .Z(n647) );
  XNOR U1988 ( .A(n644), .B(n666), .Z(n646) );
  AND U1989 ( .A(g_input[30]), .B(e_input[30]), .Z(n666) );
  XNOR U1990 ( .A(n670), .B(n667), .Z(n668) );
  XNOR U1991 ( .A(n650), .B(n648), .Z(n652) );
  XNOR U1992 ( .A(n672), .B(o_reg[27]), .Z(o[26]) );
  XNOR U1993 ( .A(n675), .B(n674), .Z(n672) );
  XNOR U1994 ( .A(n654), .B(n653), .Z(n674) );
  OR U1995 ( .A(n676), .B(n677), .Z(n653) );
  XNOR U1996 ( .A(n657), .B(n656), .Z(n654) );
  XNOR U1997 ( .A(n678), .B(n679), .Z(n656) );
  XOR U1998 ( .A(n680), .B(n681), .Z(n679) );
  AND U1999 ( .A(n682), .B(n683), .Z(n680) );
  NAND U2000 ( .A(n684), .B(n685), .Z(n683) );
  NANDN U2001 ( .B(n686), .A(n681), .Z(n682) );
  XOR U2002 ( .A(n659), .B(n691), .Z(n660) );
  AND U2003 ( .A(g_input[31]), .B(e_input[28]), .Z(n691) );
  XNOR U2004 ( .A(n695), .B(n661), .Z(n690) );
  NAND U2005 ( .A(e_input[29]), .B(g_input[30]), .Z(n661) );
  IV U2006 ( .A(n663), .Z(n695) );
  XNOR U2007 ( .A(n669), .B(n670), .Z(n665) );
  NAND U2008 ( .A(e_input[31]), .B(g_input[28]), .Z(n670) );
  XNOR U2009 ( .A(n667), .B(n699), .Z(n669) );
  AND U2010 ( .A(g_input[29]), .B(e_input[30]), .Z(n699) );
  XNOR U2011 ( .A(n703), .B(n700), .Z(n701) );
  XNOR U2012 ( .A(n673), .B(n671), .Z(n675) );
  XOR U2013 ( .A(o_reg[26]), .B(n705), .Z(o[25]) );
  XNOR U2014 ( .A(n708), .B(n707), .Z(n705) );
  XOR U2015 ( .A(n676), .B(n677), .Z(n707) );
  OR U2016 ( .A(n709), .B(n710), .Z(n677) );
  XNOR U2017 ( .A(n711), .B(n686), .Z(n688) );
  XNOR U2018 ( .A(n685), .B(n684), .Z(n686) );
  NAND U2019 ( .A(g_input[31]), .B(e_input[27]), .Z(n684) );
  XNOR U2020 ( .A(n715), .B(n712), .Z(n713) );
  XNOR U2021 ( .A(n681), .B(n687), .Z(n711) );
  XNOR U2022 ( .A(n719), .B(n722), .Z(n721) );
  XOR U2023 ( .A(n692), .B(n724), .Z(n693) );
  AND U2024 ( .A(g_input[30]), .B(e_input[28]), .Z(n724) );
  XNOR U2025 ( .A(n728), .B(n694), .Z(n723) );
  NAND U2026 ( .A(e_input[29]), .B(g_input[29]), .Z(n694) );
  IV U2027 ( .A(n696), .Z(n728) );
  XNOR U2028 ( .A(n702), .B(n703), .Z(n698) );
  NAND U2029 ( .A(e_input[31]), .B(g_input[27]), .Z(n703) );
  XNOR U2030 ( .A(n700), .B(n732), .Z(n702) );
  AND U2031 ( .A(g_input[28]), .B(e_input[30]), .Z(n732) );
  XNOR U2032 ( .A(n736), .B(n733), .Z(n734) );
  XNOR U2033 ( .A(n706), .B(n704), .Z(n708) );
  XOR U2034 ( .A(o_reg[25]), .B(n738), .Z(o[24]) );
  XNOR U2035 ( .A(n741), .B(n740), .Z(n738) );
  XOR U2036 ( .A(n709), .B(n710), .Z(n740) );
  NANDN U2037 ( .B(n742), .A(n743), .Z(n710) );
  XOR U2038 ( .A(n744), .B(n722), .Z(n717) );
  XNOR U2039 ( .A(n714), .B(n715), .Z(n722) );
  NAND U2040 ( .A(e_input[27]), .B(g_input[30]), .Z(n715) );
  XNOR U2041 ( .A(n712), .B(n745), .Z(n714) );
  AND U2042 ( .A(g_input[31]), .B(e_input[26]), .Z(n745) );
  XNOR U2043 ( .A(n749), .B(n746), .Z(n747) );
  XNOR U2044 ( .A(n720), .B(n716), .Z(n744) );
  XOR U2045 ( .A(n719), .B(n753), .Z(n720) );
  ANDN U2046 ( .A(n754), .B(n755), .Z(n753) );
  XOR U2047 ( .A(n725), .B(n760), .Z(n726) );
  AND U2048 ( .A(g_input[29]), .B(e_input[28]), .Z(n760) );
  XNOR U2049 ( .A(n764), .B(n727), .Z(n759) );
  NAND U2050 ( .A(e_input[29]), .B(g_input[28]), .Z(n727) );
  IV U2051 ( .A(n729), .Z(n764) );
  XNOR U2052 ( .A(n735), .B(n736), .Z(n731) );
  NAND U2053 ( .A(e_input[31]), .B(g_input[26]), .Z(n736) );
  XNOR U2054 ( .A(n733), .B(n768), .Z(n735) );
  AND U2055 ( .A(g_input[27]), .B(e_input[30]), .Z(n768) );
  XNOR U2056 ( .A(n772), .B(n769), .Z(n770) );
  XNOR U2057 ( .A(n739), .B(n737), .Z(n741) );
  XOR U2058 ( .A(o_reg[24]), .B(n774), .Z(o[23]) );
  XOR U2059 ( .A(n777), .B(n776), .Z(n774) );
  XOR U2060 ( .A(n781), .B(n758), .Z(n751) );
  XNOR U2061 ( .A(n748), .B(n749), .Z(n758) );
  NAND U2062 ( .A(e_input[27]), .B(g_input[29]), .Z(n749) );
  XNOR U2063 ( .A(n746), .B(n782), .Z(n748) );
  AND U2064 ( .A(g_input[30]), .B(e_input[26]), .Z(n782) );
  XNOR U2065 ( .A(n786), .B(n783), .Z(n784) );
  XNOR U2066 ( .A(n757), .B(n750), .Z(n781) );
  XNOR U2067 ( .A(n794), .B(n755), .Z(n790) );
  NAND U2068 ( .A(e_input[25]), .B(g_input[31]), .Z(n755) );
  IV U2069 ( .A(n756), .Z(n794) );
  XOR U2070 ( .A(n761), .B(n799), .Z(n762) );
  AND U2071 ( .A(g_input[28]), .B(e_input[28]), .Z(n799) );
  XNOR U2072 ( .A(n803), .B(n763), .Z(n798) );
  NAND U2073 ( .A(e_input[29]), .B(g_input[27]), .Z(n763) );
  IV U2074 ( .A(n765), .Z(n803) );
  XNOR U2075 ( .A(n771), .B(n772), .Z(n767) );
  NAND U2076 ( .A(e_input[31]), .B(g_input[25]), .Z(n772) );
  XNOR U2077 ( .A(n769), .B(n807), .Z(n771) );
  AND U2078 ( .A(g_input[26]), .B(e_input[30]), .Z(n807) );
  XNOR U2079 ( .A(n811), .B(n808), .Z(n809) );
  XNOR U2080 ( .A(n775), .B(n773), .Z(n777) );
  XNOR U2081 ( .A(n813), .B(o_reg[23]), .Z(o[22]) );
  XOR U2082 ( .A(n816), .B(n815), .Z(n813) );
  XNOR U2083 ( .A(n780), .B(n779), .Z(n815) );
  XOR U2084 ( .A(n817), .B(n818), .Z(n779) );
  XOR U2085 ( .A(n819), .B(n820), .Z(n818) );
  AND U2086 ( .A(n821), .B(n822), .Z(n819) );
  OR U2087 ( .A(n823), .B(n824), .Z(n822) );
  AND U2088 ( .A(n825), .B(n826), .Z(n821) );
  NAND U2089 ( .A(n827), .B(n828), .Z(n826) );
  NANDN U2090 ( .B(n829), .A(n820), .Z(n825) );
  XOR U2091 ( .A(n830), .B(n831), .Z(n778) );
  ANDN U2092 ( .A(n832), .B(n833), .Z(n831) );
  XNOR U2093 ( .A(n830), .B(n834), .Z(n832) );
  XOR U2094 ( .A(n835), .B(n797), .Z(n788) );
  XNOR U2095 ( .A(n785), .B(n786), .Z(n797) );
  NAND U2096 ( .A(e_input[27]), .B(g_input[28]), .Z(n786) );
  XNOR U2097 ( .A(n783), .B(n836), .Z(n785) );
  AND U2098 ( .A(g_input[29]), .B(e_input[26]), .Z(n836) );
  XNOR U2099 ( .A(n840), .B(n837), .Z(n838) );
  XNOR U2100 ( .A(n796), .B(n787), .Z(n835) );
  XOR U2101 ( .A(n791), .B(n845), .Z(n792) );
  AND U2102 ( .A(g_input[31]), .B(e_input[24]), .Z(n845) );
  XOR U2103 ( .A(n846), .B(n847), .Z(n791) );
  AND U2104 ( .A(n848), .B(n849), .Z(n847) );
  XNOR U2105 ( .A(n850), .B(n846), .Z(n848) );
  XNOR U2106 ( .A(n851), .B(n793), .Z(n844) );
  NAND U2107 ( .A(e_input[25]), .B(g_input[30]), .Z(n793) );
  IV U2108 ( .A(n795), .Z(n851) );
  XOR U2109 ( .A(n800), .B(n856), .Z(n801) );
  AND U2110 ( .A(g_input[27]), .B(e_input[28]), .Z(n856) );
  XNOR U2111 ( .A(n860), .B(n802), .Z(n855) );
  NAND U2112 ( .A(e_input[29]), .B(g_input[26]), .Z(n802) );
  IV U2113 ( .A(n804), .Z(n860) );
  XNOR U2114 ( .A(n810), .B(n811), .Z(n806) );
  NAND U2115 ( .A(e_input[31]), .B(g_input[24]), .Z(n811) );
  XNOR U2116 ( .A(n808), .B(n864), .Z(n810) );
  AND U2117 ( .A(g_input[25]), .B(e_input[30]), .Z(n864) );
  XNOR U2118 ( .A(n868), .B(n865), .Z(n866) );
  XNOR U2119 ( .A(n814), .B(n812), .Z(n816) );
  XOR U2120 ( .A(o_reg[22]), .B(n870), .Z(o[21]) );
  XNOR U2121 ( .A(n873), .B(n872), .Z(n870) );
  XOR U2122 ( .A(n834), .B(n833), .Z(n872) );
  XNOR U2123 ( .A(n874), .B(n824), .Z(n833) );
  XNOR U2124 ( .A(n829), .B(n820), .Z(n824) );
  XNOR U2125 ( .A(n828), .B(n827), .Z(n829) );
  NAND U2126 ( .A(g_input[31]), .B(e_input[23]), .Z(n827) );
  XNOR U2127 ( .A(n881), .B(n878), .Z(n879) );
  OR U2128 ( .A(n882), .B(n883), .Z(n823) );
  XOR U2129 ( .A(n887), .B(n854), .Z(n842) );
  XNOR U2130 ( .A(n839), .B(n840), .Z(n854) );
  NAND U2131 ( .A(e_input[27]), .B(g_input[27]), .Z(n840) );
  XNOR U2132 ( .A(n837), .B(n888), .Z(n839) );
  AND U2133 ( .A(g_input[28]), .B(e_input[26]), .Z(n888) );
  XNOR U2134 ( .A(n892), .B(n889), .Z(n890) );
  XNOR U2135 ( .A(n853), .B(n841), .Z(n887) );
  XOR U2136 ( .A(n846), .B(n897), .Z(n849) );
  AND U2137 ( .A(g_input[30]), .B(e_input[24]), .Z(n897) );
  XNOR U2138 ( .A(n901), .B(n850), .Z(n896) );
  NAND U2139 ( .A(e_input[25]), .B(g_input[29]), .Z(n850) );
  IV U2140 ( .A(n852), .Z(n901) );
  XOR U2141 ( .A(n857), .B(n906), .Z(n858) );
  AND U2142 ( .A(g_input[26]), .B(e_input[28]), .Z(n906) );
  XNOR U2143 ( .A(n910), .B(n859), .Z(n905) );
  NAND U2144 ( .A(e_input[29]), .B(g_input[25]), .Z(n859) );
  IV U2145 ( .A(n861), .Z(n910) );
  XNOR U2146 ( .A(n867), .B(n868), .Z(n863) );
  NAND U2147 ( .A(e_input[31]), .B(g_input[23]), .Z(n868) );
  XNOR U2148 ( .A(n865), .B(n914), .Z(n867) );
  AND U2149 ( .A(g_input[24]), .B(e_input[30]), .Z(n914) );
  XNOR U2150 ( .A(n918), .B(n915), .Z(n916) );
  XNOR U2151 ( .A(n871), .B(n869), .Z(n873) );
  XOR U2152 ( .A(o_reg[21]), .B(n920), .Z(o[20]) );
  XOR U2153 ( .A(n923), .B(n922), .Z(n920) );
  XOR U2154 ( .A(n924), .B(n883), .Z(n885) );
  XOR U2155 ( .A(n875), .B(n925), .Z(n876) );
  ANDN U2156 ( .A(n926), .B(n927), .Z(n925) );
  XNOR U2157 ( .A(n880), .B(n881), .Z(n877) );
  NAND U2158 ( .A(e_input[23]), .B(g_input[30]), .Z(n881) );
  XNOR U2159 ( .A(n878), .B(n931), .Z(n880) );
  AND U2160 ( .A(g_input[31]), .B(e_input[22]), .Z(n931) );
  XNOR U2161 ( .A(n935), .B(n932), .Z(n933) );
  NANDN U2162 ( .B(n936), .A(n937), .Z(n882) );
  XOR U2163 ( .A(n941), .B(n904), .Z(n894) );
  XNOR U2164 ( .A(n891), .B(n892), .Z(n904) );
  NAND U2165 ( .A(e_input[27]), .B(g_input[26]), .Z(n892) );
  XNOR U2166 ( .A(n889), .B(n942), .Z(n891) );
  AND U2167 ( .A(g_input[27]), .B(e_input[26]), .Z(n942) );
  XNOR U2168 ( .A(n946), .B(n943), .Z(n944) );
  XNOR U2169 ( .A(n903), .B(n893), .Z(n941) );
  XOR U2170 ( .A(n947), .B(n948), .Z(n893) );
  AND U2171 ( .A(n949), .B(n950), .Z(n948) );
  XNOR U2172 ( .A(n947), .B(n951), .Z(n949) );
  XOR U2173 ( .A(n898), .B(n953), .Z(n899) );
  AND U2174 ( .A(g_input[29]), .B(e_input[24]), .Z(n953) );
  XNOR U2175 ( .A(n957), .B(n900), .Z(n952) );
  NAND U2176 ( .A(e_input[25]), .B(g_input[28]), .Z(n900) );
  IV U2177 ( .A(n902), .Z(n957) );
  XOR U2178 ( .A(n907), .B(n962), .Z(n908) );
  AND U2179 ( .A(g_input[25]), .B(e_input[28]), .Z(n962) );
  XNOR U2180 ( .A(n966), .B(n909), .Z(n961) );
  NAND U2181 ( .A(e_input[29]), .B(g_input[24]), .Z(n909) );
  IV U2182 ( .A(n911), .Z(n966) );
  XNOR U2183 ( .A(n917), .B(n918), .Z(n913) );
  NAND U2184 ( .A(e_input[31]), .B(g_input[22]), .Z(n918) );
  XNOR U2185 ( .A(n915), .B(n970), .Z(n917) );
  AND U2186 ( .A(g_input[23]), .B(e_input[30]), .Z(n970) );
  XNOR U2187 ( .A(n974), .B(n971), .Z(n972) );
  XNOR U2188 ( .A(n921), .B(n919), .Z(n923) );
  XNOR U2189 ( .A(o_reg[2]), .B(n979), .Z(o[1]) );
  XOR U2190 ( .A(o_reg[20]), .B(n976), .Z(o[19]) );
  XOR U2191 ( .A(n980), .B(n978), .Z(n976) );
  XOR U2192 ( .A(n981), .B(n936), .Z(n939) );
  XNOR U2193 ( .A(n986), .B(n927), .Z(n982) );
  NAND U2194 ( .A(e_input[21]), .B(g_input[31]), .Z(n927) );
  IV U2195 ( .A(n928), .Z(n986) );
  XNOR U2196 ( .A(n934), .B(n935), .Z(n930) );
  NAND U2197 ( .A(e_input[23]), .B(g_input[29]), .Z(n935) );
  XNOR U2198 ( .A(n932), .B(n990), .Z(n934) );
  AND U2199 ( .A(g_input[30]), .B(e_input[22]), .Z(n990) );
  XNOR U2200 ( .A(n994), .B(n991), .Z(n992) );
  XNOR U2201 ( .A(n937), .B(n938), .Z(n981) );
  XOR U2202 ( .A(n1001), .B(n960), .Z(n950) );
  XNOR U2203 ( .A(n945), .B(n946), .Z(n960) );
  NAND U2204 ( .A(e_input[27]), .B(g_input[25]), .Z(n946) );
  XNOR U2205 ( .A(n943), .B(n1002), .Z(n945) );
  AND U2206 ( .A(g_input[26]), .B(e_input[26]), .Z(n1002) );
  XNOR U2207 ( .A(n1006), .B(n1003), .Z(n1004) );
  XNOR U2208 ( .A(n959), .B(n947), .Z(n1001) );
  XOR U2209 ( .A(n954), .B(n1011), .Z(n955) );
  AND U2210 ( .A(g_input[28]), .B(e_input[24]), .Z(n1011) );
  XNOR U2211 ( .A(n1015), .B(n956), .Z(n1010) );
  NAND U2212 ( .A(e_input[25]), .B(g_input[27]), .Z(n956) );
  IV U2213 ( .A(n958), .Z(n1015) );
  XOR U2214 ( .A(n963), .B(n1020), .Z(n964) );
  AND U2215 ( .A(g_input[24]), .B(e_input[28]), .Z(n1020) );
  XNOR U2216 ( .A(n1024), .B(n965), .Z(n1019) );
  NAND U2217 ( .A(e_input[29]), .B(g_input[23]), .Z(n965) );
  IV U2218 ( .A(n967), .Z(n1024) );
  XNOR U2219 ( .A(n973), .B(n974), .Z(n969) );
  NAND U2220 ( .A(e_input[31]), .B(g_input[21]), .Z(n974) );
  XNOR U2221 ( .A(n971), .B(n1028), .Z(n973) );
  AND U2222 ( .A(g_input[22]), .B(e_input[30]), .Z(n1028) );
  XNOR U2223 ( .A(n1032), .B(n1029), .Z(n1030) );
  XNOR U2224 ( .A(n977), .B(n975), .Z(n980) );
  XNOR U2225 ( .A(n1034), .B(o_reg[19]), .Z(o[18]) );
  XOR U2226 ( .A(n1037), .B(n1036), .Z(n1034) );
  XNOR U2227 ( .A(n997), .B(n996), .Z(n1036) );
  XNOR U2228 ( .A(n1038), .B(n1000), .Z(n996) );
  XOR U2229 ( .A(n983), .B(n1040), .Z(n984) );
  AND U2230 ( .A(g_input[31]), .B(e_input[20]), .Z(n1040) );
  XNOR U2231 ( .A(n1044), .B(n985), .Z(n1039) );
  NAND U2232 ( .A(e_input[21]), .B(g_input[30]), .Z(n985) );
  IV U2233 ( .A(n987), .Z(n1044) );
  XNOR U2234 ( .A(n993), .B(n994), .Z(n989) );
  NAND U2235 ( .A(e_input[23]), .B(g_input[28]), .Z(n994) );
  XNOR U2236 ( .A(n991), .B(n1048), .Z(n993) );
  AND U2237 ( .A(g_input[29]), .B(e_input[22]), .Z(n1048) );
  XNOR U2238 ( .A(n1052), .B(n1049), .Z(n1050) );
  XNOR U2239 ( .A(n999), .B(n995), .Z(n1038) );
  XNOR U2240 ( .A(n1056), .B(n1057), .Z(n999) );
  XOR U2241 ( .A(n1058), .B(n1059), .Z(n1057) );
  AND U2242 ( .A(n1060), .B(n1061), .Z(n1058) );
  NAND U2243 ( .A(n1062), .B(n1063), .Z(n1061) );
  NANDN U2244 ( .B(n1064), .A(n1059), .Z(n1060) );
  XOR U2245 ( .A(n1068), .B(n1018), .Z(n1008) );
  XNOR U2246 ( .A(n1005), .B(n1006), .Z(n1018) );
  NAND U2247 ( .A(e_input[27]), .B(g_input[24]), .Z(n1006) );
  XNOR U2248 ( .A(n1003), .B(n1069), .Z(n1005) );
  AND U2249 ( .A(g_input[25]), .B(e_input[26]), .Z(n1069) );
  XNOR U2250 ( .A(n1073), .B(n1070), .Z(n1071) );
  XNOR U2251 ( .A(n1017), .B(n1007), .Z(n1068) );
  XOR U2252 ( .A(n1012), .B(n1078), .Z(n1013) );
  AND U2253 ( .A(g_input[27]), .B(e_input[24]), .Z(n1078) );
  XNOR U2254 ( .A(n1082), .B(n1014), .Z(n1077) );
  NAND U2255 ( .A(e_input[25]), .B(g_input[26]), .Z(n1014) );
  IV U2256 ( .A(n1016), .Z(n1082) );
  XOR U2257 ( .A(n1021), .B(n1087), .Z(n1022) );
  AND U2258 ( .A(g_input[23]), .B(e_input[28]), .Z(n1087) );
  XNOR U2259 ( .A(n1091), .B(n1023), .Z(n1086) );
  NAND U2260 ( .A(e_input[29]), .B(g_input[22]), .Z(n1023) );
  IV U2261 ( .A(n1025), .Z(n1091) );
  XNOR U2262 ( .A(n1031), .B(n1032), .Z(n1027) );
  NAND U2263 ( .A(e_input[31]), .B(g_input[20]), .Z(n1032) );
  XNOR U2264 ( .A(n1029), .B(n1095), .Z(n1031) );
  AND U2265 ( .A(g_input[21]), .B(e_input[30]), .Z(n1095) );
  XNOR U2266 ( .A(n1099), .B(n1096), .Z(n1097) );
  XNOR U2267 ( .A(n1035), .B(n1033), .Z(n1037) );
  XOR U2268 ( .A(o_reg[18]), .B(n1101), .Z(o[17]) );
  XOR U2269 ( .A(n1104), .B(n1103), .Z(n1101) );
  XOR U2270 ( .A(n1105), .B(n1067), .Z(n1054) );
  XOR U2271 ( .A(n1041), .B(n1107), .Z(n1042) );
  AND U2272 ( .A(g_input[30]), .B(e_input[20]), .Z(n1107) );
  XNOR U2273 ( .A(n1111), .B(n1043), .Z(n1106) );
  NAND U2274 ( .A(e_input[21]), .B(g_input[29]), .Z(n1043) );
  IV U2275 ( .A(n1045), .Z(n1111) );
  XNOR U2276 ( .A(n1051), .B(n1052), .Z(n1047) );
  NAND U2277 ( .A(e_input[23]), .B(g_input[27]), .Z(n1052) );
  XNOR U2278 ( .A(n1049), .B(n1115), .Z(n1051) );
  AND U2279 ( .A(g_input[28]), .B(e_input[22]), .Z(n1115) );
  XNOR U2280 ( .A(n1119), .B(n1116), .Z(n1117) );
  XOR U2281 ( .A(n1066), .B(n1053), .Z(n1105) );
  XOR U2282 ( .A(n1123), .B(n1064), .Z(n1066) );
  XNOR U2283 ( .A(n1063), .B(n1062), .Z(n1064) );
  NAND U2284 ( .A(g_input[31]), .B(e_input[19]), .Z(n1062) );
  XNOR U2285 ( .A(n1127), .B(n1124), .Z(n1125) );
  XNOR U2286 ( .A(n1059), .B(n1065), .Z(n1123) );
  XNOR U2287 ( .A(n1131), .B(n1134), .Z(n1133) );
  XOR U2288 ( .A(n1135), .B(n1085), .Z(n1075) );
  XNOR U2289 ( .A(n1072), .B(n1073), .Z(n1085) );
  NAND U2290 ( .A(e_input[27]), .B(g_input[23]), .Z(n1073) );
  XNOR U2291 ( .A(n1070), .B(n1136), .Z(n1072) );
  AND U2292 ( .A(g_input[24]), .B(e_input[26]), .Z(n1136) );
  XNOR U2293 ( .A(n1140), .B(n1137), .Z(n1138) );
  XNOR U2294 ( .A(n1084), .B(n1074), .Z(n1135) );
  XOR U2295 ( .A(n1079), .B(n1145), .Z(n1080) );
  AND U2296 ( .A(g_input[26]), .B(e_input[24]), .Z(n1145) );
  XNOR U2297 ( .A(n1149), .B(n1081), .Z(n1144) );
  NAND U2298 ( .A(e_input[25]), .B(g_input[25]), .Z(n1081) );
  IV U2299 ( .A(n1083), .Z(n1149) );
  XOR U2300 ( .A(n1088), .B(n1154), .Z(n1089) );
  AND U2301 ( .A(g_input[22]), .B(e_input[28]), .Z(n1154) );
  XNOR U2302 ( .A(n1158), .B(n1090), .Z(n1153) );
  NAND U2303 ( .A(e_input[29]), .B(g_input[21]), .Z(n1090) );
  IV U2304 ( .A(n1092), .Z(n1158) );
  XNOR U2305 ( .A(n1098), .B(n1099), .Z(n1094) );
  NAND U2306 ( .A(e_input[31]), .B(g_input[19]), .Z(n1099) );
  XNOR U2307 ( .A(n1096), .B(n1162), .Z(n1098) );
  AND U2308 ( .A(g_input[20]), .B(e_input[30]), .Z(n1162) );
  XNOR U2309 ( .A(n1166), .B(n1163), .Z(n1164) );
  XNOR U2310 ( .A(n1102), .B(n1100), .Z(n1104) );
  XOR U2311 ( .A(o_reg[17]), .B(n1168), .Z(o[16]) );
  XOR U2312 ( .A(n1171), .B(n1170), .Z(n1168) );
  XOR U2313 ( .A(n1172), .B(n1130), .Z(n1121) );
  XOR U2314 ( .A(n1108), .B(n1174), .Z(n1109) );
  AND U2315 ( .A(g_input[29]), .B(e_input[20]), .Z(n1174) );
  XNOR U2316 ( .A(n1178), .B(n1110), .Z(n1173) );
  NAND U2317 ( .A(e_input[21]), .B(g_input[28]), .Z(n1110) );
  IV U2318 ( .A(n1112), .Z(n1178) );
  XNOR U2319 ( .A(n1118), .B(n1119), .Z(n1114) );
  NAND U2320 ( .A(e_input[23]), .B(g_input[26]), .Z(n1119) );
  XNOR U2321 ( .A(n1116), .B(n1182), .Z(n1118) );
  AND U2322 ( .A(g_input[27]), .B(e_input[22]), .Z(n1182) );
  XNOR U2323 ( .A(n1186), .B(n1183), .Z(n1184) );
  XNOR U2324 ( .A(n1129), .B(n1120), .Z(n1172) );
  XOR U2325 ( .A(n1190), .B(n1134), .Z(n1129) );
  XNOR U2326 ( .A(n1126), .B(n1127), .Z(n1134) );
  NAND U2327 ( .A(e_input[19]), .B(g_input[30]), .Z(n1127) );
  XNOR U2328 ( .A(n1124), .B(n1191), .Z(n1126) );
  AND U2329 ( .A(g_input[31]), .B(e_input[18]), .Z(n1191) );
  XNOR U2330 ( .A(n1195), .B(n1192), .Z(n1193) );
  XNOR U2331 ( .A(n1132), .B(n1128), .Z(n1190) );
  XOR U2332 ( .A(n1131), .B(n1199), .Z(n1132) );
  ANDN U2333 ( .A(n1200), .B(n1201), .Z(n1199) );
  XOR U2334 ( .A(n1205), .B(n1152), .Z(n1142) );
  XNOR U2335 ( .A(n1139), .B(n1140), .Z(n1152) );
  NAND U2336 ( .A(e_input[27]), .B(g_input[22]), .Z(n1140) );
  XNOR U2337 ( .A(n1137), .B(n1206), .Z(n1139) );
  AND U2338 ( .A(g_input[23]), .B(e_input[26]), .Z(n1206) );
  XNOR U2339 ( .A(n1210), .B(n1207), .Z(n1208) );
  XNOR U2340 ( .A(n1151), .B(n1141), .Z(n1205) );
  XOR U2341 ( .A(n1146), .B(n1215), .Z(n1147) );
  AND U2342 ( .A(g_input[25]), .B(e_input[24]), .Z(n1215) );
  XNOR U2343 ( .A(n1219), .B(n1148), .Z(n1214) );
  NAND U2344 ( .A(e_input[25]), .B(g_input[24]), .Z(n1148) );
  IV U2345 ( .A(n1150), .Z(n1219) );
  XOR U2346 ( .A(n1155), .B(n1224), .Z(n1156) );
  AND U2347 ( .A(g_input[21]), .B(e_input[28]), .Z(n1224) );
  XNOR U2348 ( .A(n1228), .B(n1157), .Z(n1223) );
  NAND U2349 ( .A(e_input[29]), .B(g_input[20]), .Z(n1157) );
  IV U2350 ( .A(n1159), .Z(n1228) );
  XNOR U2351 ( .A(n1165), .B(n1166), .Z(n1161) );
  NAND U2352 ( .A(e_input[31]), .B(g_input[18]), .Z(n1166) );
  XNOR U2353 ( .A(n1163), .B(n1232), .Z(n1165) );
  AND U2354 ( .A(g_input[19]), .B(e_input[30]), .Z(n1232) );
  XNOR U2355 ( .A(n1236), .B(n1233), .Z(n1234) );
  XNOR U2356 ( .A(n1169), .B(n1167), .Z(n1171) );
  XOR U2357 ( .A(o_reg[16]), .B(n1238), .Z(o[15]) );
  XOR U2358 ( .A(n1241), .B(n1240), .Z(n1238) );
  XOR U2359 ( .A(n1242), .B(n1198), .Z(n1188) );
  XOR U2360 ( .A(n1175), .B(n1244), .Z(n1176) );
  AND U2361 ( .A(g_input[28]), .B(e_input[20]), .Z(n1244) );
  XNOR U2362 ( .A(n1248), .B(n1177), .Z(n1243) );
  NAND U2363 ( .A(e_input[21]), .B(g_input[27]), .Z(n1177) );
  IV U2364 ( .A(n1179), .Z(n1248) );
  XNOR U2365 ( .A(n1185), .B(n1186), .Z(n1181) );
  NAND U2366 ( .A(e_input[23]), .B(g_input[25]), .Z(n1186) );
  XNOR U2367 ( .A(n1183), .B(n1252), .Z(n1185) );
  AND U2368 ( .A(g_input[26]), .B(e_input[22]), .Z(n1252) );
  XNOR U2369 ( .A(n1256), .B(n1253), .Z(n1254) );
  XNOR U2370 ( .A(n1197), .B(n1187), .Z(n1242) );
  XOR U2371 ( .A(n1260), .B(n1204), .Z(n1197) );
  XNOR U2372 ( .A(n1194), .B(n1195), .Z(n1204) );
  NAND U2373 ( .A(e_input[19]), .B(g_input[29]), .Z(n1195) );
  XNOR U2374 ( .A(n1192), .B(n1261), .Z(n1194) );
  AND U2375 ( .A(g_input[30]), .B(e_input[18]), .Z(n1261) );
  XNOR U2376 ( .A(n1265), .B(n1262), .Z(n1263) );
  XNOR U2377 ( .A(n1203), .B(n1196), .Z(n1260) );
  XNOR U2378 ( .A(n1273), .B(n1201), .Z(n1269) );
  NAND U2379 ( .A(e_input[17]), .B(g_input[31]), .Z(n1201) );
  IV U2380 ( .A(n1202), .Z(n1273) );
  XOR U2381 ( .A(n1277), .B(n1222), .Z(n1212) );
  XNOR U2382 ( .A(n1209), .B(n1210), .Z(n1222) );
  NAND U2383 ( .A(e_input[27]), .B(g_input[21]), .Z(n1210) );
  XNOR U2384 ( .A(n1207), .B(n1278), .Z(n1209) );
  AND U2385 ( .A(g_input[22]), .B(e_input[26]), .Z(n1278) );
  XNOR U2386 ( .A(n1282), .B(n1279), .Z(n1280) );
  XNOR U2387 ( .A(n1221), .B(n1211), .Z(n1277) );
  XOR U2388 ( .A(n1216), .B(n1287), .Z(n1217) );
  AND U2389 ( .A(g_input[24]), .B(e_input[24]), .Z(n1287) );
  XNOR U2390 ( .A(n1291), .B(n1218), .Z(n1286) );
  NAND U2391 ( .A(e_input[25]), .B(g_input[23]), .Z(n1218) );
  IV U2392 ( .A(n1220), .Z(n1291) );
  XOR U2393 ( .A(n1225), .B(n1296), .Z(n1226) );
  AND U2394 ( .A(g_input[20]), .B(e_input[28]), .Z(n1296) );
  XNOR U2395 ( .A(n1300), .B(n1227), .Z(n1295) );
  NAND U2396 ( .A(e_input[29]), .B(g_input[19]), .Z(n1227) );
  IV U2397 ( .A(n1229), .Z(n1300) );
  XNOR U2398 ( .A(n1235), .B(n1236), .Z(n1231) );
  NAND U2399 ( .A(e_input[31]), .B(g_input[17]), .Z(n1236) );
  XNOR U2400 ( .A(n1233), .B(n1304), .Z(n1235) );
  AND U2401 ( .A(g_input[18]), .B(e_input[30]), .Z(n1304) );
  XNOR U2402 ( .A(n1308), .B(n1305), .Z(n1306) );
  XNOR U2403 ( .A(n1239), .B(n1237), .Z(n1241) );
  XNOR U2404 ( .A(n1310), .B(o_reg[15]), .Z(o[14]) );
  XOR U2405 ( .A(n1314), .B(n1313), .Z(n1310) );
  XOR U2406 ( .A(n1315), .B(n1268), .Z(n1258) );
  XOR U2407 ( .A(n1245), .B(n1317), .Z(n1246) );
  AND U2408 ( .A(g_input[27]), .B(e_input[20]), .Z(n1317) );
  XNOR U2409 ( .A(n1321), .B(n1247), .Z(n1316) );
  NAND U2410 ( .A(e_input[21]), .B(g_input[26]), .Z(n1247) );
  IV U2411 ( .A(n1249), .Z(n1321) );
  XNOR U2412 ( .A(n1255), .B(n1256), .Z(n1251) );
  NAND U2413 ( .A(e_input[23]), .B(g_input[24]), .Z(n1256) );
  XNOR U2414 ( .A(n1253), .B(n1325), .Z(n1255) );
  AND U2415 ( .A(g_input[25]), .B(e_input[22]), .Z(n1325) );
  XNOR U2416 ( .A(n1329), .B(n1326), .Z(n1327) );
  XNOR U2417 ( .A(n1267), .B(n1257), .Z(n1315) );
  XOR U2418 ( .A(n1333), .B(n1276), .Z(n1267) );
  XNOR U2419 ( .A(n1264), .B(n1265), .Z(n1276) );
  NAND U2420 ( .A(e_input[19]), .B(g_input[28]), .Z(n1265) );
  XNOR U2421 ( .A(n1262), .B(n1334), .Z(n1264) );
  AND U2422 ( .A(g_input[29]), .B(e_input[18]), .Z(n1334) );
  XNOR U2423 ( .A(n1338), .B(n1335), .Z(n1336) );
  XNOR U2424 ( .A(n1275), .B(n1266), .Z(n1333) );
  XOR U2425 ( .A(n1270), .B(n1343), .Z(n1271) );
  AND U2426 ( .A(g_input[31]), .B(e_input[16]), .Z(n1343) );
  XNOR U2427 ( .A(n1347), .B(n1272), .Z(n1342) );
  NAND U2428 ( .A(e_input[17]), .B(g_input[30]), .Z(n1272) );
  IV U2429 ( .A(n1274), .Z(n1347) );
  XOR U2430 ( .A(n1351), .B(n1294), .Z(n1284) );
  XNOR U2431 ( .A(n1281), .B(n1282), .Z(n1294) );
  NAND U2432 ( .A(e_input[27]), .B(g_input[20]), .Z(n1282) );
  XNOR U2433 ( .A(n1279), .B(n1352), .Z(n1281) );
  AND U2434 ( .A(g_input[21]), .B(e_input[26]), .Z(n1352) );
  XNOR U2435 ( .A(n1356), .B(n1353), .Z(n1354) );
  XNOR U2436 ( .A(n1293), .B(n1283), .Z(n1351) );
  XOR U2437 ( .A(n1288), .B(n1361), .Z(n1289) );
  AND U2438 ( .A(g_input[23]), .B(e_input[24]), .Z(n1361) );
  XNOR U2439 ( .A(n1365), .B(n1290), .Z(n1360) );
  NAND U2440 ( .A(e_input[25]), .B(g_input[22]), .Z(n1290) );
  IV U2441 ( .A(n1292), .Z(n1365) );
  XOR U2442 ( .A(n1297), .B(n1370), .Z(n1298) );
  AND U2443 ( .A(g_input[19]), .B(e_input[28]), .Z(n1370) );
  XNOR U2444 ( .A(n1374), .B(n1299), .Z(n1369) );
  NAND U2445 ( .A(e_input[29]), .B(g_input[18]), .Z(n1299) );
  IV U2446 ( .A(n1301), .Z(n1374) );
  XNOR U2447 ( .A(n1307), .B(n1308), .Z(n1303) );
  NAND U2448 ( .A(e_input[31]), .B(g_input[16]), .Z(n1308) );
  XNOR U2449 ( .A(n1305), .B(n1378), .Z(n1307) );
  AND U2450 ( .A(g_input[17]), .B(e_input[30]), .Z(n1378) );
  XNOR U2451 ( .A(n1382), .B(n1379), .Z(n1380) );
  XNOR U2452 ( .A(n1312), .B(n1309), .Z(n1314) );
  XNOR U2453 ( .A(n1385), .B(n1386), .Z(n1312) );
  XOR U2454 ( .A(n1387), .B(n1388), .Z(n1386) );
  XNOR U2455 ( .A(n1389), .B(n1390), .Z(n1388) );
  AND U2456 ( .A(n1391), .B(n1392), .Z(n1389) );
  NAND U2457 ( .A(n1393), .B(n1394), .Z(n1392) );
  NANDN U2458 ( .B(n1395), .A(n1396), .Z(n1391) );
  XOR U2459 ( .A(n1397), .B(n1398), .Z(n1387) );
  ANDN U2460 ( .A(n1401), .B(n1390), .Z(n1397) );
  XOR U2461 ( .A(n1402), .B(n1403), .Z(n1385) );
  XOR U2462 ( .A(n1399), .B(n1396), .Z(n1403) );
  XOR U2463 ( .A(o_reg[14]), .B(n1384), .Z(o[13]) );
  XOR U2464 ( .A(n1407), .B(n1406), .Z(n1384) );
  XOR U2465 ( .A(n1408), .B(n1341), .Z(n1331) );
  XOR U2466 ( .A(n1318), .B(n1410), .Z(n1319) );
  AND U2467 ( .A(g_input[26]), .B(e_input[20]), .Z(n1410) );
  XNOR U2468 ( .A(n1414), .B(n1320), .Z(n1409) );
  NAND U2469 ( .A(e_input[21]), .B(g_input[25]), .Z(n1320) );
  IV U2470 ( .A(n1322), .Z(n1414) );
  XNOR U2471 ( .A(n1328), .B(n1329), .Z(n1324) );
  NAND U2472 ( .A(e_input[23]), .B(g_input[23]), .Z(n1329) );
  XNOR U2473 ( .A(n1326), .B(n1418), .Z(n1328) );
  AND U2474 ( .A(g_input[24]), .B(e_input[22]), .Z(n1418) );
  XNOR U2475 ( .A(n1422), .B(n1419), .Z(n1420) );
  XNOR U2476 ( .A(n1340), .B(n1330), .Z(n1408) );
  XOR U2477 ( .A(n1426), .B(n1350), .Z(n1340) );
  XNOR U2478 ( .A(n1337), .B(n1338), .Z(n1350) );
  NAND U2479 ( .A(e_input[19]), .B(g_input[27]), .Z(n1338) );
  XNOR U2480 ( .A(n1335), .B(n1427), .Z(n1337) );
  AND U2481 ( .A(g_input[28]), .B(e_input[18]), .Z(n1427) );
  XNOR U2482 ( .A(n1431), .B(n1428), .Z(n1429) );
  XNOR U2483 ( .A(n1349), .B(n1339), .Z(n1426) );
  XOR U2484 ( .A(n1344), .B(n1436), .Z(n1345) );
  AND U2485 ( .A(g_input[30]), .B(e_input[16]), .Z(n1436) );
  XNOR U2486 ( .A(n1440), .B(n1346), .Z(n1435) );
  NAND U2487 ( .A(e_input[17]), .B(g_input[29]), .Z(n1346) );
  IV U2488 ( .A(n1348), .Z(n1440) );
  XOR U2489 ( .A(n1444), .B(n1368), .Z(n1358) );
  XNOR U2490 ( .A(n1355), .B(n1356), .Z(n1368) );
  NAND U2491 ( .A(e_input[27]), .B(g_input[19]), .Z(n1356) );
  XNOR U2492 ( .A(n1353), .B(n1445), .Z(n1355) );
  AND U2493 ( .A(g_input[20]), .B(e_input[26]), .Z(n1445) );
  XNOR U2494 ( .A(n1449), .B(n1446), .Z(n1447) );
  XNOR U2495 ( .A(n1367), .B(n1357), .Z(n1444) );
  XOR U2496 ( .A(n1362), .B(n1454), .Z(n1363) );
  AND U2497 ( .A(g_input[22]), .B(e_input[24]), .Z(n1454) );
  XNOR U2498 ( .A(n1458), .B(n1364), .Z(n1453) );
  NAND U2499 ( .A(e_input[25]), .B(g_input[21]), .Z(n1364) );
  IV U2500 ( .A(n1366), .Z(n1458) );
  XOR U2501 ( .A(n1371), .B(n1463), .Z(n1372) );
  AND U2502 ( .A(g_input[18]), .B(e_input[28]), .Z(n1463) );
  XNOR U2503 ( .A(n1467), .B(n1373), .Z(n1462) );
  NAND U2504 ( .A(e_input[29]), .B(g_input[17]), .Z(n1373) );
  IV U2505 ( .A(n1375), .Z(n1467) );
  XNOR U2506 ( .A(n1381), .B(n1382), .Z(n1377) );
  NAND U2507 ( .A(e_input[31]), .B(g_input[15]), .Z(n1382) );
  XNOR U2508 ( .A(n1379), .B(n1471), .Z(n1381) );
  AND U2509 ( .A(g_input[16]), .B(e_input[30]), .Z(n1471) );
  XNOR U2510 ( .A(n1475), .B(n1472), .Z(n1473) );
  XNOR U2511 ( .A(n1405), .B(n1383), .Z(n1407) );
  XOR U2512 ( .A(n1478), .B(n1400), .Z(n1405) );
  XNOR U2513 ( .A(n1401), .B(n1390), .Z(n1400) );
  OR U2514 ( .A(n1479), .B(n1480), .Z(n1390) );
  XNOR U2515 ( .A(n1394), .B(n1393), .Z(n1395) );
  NAND U2516 ( .A(e_input[15]), .B(g_input[31]), .Z(n1393) );
  XNOR U2517 ( .A(n1487), .B(n1484), .Z(n1485) );
  XNOR U2518 ( .A(n1399), .B(n1404), .Z(n1478) );
  XOR U2519 ( .A(o_reg[13]), .B(n1477), .Z(o[12]) );
  XOR U2520 ( .A(n1493), .B(n1490), .Z(n1477) );
  XOR U2521 ( .A(n1494), .B(n1434), .Z(n1424) );
  XOR U2522 ( .A(n1411), .B(n1496), .Z(n1412) );
  AND U2523 ( .A(g_input[25]), .B(e_input[20]), .Z(n1496) );
  XNOR U2524 ( .A(n1500), .B(n1413), .Z(n1495) );
  NAND U2525 ( .A(e_input[21]), .B(g_input[24]), .Z(n1413) );
  IV U2526 ( .A(n1415), .Z(n1500) );
  XNOR U2527 ( .A(n1421), .B(n1422), .Z(n1417) );
  NAND U2528 ( .A(e_input[23]), .B(g_input[22]), .Z(n1422) );
  XNOR U2529 ( .A(n1419), .B(n1504), .Z(n1421) );
  AND U2530 ( .A(g_input[23]), .B(e_input[22]), .Z(n1504) );
  XNOR U2531 ( .A(n1508), .B(n1505), .Z(n1506) );
  XNOR U2532 ( .A(n1433), .B(n1423), .Z(n1494) );
  XOR U2533 ( .A(n1512), .B(n1443), .Z(n1433) );
  XNOR U2534 ( .A(n1430), .B(n1431), .Z(n1443) );
  NAND U2535 ( .A(e_input[19]), .B(g_input[26]), .Z(n1431) );
  XNOR U2536 ( .A(n1428), .B(n1513), .Z(n1430) );
  AND U2537 ( .A(g_input[27]), .B(e_input[18]), .Z(n1513) );
  XNOR U2538 ( .A(n1517), .B(n1514), .Z(n1515) );
  XNOR U2539 ( .A(n1442), .B(n1432), .Z(n1512) );
  XOR U2540 ( .A(n1437), .B(n1522), .Z(n1438) );
  AND U2541 ( .A(g_input[29]), .B(e_input[16]), .Z(n1522) );
  XNOR U2542 ( .A(n1526), .B(n1439), .Z(n1521) );
  NAND U2543 ( .A(e_input[17]), .B(g_input[28]), .Z(n1439) );
  IV U2544 ( .A(n1441), .Z(n1526) );
  XOR U2545 ( .A(n1530), .B(n1461), .Z(n1451) );
  XNOR U2546 ( .A(n1448), .B(n1449), .Z(n1461) );
  NAND U2547 ( .A(e_input[27]), .B(g_input[18]), .Z(n1449) );
  XNOR U2548 ( .A(n1446), .B(n1531), .Z(n1448) );
  AND U2549 ( .A(g_input[19]), .B(e_input[26]), .Z(n1531) );
  XNOR U2550 ( .A(n1535), .B(n1532), .Z(n1533) );
  XNOR U2551 ( .A(n1460), .B(n1450), .Z(n1530) );
  XOR U2552 ( .A(n1455), .B(n1540), .Z(n1456) );
  AND U2553 ( .A(g_input[21]), .B(e_input[24]), .Z(n1540) );
  XNOR U2554 ( .A(n1544), .B(n1457), .Z(n1539) );
  NAND U2555 ( .A(e_input[25]), .B(g_input[20]), .Z(n1457) );
  IV U2556 ( .A(n1459), .Z(n1544) );
  XOR U2557 ( .A(n1464), .B(n1549), .Z(n1465) );
  AND U2558 ( .A(g_input[17]), .B(e_input[28]), .Z(n1549) );
  XNOR U2559 ( .A(n1553), .B(n1466), .Z(n1548) );
  NAND U2560 ( .A(e_input[29]), .B(g_input[16]), .Z(n1466) );
  IV U2561 ( .A(n1468), .Z(n1553) );
  XNOR U2562 ( .A(n1474), .B(n1475), .Z(n1470) );
  NAND U2563 ( .A(e_input[31]), .B(g_input[14]), .Z(n1475) );
  XNOR U2564 ( .A(n1472), .B(n1557), .Z(n1474) );
  AND U2565 ( .A(g_input[15]), .B(e_input[30]), .Z(n1557) );
  XNOR U2566 ( .A(n1561), .B(n1558), .Z(n1559) );
  XNOR U2567 ( .A(n1489), .B(n1476), .Z(n1493) );
  XOR U2568 ( .A(n1564), .B(n1492), .Z(n1489) );
  XNOR U2569 ( .A(n1479), .B(n1480), .Z(n1492) );
  NANDN U2570 ( .B(n1565), .A(n1566), .Z(n1480) );
  XOR U2571 ( .A(n1481), .B(n1567), .Z(n1482) );
  ANDN U2572 ( .A(n1568), .B(n1569), .Z(n1567) );
  XNOR U2573 ( .A(n1486), .B(n1487), .Z(n1483) );
  NAND U2574 ( .A(g_input[30]), .B(e_input[15]), .Z(n1487) );
  XNOR U2575 ( .A(n1484), .B(n1573), .Z(n1486) );
  AND U2576 ( .A(e_input[14]), .B(g_input[31]), .Z(n1573) );
  XNOR U2577 ( .A(n1577), .B(n1574), .Z(n1575) );
  XOR U2578 ( .A(o_reg[12]), .B(n1563), .Z(o[11]) );
  XOR U2579 ( .A(n1583), .B(n1580), .Z(n1563) );
  XOR U2580 ( .A(n1584), .B(n1520), .Z(n1510) );
  XOR U2581 ( .A(n1497), .B(n1586), .Z(n1498) );
  AND U2582 ( .A(g_input[24]), .B(e_input[20]), .Z(n1586) );
  XNOR U2583 ( .A(n1590), .B(n1499), .Z(n1585) );
  NAND U2584 ( .A(e_input[21]), .B(g_input[23]), .Z(n1499) );
  IV U2585 ( .A(n1501), .Z(n1590) );
  XNOR U2586 ( .A(n1507), .B(n1508), .Z(n1503) );
  NAND U2587 ( .A(e_input[23]), .B(g_input[21]), .Z(n1508) );
  XNOR U2588 ( .A(n1505), .B(n1594), .Z(n1507) );
  AND U2589 ( .A(g_input[22]), .B(e_input[22]), .Z(n1594) );
  XNOR U2590 ( .A(n1598), .B(n1595), .Z(n1596) );
  XNOR U2591 ( .A(n1519), .B(n1509), .Z(n1584) );
  XOR U2592 ( .A(n1602), .B(n1529), .Z(n1519) );
  XNOR U2593 ( .A(n1516), .B(n1517), .Z(n1529) );
  NAND U2594 ( .A(e_input[19]), .B(g_input[25]), .Z(n1517) );
  XNOR U2595 ( .A(n1514), .B(n1603), .Z(n1516) );
  AND U2596 ( .A(g_input[26]), .B(e_input[18]), .Z(n1603) );
  XNOR U2597 ( .A(n1607), .B(n1604), .Z(n1605) );
  XNOR U2598 ( .A(n1528), .B(n1518), .Z(n1602) );
  XOR U2599 ( .A(n1523), .B(n1612), .Z(n1524) );
  AND U2600 ( .A(g_input[28]), .B(e_input[16]), .Z(n1612) );
  XNOR U2601 ( .A(n1616), .B(n1525), .Z(n1611) );
  NAND U2602 ( .A(e_input[17]), .B(g_input[27]), .Z(n1525) );
  IV U2603 ( .A(n1527), .Z(n1616) );
  XOR U2604 ( .A(n1620), .B(n1547), .Z(n1537) );
  XNOR U2605 ( .A(n1534), .B(n1535), .Z(n1547) );
  NAND U2606 ( .A(e_input[27]), .B(g_input[17]), .Z(n1535) );
  XNOR U2607 ( .A(n1532), .B(n1621), .Z(n1534) );
  AND U2608 ( .A(g_input[18]), .B(e_input[26]), .Z(n1621) );
  XNOR U2609 ( .A(n1625), .B(n1622), .Z(n1623) );
  XNOR U2610 ( .A(n1546), .B(n1536), .Z(n1620) );
  XOR U2611 ( .A(n1541), .B(n1630), .Z(n1542) );
  AND U2612 ( .A(g_input[20]), .B(e_input[24]), .Z(n1630) );
  XNOR U2613 ( .A(n1634), .B(n1543), .Z(n1629) );
  NAND U2614 ( .A(e_input[25]), .B(g_input[19]), .Z(n1543) );
  IV U2615 ( .A(n1545), .Z(n1634) );
  XOR U2616 ( .A(n1550), .B(n1639), .Z(n1551) );
  AND U2617 ( .A(g_input[16]), .B(e_input[28]), .Z(n1639) );
  XNOR U2618 ( .A(n1643), .B(n1552), .Z(n1638) );
  NAND U2619 ( .A(e_input[29]), .B(g_input[15]), .Z(n1552) );
  IV U2620 ( .A(n1554), .Z(n1643) );
  XNOR U2621 ( .A(n1560), .B(n1561), .Z(n1556) );
  NAND U2622 ( .A(e_input[31]), .B(g_input[13]), .Z(n1561) );
  XNOR U2623 ( .A(n1558), .B(n1647), .Z(n1560) );
  AND U2624 ( .A(g_input[14]), .B(e_input[30]), .Z(n1647) );
  XNOR U2625 ( .A(n1651), .B(n1648), .Z(n1649) );
  XNOR U2626 ( .A(n1579), .B(n1562), .Z(n1583) );
  XOR U2627 ( .A(n1654), .B(n1582), .Z(n1579) );
  XNOR U2628 ( .A(n1662), .B(n1569), .Z(n1658) );
  NAND U2629 ( .A(g_input[31]), .B(e_input[13]), .Z(n1569) );
  IV U2630 ( .A(n1570), .Z(n1662) );
  XNOR U2631 ( .A(n1576), .B(n1577), .Z(n1572) );
  NAND U2632 ( .A(g_input[29]), .B(e_input[15]), .Z(n1577) );
  XNOR U2633 ( .A(n1574), .B(n1666), .Z(n1576) );
  AND U2634 ( .A(e_input[14]), .B(g_input[30]), .Z(n1666) );
  XNOR U2635 ( .A(n1670), .B(n1667), .Z(n1668) );
  XNOR U2636 ( .A(n1653), .B(o_reg[11]), .Z(o[10]) );
  XOR U2637 ( .A(n1676), .B(n1673), .Z(n1653) );
  XOR U2638 ( .A(n1677), .B(n1610), .Z(n1600) );
  XOR U2639 ( .A(n1587), .B(n1679), .Z(n1588) );
  AND U2640 ( .A(g_input[23]), .B(e_input[20]), .Z(n1679) );
  XNOR U2641 ( .A(n1683), .B(n1589), .Z(n1678) );
  NAND U2642 ( .A(e_input[21]), .B(g_input[22]), .Z(n1589) );
  IV U2643 ( .A(n1591), .Z(n1683) );
  XNOR U2644 ( .A(n1597), .B(n1598), .Z(n1593) );
  NAND U2645 ( .A(e_input[23]), .B(g_input[20]), .Z(n1598) );
  XNOR U2646 ( .A(n1595), .B(n1687), .Z(n1597) );
  AND U2647 ( .A(g_input[21]), .B(e_input[22]), .Z(n1687) );
  XNOR U2648 ( .A(n1691), .B(n1688), .Z(n1689) );
  XNOR U2649 ( .A(n1609), .B(n1599), .Z(n1677) );
  XOR U2650 ( .A(n1695), .B(n1619), .Z(n1609) );
  XNOR U2651 ( .A(n1606), .B(n1607), .Z(n1619) );
  NAND U2652 ( .A(e_input[19]), .B(g_input[24]), .Z(n1607) );
  XNOR U2653 ( .A(n1604), .B(n1696), .Z(n1606) );
  AND U2654 ( .A(g_input[25]), .B(e_input[18]), .Z(n1696) );
  XNOR U2655 ( .A(n1700), .B(n1697), .Z(n1698) );
  XNOR U2656 ( .A(n1618), .B(n1608), .Z(n1695) );
  XOR U2657 ( .A(n1613), .B(n1705), .Z(n1614) );
  AND U2658 ( .A(g_input[27]), .B(e_input[16]), .Z(n1705) );
  XNOR U2659 ( .A(n1709), .B(n1615), .Z(n1704) );
  NAND U2660 ( .A(e_input[17]), .B(g_input[26]), .Z(n1615) );
  IV U2661 ( .A(n1617), .Z(n1709) );
  XOR U2662 ( .A(n1713), .B(n1637), .Z(n1627) );
  XNOR U2663 ( .A(n1624), .B(n1625), .Z(n1637) );
  NAND U2664 ( .A(e_input[27]), .B(g_input[16]), .Z(n1625) );
  XNOR U2665 ( .A(n1622), .B(n1714), .Z(n1624) );
  AND U2666 ( .A(g_input[17]), .B(e_input[26]), .Z(n1714) );
  XNOR U2667 ( .A(n1718), .B(n1715), .Z(n1716) );
  XNOR U2668 ( .A(n1636), .B(n1626), .Z(n1713) );
  XOR U2669 ( .A(n1631), .B(n1723), .Z(n1632) );
  AND U2670 ( .A(g_input[19]), .B(e_input[24]), .Z(n1723) );
  XNOR U2671 ( .A(n1727), .B(n1633), .Z(n1722) );
  NAND U2672 ( .A(e_input[25]), .B(g_input[18]), .Z(n1633) );
  IV U2673 ( .A(n1635), .Z(n1727) );
  XOR U2674 ( .A(n1640), .B(n1732), .Z(n1641) );
  AND U2675 ( .A(g_input[15]), .B(e_input[28]), .Z(n1732) );
  XNOR U2676 ( .A(n1736), .B(n1642), .Z(n1731) );
  NAND U2677 ( .A(e_input[29]), .B(g_input[14]), .Z(n1642) );
  IV U2678 ( .A(n1644), .Z(n1736) );
  XNOR U2679 ( .A(n1650), .B(n1651), .Z(n1646) );
  NAND U2680 ( .A(e_input[31]), .B(g_input[12]), .Z(n1651) );
  XNOR U2681 ( .A(n1648), .B(n1740), .Z(n1650) );
  AND U2682 ( .A(g_input[13]), .B(e_input[30]), .Z(n1740) );
  XNOR U2683 ( .A(n1744), .B(n1741), .Z(n1742) );
  XNOR U2684 ( .A(n1672), .B(n1652), .Z(n1676) );
  XOR U2685 ( .A(n1746), .B(n1747), .Z(n579) );
  XNOR U2686 ( .A(n1748), .B(n1745), .Z(n1746) );
  XNOR U2687 ( .A(n1750), .B(n1751), .Z(n580) );
  XOR U2688 ( .A(n1752), .B(n1749), .Z(n1750) );
  XNOR U2689 ( .A(n1754), .B(n1755), .Z(n581) );
  XOR U2690 ( .A(n1756), .B(n1753), .Z(n1754) );
  XNOR U2691 ( .A(n1758), .B(n1759), .Z(n582) );
  XOR U2692 ( .A(n1760), .B(n1757), .Z(n1758) );
  XNOR U2693 ( .A(n1762), .B(n1763), .Z(n583) );
  XOR U2694 ( .A(n1764), .B(n1761), .Z(n1762) );
  XNOR U2695 ( .A(n1766), .B(n1767), .Z(n584) );
  XOR U2696 ( .A(n1768), .B(n1765), .Z(n1766) );
  XNOR U2697 ( .A(n1770), .B(n1771), .Z(n585) );
  XOR U2698 ( .A(n1772), .B(n1769), .Z(n1770) );
  XNOR U2699 ( .A(n1774), .B(n1775), .Z(n615) );
  XOR U2700 ( .A(n1776), .B(n1773), .Z(n1774) );
  XNOR U2701 ( .A(n1778), .B(n1779), .Z(n979) );
  XNOR U2702 ( .A(n1780), .B(n1777), .Z(n1778) );
  XOR U2703 ( .A(n1783), .B(n1675), .Z(n1672) );
  XNOR U2704 ( .A(n1657), .B(n1656), .Z(n1675) );
  XOR U2705 ( .A(n1784), .B(n1785), .Z(n1656) );
  XOR U2706 ( .A(n1786), .B(n1787), .Z(n1785) );
  AND U2707 ( .A(n1788), .B(n1789), .Z(n1786) );
  NAND U2708 ( .A(n1790), .B(n1791), .Z(n1789) );
  NANDN U2709 ( .B(n1792), .A(n1787), .Z(n1788) );
  XOR U2710 ( .A(n1793), .B(n1794), .Z(n1655) );
  AND U2711 ( .A(n1795), .B(n1796), .Z(n1794) );
  XNOR U2712 ( .A(n1793), .B(n1797), .Z(n1795) );
  XOR U2713 ( .A(n1659), .B(n1799), .Z(n1660) );
  AND U2714 ( .A(e_input[12]), .B(g_input[31]), .Z(n1799) );
  XNOR U2715 ( .A(n1803), .B(n1661), .Z(n1798) );
  NAND U2716 ( .A(g_input[30]), .B(e_input[13]), .Z(n1661) );
  IV U2717 ( .A(n1663), .Z(n1803) );
  XNOR U2718 ( .A(n1669), .B(n1670), .Z(n1665) );
  NAND U2719 ( .A(g_input[28]), .B(e_input[15]), .Z(n1670) );
  XNOR U2720 ( .A(n1667), .B(n1807), .Z(n1669) );
  AND U2721 ( .A(e_input[14]), .B(g_input[29]), .Z(n1807) );
  XNOR U2722 ( .A(n1811), .B(n1808), .Z(n1809) );
  XOR U2723 ( .A(n1813), .B(n1703), .Z(n1693) );
  XOR U2724 ( .A(n1680), .B(n1815), .Z(n1681) );
  AND U2725 ( .A(g_input[22]), .B(e_input[20]), .Z(n1815) );
  XNOR U2726 ( .A(n1819), .B(n1682), .Z(n1814) );
  NAND U2727 ( .A(e_input[21]), .B(g_input[21]), .Z(n1682) );
  IV U2728 ( .A(n1684), .Z(n1819) );
  XNOR U2729 ( .A(n1690), .B(n1691), .Z(n1686) );
  NAND U2730 ( .A(e_input[23]), .B(g_input[19]), .Z(n1691) );
  XNOR U2731 ( .A(n1688), .B(n1823), .Z(n1690) );
  AND U2732 ( .A(g_input[20]), .B(e_input[22]), .Z(n1823) );
  XNOR U2733 ( .A(n1827), .B(n1824), .Z(n1825) );
  XNOR U2734 ( .A(n1702), .B(n1692), .Z(n1813) );
  XOR U2735 ( .A(n1831), .B(n1712), .Z(n1702) );
  XNOR U2736 ( .A(n1699), .B(n1700), .Z(n1712) );
  NAND U2737 ( .A(e_input[19]), .B(g_input[23]), .Z(n1700) );
  XNOR U2738 ( .A(n1697), .B(n1832), .Z(n1699) );
  AND U2739 ( .A(g_input[24]), .B(e_input[18]), .Z(n1832) );
  XNOR U2740 ( .A(n1836), .B(n1833), .Z(n1834) );
  XNOR U2741 ( .A(n1711), .B(n1701), .Z(n1831) );
  XOR U2742 ( .A(n1706), .B(n1841), .Z(n1707) );
  AND U2743 ( .A(g_input[26]), .B(e_input[16]), .Z(n1841) );
  XNOR U2744 ( .A(n1845), .B(n1708), .Z(n1840) );
  NAND U2745 ( .A(e_input[17]), .B(g_input[25]), .Z(n1708) );
  IV U2746 ( .A(n1710), .Z(n1845) );
  XOR U2747 ( .A(n1849), .B(n1730), .Z(n1720) );
  XNOR U2748 ( .A(n1717), .B(n1718), .Z(n1730) );
  NAND U2749 ( .A(e_input[27]), .B(g_input[15]), .Z(n1718) );
  XNOR U2750 ( .A(n1715), .B(n1850), .Z(n1717) );
  AND U2751 ( .A(g_input[16]), .B(e_input[26]), .Z(n1850) );
  XNOR U2752 ( .A(n1854), .B(n1851), .Z(n1852) );
  XNOR U2753 ( .A(n1729), .B(n1719), .Z(n1849) );
  XOR U2754 ( .A(n1724), .B(n1859), .Z(n1725) );
  AND U2755 ( .A(g_input[18]), .B(e_input[24]), .Z(n1859) );
  XNOR U2756 ( .A(n1863), .B(n1726), .Z(n1858) );
  NAND U2757 ( .A(e_input[25]), .B(g_input[17]), .Z(n1726) );
  IV U2758 ( .A(n1728), .Z(n1863) );
  XOR U2759 ( .A(n1733), .B(n1868), .Z(n1734) );
  AND U2760 ( .A(g_input[14]), .B(e_input[28]), .Z(n1868) );
  XNOR U2761 ( .A(n1872), .B(n1735), .Z(n1867) );
  NAND U2762 ( .A(e_input[29]), .B(g_input[13]), .Z(n1735) );
  IV U2763 ( .A(n1737), .Z(n1872) );
  XNOR U2764 ( .A(n1743), .B(n1744), .Z(n1739) );
  NAND U2765 ( .A(e_input[31]), .B(g_input[11]), .Z(n1744) );
  XNOR U2766 ( .A(n1741), .B(n1876), .Z(n1743) );
  AND U2767 ( .A(g_input[12]), .B(e_input[30]), .Z(n1876) );
  XNOR U2768 ( .A(n1880), .B(n1877), .Z(n1878) );
  XOR U2769 ( .A(n1881), .B(n1882), .Z(n1748) );
  XNOR U2770 ( .A(n1885), .B(n1886), .Z(n1752) );
  XNOR U2771 ( .A(n1887), .B(n1884), .Z(n1885) );
  XOR U2772 ( .A(n1888), .B(n1839), .Z(n1829) );
  XOR U2773 ( .A(n1816), .B(n1890), .Z(n1817) );
  AND U2774 ( .A(g_input[21]), .B(e_input[20]), .Z(n1890) );
  XNOR U2775 ( .A(n1894), .B(n1818), .Z(n1889) );
  NAND U2776 ( .A(e_input[21]), .B(g_input[20]), .Z(n1818) );
  IV U2777 ( .A(n1820), .Z(n1894) );
  XNOR U2778 ( .A(n1826), .B(n1827), .Z(n1822) );
  NAND U2779 ( .A(e_input[23]), .B(g_input[18]), .Z(n1827) );
  XNOR U2780 ( .A(n1824), .B(n1898), .Z(n1826) );
  AND U2781 ( .A(g_input[19]), .B(e_input[22]), .Z(n1898) );
  XNOR U2782 ( .A(n1902), .B(n1899), .Z(n1900) );
  XNOR U2783 ( .A(n1838), .B(n1828), .Z(n1888) );
  XOR U2784 ( .A(n1906), .B(n1848), .Z(n1838) );
  XNOR U2785 ( .A(n1835), .B(n1836), .Z(n1848) );
  NAND U2786 ( .A(e_input[19]), .B(g_input[22]), .Z(n1836) );
  XNOR U2787 ( .A(n1833), .B(n1907), .Z(n1835) );
  AND U2788 ( .A(g_input[23]), .B(e_input[18]), .Z(n1907) );
  XNOR U2789 ( .A(n1911), .B(n1908), .Z(n1909) );
  XNOR U2790 ( .A(n1847), .B(n1837), .Z(n1906) );
  XOR U2791 ( .A(n1842), .B(n1916), .Z(n1843) );
  AND U2792 ( .A(g_input[25]), .B(e_input[16]), .Z(n1916) );
  XNOR U2793 ( .A(n1920), .B(n1844), .Z(n1915) );
  NAND U2794 ( .A(e_input[17]), .B(g_input[24]), .Z(n1844) );
  IV U2795 ( .A(n1846), .Z(n1920) );
  XOR U2796 ( .A(n1924), .B(n1866), .Z(n1856) );
  XNOR U2797 ( .A(n1853), .B(n1854), .Z(n1866) );
  NAND U2798 ( .A(e_input[27]), .B(g_input[14]), .Z(n1854) );
  XNOR U2799 ( .A(n1851), .B(n1925), .Z(n1853) );
  AND U2800 ( .A(g_input[15]), .B(e_input[26]), .Z(n1925) );
  XNOR U2801 ( .A(n1929), .B(n1926), .Z(n1927) );
  XNOR U2802 ( .A(n1865), .B(n1855), .Z(n1924) );
  XOR U2803 ( .A(n1860), .B(n1934), .Z(n1861) );
  AND U2804 ( .A(g_input[17]), .B(e_input[24]), .Z(n1934) );
  XNOR U2805 ( .A(n1938), .B(n1862), .Z(n1933) );
  NAND U2806 ( .A(e_input[25]), .B(g_input[16]), .Z(n1862) );
  IV U2807 ( .A(n1864), .Z(n1938) );
  XOR U2808 ( .A(n1869), .B(n1943), .Z(n1870) );
  AND U2809 ( .A(g_input[13]), .B(e_input[28]), .Z(n1943) );
  XNOR U2810 ( .A(n1947), .B(n1871), .Z(n1942) );
  NAND U2811 ( .A(e_input[29]), .B(g_input[12]), .Z(n1871) );
  IV U2812 ( .A(n1873), .Z(n1947) );
  XNOR U2813 ( .A(n1879), .B(n1880), .Z(n1875) );
  NAND U2814 ( .A(e_input[31]), .B(g_input[10]), .Z(n1880) );
  XNOR U2815 ( .A(n1877), .B(n1951), .Z(n1879) );
  AND U2816 ( .A(g_input[11]), .B(e_input[30]), .Z(n1951) );
  XNOR U2817 ( .A(n1955), .B(n1952), .Z(n1953) );
  XNOR U2818 ( .A(n1957), .B(n1958), .Z(n1756) );
  XNOR U2819 ( .A(n1959), .B(n1956), .Z(n1957) );
  XOR U2820 ( .A(n1960), .B(n1914), .Z(n1904) );
  XOR U2821 ( .A(n1891), .B(n1962), .Z(n1892) );
  AND U2822 ( .A(g_input[20]), .B(e_input[20]), .Z(n1962) );
  XNOR U2823 ( .A(n1966), .B(n1893), .Z(n1961) );
  NAND U2824 ( .A(e_input[21]), .B(g_input[19]), .Z(n1893) );
  IV U2825 ( .A(n1895), .Z(n1966) );
  XNOR U2826 ( .A(n1901), .B(n1902), .Z(n1897) );
  NAND U2827 ( .A(e_input[23]), .B(g_input[17]), .Z(n1902) );
  XNOR U2828 ( .A(n1899), .B(n1970), .Z(n1901) );
  AND U2829 ( .A(g_input[18]), .B(e_input[22]), .Z(n1970) );
  XNOR U2830 ( .A(n1974), .B(n1971), .Z(n1972) );
  XNOR U2831 ( .A(n1913), .B(n1903), .Z(n1960) );
  XOR U2832 ( .A(n1978), .B(n1923), .Z(n1913) );
  XNOR U2833 ( .A(n1910), .B(n1911), .Z(n1923) );
  NAND U2834 ( .A(e_input[19]), .B(g_input[21]), .Z(n1911) );
  XNOR U2835 ( .A(n1908), .B(n1979), .Z(n1910) );
  AND U2836 ( .A(g_input[22]), .B(e_input[18]), .Z(n1979) );
  XNOR U2837 ( .A(n1983), .B(n1980), .Z(n1981) );
  XNOR U2838 ( .A(n1922), .B(n1912), .Z(n1978) );
  XOR U2839 ( .A(n1917), .B(n1988), .Z(n1918) );
  AND U2840 ( .A(g_input[24]), .B(e_input[16]), .Z(n1988) );
  XNOR U2841 ( .A(n1992), .B(n1919), .Z(n1987) );
  NAND U2842 ( .A(e_input[17]), .B(g_input[23]), .Z(n1919) );
  IV U2843 ( .A(n1921), .Z(n1992) );
  XOR U2844 ( .A(n1996), .B(n1941), .Z(n1931) );
  XNOR U2845 ( .A(n1928), .B(n1929), .Z(n1941) );
  NAND U2846 ( .A(e_input[27]), .B(g_input[13]), .Z(n1929) );
  XNOR U2847 ( .A(n1926), .B(n1997), .Z(n1928) );
  AND U2848 ( .A(g_input[14]), .B(e_input[26]), .Z(n1997) );
  XNOR U2849 ( .A(n2001), .B(n1998), .Z(n1999) );
  XNOR U2850 ( .A(n1940), .B(n1930), .Z(n1996) );
  XOR U2851 ( .A(n1935), .B(n2006), .Z(n1936) );
  AND U2852 ( .A(g_input[16]), .B(e_input[24]), .Z(n2006) );
  XNOR U2853 ( .A(n2010), .B(n1937), .Z(n2005) );
  NAND U2854 ( .A(e_input[25]), .B(g_input[15]), .Z(n1937) );
  IV U2855 ( .A(n1939), .Z(n2010) );
  XOR U2856 ( .A(n1944), .B(n2015), .Z(n1945) );
  AND U2857 ( .A(g_input[12]), .B(e_input[28]), .Z(n2015) );
  XNOR U2858 ( .A(n2019), .B(n1946), .Z(n2014) );
  NAND U2859 ( .A(e_input[29]), .B(g_input[11]), .Z(n1946) );
  IV U2860 ( .A(n1948), .Z(n2019) );
  XNOR U2861 ( .A(n1954), .B(n1955), .Z(n1950) );
  NAND U2862 ( .A(e_input[31]), .B(g_input[9]), .Z(n1955) );
  XNOR U2863 ( .A(n1952), .B(n2023), .Z(n1954) );
  AND U2864 ( .A(g_input[10]), .B(e_input[30]), .Z(n2023) );
  XNOR U2865 ( .A(n2027), .B(n2024), .Z(n2025) );
  XOR U2866 ( .A(n2029), .B(n1986), .Z(n1976) );
  XOR U2867 ( .A(n1963), .B(n2031), .Z(n1964) );
  AND U2868 ( .A(g_input[19]), .B(e_input[20]), .Z(n2031) );
  XNOR U2869 ( .A(n2035), .B(n1965), .Z(n2030) );
  NAND U2870 ( .A(e_input[21]), .B(g_input[18]), .Z(n1965) );
  IV U2871 ( .A(n1967), .Z(n2035) );
  XNOR U2872 ( .A(n1973), .B(n1974), .Z(n1969) );
  NAND U2873 ( .A(e_input[23]), .B(g_input[16]), .Z(n1974) );
  XNOR U2874 ( .A(n1971), .B(n2039), .Z(n1973) );
  AND U2875 ( .A(g_input[17]), .B(e_input[22]), .Z(n2039) );
  XNOR U2876 ( .A(n2043), .B(n2040), .Z(n2041) );
  XNOR U2877 ( .A(n1985), .B(n1975), .Z(n2029) );
  XOR U2878 ( .A(n2047), .B(n1995), .Z(n1985) );
  XNOR U2879 ( .A(n1982), .B(n1983), .Z(n1995) );
  NAND U2880 ( .A(e_input[19]), .B(g_input[20]), .Z(n1983) );
  XNOR U2881 ( .A(n1980), .B(n2048), .Z(n1982) );
  AND U2882 ( .A(g_input[21]), .B(e_input[18]), .Z(n2048) );
  XNOR U2883 ( .A(n2052), .B(n2049), .Z(n2050) );
  XNOR U2884 ( .A(n1994), .B(n1984), .Z(n2047) );
  XOR U2885 ( .A(n1989), .B(n2057), .Z(n1990) );
  AND U2886 ( .A(g_input[23]), .B(e_input[16]), .Z(n2057) );
  XNOR U2887 ( .A(n2061), .B(n1991), .Z(n2056) );
  NAND U2888 ( .A(e_input[17]), .B(g_input[22]), .Z(n1991) );
  IV U2889 ( .A(n1993), .Z(n2061) );
  XOR U2890 ( .A(n2065), .B(n2013), .Z(n2003) );
  XNOR U2891 ( .A(n2000), .B(n2001), .Z(n2013) );
  NAND U2892 ( .A(e_input[27]), .B(g_input[12]), .Z(n2001) );
  XNOR U2893 ( .A(n1998), .B(n2066), .Z(n2000) );
  AND U2894 ( .A(g_input[13]), .B(e_input[26]), .Z(n2066) );
  XNOR U2895 ( .A(n2070), .B(n2067), .Z(n2068) );
  XNOR U2896 ( .A(n2012), .B(n2002), .Z(n2065) );
  XOR U2897 ( .A(n2007), .B(n2075), .Z(n2008) );
  AND U2898 ( .A(g_input[15]), .B(e_input[24]), .Z(n2075) );
  XNOR U2899 ( .A(n2079), .B(n2009), .Z(n2074) );
  NAND U2900 ( .A(e_input[25]), .B(g_input[14]), .Z(n2009) );
  IV U2901 ( .A(n2011), .Z(n2079) );
  XOR U2902 ( .A(n2016), .B(n2084), .Z(n2017) );
  AND U2903 ( .A(g_input[11]), .B(e_input[28]), .Z(n2084) );
  XNOR U2904 ( .A(n2088), .B(n2018), .Z(n2083) );
  NAND U2905 ( .A(e_input[29]), .B(g_input[10]), .Z(n2018) );
  IV U2906 ( .A(n2020), .Z(n2088) );
  XNOR U2907 ( .A(n2026), .B(n2027), .Z(n2022) );
  NAND U2908 ( .A(e_input[31]), .B(g_input[8]), .Z(n2027) );
  XNOR U2909 ( .A(n2024), .B(n2092), .Z(n2026) );
  AND U2910 ( .A(g_input[9]), .B(e_input[30]), .Z(n2092) );
  XNOR U2911 ( .A(n2096), .B(n2093), .Z(n2094) );
  XNOR U2912 ( .A(n2097), .B(n2098), .Z(n1760) );
  XNOR U2913 ( .A(n2099), .B(n2028), .Z(n2097) );
  XNOR U2914 ( .A(n2101), .B(n2102), .Z(n1764) );
  XNOR U2915 ( .A(n2103), .B(n2100), .Z(n2101) );
  XOR U2916 ( .A(n2104), .B(n2055), .Z(n2045) );
  XOR U2917 ( .A(n2032), .B(n2106), .Z(n2033) );
  AND U2918 ( .A(g_input[18]), .B(e_input[20]), .Z(n2106) );
  XNOR U2919 ( .A(n2110), .B(n2034), .Z(n2105) );
  NAND U2920 ( .A(e_input[21]), .B(g_input[17]), .Z(n2034) );
  IV U2921 ( .A(n2036), .Z(n2110) );
  XNOR U2922 ( .A(n2042), .B(n2043), .Z(n2038) );
  NAND U2923 ( .A(e_input[23]), .B(g_input[15]), .Z(n2043) );
  XNOR U2924 ( .A(n2040), .B(n2114), .Z(n2042) );
  AND U2925 ( .A(g_input[16]), .B(e_input[22]), .Z(n2114) );
  XNOR U2926 ( .A(n2118), .B(n2115), .Z(n2116) );
  XNOR U2927 ( .A(n2054), .B(n2044), .Z(n2104) );
  XOR U2928 ( .A(n2122), .B(n2064), .Z(n2054) );
  XNOR U2929 ( .A(n2051), .B(n2052), .Z(n2064) );
  NAND U2930 ( .A(e_input[19]), .B(g_input[19]), .Z(n2052) );
  XNOR U2931 ( .A(n2049), .B(n2123), .Z(n2051) );
  AND U2932 ( .A(g_input[20]), .B(e_input[18]), .Z(n2123) );
  XNOR U2933 ( .A(n2127), .B(n2124), .Z(n2125) );
  XNOR U2934 ( .A(n2063), .B(n2053), .Z(n2122) );
  XOR U2935 ( .A(n2058), .B(n2132), .Z(n2059) );
  AND U2936 ( .A(g_input[22]), .B(e_input[16]), .Z(n2132) );
  XNOR U2937 ( .A(n2136), .B(n2060), .Z(n2131) );
  NAND U2938 ( .A(e_input[17]), .B(g_input[21]), .Z(n2060) );
  IV U2939 ( .A(n2062), .Z(n2136) );
  XOR U2940 ( .A(n2140), .B(n2082), .Z(n2072) );
  XNOR U2941 ( .A(n2069), .B(n2070), .Z(n2082) );
  NAND U2942 ( .A(e_input[27]), .B(g_input[11]), .Z(n2070) );
  XNOR U2943 ( .A(n2067), .B(n2141), .Z(n2069) );
  AND U2944 ( .A(g_input[12]), .B(e_input[26]), .Z(n2141) );
  XNOR U2945 ( .A(n2145), .B(n2142), .Z(n2143) );
  XNOR U2946 ( .A(n2081), .B(n2071), .Z(n2140) );
  XOR U2947 ( .A(n2076), .B(n2150), .Z(n2077) );
  AND U2948 ( .A(g_input[14]), .B(e_input[24]), .Z(n2150) );
  XNOR U2949 ( .A(n2154), .B(n2078), .Z(n2149) );
  NAND U2950 ( .A(e_input[25]), .B(g_input[13]), .Z(n2078) );
  IV U2951 ( .A(n2080), .Z(n2154) );
  XOR U2952 ( .A(n2085), .B(n2159), .Z(n2086) );
  AND U2953 ( .A(g_input[10]), .B(e_input[28]), .Z(n2159) );
  XNOR U2954 ( .A(n2163), .B(n2087), .Z(n2158) );
  NAND U2955 ( .A(e_input[29]), .B(g_input[9]), .Z(n2087) );
  IV U2956 ( .A(n2089), .Z(n2163) );
  XNOR U2957 ( .A(n2095), .B(n2096), .Z(n2091) );
  NAND U2958 ( .A(e_input[31]), .B(g_input[7]), .Z(n2096) );
  XNOR U2959 ( .A(n2093), .B(n2167), .Z(n2095) );
  AND U2960 ( .A(g_input[8]), .B(e_input[30]), .Z(n2167) );
  XNOR U2961 ( .A(n2171), .B(n2168), .Z(n2169) );
  XNOR U2962 ( .A(n2173), .B(n2174), .Z(n1768) );
  XNOR U2963 ( .A(n2175), .B(n2172), .Z(n2173) );
  XOR U2964 ( .A(n2176), .B(n2130), .Z(n2120) );
  XOR U2965 ( .A(n2107), .B(n2178), .Z(n2108) );
  AND U2966 ( .A(g_input[17]), .B(e_input[20]), .Z(n2178) );
  XNOR U2967 ( .A(n2182), .B(n2109), .Z(n2177) );
  NAND U2968 ( .A(e_input[21]), .B(g_input[16]), .Z(n2109) );
  IV U2969 ( .A(n2111), .Z(n2182) );
  XNOR U2970 ( .A(n2117), .B(n2118), .Z(n2113) );
  NAND U2971 ( .A(e_input[23]), .B(g_input[14]), .Z(n2118) );
  XNOR U2972 ( .A(n2115), .B(n2186), .Z(n2117) );
  AND U2973 ( .A(g_input[15]), .B(e_input[22]), .Z(n2186) );
  XNOR U2974 ( .A(n2190), .B(n2187), .Z(n2188) );
  XNOR U2975 ( .A(n2129), .B(n2119), .Z(n2176) );
  XOR U2976 ( .A(n2194), .B(n2139), .Z(n2129) );
  XNOR U2977 ( .A(n2126), .B(n2127), .Z(n2139) );
  NAND U2978 ( .A(e_input[19]), .B(g_input[18]), .Z(n2127) );
  XNOR U2979 ( .A(n2124), .B(n2195), .Z(n2126) );
  AND U2980 ( .A(g_input[19]), .B(e_input[18]), .Z(n2195) );
  XNOR U2981 ( .A(n2199), .B(n2196), .Z(n2197) );
  XNOR U2982 ( .A(n2138), .B(n2128), .Z(n2194) );
  XOR U2983 ( .A(n2133), .B(n2204), .Z(n2134) );
  AND U2984 ( .A(g_input[21]), .B(e_input[16]), .Z(n2204) );
  XNOR U2985 ( .A(n2208), .B(n2135), .Z(n2203) );
  NAND U2986 ( .A(e_input[17]), .B(g_input[20]), .Z(n2135) );
  IV U2987 ( .A(n2137), .Z(n2208) );
  XOR U2988 ( .A(n2212), .B(n2157), .Z(n2147) );
  XNOR U2989 ( .A(n2144), .B(n2145), .Z(n2157) );
  NAND U2990 ( .A(e_input[27]), .B(g_input[10]), .Z(n2145) );
  XNOR U2991 ( .A(n2142), .B(n2213), .Z(n2144) );
  AND U2992 ( .A(g_input[11]), .B(e_input[26]), .Z(n2213) );
  XNOR U2993 ( .A(n2217), .B(n2214), .Z(n2215) );
  XNOR U2994 ( .A(n2156), .B(n2146), .Z(n2212) );
  XOR U2995 ( .A(n2151), .B(n2222), .Z(n2152) );
  AND U2996 ( .A(g_input[13]), .B(e_input[24]), .Z(n2222) );
  XNOR U2997 ( .A(n2226), .B(n2153), .Z(n2221) );
  NAND U2998 ( .A(e_input[25]), .B(g_input[12]), .Z(n2153) );
  IV U2999 ( .A(n2155), .Z(n2226) );
  XOR U3000 ( .A(n2160), .B(n2231), .Z(n2161) );
  AND U3001 ( .A(g_input[9]), .B(e_input[28]), .Z(n2231) );
  XNOR U3002 ( .A(n2235), .B(n2162), .Z(n2230) );
  NAND U3003 ( .A(e_input[29]), .B(g_input[8]), .Z(n2162) );
  IV U3004 ( .A(n2164), .Z(n2235) );
  XNOR U3005 ( .A(n2170), .B(n2171), .Z(n2166) );
  NAND U3006 ( .A(e_input[31]), .B(g_input[6]), .Z(n2171) );
  XNOR U3007 ( .A(n2168), .B(n2239), .Z(n2170) );
  AND U3008 ( .A(g_input[7]), .B(e_input[30]), .Z(n2239) );
  XNOR U3009 ( .A(n2243), .B(n2240), .Z(n2241) );
  XNOR U3010 ( .A(n2245), .B(n2246), .Z(n1772) );
  XNOR U3011 ( .A(n2247), .B(n2244), .Z(n2245) );
  XOR U3012 ( .A(n2248), .B(n2202), .Z(n2192) );
  XOR U3013 ( .A(n2179), .B(n2250), .Z(n2180) );
  AND U3014 ( .A(g_input[16]), .B(e_input[20]), .Z(n2250) );
  XNOR U3015 ( .A(n2254), .B(n2181), .Z(n2249) );
  NAND U3016 ( .A(e_input[21]), .B(g_input[15]), .Z(n2181) );
  IV U3017 ( .A(n2183), .Z(n2254) );
  XNOR U3018 ( .A(n2189), .B(n2190), .Z(n2185) );
  NAND U3019 ( .A(e_input[23]), .B(g_input[13]), .Z(n2190) );
  XNOR U3020 ( .A(n2187), .B(n2258), .Z(n2189) );
  AND U3021 ( .A(g_input[14]), .B(e_input[22]), .Z(n2258) );
  XNOR U3022 ( .A(n2262), .B(n2259), .Z(n2260) );
  XNOR U3023 ( .A(n2201), .B(n2191), .Z(n2248) );
  XOR U3024 ( .A(n2266), .B(n2211), .Z(n2201) );
  XNOR U3025 ( .A(n2198), .B(n2199), .Z(n2211) );
  NAND U3026 ( .A(e_input[19]), .B(g_input[17]), .Z(n2199) );
  XNOR U3027 ( .A(n2196), .B(n2267), .Z(n2198) );
  AND U3028 ( .A(g_input[18]), .B(e_input[18]), .Z(n2267) );
  XNOR U3029 ( .A(n2271), .B(n2268), .Z(n2269) );
  XNOR U3030 ( .A(n2210), .B(n2200), .Z(n2266) );
  XOR U3031 ( .A(n2205), .B(n2276), .Z(n2206) );
  AND U3032 ( .A(g_input[20]), .B(e_input[16]), .Z(n2276) );
  XNOR U3033 ( .A(n2280), .B(n2207), .Z(n2275) );
  NAND U3034 ( .A(e_input[17]), .B(g_input[19]), .Z(n2207) );
  IV U3035 ( .A(n2209), .Z(n2280) );
  XOR U3036 ( .A(n2284), .B(n2229), .Z(n2219) );
  XNOR U3037 ( .A(n2216), .B(n2217), .Z(n2229) );
  NAND U3038 ( .A(e_input[27]), .B(g_input[9]), .Z(n2217) );
  XNOR U3039 ( .A(n2214), .B(n2285), .Z(n2216) );
  AND U3040 ( .A(g_input[10]), .B(e_input[26]), .Z(n2285) );
  XNOR U3041 ( .A(n2289), .B(n2286), .Z(n2287) );
  XNOR U3042 ( .A(n2228), .B(n2218), .Z(n2284) );
  XOR U3043 ( .A(n2223), .B(n2294), .Z(n2224) );
  AND U3044 ( .A(g_input[12]), .B(e_input[24]), .Z(n2294) );
  XNOR U3045 ( .A(n2298), .B(n2225), .Z(n2293) );
  NAND U3046 ( .A(e_input[25]), .B(g_input[11]), .Z(n2225) );
  IV U3047 ( .A(n2227), .Z(n2298) );
  XOR U3048 ( .A(n2232), .B(n2303), .Z(n2233) );
  AND U3049 ( .A(g_input[8]), .B(e_input[28]), .Z(n2303) );
  XNOR U3050 ( .A(n2307), .B(n2234), .Z(n2302) );
  NAND U3051 ( .A(e_input[29]), .B(g_input[7]), .Z(n2234) );
  IV U3052 ( .A(n2236), .Z(n2307) );
  XNOR U3053 ( .A(n2242), .B(n2243), .Z(n2238) );
  NAND U3054 ( .A(e_input[31]), .B(g_input[5]), .Z(n2243) );
  XNOR U3055 ( .A(n2240), .B(n2311), .Z(n2242) );
  AND U3056 ( .A(g_input[6]), .B(e_input[30]), .Z(n2311) );
  XNOR U3057 ( .A(n2315), .B(n2312), .Z(n2313) );
  XOR U3058 ( .A(n2317), .B(n2274), .Z(n2264) );
  XOR U3059 ( .A(n2251), .B(n2319), .Z(n2252) );
  AND U3060 ( .A(g_input[15]), .B(e_input[20]), .Z(n2319) );
  XNOR U3061 ( .A(n2323), .B(n2253), .Z(n2318) );
  NAND U3062 ( .A(e_input[21]), .B(g_input[14]), .Z(n2253) );
  IV U3063 ( .A(n2255), .Z(n2323) );
  XNOR U3064 ( .A(n2261), .B(n2262), .Z(n2257) );
  NAND U3065 ( .A(e_input[23]), .B(g_input[12]), .Z(n2262) );
  XNOR U3066 ( .A(n2259), .B(n2327), .Z(n2261) );
  AND U3067 ( .A(g_input[13]), .B(e_input[22]), .Z(n2327) );
  XNOR U3068 ( .A(n2331), .B(n2328), .Z(n2329) );
  XNOR U3069 ( .A(n2273), .B(n2263), .Z(n2317) );
  XOR U3070 ( .A(n2335), .B(n2283), .Z(n2273) );
  XNOR U3071 ( .A(n2270), .B(n2271), .Z(n2283) );
  NAND U3072 ( .A(e_input[19]), .B(g_input[16]), .Z(n2271) );
  XNOR U3073 ( .A(n2268), .B(n2336), .Z(n2270) );
  AND U3074 ( .A(g_input[17]), .B(e_input[18]), .Z(n2336) );
  XNOR U3075 ( .A(n2340), .B(n2337), .Z(n2338) );
  XNOR U3076 ( .A(n2282), .B(n2272), .Z(n2335) );
  XOR U3077 ( .A(n2277), .B(n2345), .Z(n2278) );
  AND U3078 ( .A(g_input[19]), .B(e_input[16]), .Z(n2345) );
  XNOR U3079 ( .A(n2349), .B(n2279), .Z(n2344) );
  NAND U3080 ( .A(e_input[17]), .B(g_input[18]), .Z(n2279) );
  IV U3081 ( .A(n2281), .Z(n2349) );
  XOR U3082 ( .A(n2353), .B(n2301), .Z(n2291) );
  XNOR U3083 ( .A(n2288), .B(n2289), .Z(n2301) );
  NAND U3084 ( .A(e_input[27]), .B(g_input[8]), .Z(n2289) );
  XNOR U3085 ( .A(n2286), .B(n2354), .Z(n2288) );
  AND U3086 ( .A(g_input[9]), .B(e_input[26]), .Z(n2354) );
  XNOR U3087 ( .A(n2358), .B(n2355), .Z(n2356) );
  XNOR U3088 ( .A(n2300), .B(n2290), .Z(n2353) );
  XOR U3089 ( .A(n2295), .B(n2363), .Z(n2296) );
  AND U3090 ( .A(g_input[11]), .B(e_input[24]), .Z(n2363) );
  XNOR U3091 ( .A(n2367), .B(n2297), .Z(n2362) );
  NAND U3092 ( .A(e_input[25]), .B(g_input[10]), .Z(n2297) );
  IV U3093 ( .A(n2299), .Z(n2367) );
  XOR U3094 ( .A(n2304), .B(n2372), .Z(n2305) );
  AND U3095 ( .A(g_input[7]), .B(e_input[28]), .Z(n2372) );
  XNOR U3096 ( .A(n2376), .B(n2306), .Z(n2371) );
  NAND U3097 ( .A(e_input[29]), .B(g_input[6]), .Z(n2306) );
  IV U3098 ( .A(n2308), .Z(n2376) );
  XNOR U3099 ( .A(n2314), .B(n2315), .Z(n2310) );
  NAND U3100 ( .A(e_input[31]), .B(g_input[4]), .Z(n2315) );
  XNOR U3101 ( .A(n2312), .B(n2380), .Z(n2314) );
  AND U3102 ( .A(g_input[5]), .B(e_input[30]), .Z(n2380) );
  XNOR U3103 ( .A(n2384), .B(n2381), .Z(n2382) );
  XNOR U3104 ( .A(n2385), .B(n2386), .Z(n1776) );
  XNOR U3105 ( .A(n2387), .B(n2316), .Z(n2385) );
  XNOR U3106 ( .A(n2389), .B(n2390), .Z(n1780) );
  XNOR U3107 ( .A(n2391), .B(n2388), .Z(n2389) );
  XOR U3108 ( .A(n2392), .B(n2343), .Z(n2333) );
  XOR U3109 ( .A(n2320), .B(n2394), .Z(n2321) );
  AND U3110 ( .A(g_input[14]), .B(e_input[20]), .Z(n2394) );
  XNOR U3111 ( .A(n2398), .B(n2322), .Z(n2393) );
  NAND U3112 ( .A(e_input[21]), .B(g_input[13]), .Z(n2322) );
  IV U3113 ( .A(n2324), .Z(n2398) );
  XNOR U3114 ( .A(n2330), .B(n2331), .Z(n2326) );
  NAND U3115 ( .A(e_input[23]), .B(g_input[11]), .Z(n2331) );
  XNOR U3116 ( .A(n2328), .B(n2402), .Z(n2330) );
  AND U3117 ( .A(g_input[12]), .B(e_input[22]), .Z(n2402) );
  XNOR U3118 ( .A(n2406), .B(n2403), .Z(n2404) );
  XNOR U3119 ( .A(n2342), .B(n2332), .Z(n2392) );
  XOR U3120 ( .A(n2410), .B(n2352), .Z(n2342) );
  XNOR U3121 ( .A(n2339), .B(n2340), .Z(n2352) );
  NAND U3122 ( .A(e_input[19]), .B(g_input[15]), .Z(n2340) );
  XNOR U3123 ( .A(n2337), .B(n2411), .Z(n2339) );
  AND U3124 ( .A(g_input[16]), .B(e_input[18]), .Z(n2411) );
  XNOR U3125 ( .A(n2415), .B(n2412), .Z(n2413) );
  XNOR U3126 ( .A(n2351), .B(n2341), .Z(n2410) );
  XOR U3127 ( .A(n2346), .B(n2420), .Z(n2347) );
  AND U3128 ( .A(g_input[18]), .B(e_input[16]), .Z(n2420) );
  XNOR U3129 ( .A(n2424), .B(n2348), .Z(n2419) );
  NAND U3130 ( .A(e_input[17]), .B(g_input[17]), .Z(n2348) );
  IV U3131 ( .A(n2350), .Z(n2424) );
  XOR U3132 ( .A(n2428), .B(n2370), .Z(n2360) );
  XNOR U3133 ( .A(n2357), .B(n2358), .Z(n2370) );
  NAND U3134 ( .A(e_input[27]), .B(g_input[7]), .Z(n2358) );
  XNOR U3135 ( .A(n2355), .B(n2429), .Z(n2357) );
  AND U3136 ( .A(g_input[8]), .B(e_input[26]), .Z(n2429) );
  XNOR U3137 ( .A(n2433), .B(n2430), .Z(n2431) );
  XNOR U3138 ( .A(n2369), .B(n2359), .Z(n2428) );
  XOR U3139 ( .A(n2364), .B(n2438), .Z(n2365) );
  AND U3140 ( .A(g_input[10]), .B(e_input[24]), .Z(n2438) );
  XNOR U3141 ( .A(n2442), .B(n2366), .Z(n2437) );
  NAND U3142 ( .A(e_input[25]), .B(g_input[9]), .Z(n2366) );
  IV U3143 ( .A(n2368), .Z(n2442) );
  XOR U3144 ( .A(n2373), .B(n2447), .Z(n2374) );
  AND U3145 ( .A(g_input[6]), .B(e_input[28]), .Z(n2447) );
  XNOR U3146 ( .A(n2451), .B(n2375), .Z(n2446) );
  NAND U3147 ( .A(e_input[29]), .B(g_input[5]), .Z(n2375) );
  IV U3148 ( .A(n2377), .Z(n2451) );
  XNOR U3149 ( .A(n2383), .B(n2384), .Z(n2379) );
  NAND U3150 ( .A(e_input[31]), .B(g_input[3]), .Z(n2384) );
  XNOR U3151 ( .A(n2381), .B(n2455), .Z(n2383) );
  AND U3152 ( .A(g_input[4]), .B(e_input[30]), .Z(n2455) );
  XNOR U3153 ( .A(n2459), .B(n2456), .Z(n2457) );
  XNOR U3154 ( .A(n2463), .B(n1792), .Z(n1796) );
  XNOR U3155 ( .A(n1791), .B(n1790), .Z(n1792) );
  NAND U3156 ( .A(e_input[11]), .B(g_input[31]), .Z(n1790) );
  XNOR U3157 ( .A(n2467), .B(n2464), .Z(n2465) );
  XNOR U3158 ( .A(n1787), .B(n1793), .Z(n2463) );
  XNOR U3159 ( .A(n2471), .B(n2474), .Z(n2473) );
  XOR U3160 ( .A(n1800), .B(n2476), .Z(n1801) );
  AND U3161 ( .A(e_input[12]), .B(g_input[30]), .Z(n2476) );
  XNOR U3162 ( .A(n2480), .B(n1802), .Z(n2475) );
  NAND U3163 ( .A(g_input[29]), .B(e_input[13]), .Z(n1802) );
  IV U3164 ( .A(n1804), .Z(n2480) );
  XOR U3165 ( .A(n2481), .B(n2482), .Z(n1804) );
  AND U3166 ( .A(n2483), .B(n2484), .Z(n2482) );
  XNOR U3167 ( .A(n2481), .B(n2485), .Z(n2483) );
  XNOR U3168 ( .A(n1810), .B(n1811), .Z(n1806) );
  NAND U3169 ( .A(g_input[27]), .B(e_input[15]), .Z(n1811) );
  XNOR U3170 ( .A(n1808), .B(n2486), .Z(n1810) );
  AND U3171 ( .A(e_input[14]), .B(g_input[28]), .Z(n2486) );
  XNOR U3172 ( .A(n2490), .B(n2487), .Z(n2488) );
  XOR U3173 ( .A(n2491), .B(n2474), .Z(n2469) );
  XNOR U3174 ( .A(n2466), .B(n2467), .Z(n2474) );
  NAND U3175 ( .A(g_input[30]), .B(e_input[11]), .Z(n2467) );
  XNOR U3176 ( .A(n2464), .B(n2492), .Z(n2466) );
  AND U3177 ( .A(e_input[10]), .B(g_input[31]), .Z(n2492) );
  XNOR U3178 ( .A(n2496), .B(n2493), .Z(n2494) );
  XNOR U3179 ( .A(n2472), .B(n2468), .Z(n2491) );
  XOR U3180 ( .A(n2471), .B(n2500), .Z(n2472) );
  ANDN U3181 ( .A(n2501), .B(n2502), .Z(n2500) );
  XOR U3182 ( .A(n2477), .B(n2507), .Z(n2478) );
  AND U3183 ( .A(e_input[12]), .B(g_input[29]), .Z(n2507) );
  XNOR U3184 ( .A(n2511), .B(n2479), .Z(n2506) );
  NAND U3185 ( .A(g_input[28]), .B(e_input[13]), .Z(n2479) );
  IV U3186 ( .A(n2481), .Z(n2511) );
  XNOR U3187 ( .A(n2489), .B(n2490), .Z(n2485) );
  NAND U3188 ( .A(g_input[26]), .B(e_input[15]), .Z(n2490) );
  XNOR U3189 ( .A(n2487), .B(n2515), .Z(n2489) );
  AND U3190 ( .A(e_input[14]), .B(g_input[27]), .Z(n2515) );
  XNOR U3191 ( .A(n2519), .B(n2516), .Z(n2517) );
  XOR U3192 ( .A(n2520), .B(n2505), .Z(n2498) );
  XNOR U3193 ( .A(n2495), .B(n2496), .Z(n2505) );
  NAND U3194 ( .A(g_input[29]), .B(e_input[11]), .Z(n2496) );
  XNOR U3195 ( .A(n2493), .B(n2521), .Z(n2495) );
  AND U3196 ( .A(e_input[10]), .B(g_input[30]), .Z(n2521) );
  XNOR U3197 ( .A(n2525), .B(n2522), .Z(n2523) );
  XNOR U3198 ( .A(n2504), .B(n2497), .Z(n2520) );
  XNOR U3199 ( .A(n2533), .B(n2502), .Z(n2529) );
  NAND U3200 ( .A(g_input[31]), .B(e_input[9]), .Z(n2502) );
  IV U3201 ( .A(n2503), .Z(n2533) );
  XOR U3202 ( .A(n2508), .B(n2538), .Z(n2509) );
  AND U3203 ( .A(e_input[12]), .B(g_input[28]), .Z(n2538) );
  XNOR U3204 ( .A(n2542), .B(n2510), .Z(n2537) );
  NAND U3205 ( .A(g_input[27]), .B(e_input[13]), .Z(n2510) );
  IV U3206 ( .A(n2512), .Z(n2542) );
  XNOR U3207 ( .A(n2518), .B(n2519), .Z(n2514) );
  NAND U3208 ( .A(g_input[25]), .B(e_input[15]), .Z(n2519) );
  XNOR U3209 ( .A(n2516), .B(n2546), .Z(n2518) );
  AND U3210 ( .A(e_input[14]), .B(g_input[26]), .Z(n2546) );
  XNOR U3211 ( .A(n2550), .B(n2547), .Z(n2548) );
  XNOR U3212 ( .A(n2552), .B(n2553), .Z(n2099) );
  XOR U3213 ( .A(n2554), .B(n2555), .Z(n2553) );
  AND U3214 ( .A(n2556), .B(n2557), .Z(n2554) );
  OR U3215 ( .A(n2558), .B(n2559), .Z(n2557) );
  AND U3216 ( .A(n2560), .B(n2561), .Z(n2556) );
  NAND U3217 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U3218 ( .B(n2564), .A(n2555), .Z(n2560) );
  XOR U3219 ( .A(n2565), .B(n2536), .Z(n2527) );
  XNOR U3220 ( .A(n2524), .B(n2525), .Z(n2536) );
  NAND U3221 ( .A(g_input[28]), .B(e_input[11]), .Z(n2525) );
  XNOR U3222 ( .A(n2522), .B(n2566), .Z(n2524) );
  AND U3223 ( .A(e_input[10]), .B(g_input[29]), .Z(n2566) );
  XNOR U3224 ( .A(n2570), .B(n2567), .Z(n2568) );
  XNOR U3225 ( .A(n2535), .B(n2526), .Z(n2565) );
  XOR U3226 ( .A(n2530), .B(n2575), .Z(n2531) );
  AND U3227 ( .A(e_input[8]), .B(g_input[31]), .Z(n2575) );
  XOR U3228 ( .A(n2576), .B(n2577), .Z(n2530) );
  AND U3229 ( .A(n2578), .B(n2579), .Z(n2577) );
  XNOR U3230 ( .A(n2580), .B(n2576), .Z(n2578) );
  XNOR U3231 ( .A(n2581), .B(n2532), .Z(n2574) );
  NAND U3232 ( .A(g_input[30]), .B(e_input[9]), .Z(n2532) );
  IV U3233 ( .A(n2534), .Z(n2581) );
  XOR U3234 ( .A(n2539), .B(n2586), .Z(n2540) );
  AND U3235 ( .A(e_input[12]), .B(g_input[27]), .Z(n2586) );
  XNOR U3236 ( .A(n2590), .B(n2541), .Z(n2585) );
  NAND U3237 ( .A(g_input[26]), .B(e_input[13]), .Z(n2541) );
  IV U3238 ( .A(n2543), .Z(n2590) );
  XNOR U3239 ( .A(n2549), .B(n2550), .Z(n2545) );
  NAND U3240 ( .A(g_input[24]), .B(e_input[15]), .Z(n2550) );
  XNOR U3241 ( .A(n2547), .B(n2594), .Z(n2549) );
  AND U3242 ( .A(e_input[14]), .B(g_input[25]), .Z(n2594) );
  XNOR U3243 ( .A(n2598), .B(n2595), .Z(n2596) );
  XOR U3244 ( .A(n2600), .B(n2584), .Z(n2572) );
  XNOR U3245 ( .A(n2569), .B(n2570), .Z(n2584) );
  NAND U3246 ( .A(g_input[27]), .B(e_input[11]), .Z(n2570) );
  XNOR U3247 ( .A(n2567), .B(n2601), .Z(n2569) );
  AND U3248 ( .A(e_input[10]), .B(g_input[28]), .Z(n2601) );
  XNOR U3249 ( .A(n2605), .B(n2602), .Z(n2603) );
  XNOR U3250 ( .A(n2583), .B(n2571), .Z(n2600) );
  XOR U3251 ( .A(n2576), .B(n2610), .Z(n2579) );
  AND U3252 ( .A(e_input[8]), .B(g_input[30]), .Z(n2610) );
  XNOR U3253 ( .A(n2614), .B(n2580), .Z(n2609) );
  NAND U3254 ( .A(g_input[29]), .B(e_input[9]), .Z(n2580) );
  IV U3255 ( .A(n2582), .Z(n2614) );
  XOR U3256 ( .A(n2587), .B(n2619), .Z(n2588) );
  AND U3257 ( .A(e_input[12]), .B(g_input[26]), .Z(n2619) );
  XNOR U3258 ( .A(n2623), .B(n2589), .Z(n2618) );
  NAND U3259 ( .A(g_input[25]), .B(e_input[13]), .Z(n2589) );
  IV U3260 ( .A(n2591), .Z(n2623) );
  XNOR U3261 ( .A(n2597), .B(n2598), .Z(n2593) );
  NAND U3262 ( .A(g_input[23]), .B(e_input[15]), .Z(n2598) );
  XNOR U3263 ( .A(n2595), .B(n2627), .Z(n2597) );
  AND U3264 ( .A(e_input[14]), .B(g_input[24]), .Z(n2627) );
  XNOR U3265 ( .A(n2631), .B(n2628), .Z(n2629) );
  XOR U3266 ( .A(n2632), .B(n2559), .Z(n2103) );
  XNOR U3267 ( .A(n2564), .B(n2555), .Z(n2559) );
  XNOR U3268 ( .A(n2563), .B(n2562), .Z(n2564) );
  NAND U3269 ( .A(e_input[7]), .B(g_input[31]), .Z(n2562) );
  XNOR U3270 ( .A(n2639), .B(n2636), .Z(n2637) );
  OR U3271 ( .A(n2640), .B(n2641), .Z(n2558) );
  XOR U3272 ( .A(n2643), .B(n2617), .Z(n2607) );
  XNOR U3273 ( .A(n2604), .B(n2605), .Z(n2617) );
  NAND U3274 ( .A(g_input[26]), .B(e_input[11]), .Z(n2605) );
  XNOR U3275 ( .A(n2602), .B(n2644), .Z(n2604) );
  AND U3276 ( .A(e_input[10]), .B(g_input[27]), .Z(n2644) );
  XNOR U3277 ( .A(n2648), .B(n2645), .Z(n2646) );
  XNOR U3278 ( .A(n2616), .B(n2606), .Z(n2643) );
  XOR U3279 ( .A(n2611), .B(n2653), .Z(n2612) );
  AND U3280 ( .A(e_input[8]), .B(g_input[29]), .Z(n2653) );
  XNOR U3281 ( .A(n2657), .B(n2613), .Z(n2652) );
  NAND U3282 ( .A(g_input[28]), .B(e_input[9]), .Z(n2613) );
  IV U3283 ( .A(n2615), .Z(n2657) );
  XOR U3284 ( .A(n2620), .B(n2662), .Z(n2621) );
  AND U3285 ( .A(e_input[12]), .B(g_input[25]), .Z(n2662) );
  XNOR U3286 ( .A(n2666), .B(n2622), .Z(n2661) );
  NAND U3287 ( .A(g_input[24]), .B(e_input[13]), .Z(n2622) );
  IV U3288 ( .A(n2624), .Z(n2666) );
  XNOR U3289 ( .A(n2630), .B(n2631), .Z(n2626) );
  NAND U3290 ( .A(g_input[22]), .B(e_input[15]), .Z(n2631) );
  XNOR U3291 ( .A(n2628), .B(n2670), .Z(n2630) );
  AND U3292 ( .A(e_input[14]), .B(g_input[23]), .Z(n2670) );
  XNOR U3293 ( .A(n2674), .B(n2671), .Z(n2672) );
  XOR U3294 ( .A(n2675), .B(n2641), .Z(n2175) );
  XOR U3295 ( .A(n2633), .B(n2676), .Z(n2634) );
  ANDN U3296 ( .A(n2677), .B(n2678), .Z(n2676) );
  XNOR U3297 ( .A(n2638), .B(n2639), .Z(n2635) );
  NAND U3298 ( .A(g_input[30]), .B(e_input[7]), .Z(n2639) );
  XNOR U3299 ( .A(n2636), .B(n2682), .Z(n2638) );
  AND U3300 ( .A(e_input[6]), .B(g_input[31]), .Z(n2682) );
  XNOR U3301 ( .A(n2686), .B(n2683), .Z(n2684) );
  NANDN U3302 ( .B(n2687), .A(n2688), .Z(n2640) );
  XOR U3303 ( .A(n2690), .B(n2660), .Z(n2650) );
  XNOR U3304 ( .A(n2647), .B(n2648), .Z(n2660) );
  NAND U3305 ( .A(g_input[25]), .B(e_input[11]), .Z(n2648) );
  XNOR U3306 ( .A(n2645), .B(n2691), .Z(n2647) );
  AND U3307 ( .A(e_input[10]), .B(g_input[26]), .Z(n2691) );
  XNOR U3308 ( .A(n2695), .B(n2692), .Z(n2693) );
  XNOR U3309 ( .A(n2659), .B(n2649), .Z(n2690) );
  XOR U3310 ( .A(n2654), .B(n2700), .Z(n2655) );
  AND U3311 ( .A(e_input[8]), .B(g_input[28]), .Z(n2700) );
  XNOR U3312 ( .A(n2704), .B(n2656), .Z(n2699) );
  NAND U3313 ( .A(g_input[27]), .B(e_input[9]), .Z(n2656) );
  IV U3314 ( .A(n2658), .Z(n2704) );
  XOR U3315 ( .A(n2663), .B(n2709), .Z(n2664) );
  AND U3316 ( .A(e_input[12]), .B(g_input[24]), .Z(n2709) );
  XNOR U3317 ( .A(n2713), .B(n2665), .Z(n2708) );
  NAND U3318 ( .A(g_input[23]), .B(e_input[13]), .Z(n2665) );
  IV U3319 ( .A(n2667), .Z(n2713) );
  XNOR U3320 ( .A(n2673), .B(n2674), .Z(n2669) );
  NAND U3321 ( .A(g_input[21]), .B(e_input[15]), .Z(n2674) );
  XNOR U3322 ( .A(n2671), .B(n2717), .Z(n2673) );
  AND U3323 ( .A(e_input[14]), .B(g_input[22]), .Z(n2717) );
  XNOR U3324 ( .A(n2721), .B(n2718), .Z(n2719) );
  XOR U3325 ( .A(n2722), .B(n2687), .Z(n2247) );
  XNOR U3326 ( .A(n2727), .B(n2678), .Z(n2723) );
  NAND U3327 ( .A(g_input[31]), .B(e_input[5]), .Z(n2678) );
  IV U3328 ( .A(n2679), .Z(n2727) );
  XNOR U3329 ( .A(n2685), .B(n2686), .Z(n2681) );
  NAND U3330 ( .A(g_input[29]), .B(e_input[7]), .Z(n2686) );
  XNOR U3331 ( .A(n2683), .B(n2731), .Z(n2685) );
  AND U3332 ( .A(e_input[6]), .B(g_input[30]), .Z(n2731) );
  XNOR U3333 ( .A(n2735), .B(n2732), .Z(n2733) );
  XNOR U3334 ( .A(n2688), .B(n2689), .Z(n2722) );
  XOR U3335 ( .A(n2740), .B(n2738), .Z(n2387) );
  XOR U3336 ( .A(n2724), .B(n2742), .Z(n2725) );
  AND U3337 ( .A(e_input[4]), .B(g_input[31]), .Z(n2742) );
  XNOR U3338 ( .A(n2746), .B(n2726), .Z(n2741) );
  NAND U3339 ( .A(g_input[30]), .B(e_input[5]), .Z(n2726) );
  IV U3340 ( .A(n2728), .Z(n2746) );
  XNOR U3341 ( .A(n2734), .B(n2735), .Z(n2730) );
  NAND U3342 ( .A(g_input[28]), .B(e_input[7]), .Z(n2735) );
  XNOR U3343 ( .A(n2732), .B(n2750), .Z(n2734) );
  AND U3344 ( .A(e_input[6]), .B(g_input[29]), .Z(n2750) );
  XNOR U3345 ( .A(n2754), .B(n2751), .Z(n2752) );
  XNOR U3346 ( .A(n2737), .B(n2739), .Z(n2740) );
  XNOR U3347 ( .A(n2755), .B(n2756), .Z(n2737) );
  XOR U3348 ( .A(n2757), .B(n2758), .Z(n2756) );
  AND U3349 ( .A(n2759), .B(n2760), .Z(n2757) );
  NAND U3350 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U3351 ( .B(n2763), .A(n2758), .Z(n2759) );
  XOR U3352 ( .A(n2767), .B(n2707), .Z(n2697) );
  XNOR U3353 ( .A(n2694), .B(n2695), .Z(n2707) );
  NAND U3354 ( .A(g_input[24]), .B(e_input[11]), .Z(n2695) );
  XNOR U3355 ( .A(n2692), .B(n2768), .Z(n2694) );
  AND U3356 ( .A(e_input[10]), .B(g_input[25]), .Z(n2768) );
  XNOR U3357 ( .A(n2772), .B(n2769), .Z(n2770) );
  XNOR U3358 ( .A(n2706), .B(n2696), .Z(n2767) );
  XOR U3359 ( .A(n2701), .B(n2777), .Z(n2702) );
  AND U3360 ( .A(e_input[8]), .B(g_input[27]), .Z(n2777) );
  XNOR U3361 ( .A(n2781), .B(n2703), .Z(n2776) );
  NAND U3362 ( .A(g_input[26]), .B(e_input[9]), .Z(n2703) );
  IV U3363 ( .A(n2705), .Z(n2781) );
  XOR U3364 ( .A(n2710), .B(n2786), .Z(n2711) );
  AND U3365 ( .A(e_input[12]), .B(g_input[23]), .Z(n2786) );
  XNOR U3366 ( .A(n2790), .B(n2712), .Z(n2785) );
  NAND U3367 ( .A(g_input[22]), .B(e_input[13]), .Z(n2712) );
  IV U3368 ( .A(n2714), .Z(n2790) );
  XNOR U3369 ( .A(n2720), .B(n2721), .Z(n2716) );
  NAND U3370 ( .A(g_input[20]), .B(e_input[15]), .Z(n2721) );
  XNOR U3371 ( .A(n2718), .B(n2794), .Z(n2720) );
  AND U3372 ( .A(e_input[14]), .B(g_input[21]), .Z(n2794) );
  XNOR U3373 ( .A(n2798), .B(n2795), .Z(n2796) );
  XOR U3374 ( .A(n2800), .B(n2784), .Z(n2774) );
  XNOR U3375 ( .A(n2771), .B(n2772), .Z(n2784) );
  NAND U3376 ( .A(g_input[23]), .B(e_input[11]), .Z(n2772) );
  XNOR U3377 ( .A(n2769), .B(n2801), .Z(n2771) );
  AND U3378 ( .A(e_input[10]), .B(g_input[24]), .Z(n2801) );
  XNOR U3379 ( .A(n2805), .B(n2802), .Z(n2803) );
  XNOR U3380 ( .A(n2783), .B(n2773), .Z(n2800) );
  XOR U3381 ( .A(n2778), .B(n2810), .Z(n2779) );
  AND U3382 ( .A(e_input[8]), .B(g_input[26]), .Z(n2810) );
  XNOR U3383 ( .A(n2814), .B(n2780), .Z(n2809) );
  NAND U3384 ( .A(g_input[25]), .B(e_input[9]), .Z(n2780) );
  IV U3385 ( .A(n2782), .Z(n2814) );
  XOR U3386 ( .A(n2787), .B(n2819), .Z(n2788) );
  AND U3387 ( .A(e_input[12]), .B(g_input[22]), .Z(n2819) );
  XNOR U3388 ( .A(n2823), .B(n2789), .Z(n2818) );
  NAND U3389 ( .A(g_input[21]), .B(e_input[13]), .Z(n2789) );
  IV U3390 ( .A(n2791), .Z(n2823) );
  XNOR U3391 ( .A(n2797), .B(n2798), .Z(n2793) );
  NAND U3392 ( .A(g_input[19]), .B(e_input[15]), .Z(n2798) );
  XNOR U3393 ( .A(n2795), .B(n2827), .Z(n2797) );
  AND U3394 ( .A(e_input[14]), .B(g_input[20]), .Z(n2827) );
  XNOR U3395 ( .A(n2831), .B(n2828), .Z(n2829) );
  XOR U3396 ( .A(n2832), .B(n2766), .Z(n2391) );
  XOR U3397 ( .A(n2743), .B(n2834), .Z(n2744) );
  AND U3398 ( .A(e_input[4]), .B(g_input[30]), .Z(n2834) );
  XNOR U3399 ( .A(n2838), .B(n2745), .Z(n2833) );
  NAND U3400 ( .A(g_input[29]), .B(e_input[5]), .Z(n2745) );
  IV U3401 ( .A(n2747), .Z(n2838) );
  XNOR U3402 ( .A(n2753), .B(n2754), .Z(n2749) );
  NAND U3403 ( .A(g_input[27]), .B(e_input[7]), .Z(n2754) );
  XNOR U3404 ( .A(n2751), .B(n2842), .Z(n2753) );
  AND U3405 ( .A(e_input[6]), .B(g_input[28]), .Z(n2842) );
  XNOR U3406 ( .A(n2846), .B(n2843), .Z(n2844) );
  XOR U3407 ( .A(n2765), .B(n2799), .Z(n2832) );
  XOR U3408 ( .A(n2847), .B(n2763), .Z(n2765) );
  XNOR U3409 ( .A(n2762), .B(n2761), .Z(n2763) );
  NAND U3410 ( .A(e_input[3]), .B(g_input[31]), .Z(n2761) );
  XNOR U3411 ( .A(n2851), .B(n2848), .Z(n2849) );
  XNOR U3412 ( .A(n2758), .B(n2764), .Z(n2847) );
  XNOR U3413 ( .A(n2855), .B(n2858), .Z(n2857) );
  XNOR U3414 ( .A(o_reg[1]), .B(n1782), .Z(o[0]) );
  XNOR U3415 ( .A(n2862), .B(n2461), .Z(n1782) );
  XNOR U3416 ( .A(n2863), .B(n2861), .Z(n2461) );
  XOR U3417 ( .A(n2864), .B(n2817), .Z(n2807) );
  XNOR U3418 ( .A(n2804), .B(n2805), .Z(n2817) );
  NAND U3419 ( .A(g_input[22]), .B(e_input[11]), .Z(n2805) );
  XNOR U3420 ( .A(n2802), .B(n2865), .Z(n2804) );
  AND U3421 ( .A(e_input[10]), .B(g_input[23]), .Z(n2865) );
  XNOR U3422 ( .A(n2869), .B(n2866), .Z(n2867) );
  XNOR U3423 ( .A(n2816), .B(n2806), .Z(n2864) );
  XOR U3424 ( .A(n2811), .B(n2874), .Z(n2812) );
  AND U3425 ( .A(e_input[8]), .B(g_input[25]), .Z(n2874) );
  XNOR U3426 ( .A(n2878), .B(n2813), .Z(n2873) );
  NAND U3427 ( .A(g_input[24]), .B(e_input[9]), .Z(n2813) );
  IV U3428 ( .A(n2815), .Z(n2878) );
  XOR U3429 ( .A(n2820), .B(n2883), .Z(n2821) );
  AND U3430 ( .A(e_input[12]), .B(g_input[21]), .Z(n2883) );
  XNOR U3431 ( .A(n2887), .B(n2822), .Z(n2882) );
  NAND U3432 ( .A(g_input[20]), .B(e_input[13]), .Z(n2822) );
  IV U3433 ( .A(n2824), .Z(n2887) );
  XNOR U3434 ( .A(n2830), .B(n2831), .Z(n2826) );
  NAND U3435 ( .A(g_input[18]), .B(e_input[15]), .Z(n2831) );
  XNOR U3436 ( .A(n2828), .B(n2891), .Z(n2830) );
  AND U3437 ( .A(e_input[14]), .B(g_input[19]), .Z(n2891) );
  XNOR U3438 ( .A(n2895), .B(n2892), .Z(n2893) );
  XNOR U3439 ( .A(n2860), .B(n2460), .Z(n2863) );
  XOR U3440 ( .A(n2899), .B(n2854), .Z(n2860) );
  XOR U3441 ( .A(n2835), .B(n2901), .Z(n2836) );
  AND U3442 ( .A(e_input[4]), .B(g_input[29]), .Z(n2901) );
  XNOR U3443 ( .A(n2905), .B(n2837), .Z(n2900) );
  NAND U3444 ( .A(g_input[28]), .B(e_input[5]), .Z(n2837) );
  IV U3445 ( .A(n2839), .Z(n2905) );
  XNOR U3446 ( .A(n2845), .B(n2846), .Z(n2841) );
  NAND U3447 ( .A(g_input[26]), .B(e_input[7]), .Z(n2846) );
  XNOR U3448 ( .A(n2843), .B(n2909), .Z(n2845) );
  AND U3449 ( .A(e_input[6]), .B(g_input[27]), .Z(n2909) );
  XNOR U3450 ( .A(n2913), .B(n2910), .Z(n2911) );
  XNOR U3451 ( .A(n2853), .B(n2859), .Z(n2899) );
  XOR U3452 ( .A(n2917), .B(n2858), .Z(n2853) );
  XNOR U3453 ( .A(n2850), .B(n2851), .Z(n2858) );
  NAND U3454 ( .A(g_input[30]), .B(e_input[3]), .Z(n2851) );
  XNOR U3455 ( .A(n2848), .B(n2918), .Z(n2850) );
  AND U3456 ( .A(e_input[2]), .B(g_input[31]), .Z(n2918) );
  XNOR U3457 ( .A(n2922), .B(n2919), .Z(n2920) );
  XNOR U3458 ( .A(n2856), .B(n2852), .Z(n2917) );
  XOR U3459 ( .A(n2855), .B(n2926), .Z(n2856) );
  ANDN U3460 ( .A(n2927), .B(n2928), .Z(n2926) );
  AND U3461 ( .A(n2932), .B(o_reg[0]), .Z(n1781) );
  XOR U3462 ( .A(n2897), .B(n2898), .Z(n2932) );
  XNOR U3463 ( .A(n2935), .B(n2916), .Z(n2897) );
  XOR U3464 ( .A(n2936), .B(n2881), .Z(n2871) );
  XNOR U3465 ( .A(n2868), .B(n2869), .Z(n2881) );
  NAND U3466 ( .A(g_input[21]), .B(e_input[11]), .Z(n2869) );
  XNOR U3467 ( .A(n2866), .B(n2937), .Z(n2868) );
  AND U3468 ( .A(e_input[10]), .B(g_input[22]), .Z(n2937) );
  XNOR U3469 ( .A(n2941), .B(n2938), .Z(n2939) );
  XNOR U3470 ( .A(n2880), .B(n2870), .Z(n2936) );
  XOR U3471 ( .A(n2875), .B(n2946), .Z(n2876) );
  AND U3472 ( .A(e_input[8]), .B(g_input[24]), .Z(n2946) );
  XNOR U3473 ( .A(n2950), .B(n2877), .Z(n2945) );
  NAND U3474 ( .A(g_input[23]), .B(e_input[9]), .Z(n2877) );
  IV U3475 ( .A(n2879), .Z(n2950) );
  XOR U3476 ( .A(n2884), .B(n2955), .Z(n2885) );
  AND U3477 ( .A(e_input[12]), .B(g_input[20]), .Z(n2955) );
  XNOR U3478 ( .A(n2959), .B(n2886), .Z(n2954) );
  NAND U3479 ( .A(g_input[19]), .B(e_input[13]), .Z(n2886) );
  IV U3480 ( .A(n2888), .Z(n2959) );
  XNOR U3481 ( .A(n2894), .B(n2895), .Z(n2890) );
  NAND U3482 ( .A(g_input[17]), .B(e_input[15]), .Z(n2895) );
  XNOR U3483 ( .A(n2892), .B(n2963), .Z(n2894) );
  AND U3484 ( .A(e_input[14]), .B(g_input[18]), .Z(n2963) );
  XNOR U3485 ( .A(n2967), .B(n2964), .Z(n2965) );
  XNOR U3486 ( .A(n2915), .B(n2896), .Z(n2935) );
  XNOR U3487 ( .A(n2968), .B(n2969), .Z(n2896) );
  XOR U3488 ( .A(n2970), .B(n2925), .Z(n2915) );
  XOR U3489 ( .A(n2902), .B(n2972), .Z(n2903) );
  AND U3490 ( .A(e_input[4]), .B(g_input[28]), .Z(n2972) );
  XNOR U3491 ( .A(n2976), .B(n2904), .Z(n2971) );
  NAND U3492 ( .A(g_input[27]), .B(e_input[5]), .Z(n2904) );
  IV U3493 ( .A(n2906), .Z(n2976) );
  XNOR U3494 ( .A(n2912), .B(n2913), .Z(n2908) );
  NAND U3495 ( .A(g_input[25]), .B(e_input[7]), .Z(n2913) );
  XNOR U3496 ( .A(n2910), .B(n2980), .Z(n2912) );
  AND U3497 ( .A(e_input[6]), .B(g_input[26]), .Z(n2980) );
  XNOR U3498 ( .A(n2984), .B(n2981), .Z(n2982) );
  XNOR U3499 ( .A(n2924), .B(n2914), .Z(n2970) );
  XOR U3500 ( .A(n2985), .B(n2986), .Z(n2914) );
  AND U3501 ( .A(n2987), .B(n2988), .Z(n2986) );
  XNOR U3502 ( .A(n2989), .B(n2990), .Z(n2988) );
  XOR U3503 ( .A(n2985), .B(n2991), .Z(n2990) );
  XOR U3504 ( .A(n2943), .B(n2992), .Z(n2987) );
  XNOR U3505 ( .A(n2985), .B(n2944), .Z(n2992) );
  XOR U3506 ( .A(n2956), .B(n2994), .Z(n2957) );
  AND U3507 ( .A(e_input[12]), .B(g_input[19]), .Z(n2994) );
  XNOR U3508 ( .A(n2998), .B(n2958), .Z(n2993) );
  NAND U3509 ( .A(g_input[18]), .B(e_input[13]), .Z(n2958) );
  IV U3510 ( .A(n2960), .Z(n2998) );
  XNOR U3511 ( .A(n2966), .B(n2967), .Z(n2962) );
  NAND U3512 ( .A(e_input[15]), .B(g_input[16]), .Z(n2967) );
  XNOR U3513 ( .A(n2964), .B(n3002), .Z(n2966) );
  AND U3514 ( .A(e_input[14]), .B(g_input[17]), .Z(n3002) );
  XNOR U3515 ( .A(n3006), .B(n3003), .Z(n3004) );
  XOR U3516 ( .A(n3007), .B(n2953), .Z(n2943) );
  XNOR U3517 ( .A(n2940), .B(n2941), .Z(n2953) );
  NAND U3518 ( .A(g_input[20]), .B(e_input[11]), .Z(n2941) );
  XNOR U3519 ( .A(n2938), .B(n3008), .Z(n2940) );
  AND U3520 ( .A(e_input[10]), .B(g_input[21]), .Z(n3008) );
  XNOR U3521 ( .A(n3012), .B(n3009), .Z(n3010) );
  XNOR U3522 ( .A(n2952), .B(n2942), .Z(n3007) );
  XOR U3523 ( .A(n2947), .B(n3017), .Z(n2948) );
  AND U3524 ( .A(e_input[8]), .B(g_input[23]), .Z(n3017) );
  XNOR U3525 ( .A(n3021), .B(n2949), .Z(n3016) );
  NAND U3526 ( .A(g_input[22]), .B(e_input[9]), .Z(n2949) );
  IV U3527 ( .A(n2951), .Z(n3021) );
  XOR U3528 ( .A(n3025), .B(n3026), .Z(n2985) );
  AND U3529 ( .A(n3027), .B(n3028), .Z(n3026) );
  XNOR U3530 ( .A(n3029), .B(n3030), .Z(n3028) );
  XOR U3531 ( .A(n3025), .B(n3031), .Z(n3030) );
  XOR U3532 ( .A(n3014), .B(n3032), .Z(n3027) );
  XNOR U3533 ( .A(n3025), .B(n3015), .Z(n3032) );
  XOR U3534 ( .A(n2995), .B(n3034), .Z(n2996) );
  AND U3535 ( .A(e_input[12]), .B(g_input[18]), .Z(n3034) );
  XNOR U3536 ( .A(n3038), .B(n2997), .Z(n3033) );
  NAND U3537 ( .A(g_input[17]), .B(e_input[13]), .Z(n2997) );
  IV U3538 ( .A(n2999), .Z(n3038) );
  XNOR U3539 ( .A(n3005), .B(n3006), .Z(n3001) );
  NAND U3540 ( .A(e_input[15]), .B(g_input[15]), .Z(n3006) );
  XNOR U3541 ( .A(n3003), .B(n3042), .Z(n3005) );
  AND U3542 ( .A(g_input[16]), .B(e_input[14]), .Z(n3042) );
  XNOR U3543 ( .A(n3046), .B(n3043), .Z(n3044) );
  XOR U3544 ( .A(n3047), .B(n3024), .Z(n3014) );
  XNOR U3545 ( .A(n3011), .B(n3012), .Z(n3024) );
  NAND U3546 ( .A(g_input[19]), .B(e_input[11]), .Z(n3012) );
  XNOR U3547 ( .A(n3009), .B(n3048), .Z(n3011) );
  AND U3548 ( .A(e_input[10]), .B(g_input[20]), .Z(n3048) );
  XNOR U3549 ( .A(n3052), .B(n3049), .Z(n3050) );
  XNOR U3550 ( .A(n3023), .B(n3013), .Z(n3047) );
  XOR U3551 ( .A(n3018), .B(n3057), .Z(n3019) );
  AND U3552 ( .A(e_input[8]), .B(g_input[22]), .Z(n3057) );
  XNOR U3553 ( .A(n3061), .B(n3020), .Z(n3056) );
  NAND U3554 ( .A(g_input[21]), .B(e_input[9]), .Z(n3020) );
  IV U3555 ( .A(n3022), .Z(n3061) );
  XOR U3556 ( .A(n3065), .B(n3066), .Z(n3025) );
  AND U3557 ( .A(n3067), .B(n3068), .Z(n3066) );
  XNOR U3558 ( .A(n3069), .B(n3070), .Z(n3068) );
  XOR U3559 ( .A(n3065), .B(n3071), .Z(n3070) );
  XOR U3560 ( .A(n3054), .B(n3072), .Z(n3067) );
  XNOR U3561 ( .A(n3065), .B(n3055), .Z(n3072) );
  XOR U3562 ( .A(n3035), .B(n3074), .Z(n3036) );
  AND U3563 ( .A(e_input[12]), .B(g_input[17]), .Z(n3074) );
  XNOR U3564 ( .A(n3078), .B(n3037), .Z(n3073) );
  NAND U3565 ( .A(e_input[13]), .B(g_input[16]), .Z(n3037) );
  IV U3566 ( .A(n3039), .Z(n3078) );
  XNOR U3567 ( .A(n3045), .B(n3046), .Z(n3041) );
  NAND U3568 ( .A(e_input[15]), .B(g_input[14]), .Z(n3046) );
  XNOR U3569 ( .A(n3043), .B(n3082), .Z(n3045) );
  AND U3570 ( .A(g_input[15]), .B(e_input[14]), .Z(n3082) );
  XNOR U3571 ( .A(n3086), .B(n3083), .Z(n3084) );
  XOR U3572 ( .A(n3087), .B(n3064), .Z(n3054) );
  XNOR U3573 ( .A(n3051), .B(n3052), .Z(n3064) );
  NAND U3574 ( .A(g_input[18]), .B(e_input[11]), .Z(n3052) );
  XNOR U3575 ( .A(n3049), .B(n3088), .Z(n3051) );
  AND U3576 ( .A(e_input[10]), .B(g_input[19]), .Z(n3088) );
  XNOR U3577 ( .A(n3092), .B(n3089), .Z(n3090) );
  XNOR U3578 ( .A(n3063), .B(n3053), .Z(n3087) );
  XOR U3579 ( .A(n3058), .B(n3097), .Z(n3059) );
  AND U3580 ( .A(e_input[8]), .B(g_input[21]), .Z(n3097) );
  XNOR U3581 ( .A(n3101), .B(n3060), .Z(n3096) );
  NAND U3582 ( .A(g_input[20]), .B(e_input[9]), .Z(n3060) );
  IV U3583 ( .A(n3062), .Z(n3101) );
  XOR U3584 ( .A(n3105), .B(n3106), .Z(n3065) );
  AND U3585 ( .A(n3107), .B(n3108), .Z(n3106) );
  XNOR U3586 ( .A(n3109), .B(n3110), .Z(n3108) );
  XOR U3587 ( .A(n3105), .B(n3111), .Z(n3110) );
  XOR U3588 ( .A(n3094), .B(n3112), .Z(n3107) );
  XNOR U3589 ( .A(n3105), .B(n3095), .Z(n3112) );
  XOR U3590 ( .A(n3075), .B(n3114), .Z(n3076) );
  AND U3591 ( .A(g_input[16]), .B(e_input[12]), .Z(n3114) );
  XNOR U3592 ( .A(n3118), .B(n3077), .Z(n3113) );
  NAND U3593 ( .A(e_input[13]), .B(g_input[15]), .Z(n3077) );
  IV U3594 ( .A(n3079), .Z(n3118) );
  XNOR U3595 ( .A(n3085), .B(n3086), .Z(n3081) );
  NAND U3596 ( .A(e_input[15]), .B(g_input[13]), .Z(n3086) );
  XNOR U3597 ( .A(n3083), .B(n3122), .Z(n3085) );
  AND U3598 ( .A(g_input[14]), .B(e_input[14]), .Z(n3122) );
  XNOR U3599 ( .A(n3126), .B(n3123), .Z(n3124) );
  XOR U3600 ( .A(n3127), .B(n3104), .Z(n3094) );
  XNOR U3601 ( .A(n3091), .B(n3092), .Z(n3104) );
  NAND U3602 ( .A(g_input[17]), .B(e_input[11]), .Z(n3092) );
  XNOR U3603 ( .A(n3089), .B(n3128), .Z(n3091) );
  AND U3604 ( .A(e_input[10]), .B(g_input[18]), .Z(n3128) );
  XNOR U3605 ( .A(n3132), .B(n3129), .Z(n3130) );
  XNOR U3606 ( .A(n3103), .B(n3093), .Z(n3127) );
  XOR U3607 ( .A(n3098), .B(n3137), .Z(n3099) );
  AND U3608 ( .A(e_input[8]), .B(g_input[20]), .Z(n3137) );
  XNOR U3609 ( .A(n3141), .B(n3100), .Z(n3136) );
  NAND U3610 ( .A(g_input[19]), .B(e_input[9]), .Z(n3100) );
  IV U3611 ( .A(n3102), .Z(n3141) );
  XOR U3612 ( .A(n3145), .B(n3146), .Z(n3105) );
  AND U3613 ( .A(n3147), .B(n3148), .Z(n3146) );
  XNOR U3614 ( .A(n3149), .B(n3150), .Z(n3148) );
  XOR U3615 ( .A(n3145), .B(n3151), .Z(n3150) );
  XOR U3616 ( .A(n3134), .B(n3152), .Z(n3147) );
  XNOR U3617 ( .A(n3145), .B(n3135), .Z(n3152) );
  XOR U3618 ( .A(n3115), .B(n3154), .Z(n3116) );
  AND U3619 ( .A(g_input[15]), .B(e_input[12]), .Z(n3154) );
  XNOR U3620 ( .A(n3158), .B(n3117), .Z(n3153) );
  NAND U3621 ( .A(e_input[13]), .B(g_input[14]), .Z(n3117) );
  IV U3622 ( .A(n3119), .Z(n3158) );
  XNOR U3623 ( .A(n3125), .B(n3126), .Z(n3121) );
  NAND U3624 ( .A(e_input[15]), .B(g_input[12]), .Z(n3126) );
  XNOR U3625 ( .A(n3123), .B(n3162), .Z(n3125) );
  AND U3626 ( .A(g_input[13]), .B(e_input[14]), .Z(n3162) );
  XNOR U3627 ( .A(n3166), .B(n3163), .Z(n3164) );
  XOR U3628 ( .A(n3167), .B(n3144), .Z(n3134) );
  XNOR U3629 ( .A(n3131), .B(n3132), .Z(n3144) );
  NAND U3630 ( .A(e_input[11]), .B(g_input[16]), .Z(n3132) );
  XNOR U3631 ( .A(n3129), .B(n3168), .Z(n3131) );
  AND U3632 ( .A(e_input[10]), .B(g_input[17]), .Z(n3168) );
  XNOR U3633 ( .A(n3172), .B(n3169), .Z(n3170) );
  XNOR U3634 ( .A(n3143), .B(n3133), .Z(n3167) );
  XOR U3635 ( .A(n3138), .B(n3177), .Z(n3139) );
  AND U3636 ( .A(e_input[8]), .B(g_input[19]), .Z(n3177) );
  XNOR U3637 ( .A(n3181), .B(n3140), .Z(n3176) );
  NAND U3638 ( .A(g_input[18]), .B(e_input[9]), .Z(n3140) );
  IV U3639 ( .A(n3142), .Z(n3181) );
  XOR U3640 ( .A(n3185), .B(n3186), .Z(n3145) );
  AND U3641 ( .A(n3187), .B(n3188), .Z(n3186) );
  XNOR U3642 ( .A(n3189), .B(n3190), .Z(n3188) );
  XOR U3643 ( .A(n3185), .B(n3191), .Z(n3190) );
  XOR U3644 ( .A(n3174), .B(n3192), .Z(n3187) );
  XNOR U3645 ( .A(n3185), .B(n3175), .Z(n3192) );
  XOR U3646 ( .A(n3155), .B(n3194), .Z(n3156) );
  AND U3647 ( .A(g_input[14]), .B(e_input[12]), .Z(n3194) );
  XNOR U3648 ( .A(n3198), .B(n3157), .Z(n3193) );
  NAND U3649 ( .A(e_input[13]), .B(g_input[13]), .Z(n3157) );
  IV U3650 ( .A(n3159), .Z(n3198) );
  XNOR U3651 ( .A(n3165), .B(n3166), .Z(n3161) );
  NAND U3652 ( .A(e_input[15]), .B(g_input[11]), .Z(n3166) );
  XNOR U3653 ( .A(n3163), .B(n3202), .Z(n3165) );
  AND U3654 ( .A(g_input[12]), .B(e_input[14]), .Z(n3202) );
  XNOR U3655 ( .A(n3206), .B(n3203), .Z(n3204) );
  XOR U3656 ( .A(n3207), .B(n3184), .Z(n3174) );
  XNOR U3657 ( .A(n3171), .B(n3172), .Z(n3184) );
  NAND U3658 ( .A(e_input[11]), .B(g_input[15]), .Z(n3172) );
  XNOR U3659 ( .A(n3169), .B(n3208), .Z(n3171) );
  AND U3660 ( .A(g_input[16]), .B(e_input[10]), .Z(n3208) );
  XNOR U3661 ( .A(n3212), .B(n3209), .Z(n3210) );
  XNOR U3662 ( .A(n3183), .B(n3173), .Z(n3207) );
  XOR U3663 ( .A(n3178), .B(n3217), .Z(n3179) );
  AND U3664 ( .A(e_input[8]), .B(g_input[18]), .Z(n3217) );
  XNOR U3665 ( .A(n3221), .B(n3180), .Z(n3216) );
  NAND U3666 ( .A(g_input[17]), .B(e_input[9]), .Z(n3180) );
  IV U3667 ( .A(n3182), .Z(n3221) );
  XOR U3668 ( .A(n3225), .B(n3226), .Z(n3185) );
  AND U3669 ( .A(n3227), .B(n3228), .Z(n3226) );
  XNOR U3670 ( .A(n3229), .B(n3230), .Z(n3228) );
  XOR U3671 ( .A(n3225), .B(n3231), .Z(n3230) );
  XOR U3672 ( .A(n3214), .B(n3232), .Z(n3227) );
  XNOR U3673 ( .A(n3225), .B(n3215), .Z(n3232) );
  XOR U3674 ( .A(n3195), .B(n3234), .Z(n3196) );
  AND U3675 ( .A(g_input[13]), .B(e_input[12]), .Z(n3234) );
  XNOR U3676 ( .A(n3238), .B(n3197), .Z(n3233) );
  NAND U3677 ( .A(e_input[13]), .B(g_input[12]), .Z(n3197) );
  IV U3678 ( .A(n3199), .Z(n3238) );
  XNOR U3679 ( .A(n3205), .B(n3206), .Z(n3201) );
  NAND U3680 ( .A(e_input[15]), .B(g_input[10]), .Z(n3206) );
  XNOR U3681 ( .A(n3203), .B(n3242), .Z(n3205) );
  AND U3682 ( .A(g_input[11]), .B(e_input[14]), .Z(n3242) );
  XNOR U3683 ( .A(n3246), .B(n3243), .Z(n3244) );
  XOR U3684 ( .A(n3247), .B(n3224), .Z(n3214) );
  XNOR U3685 ( .A(n3211), .B(n3212), .Z(n3224) );
  NAND U3686 ( .A(e_input[11]), .B(g_input[14]), .Z(n3212) );
  XNOR U3687 ( .A(n3209), .B(n3248), .Z(n3211) );
  AND U3688 ( .A(g_input[15]), .B(e_input[10]), .Z(n3248) );
  XNOR U3689 ( .A(n3252), .B(n3249), .Z(n3250) );
  XNOR U3690 ( .A(n3223), .B(n3213), .Z(n3247) );
  XOR U3691 ( .A(n3218), .B(n3257), .Z(n3219) );
  AND U3692 ( .A(e_input[8]), .B(g_input[17]), .Z(n3257) );
  XNOR U3693 ( .A(n3261), .B(n3220), .Z(n3256) );
  NAND U3694 ( .A(e_input[9]), .B(g_input[16]), .Z(n3220) );
  IV U3695 ( .A(n3222), .Z(n3261) );
  XOR U3696 ( .A(n3265), .B(n3266), .Z(n3225) );
  AND U3697 ( .A(n3267), .B(n3268), .Z(n3266) );
  XNOR U3698 ( .A(n3269), .B(n3270), .Z(n3268) );
  XOR U3699 ( .A(n3265), .B(n3271), .Z(n3270) );
  XOR U3700 ( .A(n3254), .B(n3272), .Z(n3267) );
  XNOR U3701 ( .A(n3265), .B(n3255), .Z(n3272) );
  XOR U3702 ( .A(n3235), .B(n3274), .Z(n3236) );
  AND U3703 ( .A(g_input[12]), .B(e_input[12]), .Z(n3274) );
  XNOR U3704 ( .A(n3278), .B(n3237), .Z(n3273) );
  NAND U3705 ( .A(e_input[13]), .B(g_input[11]), .Z(n3237) );
  IV U3706 ( .A(n3239), .Z(n3278) );
  XNOR U3707 ( .A(n3245), .B(n3246), .Z(n3241) );
  NAND U3708 ( .A(e_input[15]), .B(g_input[9]), .Z(n3246) );
  XNOR U3709 ( .A(n3243), .B(n3282), .Z(n3245) );
  AND U3710 ( .A(g_input[10]), .B(e_input[14]), .Z(n3282) );
  XNOR U3711 ( .A(n3286), .B(n3283), .Z(n3284) );
  XOR U3712 ( .A(n3287), .B(n3264), .Z(n3254) );
  XNOR U3713 ( .A(n3251), .B(n3252), .Z(n3264) );
  NAND U3714 ( .A(e_input[11]), .B(g_input[13]), .Z(n3252) );
  XNOR U3715 ( .A(n3249), .B(n3288), .Z(n3251) );
  AND U3716 ( .A(g_input[14]), .B(e_input[10]), .Z(n3288) );
  XNOR U3717 ( .A(n3292), .B(n3289), .Z(n3290) );
  XNOR U3718 ( .A(n3263), .B(n3253), .Z(n3287) );
  XOR U3719 ( .A(n3258), .B(n3297), .Z(n3259) );
  AND U3720 ( .A(g_input[16]), .B(e_input[8]), .Z(n3297) );
  XNOR U3721 ( .A(n3301), .B(n3260), .Z(n3296) );
  NAND U3722 ( .A(e_input[9]), .B(g_input[15]), .Z(n3260) );
  IV U3723 ( .A(n3262), .Z(n3301) );
  XOR U3724 ( .A(n3305), .B(n3306), .Z(n3265) );
  AND U3725 ( .A(n3307), .B(n3308), .Z(n3306) );
  XNOR U3726 ( .A(n3309), .B(n3310), .Z(n3308) );
  XOR U3727 ( .A(n3305), .B(n3311), .Z(n3310) );
  XOR U3728 ( .A(n3294), .B(n3312), .Z(n3307) );
  XNOR U3729 ( .A(n3305), .B(n3295), .Z(n3312) );
  XOR U3730 ( .A(n3275), .B(n3314), .Z(n3276) );
  AND U3731 ( .A(g_input[11]), .B(e_input[12]), .Z(n3314) );
  XNOR U3732 ( .A(n3318), .B(n3277), .Z(n3313) );
  NAND U3733 ( .A(e_input[13]), .B(g_input[10]), .Z(n3277) );
  IV U3734 ( .A(n3279), .Z(n3318) );
  XNOR U3735 ( .A(n3285), .B(n3286), .Z(n3281) );
  NAND U3736 ( .A(e_input[15]), .B(g_input[8]), .Z(n3286) );
  XNOR U3737 ( .A(n3283), .B(n3322), .Z(n3285) );
  AND U3738 ( .A(g_input[9]), .B(e_input[14]), .Z(n3322) );
  XNOR U3739 ( .A(n3326), .B(n3323), .Z(n3324) );
  XOR U3740 ( .A(n3327), .B(n3304), .Z(n3294) );
  XNOR U3741 ( .A(n3291), .B(n3292), .Z(n3304) );
  NAND U3742 ( .A(e_input[11]), .B(g_input[12]), .Z(n3292) );
  XNOR U3743 ( .A(n3289), .B(n3328), .Z(n3291) );
  AND U3744 ( .A(g_input[13]), .B(e_input[10]), .Z(n3328) );
  XNOR U3745 ( .A(n3332), .B(n3329), .Z(n3330) );
  XNOR U3746 ( .A(n3303), .B(n3293), .Z(n3327) );
  XOR U3747 ( .A(n3298), .B(n3337), .Z(n3299) );
  AND U3748 ( .A(g_input[15]), .B(e_input[8]), .Z(n3337) );
  XNOR U3749 ( .A(n3341), .B(n3300), .Z(n3336) );
  NAND U3750 ( .A(e_input[9]), .B(g_input[14]), .Z(n3300) );
  IV U3751 ( .A(n3302), .Z(n3341) );
  XOR U3752 ( .A(n3345), .B(n3346), .Z(n3305) );
  AND U3753 ( .A(n3347), .B(n3348), .Z(n3346) );
  XNOR U3754 ( .A(n3349), .B(n3350), .Z(n3348) );
  XOR U3755 ( .A(n3345), .B(n3351), .Z(n3350) );
  XOR U3756 ( .A(n3334), .B(n3352), .Z(n3347) );
  XNOR U3757 ( .A(n3345), .B(n3335), .Z(n3352) );
  XOR U3758 ( .A(n3315), .B(n3354), .Z(n3316) );
  AND U3759 ( .A(g_input[10]), .B(e_input[12]), .Z(n3354) );
  XNOR U3760 ( .A(n3358), .B(n3317), .Z(n3353) );
  NAND U3761 ( .A(e_input[13]), .B(g_input[9]), .Z(n3317) );
  IV U3762 ( .A(n3319), .Z(n3358) );
  XNOR U3763 ( .A(n3325), .B(n3326), .Z(n3321) );
  NAND U3764 ( .A(e_input[15]), .B(g_input[7]), .Z(n3326) );
  XNOR U3765 ( .A(n3323), .B(n3362), .Z(n3325) );
  AND U3766 ( .A(g_input[8]), .B(e_input[14]), .Z(n3362) );
  XNOR U3767 ( .A(n3366), .B(n3363), .Z(n3364) );
  XOR U3768 ( .A(n3367), .B(n3344), .Z(n3334) );
  XNOR U3769 ( .A(n3331), .B(n3332), .Z(n3344) );
  NAND U3770 ( .A(e_input[11]), .B(g_input[11]), .Z(n3332) );
  XNOR U3771 ( .A(n3329), .B(n3368), .Z(n3331) );
  AND U3772 ( .A(g_input[12]), .B(e_input[10]), .Z(n3368) );
  XNOR U3773 ( .A(n3372), .B(n3369), .Z(n3370) );
  XNOR U3774 ( .A(n3343), .B(n3333), .Z(n3367) );
  XOR U3775 ( .A(n3338), .B(n3377), .Z(n3339) );
  AND U3776 ( .A(g_input[14]), .B(e_input[8]), .Z(n3377) );
  XNOR U3777 ( .A(n3381), .B(n3340), .Z(n3376) );
  NAND U3778 ( .A(e_input[9]), .B(g_input[13]), .Z(n3340) );
  IV U3779 ( .A(n3342), .Z(n3381) );
  XOR U3780 ( .A(n3385), .B(n3386), .Z(n3345) );
  AND U3781 ( .A(n3387), .B(n3388), .Z(n3386) );
  XNOR U3782 ( .A(n3389), .B(n3390), .Z(n3388) );
  XOR U3783 ( .A(n3385), .B(n3391), .Z(n3390) );
  XOR U3784 ( .A(n3374), .B(n3392), .Z(n3387) );
  XNOR U3785 ( .A(n3385), .B(n3375), .Z(n3392) );
  XOR U3786 ( .A(n3355), .B(n3394), .Z(n3356) );
  AND U3787 ( .A(g_input[9]), .B(e_input[12]), .Z(n3394) );
  XNOR U3788 ( .A(n3398), .B(n3357), .Z(n3393) );
  NAND U3789 ( .A(e_input[13]), .B(g_input[8]), .Z(n3357) );
  IV U3790 ( .A(n3359), .Z(n3398) );
  XNOR U3791 ( .A(n3365), .B(n3366), .Z(n3361) );
  NAND U3792 ( .A(e_input[15]), .B(g_input[6]), .Z(n3366) );
  XNOR U3793 ( .A(n3363), .B(n3402), .Z(n3365) );
  AND U3794 ( .A(g_input[7]), .B(e_input[14]), .Z(n3402) );
  XNOR U3795 ( .A(n3406), .B(n3403), .Z(n3404) );
  XOR U3796 ( .A(n3407), .B(n3384), .Z(n3374) );
  XNOR U3797 ( .A(n3371), .B(n3372), .Z(n3384) );
  NAND U3798 ( .A(e_input[11]), .B(g_input[10]), .Z(n3372) );
  XNOR U3799 ( .A(n3369), .B(n3408), .Z(n3371) );
  AND U3800 ( .A(g_input[11]), .B(e_input[10]), .Z(n3408) );
  XNOR U3801 ( .A(n3412), .B(n3409), .Z(n3410) );
  XNOR U3802 ( .A(n3383), .B(n3373), .Z(n3407) );
  XOR U3803 ( .A(n3378), .B(n3417), .Z(n3379) );
  AND U3804 ( .A(g_input[13]), .B(e_input[8]), .Z(n3417) );
  XNOR U3805 ( .A(n3421), .B(n3380), .Z(n3416) );
  NAND U3806 ( .A(e_input[9]), .B(g_input[12]), .Z(n3380) );
  IV U3807 ( .A(n3382), .Z(n3421) );
  XOR U3808 ( .A(n3425), .B(n3426), .Z(n3385) );
  AND U3809 ( .A(n3427), .B(n3428), .Z(n3426) );
  XNOR U3810 ( .A(n3429), .B(n3430), .Z(n3428) );
  XOR U3811 ( .A(n3425), .B(n3431), .Z(n3430) );
  XOR U3812 ( .A(n3414), .B(n3432), .Z(n3427) );
  XNOR U3813 ( .A(n3425), .B(n3415), .Z(n3432) );
  XOR U3814 ( .A(n3395), .B(n3434), .Z(n3396) );
  AND U3815 ( .A(g_input[8]), .B(e_input[12]), .Z(n3434) );
  XNOR U3816 ( .A(n3438), .B(n3397), .Z(n3433) );
  NAND U3817 ( .A(e_input[13]), .B(g_input[7]), .Z(n3397) );
  IV U3818 ( .A(n3399), .Z(n3438) );
  XNOR U3819 ( .A(n3405), .B(n3406), .Z(n3401) );
  NAND U3820 ( .A(e_input[15]), .B(g_input[5]), .Z(n3406) );
  XNOR U3821 ( .A(n3403), .B(n3442), .Z(n3405) );
  AND U3822 ( .A(g_input[6]), .B(e_input[14]), .Z(n3442) );
  XNOR U3823 ( .A(n3446), .B(n3443), .Z(n3444) );
  XOR U3824 ( .A(n3447), .B(n3424), .Z(n3414) );
  XNOR U3825 ( .A(n3411), .B(n3412), .Z(n3424) );
  NAND U3826 ( .A(e_input[11]), .B(g_input[9]), .Z(n3412) );
  XNOR U3827 ( .A(n3409), .B(n3448), .Z(n3411) );
  AND U3828 ( .A(g_input[10]), .B(e_input[10]), .Z(n3448) );
  XNOR U3829 ( .A(n3452), .B(n3449), .Z(n3450) );
  XNOR U3830 ( .A(n3423), .B(n3413), .Z(n3447) );
  XOR U3831 ( .A(n3418), .B(n3457), .Z(n3419) );
  AND U3832 ( .A(g_input[12]), .B(e_input[8]), .Z(n3457) );
  XNOR U3833 ( .A(n3461), .B(n3420), .Z(n3456) );
  NAND U3834 ( .A(e_input[9]), .B(g_input[11]), .Z(n3420) );
  IV U3835 ( .A(n3422), .Z(n3461) );
  XOR U3836 ( .A(n3465), .B(n3466), .Z(n3425) );
  AND U3837 ( .A(n3467), .B(n3468), .Z(n3466) );
  XNOR U3838 ( .A(n3469), .B(n3470), .Z(n3468) );
  XOR U3839 ( .A(n3465), .B(n3471), .Z(n3470) );
  XOR U3840 ( .A(n3454), .B(n3472), .Z(n3467) );
  XNOR U3841 ( .A(n3465), .B(n3455), .Z(n3472) );
  XOR U3842 ( .A(n3435), .B(n3474), .Z(n3436) );
  AND U3843 ( .A(g_input[7]), .B(e_input[12]), .Z(n3474) );
  XNOR U3844 ( .A(n3478), .B(n3437), .Z(n3473) );
  NAND U3845 ( .A(e_input[13]), .B(g_input[6]), .Z(n3437) );
  IV U3846 ( .A(n3439), .Z(n3478) );
  XNOR U3847 ( .A(n3445), .B(n3446), .Z(n3441) );
  NAND U3848 ( .A(e_input[15]), .B(g_input[4]), .Z(n3446) );
  XNOR U3849 ( .A(n3443), .B(n3482), .Z(n3445) );
  AND U3850 ( .A(g_input[5]), .B(e_input[14]), .Z(n3482) );
  XNOR U3851 ( .A(n3486), .B(n3483), .Z(n3484) );
  XOR U3852 ( .A(n3487), .B(n3464), .Z(n3454) );
  XNOR U3853 ( .A(n3451), .B(n3452), .Z(n3464) );
  NAND U3854 ( .A(e_input[11]), .B(g_input[8]), .Z(n3452) );
  XNOR U3855 ( .A(n3449), .B(n3488), .Z(n3451) );
  AND U3856 ( .A(g_input[9]), .B(e_input[10]), .Z(n3488) );
  XNOR U3857 ( .A(n3492), .B(n3489), .Z(n3490) );
  XNOR U3858 ( .A(n3463), .B(n3453), .Z(n3487) );
  XOR U3859 ( .A(n3458), .B(n3497), .Z(n3459) );
  AND U3860 ( .A(g_input[11]), .B(e_input[8]), .Z(n3497) );
  XNOR U3861 ( .A(n3501), .B(n3460), .Z(n3496) );
  NAND U3862 ( .A(e_input[9]), .B(g_input[10]), .Z(n3460) );
  IV U3863 ( .A(n3462), .Z(n3501) );
  XOR U3864 ( .A(n3505), .B(n3506), .Z(n3465) );
  AND U3865 ( .A(n3507), .B(n3508), .Z(n3506) );
  XNOR U3866 ( .A(n3509), .B(n3510), .Z(n3508) );
  XOR U3867 ( .A(n3505), .B(n3511), .Z(n3510) );
  XOR U3868 ( .A(n3494), .B(n3512), .Z(n3507) );
  XNOR U3869 ( .A(n3505), .B(n3495), .Z(n3512) );
  XOR U3870 ( .A(n3475), .B(n3514), .Z(n3476) );
  AND U3871 ( .A(g_input[6]), .B(e_input[12]), .Z(n3514) );
  XNOR U3872 ( .A(n3518), .B(n3477), .Z(n3513) );
  NAND U3873 ( .A(e_input[13]), .B(g_input[5]), .Z(n3477) );
  IV U3874 ( .A(n3479), .Z(n3518) );
  XNOR U3875 ( .A(n3485), .B(n3486), .Z(n3481) );
  NAND U3876 ( .A(e_input[15]), .B(g_input[3]), .Z(n3486) );
  XNOR U3877 ( .A(n3483), .B(n3522), .Z(n3485) );
  AND U3878 ( .A(g_input[4]), .B(e_input[14]), .Z(n3522) );
  XNOR U3879 ( .A(n3526), .B(n3523), .Z(n3524) );
  XOR U3880 ( .A(n3527), .B(n3504), .Z(n3494) );
  XNOR U3881 ( .A(n3491), .B(n3492), .Z(n3504) );
  NAND U3882 ( .A(e_input[11]), .B(g_input[7]), .Z(n3492) );
  XNOR U3883 ( .A(n3489), .B(n3528), .Z(n3491) );
  AND U3884 ( .A(g_input[8]), .B(e_input[10]), .Z(n3528) );
  XNOR U3885 ( .A(n3532), .B(n3529), .Z(n3530) );
  XNOR U3886 ( .A(n3503), .B(n3493), .Z(n3527) );
  XOR U3887 ( .A(n3498), .B(n3537), .Z(n3499) );
  AND U3888 ( .A(g_input[10]), .B(e_input[8]), .Z(n3537) );
  XNOR U3889 ( .A(n3541), .B(n3500), .Z(n3536) );
  NAND U3890 ( .A(e_input[9]), .B(g_input[9]), .Z(n3500) );
  IV U3891 ( .A(n3502), .Z(n3541) );
  XOR U3892 ( .A(n3545), .B(n3546), .Z(n3505) );
  AND U3893 ( .A(n3547), .B(n3548), .Z(n3546) );
  XNOR U3894 ( .A(n3549), .B(n3550), .Z(n3548) );
  XOR U3895 ( .A(n3545), .B(n3551), .Z(n3550) );
  XOR U3896 ( .A(n3534), .B(n3552), .Z(n3547) );
  XNOR U3897 ( .A(n3545), .B(n3535), .Z(n3552) );
  XOR U3898 ( .A(n3515), .B(n3554), .Z(n3516) );
  AND U3899 ( .A(g_input[5]), .B(e_input[12]), .Z(n3554) );
  XNOR U3900 ( .A(n3558), .B(n3517), .Z(n3553) );
  NAND U3901 ( .A(e_input[13]), .B(g_input[4]), .Z(n3517) );
  IV U3902 ( .A(n3519), .Z(n3558) );
  XNOR U3903 ( .A(n3525), .B(n3526), .Z(n3521) );
  NAND U3904 ( .A(e_input[15]), .B(g_input[2]), .Z(n3526) );
  XNOR U3905 ( .A(n3523), .B(n3562), .Z(n3525) );
  AND U3906 ( .A(g_input[3]), .B(e_input[14]), .Z(n3562) );
  XNOR U3907 ( .A(n3566), .B(n3563), .Z(n3564) );
  XOR U3908 ( .A(n3567), .B(n3544), .Z(n3534) );
  XNOR U3909 ( .A(n3531), .B(n3532), .Z(n3544) );
  NAND U3910 ( .A(e_input[11]), .B(g_input[6]), .Z(n3532) );
  XNOR U3911 ( .A(n3529), .B(n3568), .Z(n3531) );
  AND U3912 ( .A(g_input[7]), .B(e_input[10]), .Z(n3568) );
  XNOR U3913 ( .A(n3572), .B(n3569), .Z(n3570) );
  XNOR U3914 ( .A(n3543), .B(n3533), .Z(n3567) );
  XOR U3915 ( .A(n3538), .B(n3577), .Z(n3539) );
  AND U3916 ( .A(g_input[9]), .B(e_input[8]), .Z(n3577) );
  XNOR U3917 ( .A(n3581), .B(n3540), .Z(n3576) );
  NAND U3918 ( .A(e_input[9]), .B(g_input[8]), .Z(n3540) );
  IV U3919 ( .A(n3542), .Z(n3581) );
  XOR U3920 ( .A(n3586), .B(n3584), .Z(n3574) );
  XNOR U3921 ( .A(n3571), .B(n3572), .Z(n3584) );
  NAND U3922 ( .A(e_input[11]), .B(g_input[5]), .Z(n3572) );
  XNOR U3923 ( .A(n3569), .B(n3587), .Z(n3571) );
  AND U3924 ( .A(g_input[6]), .B(e_input[10]), .Z(n3587) );
  XNOR U3925 ( .A(n3591), .B(n3588), .Z(n3590) );
  XNOR U3926 ( .A(n3583), .B(n3573), .Z(n3586) );
  XOR U3927 ( .A(n3592), .B(n3593), .Z(n3573) );
  XOR U3928 ( .A(n3578), .B(n3595), .Z(n3579) );
  AND U3929 ( .A(g_input[8]), .B(e_input[8]), .Z(n3595) );
  XNOR U3930 ( .A(n3599), .B(n3596), .Z(n3598) );
  XNOR U3931 ( .A(n3600), .B(n3580), .Z(n3594) );
  NAND U3932 ( .A(e_input[9]), .B(g_input[7]), .Z(n3580) );
  IV U3933 ( .A(n3582), .Z(n3600) );
  XOR U3934 ( .A(n3601), .B(n3602), .Z(n3582) );
  AND U3935 ( .A(n3603), .B(n3604), .Z(n3602) );
  XOR U3936 ( .A(n3597), .B(n3605), .Z(n3604) );
  XNOR U3937 ( .A(n3599), .B(n3601), .Z(n3605) );
  NAND U3938 ( .A(e_input[9]), .B(g_input[6]), .Z(n3599) );
  XOR U3939 ( .A(n3596), .B(n3606), .Z(n3597) );
  AND U3940 ( .A(g_input[7]), .B(e_input[8]), .Z(n3606) );
  XNOR U3941 ( .A(n3610), .B(n3607), .Z(n3609) );
  XOR U3942 ( .A(n3589), .B(n3611), .Z(n3603) );
  XNOR U3943 ( .A(n3591), .B(n3601), .Z(n3611) );
  NAND U3944 ( .A(e_input[11]), .B(g_input[4]), .Z(n3591) );
  XOR U3945 ( .A(n3588), .B(n3612), .Z(n3589) );
  AND U3946 ( .A(g_input[5]), .B(e_input[10]), .Z(n3612) );
  XNOR U3947 ( .A(n3616), .B(n3613), .Z(n3615) );
  XOR U3948 ( .A(n3617), .B(n3618), .Z(n3601) );
  AND U3949 ( .A(n3619), .B(n3620), .Z(n3618) );
  XOR U3950 ( .A(n3608), .B(n3621), .Z(n3620) );
  XNOR U3951 ( .A(n3610), .B(n3617), .Z(n3621) );
  NAND U3952 ( .A(e_input[9]), .B(g_input[5]), .Z(n3610) );
  XOR U3953 ( .A(n3607), .B(n3622), .Z(n3608) );
  AND U3954 ( .A(g_input[6]), .B(e_input[8]), .Z(n3622) );
  XNOR U3955 ( .A(n3626), .B(n3623), .Z(n3625) );
  XOR U3956 ( .A(n3614), .B(n3627), .Z(n3619) );
  XNOR U3957 ( .A(n3616), .B(n3617), .Z(n3627) );
  NAND U3958 ( .A(e_input[11]), .B(g_input[3]), .Z(n3616) );
  XOR U3959 ( .A(n3613), .B(n3628), .Z(n3614) );
  AND U3960 ( .A(g_input[4]), .B(e_input[10]), .Z(n3628) );
  XNOR U3961 ( .A(n3632), .B(n3629), .Z(n3631) );
  XOR U3962 ( .A(n3633), .B(n3634), .Z(n3617) );
  AND U3963 ( .A(n3635), .B(n3636), .Z(n3634) );
  XOR U3964 ( .A(n3624), .B(n3637), .Z(n3636) );
  XNOR U3965 ( .A(n3626), .B(n3633), .Z(n3637) );
  NAND U3966 ( .A(e_input[9]), .B(g_input[4]), .Z(n3626) );
  XOR U3967 ( .A(n3623), .B(n3638), .Z(n3624) );
  AND U3968 ( .A(g_input[5]), .B(e_input[8]), .Z(n3638) );
  XOR U3969 ( .A(n3630), .B(n3642), .Z(n3635) );
  XNOR U3970 ( .A(n3632), .B(n3633), .Z(n3642) );
  NAND U3971 ( .A(e_input[11]), .B(g_input[2]), .Z(n3632) );
  XOR U3972 ( .A(n3629), .B(n3643), .Z(n3630) );
  AND U3973 ( .A(g_input[3]), .B(e_input[10]), .Z(n3643) );
  XNOR U3974 ( .A(n3647), .B(n3644), .Z(n3645) );
  NAND U3975 ( .A(e_input[11]), .B(g_input[1]), .Z(n3647) );
  XOR U3976 ( .A(n3644), .B(n3649), .Z(n3646) );
  AND U3977 ( .A(g_input[2]), .B(e_input[10]), .Z(n3649) );
  AND U3978 ( .A(n3650), .B(g_input[0]), .Z(n3644) );
  NANDN U3979 ( .B(e_input[11]), .A(n3651), .Z(n3650) );
  NAND U3980 ( .A(g_input[1]), .B(e_input[10]), .Z(n3651) );
  XOR U3981 ( .A(n3639), .B(n3653), .Z(n3640) );
  AND U3982 ( .A(g_input[4]), .B(e_input[8]), .Z(n3653) );
  XOR U3983 ( .A(n3656), .B(n3654), .Z(n3655) );
  AND U3984 ( .A(g_input[3]), .B(e_input[8]), .Z(n3656) );
  AND U3985 ( .A(g_input[2]), .B(e_input[9]), .Z(n3657) );
  XNOR U3986 ( .A(n3661), .B(n3658), .Z(n3659) );
  XNOR U3987 ( .A(n3662), .B(n3641), .Z(n3652) );
  NAND U3988 ( .A(e_input[9]), .B(g_input[3]), .Z(n3641) );
  IV U3989 ( .A(n3648), .Z(n3662) );
  NAND U3990 ( .A(e_input[9]), .B(g_input[1]), .Z(n3661) );
  XOR U3991 ( .A(n3658), .B(n3663), .Z(n3660) );
  AND U3992 ( .A(g_input[2]), .B(e_input[8]), .Z(n3663) );
  AND U3993 ( .A(n3664), .B(g_input[0]), .Z(n3658) );
  NANDN U3994 ( .B(e_input[9]), .A(n3665), .Z(n3664) );
  NAND U3995 ( .A(g_input[1]), .B(e_input[8]), .Z(n3665) );
  XOR U3996 ( .A(n3555), .B(n3667), .Z(n3556) );
  AND U3997 ( .A(g_input[4]), .B(e_input[12]), .Z(n3667) );
  XOR U3998 ( .A(n3670), .B(n3668), .Z(n3669) );
  AND U3999 ( .A(g_input[3]), .B(e_input[12]), .Z(n3670) );
  AND U4000 ( .A(g_input[2]), .B(e_input[13]), .Z(n3671) );
  XNOR U4001 ( .A(n3675), .B(n3672), .Z(n3673) );
  XNOR U4002 ( .A(n3676), .B(n3557), .Z(n3666) );
  NAND U4003 ( .A(e_input[13]), .B(g_input[3]), .Z(n3557) );
  IV U4004 ( .A(n3559), .Z(n3676) );
  NAND U4005 ( .A(e_input[13]), .B(g_input[1]), .Z(n3675) );
  XOR U4006 ( .A(n3672), .B(n3677), .Z(n3674) );
  AND U4007 ( .A(g_input[2]), .B(e_input[12]), .Z(n3677) );
  AND U4008 ( .A(n3678), .B(g_input[0]), .Z(n3672) );
  NANDN U4009 ( .B(e_input[13]), .A(n3679), .Z(n3678) );
  NAND U4010 ( .A(g_input[1]), .B(e_input[12]), .Z(n3679) );
  XNOR U4011 ( .A(n3565), .B(n3566), .Z(n3561) );
  NAND U4012 ( .A(e_input[15]), .B(g_input[1]), .Z(n3566) );
  XNOR U4013 ( .A(n3563), .B(n3680), .Z(n3565) );
  AND U4014 ( .A(g_input[2]), .B(e_input[14]), .Z(n3680) );
  AND U4015 ( .A(n3681), .B(g_input[0]), .Z(n3563) );
  NANDN U4016 ( .B(e_input[15]), .A(n3682), .Z(n3681) );
  NAND U4017 ( .A(g_input[1]), .B(e_input[14]), .Z(n3682) );
  XOR U4018 ( .A(n3683), .B(n3684), .Z(n2969) );
  XNOR U4019 ( .A(n3685), .B(n3585), .Z(n3683) );
  XOR U4020 ( .A(n3686), .B(n3687), .Z(n3585) );
  XOR U4021 ( .A(n3688), .B(n2931), .Z(n2924) );
  XNOR U4022 ( .A(n2921), .B(n2922), .Z(n2931) );
  NAND U4023 ( .A(g_input[29]), .B(e_input[3]), .Z(n2922) );
  XNOR U4024 ( .A(n2919), .B(n3689), .Z(n2921) );
  AND U4025 ( .A(e_input[2]), .B(g_input[30]), .Z(n3689) );
  XNOR U4026 ( .A(n3693), .B(n3690), .Z(n3691) );
  XNOR U4027 ( .A(n2930), .B(n2923), .Z(n3688) );
  XOR U4028 ( .A(n2973), .B(n3696), .Z(n2974) );
  AND U4029 ( .A(e_input[4]), .B(g_input[27]), .Z(n3696) );
  XNOR U4030 ( .A(n3700), .B(n2975), .Z(n3695) );
  NAND U4031 ( .A(g_input[26]), .B(e_input[5]), .Z(n2975) );
  IV U4032 ( .A(n2977), .Z(n3700) );
  XNOR U4033 ( .A(n2983), .B(n2984), .Z(n2979) );
  NAND U4034 ( .A(g_input[24]), .B(e_input[7]), .Z(n2984) );
  XNOR U4035 ( .A(n2981), .B(n3704), .Z(n2983) );
  AND U4036 ( .A(e_input[6]), .B(g_input[25]), .Z(n3704) );
  XNOR U4037 ( .A(n3708), .B(n3705), .Z(n3706) );
  XOR U4038 ( .A(n3709), .B(n3710), .Z(n2991) );
  XNOR U4039 ( .A(n3711), .B(n3694), .Z(n3709) );
  XOR U4040 ( .A(n3697), .B(n3714), .Z(n3698) );
  AND U4041 ( .A(e_input[4]), .B(g_input[26]), .Z(n3714) );
  XNOR U4042 ( .A(n3718), .B(n3699), .Z(n3713) );
  NAND U4043 ( .A(g_input[25]), .B(e_input[5]), .Z(n3699) );
  IV U4044 ( .A(n3701), .Z(n3718) );
  XNOR U4045 ( .A(n3707), .B(n3708), .Z(n3703) );
  NAND U4046 ( .A(g_input[23]), .B(e_input[7]), .Z(n3708) );
  XNOR U4047 ( .A(n3705), .B(n3722), .Z(n3707) );
  AND U4048 ( .A(e_input[6]), .B(g_input[24]), .Z(n3722) );
  XNOR U4049 ( .A(n3726), .B(n3723), .Z(n3724) );
  XOR U4050 ( .A(n3727), .B(n3728), .Z(n3031) );
  XNOR U4051 ( .A(n3729), .B(n3712), .Z(n3727) );
  XOR U4052 ( .A(n3715), .B(n3732), .Z(n3716) );
  AND U4053 ( .A(e_input[4]), .B(g_input[25]), .Z(n3732) );
  XNOR U4054 ( .A(n3736), .B(n3717), .Z(n3731) );
  NAND U4055 ( .A(g_input[24]), .B(e_input[5]), .Z(n3717) );
  IV U4056 ( .A(n3719), .Z(n3736) );
  XNOR U4057 ( .A(n3725), .B(n3726), .Z(n3721) );
  NAND U4058 ( .A(g_input[22]), .B(e_input[7]), .Z(n3726) );
  XNOR U4059 ( .A(n3723), .B(n3740), .Z(n3725) );
  AND U4060 ( .A(e_input[6]), .B(g_input[23]), .Z(n3740) );
  XNOR U4061 ( .A(n3744), .B(n3741), .Z(n3742) );
  XOR U4062 ( .A(n3745), .B(n3746), .Z(n3071) );
  XNOR U4063 ( .A(n3747), .B(n3730), .Z(n3745) );
  XOR U4064 ( .A(n3733), .B(n3750), .Z(n3734) );
  AND U4065 ( .A(e_input[4]), .B(g_input[24]), .Z(n3750) );
  XNOR U4066 ( .A(n3754), .B(n3735), .Z(n3749) );
  NAND U4067 ( .A(g_input[23]), .B(e_input[5]), .Z(n3735) );
  IV U4068 ( .A(n3737), .Z(n3754) );
  XNOR U4069 ( .A(n3743), .B(n3744), .Z(n3739) );
  NAND U4070 ( .A(g_input[21]), .B(e_input[7]), .Z(n3744) );
  XNOR U4071 ( .A(n3741), .B(n3758), .Z(n3743) );
  AND U4072 ( .A(e_input[6]), .B(g_input[22]), .Z(n3758) );
  XNOR U4073 ( .A(n3762), .B(n3759), .Z(n3760) );
  XOR U4074 ( .A(n3763), .B(n3764), .Z(n3111) );
  XNOR U4075 ( .A(n3765), .B(n3748), .Z(n3763) );
  XOR U4076 ( .A(n3751), .B(n3768), .Z(n3752) );
  AND U4077 ( .A(e_input[4]), .B(g_input[23]), .Z(n3768) );
  XNOR U4078 ( .A(n3772), .B(n3753), .Z(n3767) );
  NAND U4079 ( .A(g_input[22]), .B(e_input[5]), .Z(n3753) );
  IV U4080 ( .A(n3755), .Z(n3772) );
  XNOR U4081 ( .A(n3761), .B(n3762), .Z(n3757) );
  NAND U4082 ( .A(g_input[20]), .B(e_input[7]), .Z(n3762) );
  XNOR U4083 ( .A(n3759), .B(n3776), .Z(n3761) );
  AND U4084 ( .A(e_input[6]), .B(g_input[21]), .Z(n3776) );
  XNOR U4085 ( .A(n3780), .B(n3777), .Z(n3778) );
  XOR U4086 ( .A(n3781), .B(n3782), .Z(n3151) );
  XNOR U4087 ( .A(n3783), .B(n3766), .Z(n3781) );
  XOR U4088 ( .A(n3769), .B(n3786), .Z(n3770) );
  AND U4089 ( .A(e_input[4]), .B(g_input[22]), .Z(n3786) );
  XNOR U4090 ( .A(n3790), .B(n3771), .Z(n3785) );
  NAND U4091 ( .A(g_input[21]), .B(e_input[5]), .Z(n3771) );
  IV U4092 ( .A(n3773), .Z(n3790) );
  XNOR U4093 ( .A(n3779), .B(n3780), .Z(n3775) );
  NAND U4094 ( .A(g_input[19]), .B(e_input[7]), .Z(n3780) );
  XNOR U4095 ( .A(n3777), .B(n3794), .Z(n3779) );
  AND U4096 ( .A(e_input[6]), .B(g_input[20]), .Z(n3794) );
  XNOR U4097 ( .A(n3798), .B(n3795), .Z(n3796) );
  XOR U4098 ( .A(n3799), .B(n3800), .Z(n3191) );
  XNOR U4099 ( .A(n3801), .B(n3784), .Z(n3799) );
  XOR U4100 ( .A(n3787), .B(n3804), .Z(n3788) );
  AND U4101 ( .A(e_input[4]), .B(g_input[21]), .Z(n3804) );
  XNOR U4102 ( .A(n3808), .B(n3789), .Z(n3803) );
  NAND U4103 ( .A(g_input[20]), .B(e_input[5]), .Z(n3789) );
  IV U4104 ( .A(n3791), .Z(n3808) );
  XNOR U4105 ( .A(n3797), .B(n3798), .Z(n3793) );
  NAND U4106 ( .A(g_input[18]), .B(e_input[7]), .Z(n3798) );
  XNOR U4107 ( .A(n3795), .B(n3812), .Z(n3797) );
  AND U4108 ( .A(e_input[6]), .B(g_input[19]), .Z(n3812) );
  XNOR U4109 ( .A(n3816), .B(n3813), .Z(n3814) );
  XOR U4110 ( .A(n3817), .B(n3818), .Z(n3231) );
  XNOR U4111 ( .A(n3819), .B(n3802), .Z(n3817) );
  XOR U4112 ( .A(n3805), .B(n3822), .Z(n3806) );
  AND U4113 ( .A(e_input[4]), .B(g_input[20]), .Z(n3822) );
  XNOR U4114 ( .A(n3826), .B(n3807), .Z(n3821) );
  NAND U4115 ( .A(g_input[19]), .B(e_input[5]), .Z(n3807) );
  IV U4116 ( .A(n3809), .Z(n3826) );
  XNOR U4117 ( .A(n3815), .B(n3816), .Z(n3811) );
  NAND U4118 ( .A(g_input[17]), .B(e_input[7]), .Z(n3816) );
  XNOR U4119 ( .A(n3813), .B(n3830), .Z(n3815) );
  AND U4120 ( .A(e_input[6]), .B(g_input[18]), .Z(n3830) );
  XNOR U4121 ( .A(n3834), .B(n3831), .Z(n3832) );
  XOR U4122 ( .A(n3835), .B(n3836), .Z(n3271) );
  XNOR U4123 ( .A(n3837), .B(n3820), .Z(n3835) );
  XOR U4124 ( .A(n3823), .B(n3840), .Z(n3824) );
  AND U4125 ( .A(e_input[4]), .B(g_input[19]), .Z(n3840) );
  XNOR U4126 ( .A(n3844), .B(n3825), .Z(n3839) );
  NAND U4127 ( .A(g_input[18]), .B(e_input[5]), .Z(n3825) );
  IV U4128 ( .A(n3827), .Z(n3844) );
  XNOR U4129 ( .A(n3833), .B(n3834), .Z(n3829) );
  NAND U4130 ( .A(g_input[16]), .B(e_input[7]), .Z(n3834) );
  XNOR U4131 ( .A(n3831), .B(n3848), .Z(n3833) );
  AND U4132 ( .A(e_input[6]), .B(g_input[17]), .Z(n3848) );
  XNOR U4133 ( .A(n3852), .B(n3849), .Z(n3850) );
  XOR U4134 ( .A(n3853), .B(n3854), .Z(n3311) );
  XNOR U4135 ( .A(n3855), .B(n3838), .Z(n3853) );
  XOR U4136 ( .A(n3841), .B(n3858), .Z(n3842) );
  AND U4137 ( .A(e_input[4]), .B(g_input[18]), .Z(n3858) );
  XNOR U4138 ( .A(n3862), .B(n3843), .Z(n3857) );
  NAND U4139 ( .A(g_input[17]), .B(e_input[5]), .Z(n3843) );
  IV U4140 ( .A(n3845), .Z(n3862) );
  XNOR U4141 ( .A(n3851), .B(n3852), .Z(n3847) );
  NAND U4142 ( .A(g_input[15]), .B(e_input[7]), .Z(n3852) );
  XNOR U4143 ( .A(n3849), .B(n3866), .Z(n3851) );
  AND U4144 ( .A(e_input[6]), .B(g_input[16]), .Z(n3866) );
  XNOR U4145 ( .A(n3870), .B(n3867), .Z(n3868) );
  XOR U4146 ( .A(n3871), .B(n3872), .Z(n3351) );
  XNOR U4147 ( .A(n3873), .B(n3856), .Z(n3871) );
  XOR U4148 ( .A(n3859), .B(n3876), .Z(n3860) );
  AND U4149 ( .A(e_input[4]), .B(g_input[17]), .Z(n3876) );
  XNOR U4150 ( .A(n3880), .B(n3861), .Z(n3875) );
  NAND U4151 ( .A(g_input[16]), .B(e_input[5]), .Z(n3861) );
  IV U4152 ( .A(n3863), .Z(n3880) );
  XNOR U4153 ( .A(n3869), .B(n3870), .Z(n3865) );
  NAND U4154 ( .A(g_input[14]), .B(e_input[7]), .Z(n3870) );
  XNOR U4155 ( .A(n3867), .B(n3884), .Z(n3869) );
  AND U4156 ( .A(e_input[6]), .B(g_input[15]), .Z(n3884) );
  XNOR U4157 ( .A(n3888), .B(n3885), .Z(n3886) );
  XOR U4158 ( .A(n3889), .B(n3890), .Z(n3391) );
  XNOR U4159 ( .A(n3891), .B(n3874), .Z(n3889) );
  XOR U4160 ( .A(n3877), .B(n3894), .Z(n3878) );
  AND U4161 ( .A(e_input[4]), .B(g_input[16]), .Z(n3894) );
  XNOR U4162 ( .A(n3898), .B(n3879), .Z(n3893) );
  NAND U4163 ( .A(g_input[15]), .B(e_input[5]), .Z(n3879) );
  IV U4164 ( .A(n3881), .Z(n3898) );
  XNOR U4165 ( .A(n3887), .B(n3888), .Z(n3883) );
  NAND U4166 ( .A(g_input[13]), .B(e_input[7]), .Z(n3888) );
  XNOR U4167 ( .A(n3885), .B(n3902), .Z(n3887) );
  AND U4168 ( .A(e_input[6]), .B(g_input[14]), .Z(n3902) );
  XNOR U4169 ( .A(n3906), .B(n3903), .Z(n3904) );
  XOR U4170 ( .A(n3907), .B(n3908), .Z(n3431) );
  XNOR U4171 ( .A(n3909), .B(n3892), .Z(n3907) );
  XOR U4172 ( .A(n3895), .B(n3912), .Z(n3896) );
  AND U4173 ( .A(e_input[4]), .B(g_input[15]), .Z(n3912) );
  XNOR U4174 ( .A(n3916), .B(n3897), .Z(n3911) );
  NAND U4175 ( .A(g_input[14]), .B(e_input[5]), .Z(n3897) );
  IV U4176 ( .A(n3899), .Z(n3916) );
  XNOR U4177 ( .A(n3905), .B(n3906), .Z(n3901) );
  NAND U4178 ( .A(g_input[12]), .B(e_input[7]), .Z(n3906) );
  XNOR U4179 ( .A(n3903), .B(n3920), .Z(n3905) );
  AND U4180 ( .A(e_input[6]), .B(g_input[13]), .Z(n3920) );
  XNOR U4181 ( .A(n3924), .B(n3921), .Z(n3922) );
  XOR U4182 ( .A(n3925), .B(n3926), .Z(n3471) );
  XNOR U4183 ( .A(n3927), .B(n3910), .Z(n3925) );
  XOR U4184 ( .A(n3913), .B(n3930), .Z(n3914) );
  AND U4185 ( .A(e_input[4]), .B(g_input[14]), .Z(n3930) );
  XNOR U4186 ( .A(n3934), .B(n3915), .Z(n3929) );
  NAND U4187 ( .A(g_input[13]), .B(e_input[5]), .Z(n3915) );
  IV U4188 ( .A(n3917), .Z(n3934) );
  XNOR U4189 ( .A(n3923), .B(n3924), .Z(n3919) );
  NAND U4190 ( .A(g_input[11]), .B(e_input[7]), .Z(n3924) );
  XNOR U4191 ( .A(n3921), .B(n3938), .Z(n3923) );
  AND U4192 ( .A(e_input[6]), .B(g_input[12]), .Z(n3938) );
  XNOR U4193 ( .A(n3942), .B(n3939), .Z(n3940) );
  XOR U4194 ( .A(n3943), .B(n3944), .Z(n3511) );
  XNOR U4195 ( .A(n3945), .B(n3928), .Z(n3943) );
  XOR U4196 ( .A(n3931), .B(n3948), .Z(n3932) );
  AND U4197 ( .A(e_input[4]), .B(g_input[13]), .Z(n3948) );
  XNOR U4198 ( .A(n3952), .B(n3933), .Z(n3947) );
  NAND U4199 ( .A(g_input[12]), .B(e_input[5]), .Z(n3933) );
  IV U4200 ( .A(n3935), .Z(n3952) );
  XNOR U4201 ( .A(n3941), .B(n3942), .Z(n3937) );
  NAND U4202 ( .A(g_input[10]), .B(e_input[7]), .Z(n3942) );
  XNOR U4203 ( .A(n3939), .B(n3956), .Z(n3941) );
  AND U4204 ( .A(e_input[6]), .B(g_input[11]), .Z(n3956) );
  XNOR U4205 ( .A(n3960), .B(n3957), .Z(n3958) );
  XOR U4206 ( .A(n3961), .B(n3962), .Z(n3551) );
  XNOR U4207 ( .A(n3963), .B(n3946), .Z(n3961) );
  XOR U4208 ( .A(n3949), .B(n3966), .Z(n3950) );
  AND U4209 ( .A(e_input[4]), .B(g_input[12]), .Z(n3966) );
  XNOR U4210 ( .A(n3970), .B(n3951), .Z(n3965) );
  NAND U4211 ( .A(g_input[11]), .B(e_input[5]), .Z(n3951) );
  IV U4212 ( .A(n3953), .Z(n3970) );
  XNOR U4213 ( .A(n3959), .B(n3960), .Z(n3955) );
  NAND U4214 ( .A(g_input[9]), .B(e_input[7]), .Z(n3960) );
  XNOR U4215 ( .A(n3957), .B(n3974), .Z(n3959) );
  AND U4216 ( .A(e_input[6]), .B(g_input[10]), .Z(n3974) );
  XNOR U4217 ( .A(n3978), .B(n3975), .Z(n3976) );
  XOR U4218 ( .A(n3979), .B(n3980), .Z(n3685) );
  XNOR U4219 ( .A(n3981), .B(n3964), .Z(n3979) );
  XOR U4220 ( .A(n3982), .B(n3983), .Z(n3964) );
  AND U4221 ( .A(n3984), .B(n3985), .Z(n3983) );
  XOR U4222 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U4223 ( .A(n3982), .B(n3988), .Z(n3987) );
  XOR U4224 ( .A(n3972), .B(n3989), .Z(n3984) );
  XOR U4225 ( .A(n3982), .B(n3973), .Z(n3989) );
  NAND U4226 ( .A(e_input[7]), .B(g_input[8]), .Z(n3978) );
  XOR U4227 ( .A(n3975), .B(n3990), .Z(n3977) );
  AND U4228 ( .A(e_input[6]), .B(g_input[9]), .Z(n3990) );
  XNOR U4229 ( .A(n3994), .B(n3991), .Z(n3992) );
  XOR U4230 ( .A(n3967), .B(n3996), .Z(n3968) );
  AND U4231 ( .A(e_input[4]), .B(g_input[11]), .Z(n3996) );
  XNOR U4232 ( .A(n4000), .B(n3969), .Z(n3995) );
  NAND U4233 ( .A(g_input[10]), .B(e_input[5]), .Z(n3969) );
  IV U4234 ( .A(n3971), .Z(n4000) );
  XOR U4235 ( .A(n4004), .B(n4005), .Z(n3982) );
  AND U4236 ( .A(n4006), .B(n4007), .Z(n4005) );
  XOR U4237 ( .A(n4008), .B(n4009), .Z(n4007) );
  XOR U4238 ( .A(n4004), .B(n4010), .Z(n4009) );
  XOR U4239 ( .A(n4002), .B(n4011), .Z(n4006) );
  XOR U4240 ( .A(n4004), .B(n4003), .Z(n4011) );
  NAND U4241 ( .A(e_input[7]), .B(g_input[7]), .Z(n3994) );
  XOR U4242 ( .A(n3991), .B(n4012), .Z(n3993) );
  AND U4243 ( .A(g_input[8]), .B(e_input[6]), .Z(n4012) );
  XNOR U4244 ( .A(n4016), .B(n4013), .Z(n4014) );
  XOR U4245 ( .A(n3997), .B(n4018), .Z(n3998) );
  AND U4246 ( .A(e_input[4]), .B(g_input[10]), .Z(n4018) );
  XNOR U4247 ( .A(n4022), .B(n3999), .Z(n4017) );
  NAND U4248 ( .A(g_input[9]), .B(e_input[5]), .Z(n3999) );
  IV U4249 ( .A(n4001), .Z(n4022) );
  XOR U4250 ( .A(n4026), .B(n4027), .Z(n4004) );
  AND U4251 ( .A(n4028), .B(n4029), .Z(n4027) );
  XOR U4252 ( .A(n4030), .B(n4031), .Z(n4029) );
  XOR U4253 ( .A(n4026), .B(n4032), .Z(n4031) );
  XOR U4254 ( .A(n4024), .B(n4033), .Z(n4028) );
  XOR U4255 ( .A(n4026), .B(n4025), .Z(n4033) );
  NAND U4256 ( .A(e_input[7]), .B(g_input[6]), .Z(n4016) );
  XOR U4257 ( .A(n4013), .B(n4034), .Z(n4015) );
  AND U4258 ( .A(g_input[7]), .B(e_input[6]), .Z(n4034) );
  XNOR U4259 ( .A(n4038), .B(n4035), .Z(n4036) );
  XOR U4260 ( .A(n4019), .B(n4040), .Z(n4020) );
  AND U4261 ( .A(e_input[4]), .B(g_input[9]), .Z(n4040) );
  XNOR U4262 ( .A(n4044), .B(n4021), .Z(n4039) );
  NAND U4263 ( .A(e_input[5]), .B(g_input[8]), .Z(n4021) );
  IV U4264 ( .A(n4023), .Z(n4044) );
  XOR U4265 ( .A(n4048), .B(n4049), .Z(n4026) );
  AND U4266 ( .A(n4050), .B(n4051), .Z(n4049) );
  XOR U4267 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U4268 ( .A(n4048), .B(n4054), .Z(n4053) );
  XOR U4269 ( .A(n4046), .B(n4055), .Z(n4050) );
  XOR U4270 ( .A(n4048), .B(n4047), .Z(n4055) );
  NAND U4271 ( .A(e_input[7]), .B(g_input[5]), .Z(n4038) );
  XOR U4272 ( .A(n4035), .B(n4056), .Z(n4037) );
  AND U4273 ( .A(g_input[6]), .B(e_input[6]), .Z(n4056) );
  XNOR U4274 ( .A(n4060), .B(n4057), .Z(n4058) );
  XOR U4275 ( .A(n4041), .B(n4062), .Z(n4042) );
  AND U4276 ( .A(g_input[8]), .B(e_input[4]), .Z(n4062) );
  XNOR U4277 ( .A(n4066), .B(n4043), .Z(n4061) );
  NAND U4278 ( .A(e_input[5]), .B(g_input[7]), .Z(n4043) );
  IV U4279 ( .A(n4045), .Z(n4066) );
  XOR U4280 ( .A(n4070), .B(n4071), .Z(n4048) );
  AND U4281 ( .A(n4072), .B(n4073), .Z(n4071) );
  XOR U4282 ( .A(n4074), .B(n4075), .Z(n4073) );
  XOR U4283 ( .A(n4070), .B(n4076), .Z(n4075) );
  XOR U4284 ( .A(n4068), .B(n4077), .Z(n4072) );
  XOR U4285 ( .A(n4070), .B(n4069), .Z(n4077) );
  NAND U4286 ( .A(e_input[7]), .B(g_input[4]), .Z(n4060) );
  XOR U4287 ( .A(n4057), .B(n4078), .Z(n4059) );
  AND U4288 ( .A(g_input[5]), .B(e_input[6]), .Z(n4078) );
  XNOR U4289 ( .A(n4082), .B(n4079), .Z(n4080) );
  XOR U4290 ( .A(n4063), .B(n4084), .Z(n4064) );
  AND U4291 ( .A(g_input[7]), .B(e_input[4]), .Z(n4084) );
  XNOR U4292 ( .A(n4088), .B(n4065), .Z(n4083) );
  NAND U4293 ( .A(e_input[5]), .B(g_input[6]), .Z(n4065) );
  IV U4294 ( .A(n4067), .Z(n4088) );
  XOR U4295 ( .A(n4092), .B(n4093), .Z(n4070) );
  AND U4296 ( .A(n4094), .B(n4095), .Z(n4093) );
  XOR U4297 ( .A(n4096), .B(n4097), .Z(n4095) );
  XOR U4298 ( .A(n4092), .B(n4098), .Z(n4097) );
  XOR U4299 ( .A(n4090), .B(n4099), .Z(n4094) );
  XOR U4300 ( .A(n4092), .B(n4091), .Z(n4099) );
  NAND U4301 ( .A(e_input[7]), .B(g_input[3]), .Z(n4082) );
  XOR U4302 ( .A(n4079), .B(n4100), .Z(n4081) );
  AND U4303 ( .A(g_input[4]), .B(e_input[6]), .Z(n4100) );
  XNOR U4304 ( .A(n4104), .B(n4101), .Z(n4102) );
  XOR U4305 ( .A(n4085), .B(n4106), .Z(n4086) );
  AND U4306 ( .A(g_input[6]), .B(e_input[4]), .Z(n4106) );
  XNOR U4307 ( .A(n4110), .B(n4087), .Z(n4105) );
  NAND U4308 ( .A(e_input[5]), .B(g_input[5]), .Z(n4087) );
  IV U4309 ( .A(n4089), .Z(n4110) );
  XOR U4310 ( .A(n4114), .B(n4115), .Z(n4092) );
  AND U4311 ( .A(n4116), .B(n4117), .Z(n4115) );
  XOR U4312 ( .A(n4118), .B(n4119), .Z(n4117) );
  XOR U4313 ( .A(n4114), .B(n4120), .Z(n4119) );
  XOR U4314 ( .A(n4112), .B(n4121), .Z(n4116) );
  XOR U4315 ( .A(n4114), .B(n4113), .Z(n4121) );
  NAND U4316 ( .A(e_input[7]), .B(g_input[2]), .Z(n4104) );
  XOR U4317 ( .A(n4101), .B(n4122), .Z(n4103) );
  AND U4318 ( .A(g_input[3]), .B(e_input[6]), .Z(n4122) );
  XNOR U4319 ( .A(n4126), .B(n4123), .Z(n4124) );
  XOR U4320 ( .A(n4107), .B(n4128), .Z(n4108) );
  AND U4321 ( .A(g_input[5]), .B(e_input[4]), .Z(n4128) );
  XNOR U4322 ( .A(n4132), .B(n4109), .Z(n4127) );
  NAND U4323 ( .A(e_input[5]), .B(g_input[4]), .Z(n4109) );
  IV U4324 ( .A(n4111), .Z(n4132) );
  XNOR U4325 ( .A(n4137), .B(n4138), .Z(n3687) );
  XNOR U4326 ( .A(n4139), .B(n4136), .Z(n4137) );
  XOR U4327 ( .A(n4129), .B(n4141), .Z(n4130) );
  AND U4328 ( .A(g_input[4]), .B(e_input[4]), .Z(n4141) );
  XOR U4329 ( .A(n4144), .B(n4142), .Z(n4143) );
  AND U4330 ( .A(g_input[3]), .B(e_input[4]), .Z(n4144) );
  AND U4331 ( .A(g_input[2]), .B(e_input[5]), .Z(n4145) );
  XNOR U4332 ( .A(n4149), .B(n4146), .Z(n4147) );
  XNOR U4333 ( .A(n4150), .B(n4131), .Z(n4140) );
  NAND U4334 ( .A(e_input[5]), .B(g_input[3]), .Z(n4131) );
  IV U4335 ( .A(n4133), .Z(n4150) );
  NAND U4336 ( .A(e_input[5]), .B(g_input[1]), .Z(n4149) );
  XOR U4337 ( .A(n4146), .B(n4151), .Z(n4148) );
  AND U4338 ( .A(g_input[2]), .B(e_input[4]), .Z(n4151) );
  AND U4339 ( .A(n4152), .B(g_input[0]), .Z(n4146) );
  NANDN U4340 ( .B(e_input[5]), .A(n4153), .Z(n4152) );
  NAND U4341 ( .A(g_input[1]), .B(e_input[4]), .Z(n4153) );
  XNOR U4342 ( .A(n4125), .B(n4126), .Z(n4135) );
  NAND U4343 ( .A(e_input[7]), .B(g_input[1]), .Z(n4126) );
  XNOR U4344 ( .A(n4123), .B(n4154), .Z(n4125) );
  AND U4345 ( .A(g_input[2]), .B(e_input[6]), .Z(n4154) );
  AND U4346 ( .A(n4155), .B(g_input[0]), .Z(n4123) );
  NANDN U4347 ( .B(e_input[7]), .A(n4156), .Z(n4155) );
  NAND U4348 ( .A(g_input[1]), .B(e_input[6]), .Z(n4156) );
  XOR U4349 ( .A(n4157), .B(n4158), .Z(n4136) );
  XNOR U4350 ( .A(n4163), .B(n2928), .Z(n4159) );
  NAND U4351 ( .A(g_input[31]), .B(e_input[1]), .Z(n2928) );
  IV U4352 ( .A(n2929), .Z(n4163) );
  XNOR U4353 ( .A(n3692), .B(n3693), .Z(n3710) );
  NAND U4354 ( .A(g_input[28]), .B(e_input[3]), .Z(n3693) );
  XNOR U4355 ( .A(n3690), .B(n4165), .Z(n3692) );
  AND U4356 ( .A(e_input[2]), .B(g_input[29]), .Z(n4165) );
  XNOR U4357 ( .A(n4169), .B(n4166), .Z(n4167) );
  XOR U4358 ( .A(n4160), .B(n4171), .Z(n4161) );
  AND U4359 ( .A(e_input[0]), .B(g_input[31]), .Z(n4171) );
  XNOR U4360 ( .A(n4175), .B(n4162), .Z(n4170) );
  NAND U4361 ( .A(g_input[30]), .B(e_input[1]), .Z(n4162) );
  IV U4362 ( .A(n4164), .Z(n4175) );
  XNOR U4363 ( .A(n4168), .B(n4169), .Z(n3728) );
  NAND U4364 ( .A(g_input[27]), .B(e_input[3]), .Z(n4169) );
  XNOR U4365 ( .A(n4166), .B(n4177), .Z(n4168) );
  AND U4366 ( .A(e_input[2]), .B(g_input[28]), .Z(n4177) );
  XNOR U4367 ( .A(n4181), .B(n4178), .Z(n4179) );
  XOR U4368 ( .A(n4172), .B(n4183), .Z(n4173) );
  AND U4369 ( .A(e_input[0]), .B(g_input[30]), .Z(n4183) );
  XNOR U4370 ( .A(n4187), .B(n4174), .Z(n4182) );
  NAND U4371 ( .A(g_input[29]), .B(e_input[1]), .Z(n4174) );
  IV U4372 ( .A(n4176), .Z(n4187) );
  XNOR U4373 ( .A(n4180), .B(n4181), .Z(n3746) );
  NAND U4374 ( .A(g_input[26]), .B(e_input[3]), .Z(n4181) );
  XNOR U4375 ( .A(n4178), .B(n4189), .Z(n4180) );
  AND U4376 ( .A(e_input[2]), .B(g_input[27]), .Z(n4189) );
  XNOR U4377 ( .A(n4193), .B(n4190), .Z(n4191) );
  XOR U4378 ( .A(n4184), .B(n4195), .Z(n4185) );
  AND U4379 ( .A(e_input[0]), .B(g_input[29]), .Z(n4195) );
  XNOR U4380 ( .A(n4199), .B(n4186), .Z(n4194) );
  NAND U4381 ( .A(g_input[28]), .B(e_input[1]), .Z(n4186) );
  IV U4382 ( .A(n4188), .Z(n4199) );
  XNOR U4383 ( .A(n4192), .B(n4193), .Z(n3764) );
  NAND U4384 ( .A(g_input[25]), .B(e_input[3]), .Z(n4193) );
  XNOR U4385 ( .A(n4190), .B(n4201), .Z(n4192) );
  AND U4386 ( .A(e_input[2]), .B(g_input[26]), .Z(n4201) );
  XNOR U4387 ( .A(n4205), .B(n4202), .Z(n4203) );
  XOR U4388 ( .A(n4196), .B(n4207), .Z(n4197) );
  AND U4389 ( .A(e_input[0]), .B(g_input[28]), .Z(n4207) );
  XNOR U4390 ( .A(n4211), .B(n4198), .Z(n4206) );
  NAND U4391 ( .A(g_input[27]), .B(e_input[1]), .Z(n4198) );
  IV U4392 ( .A(n4200), .Z(n4211) );
  XNOR U4393 ( .A(n4204), .B(n4205), .Z(n3782) );
  NAND U4394 ( .A(g_input[24]), .B(e_input[3]), .Z(n4205) );
  XNOR U4395 ( .A(n4202), .B(n4213), .Z(n4204) );
  AND U4396 ( .A(e_input[2]), .B(g_input[25]), .Z(n4213) );
  XNOR U4397 ( .A(n4217), .B(n4214), .Z(n4215) );
  XOR U4398 ( .A(n4208), .B(n4219), .Z(n4209) );
  AND U4399 ( .A(e_input[0]), .B(g_input[27]), .Z(n4219) );
  XNOR U4400 ( .A(n4223), .B(n4210), .Z(n4218) );
  NAND U4401 ( .A(g_input[26]), .B(e_input[1]), .Z(n4210) );
  IV U4402 ( .A(n4212), .Z(n4223) );
  XNOR U4403 ( .A(n4216), .B(n4217), .Z(n3800) );
  NAND U4404 ( .A(g_input[23]), .B(e_input[3]), .Z(n4217) );
  XNOR U4405 ( .A(n4214), .B(n4225), .Z(n4216) );
  AND U4406 ( .A(e_input[2]), .B(g_input[24]), .Z(n4225) );
  XNOR U4407 ( .A(n4229), .B(n4226), .Z(n4227) );
  XOR U4408 ( .A(n4220), .B(n4231), .Z(n4221) );
  AND U4409 ( .A(e_input[0]), .B(g_input[26]), .Z(n4231) );
  XNOR U4410 ( .A(n4235), .B(n4222), .Z(n4230) );
  NAND U4411 ( .A(g_input[25]), .B(e_input[1]), .Z(n4222) );
  IV U4412 ( .A(n4224), .Z(n4235) );
  XNOR U4413 ( .A(n4228), .B(n4229), .Z(n3818) );
  NAND U4414 ( .A(g_input[22]), .B(e_input[3]), .Z(n4229) );
  XNOR U4415 ( .A(n4226), .B(n4237), .Z(n4228) );
  AND U4416 ( .A(e_input[2]), .B(g_input[23]), .Z(n4237) );
  XNOR U4417 ( .A(n4241), .B(n4238), .Z(n4239) );
  XOR U4418 ( .A(n4232), .B(n4243), .Z(n4233) );
  AND U4419 ( .A(e_input[0]), .B(g_input[25]), .Z(n4243) );
  XNOR U4420 ( .A(n4247), .B(n4234), .Z(n4242) );
  NAND U4421 ( .A(g_input[24]), .B(e_input[1]), .Z(n4234) );
  IV U4422 ( .A(n4236), .Z(n4247) );
  XNOR U4423 ( .A(n4240), .B(n4241), .Z(n3836) );
  NAND U4424 ( .A(g_input[21]), .B(e_input[3]), .Z(n4241) );
  XNOR U4425 ( .A(n4238), .B(n4249), .Z(n4240) );
  AND U4426 ( .A(e_input[2]), .B(g_input[22]), .Z(n4249) );
  XNOR U4427 ( .A(n4253), .B(n4250), .Z(n4251) );
  XOR U4428 ( .A(n4244), .B(n4255), .Z(n4245) );
  AND U4429 ( .A(e_input[0]), .B(g_input[24]), .Z(n4255) );
  XNOR U4430 ( .A(n4259), .B(n4246), .Z(n4254) );
  NAND U4431 ( .A(g_input[23]), .B(e_input[1]), .Z(n4246) );
  IV U4432 ( .A(n4248), .Z(n4259) );
  XNOR U4433 ( .A(n4252), .B(n4253), .Z(n3854) );
  NAND U4434 ( .A(g_input[20]), .B(e_input[3]), .Z(n4253) );
  XNOR U4435 ( .A(n4250), .B(n4261), .Z(n4252) );
  AND U4436 ( .A(e_input[2]), .B(g_input[21]), .Z(n4261) );
  XNOR U4437 ( .A(n4265), .B(n4262), .Z(n4263) );
  XOR U4438 ( .A(n4256), .B(n4267), .Z(n4257) );
  AND U4439 ( .A(e_input[0]), .B(g_input[23]), .Z(n4267) );
  XNOR U4440 ( .A(n4271), .B(n4258), .Z(n4266) );
  NAND U4441 ( .A(g_input[22]), .B(e_input[1]), .Z(n4258) );
  IV U4442 ( .A(n4260), .Z(n4271) );
  XNOR U4443 ( .A(n4264), .B(n4265), .Z(n3872) );
  NAND U4444 ( .A(g_input[19]), .B(e_input[3]), .Z(n4265) );
  XNOR U4445 ( .A(n4262), .B(n4273), .Z(n4264) );
  AND U4446 ( .A(e_input[2]), .B(g_input[20]), .Z(n4273) );
  XNOR U4447 ( .A(n4277), .B(n4274), .Z(n4275) );
  XOR U4448 ( .A(n4268), .B(n4279), .Z(n4269) );
  AND U4449 ( .A(e_input[0]), .B(g_input[22]), .Z(n4279) );
  XNOR U4450 ( .A(n4283), .B(n4270), .Z(n4278) );
  NAND U4451 ( .A(g_input[21]), .B(e_input[1]), .Z(n4270) );
  IV U4452 ( .A(n4272), .Z(n4283) );
  XNOR U4453 ( .A(n4276), .B(n4277), .Z(n3890) );
  NAND U4454 ( .A(g_input[18]), .B(e_input[3]), .Z(n4277) );
  XNOR U4455 ( .A(n4274), .B(n4285), .Z(n4276) );
  AND U4456 ( .A(e_input[2]), .B(g_input[19]), .Z(n4285) );
  XNOR U4457 ( .A(n4289), .B(n4286), .Z(n4287) );
  XOR U4458 ( .A(n4280), .B(n4291), .Z(n4281) );
  AND U4459 ( .A(e_input[0]), .B(g_input[21]), .Z(n4291) );
  XNOR U4460 ( .A(n4295), .B(n4282), .Z(n4290) );
  NAND U4461 ( .A(g_input[20]), .B(e_input[1]), .Z(n4282) );
  IV U4462 ( .A(n4284), .Z(n4295) );
  XNOR U4463 ( .A(n4288), .B(n4289), .Z(n3908) );
  NAND U4464 ( .A(g_input[17]), .B(e_input[3]), .Z(n4289) );
  XNOR U4465 ( .A(n4286), .B(n4297), .Z(n4288) );
  AND U4466 ( .A(e_input[2]), .B(g_input[18]), .Z(n4297) );
  XNOR U4467 ( .A(n4301), .B(n4298), .Z(n4299) );
  XOR U4468 ( .A(n4292), .B(n4303), .Z(n4293) );
  AND U4469 ( .A(e_input[0]), .B(g_input[20]), .Z(n4303) );
  XNOR U4470 ( .A(n4307), .B(n4294), .Z(n4302) );
  NAND U4471 ( .A(g_input[19]), .B(e_input[1]), .Z(n4294) );
  IV U4472 ( .A(n4296), .Z(n4307) );
  XNOR U4473 ( .A(n4300), .B(n4301), .Z(n3926) );
  NAND U4474 ( .A(g_input[16]), .B(e_input[3]), .Z(n4301) );
  XNOR U4475 ( .A(n4298), .B(n4309), .Z(n4300) );
  AND U4476 ( .A(e_input[2]), .B(g_input[17]), .Z(n4309) );
  XNOR U4477 ( .A(n4313), .B(n4310), .Z(n4311) );
  XOR U4478 ( .A(n4304), .B(n4315), .Z(n4305) );
  AND U4479 ( .A(e_input[0]), .B(g_input[19]), .Z(n4315) );
  XNOR U4480 ( .A(n4319), .B(n4306), .Z(n4314) );
  NAND U4481 ( .A(g_input[18]), .B(e_input[1]), .Z(n4306) );
  IV U4482 ( .A(n4308), .Z(n4319) );
  XNOR U4483 ( .A(n4312), .B(n4313), .Z(n3944) );
  NAND U4484 ( .A(g_input[15]), .B(e_input[3]), .Z(n4313) );
  XNOR U4485 ( .A(n4310), .B(n4321), .Z(n4312) );
  AND U4486 ( .A(e_input[2]), .B(g_input[16]), .Z(n4321) );
  XNOR U4487 ( .A(n4325), .B(n4322), .Z(n4323) );
  XOR U4488 ( .A(n4316), .B(n4327), .Z(n4317) );
  AND U4489 ( .A(e_input[0]), .B(g_input[18]), .Z(n4327) );
  XNOR U4490 ( .A(n4331), .B(n4318), .Z(n4326) );
  NAND U4491 ( .A(g_input[17]), .B(e_input[1]), .Z(n4318) );
  IV U4492 ( .A(n4320), .Z(n4331) );
  XNOR U4493 ( .A(n4324), .B(n4325), .Z(n3962) );
  NAND U4494 ( .A(g_input[14]), .B(e_input[3]), .Z(n4325) );
  XNOR U4495 ( .A(n4322), .B(n4333), .Z(n4324) );
  AND U4496 ( .A(e_input[2]), .B(g_input[15]), .Z(n4333) );
  XNOR U4497 ( .A(n4337), .B(n4334), .Z(n4335) );
  XOR U4498 ( .A(n4328), .B(n4339), .Z(n4329) );
  AND U4499 ( .A(e_input[0]), .B(g_input[17]), .Z(n4339) );
  XNOR U4500 ( .A(n4343), .B(n4330), .Z(n4338) );
  NAND U4501 ( .A(g_input[16]), .B(e_input[1]), .Z(n4330) );
  IV U4502 ( .A(n4332), .Z(n4343) );
  XNOR U4503 ( .A(n4336), .B(n4337), .Z(n3980) );
  NAND U4504 ( .A(g_input[13]), .B(e_input[3]), .Z(n4337) );
  XNOR U4505 ( .A(n4334), .B(n4345), .Z(n4336) );
  AND U4506 ( .A(e_input[2]), .B(g_input[14]), .Z(n4345) );
  XNOR U4507 ( .A(n4349), .B(n4346), .Z(n4347) );
  XOR U4508 ( .A(n4340), .B(n4351), .Z(n4341) );
  AND U4509 ( .A(e_input[0]), .B(g_input[16]), .Z(n4351) );
  XNOR U4510 ( .A(n4355), .B(n4342), .Z(n4350) );
  NAND U4511 ( .A(g_input[15]), .B(e_input[1]), .Z(n4342) );
  IV U4512 ( .A(n4344), .Z(n4355) );
  NAND U4513 ( .A(g_input[12]), .B(e_input[3]), .Z(n4349) );
  XOR U4514 ( .A(n4346), .B(n4357), .Z(n4348) );
  AND U4515 ( .A(e_input[2]), .B(g_input[13]), .Z(n4357) );
  XNOR U4516 ( .A(n4361), .B(n4358), .Z(n4359) );
  XOR U4517 ( .A(n4352), .B(n4363), .Z(n4353) );
  AND U4518 ( .A(e_input[0]), .B(g_input[15]), .Z(n4363) );
  XNOR U4519 ( .A(n4367), .B(n4354), .Z(n4362) );
  NAND U4520 ( .A(g_input[14]), .B(e_input[1]), .Z(n4354) );
  IV U4521 ( .A(n4356), .Z(n4367) );
  NAND U4522 ( .A(g_input[11]), .B(e_input[3]), .Z(n4361) );
  XOR U4523 ( .A(n4358), .B(n4369), .Z(n4360) );
  AND U4524 ( .A(e_input[2]), .B(g_input[12]), .Z(n4369) );
  XNOR U4525 ( .A(n4373), .B(n4370), .Z(n4371) );
  XOR U4526 ( .A(n4364), .B(n4375), .Z(n4365) );
  AND U4527 ( .A(e_input[0]), .B(g_input[14]), .Z(n4375) );
  XNOR U4528 ( .A(n4379), .B(n4366), .Z(n4374) );
  NAND U4529 ( .A(g_input[13]), .B(e_input[1]), .Z(n4366) );
  IV U4530 ( .A(n4368), .Z(n4379) );
  NAND U4531 ( .A(g_input[10]), .B(e_input[3]), .Z(n4373) );
  XOR U4532 ( .A(n4370), .B(n4381), .Z(n4372) );
  AND U4533 ( .A(e_input[2]), .B(g_input[11]), .Z(n4381) );
  XNOR U4534 ( .A(n4385), .B(n4382), .Z(n4383) );
  XOR U4535 ( .A(n4376), .B(n4387), .Z(n4377) );
  AND U4536 ( .A(e_input[0]), .B(g_input[13]), .Z(n4387) );
  XNOR U4537 ( .A(n4391), .B(n4378), .Z(n4386) );
  NAND U4538 ( .A(g_input[12]), .B(e_input[1]), .Z(n4378) );
  IV U4539 ( .A(n4380), .Z(n4391) );
  NAND U4540 ( .A(g_input[9]), .B(e_input[3]), .Z(n4385) );
  XOR U4541 ( .A(n4382), .B(n4393), .Z(n4384) );
  AND U4542 ( .A(e_input[2]), .B(g_input[10]), .Z(n4393) );
  XNOR U4543 ( .A(n4397), .B(n4394), .Z(n4395) );
  XOR U4544 ( .A(n4388), .B(n4399), .Z(n4389) );
  AND U4545 ( .A(e_input[0]), .B(g_input[12]), .Z(n4399) );
  XNOR U4546 ( .A(n4403), .B(n4390), .Z(n4398) );
  NAND U4547 ( .A(g_input[11]), .B(e_input[1]), .Z(n4390) );
  IV U4548 ( .A(n4392), .Z(n4403) );
  NAND U4549 ( .A(g_input[8]), .B(e_input[3]), .Z(n4397) );
  XOR U4550 ( .A(n4394), .B(n4405), .Z(n4396) );
  AND U4551 ( .A(e_input[2]), .B(g_input[9]), .Z(n4405) );
  XNOR U4552 ( .A(n4409), .B(n4406), .Z(n4407) );
  XOR U4553 ( .A(n4400), .B(n4411), .Z(n4401) );
  AND U4554 ( .A(e_input[0]), .B(g_input[11]), .Z(n4411) );
  XNOR U4555 ( .A(n4415), .B(n4402), .Z(n4410) );
  NAND U4556 ( .A(g_input[10]), .B(e_input[1]), .Z(n4402) );
  IV U4557 ( .A(n4404), .Z(n4415) );
  NAND U4558 ( .A(g_input[7]), .B(e_input[3]), .Z(n4409) );
  XOR U4559 ( .A(n4406), .B(n4417), .Z(n4408) );
  AND U4560 ( .A(e_input[2]), .B(g_input[8]), .Z(n4417) );
  XNOR U4561 ( .A(n4421), .B(n4418), .Z(n4419) );
  XOR U4562 ( .A(n4412), .B(n4423), .Z(n4413) );
  AND U4563 ( .A(e_input[0]), .B(g_input[10]), .Z(n4423) );
  XNOR U4564 ( .A(n4427), .B(n4414), .Z(n4422) );
  NAND U4565 ( .A(g_input[9]), .B(e_input[1]), .Z(n4414) );
  IV U4566 ( .A(n4416), .Z(n4427) );
  NAND U4567 ( .A(g_input[6]), .B(e_input[3]), .Z(n4421) );
  XOR U4568 ( .A(n4418), .B(n4429), .Z(n4420) );
  AND U4569 ( .A(e_input[2]), .B(g_input[7]), .Z(n4429) );
  XNOR U4570 ( .A(n4433), .B(n4430), .Z(n4431) );
  XOR U4571 ( .A(n4424), .B(n4435), .Z(n4425) );
  AND U4572 ( .A(e_input[0]), .B(g_input[9]), .Z(n4435) );
  XNOR U4573 ( .A(n4439), .B(n4426), .Z(n4434) );
  NAND U4574 ( .A(g_input[8]), .B(e_input[1]), .Z(n4426) );
  IV U4575 ( .A(n4428), .Z(n4439) );
  XNOR U4576 ( .A(n4432), .B(n4433), .Z(n4138) );
  NAND U4577 ( .A(g_input[5]), .B(e_input[3]), .Z(n4433) );
  XNOR U4578 ( .A(n4430), .B(n4441), .Z(n4432) );
  AND U4579 ( .A(e_input[2]), .B(g_input[6]), .Z(n4441) );
  XNOR U4580 ( .A(n4445), .B(n4442), .Z(n4444) );
  XOR U4581 ( .A(n4436), .B(n4447), .Z(n4437) );
  AND U4582 ( .A(e_input[0]), .B(g_input[8]), .Z(n4447) );
  XNOR U4583 ( .A(n4451), .B(n4448), .Z(n4450) );
  XNOR U4584 ( .A(n4452), .B(n4438), .Z(n4446) );
  NAND U4585 ( .A(g_input[7]), .B(e_input[1]), .Z(n4438) );
  IV U4586 ( .A(n4440), .Z(n4452) );
  XOR U4587 ( .A(n4453), .B(n4454), .Z(n4440) );
  AND U4588 ( .A(n4455), .B(n4456), .Z(n4454) );
  XOR U4589 ( .A(n4449), .B(n4457), .Z(n4456) );
  XNOR U4590 ( .A(n4451), .B(n4453), .Z(n4457) );
  NAND U4591 ( .A(g_input[6]), .B(e_input[1]), .Z(n4451) );
  XOR U4592 ( .A(n4448), .B(n4458), .Z(n4449) );
  AND U4593 ( .A(e_input[0]), .B(g_input[7]), .Z(n4458) );
  XNOR U4594 ( .A(n4462), .B(n4459), .Z(n4461) );
  XOR U4595 ( .A(n4443), .B(n4463), .Z(n4455) );
  XNOR U4596 ( .A(n4445), .B(n4453), .Z(n4463) );
  NAND U4597 ( .A(e_input[3]), .B(g_input[4]), .Z(n4445) );
  XOR U4598 ( .A(n4442), .B(n4464), .Z(n4443) );
  AND U4599 ( .A(e_input[2]), .B(g_input[5]), .Z(n4464) );
  XNOR U4600 ( .A(n4468), .B(n4465), .Z(n4467) );
  XOR U4601 ( .A(n4469), .B(n4470), .Z(n4453) );
  AND U4602 ( .A(n4471), .B(n4472), .Z(n4470) );
  XOR U4603 ( .A(n4460), .B(n4473), .Z(n4472) );
  XNOR U4604 ( .A(n4462), .B(n4469), .Z(n4473) );
  NAND U4605 ( .A(g_input[5]), .B(e_input[1]), .Z(n4462) );
  XOR U4606 ( .A(n4459), .B(n4474), .Z(n4460) );
  AND U4607 ( .A(e_input[0]), .B(g_input[6]), .Z(n4474) );
  XNOR U4608 ( .A(n4478), .B(n4475), .Z(n4477) );
  XOR U4609 ( .A(n4466), .B(n4479), .Z(n4471) );
  XNOR U4610 ( .A(n4468), .B(n4469), .Z(n4479) );
  NAND U4611 ( .A(e_input[3]), .B(g_input[3]), .Z(n4468) );
  XOR U4612 ( .A(n4465), .B(n4480), .Z(n4466) );
  AND U4613 ( .A(g_input[4]), .B(e_input[2]), .Z(n4480) );
  XNOR U4614 ( .A(n4484), .B(n4481), .Z(n4483) );
  XOR U4615 ( .A(n4485), .B(n4486), .Z(n4469) );
  AND U4616 ( .A(n4487), .B(n4488), .Z(n4486) );
  XOR U4617 ( .A(n4476), .B(n4489), .Z(n4488) );
  XNOR U4618 ( .A(n4478), .B(n4485), .Z(n4489) );
  NAND U4619 ( .A(g_input[4]), .B(e_input[1]), .Z(n4478) );
  XOR U4620 ( .A(n4475), .B(n4490), .Z(n4476) );
  AND U4621 ( .A(e_input[0]), .B(g_input[5]), .Z(n4490) );
  XOR U4622 ( .A(n4482), .B(n4494), .Z(n4487) );
  XNOR U4623 ( .A(n4484), .B(n4485), .Z(n4494) );
  NAND U4624 ( .A(e_input[3]), .B(g_input[2]), .Z(n4484) );
  XOR U4625 ( .A(n4481), .B(n4495), .Z(n4482) );
  AND U4626 ( .A(g_input[3]), .B(e_input[2]), .Z(n4495) );
  XNOR U4627 ( .A(n4499), .B(n4496), .Z(n4497) );
  NAND U4628 ( .A(e_input[3]), .B(g_input[1]), .Z(n4499) );
  XOR U4629 ( .A(n4496), .B(n4501), .Z(n4498) );
  AND U4630 ( .A(g_input[2]), .B(e_input[2]), .Z(n4501) );
  AND U4631 ( .A(n4502), .B(g_input[0]), .Z(n4496) );
  NANDN U4632 ( .B(e_input[3]), .A(n4503), .Z(n4502) );
  NAND U4633 ( .A(g_input[1]), .B(e_input[2]), .Z(n4503) );
  XOR U4634 ( .A(n4491), .B(n4505), .Z(n4492) );
  AND U4635 ( .A(e_input[0]), .B(g_input[4]), .Z(n4505) );
  XOR U4636 ( .A(n4508), .B(n4506), .Z(n4507) );
  AND U4637 ( .A(e_input[0]), .B(g_input[3]), .Z(n4508) );
  AND U4638 ( .A(e_input[1]), .B(g_input[2]), .Z(n4509) );
  XNOR U4639 ( .A(n4513), .B(n4510), .Z(n4511) );
  XNOR U4640 ( .A(n4514), .B(n4493), .Z(n4504) );
  NAND U4641 ( .A(g_input[3]), .B(e_input[1]), .Z(n4493) );
  IV U4642 ( .A(n4500), .Z(n4514) );
  NAND U4643 ( .A(g_input[1]), .B(e_input[1]), .Z(n4513) );
  XOR U4644 ( .A(n4510), .B(n4515), .Z(n4512) );
  AND U4645 ( .A(e_input[0]), .B(g_input[2]), .Z(n4515) );
  AND U4646 ( .A(n4516), .B(g_input[0]), .Z(n4510) );
  NANDN U4647 ( .B(e_input[1]), .A(n4517), .Z(n4516) );
  NAND U4648 ( .A(g_input[1]), .B(e_input[0]), .Z(n4517) );
  XOR U4649 ( .A(n4518), .B(n2418), .Z(n2408) );
  XOR U4650 ( .A(n2395), .B(n4520), .Z(n2396) );
  AND U4651 ( .A(g_input[13]), .B(e_input[20]), .Z(n4520) );
  XNOR U4652 ( .A(n4524), .B(n2397), .Z(n4519) );
  NAND U4653 ( .A(e_input[21]), .B(g_input[12]), .Z(n2397) );
  IV U4654 ( .A(n2399), .Z(n4524) );
  XNOR U4655 ( .A(n2405), .B(n2406), .Z(n2401) );
  NAND U4656 ( .A(e_input[23]), .B(g_input[10]), .Z(n2406) );
  XNOR U4657 ( .A(n2403), .B(n4528), .Z(n2405) );
  AND U4658 ( .A(g_input[11]), .B(e_input[22]), .Z(n4528) );
  XNOR U4659 ( .A(n4532), .B(n4529), .Z(n4530) );
  XNOR U4660 ( .A(n2417), .B(n2407), .Z(n4518) );
  XOR U4661 ( .A(n4534), .B(n4535), .Z(n2934) );
  XNOR U4662 ( .A(n4536), .B(n4533), .Z(n4534) );
  XOR U4663 ( .A(n4539), .B(n4540), .Z(n4533) );
  XOR U4664 ( .A(n4541), .B(n2427), .Z(n2417) );
  XNOR U4665 ( .A(n2414), .B(n2415), .Z(n2427) );
  NAND U4666 ( .A(e_input[19]), .B(g_input[14]), .Z(n2415) );
  XNOR U4667 ( .A(n2412), .B(n4542), .Z(n2414) );
  AND U4668 ( .A(g_input[15]), .B(e_input[18]), .Z(n4542) );
  XNOR U4669 ( .A(n4546), .B(n4543), .Z(n4544) );
  XNOR U4670 ( .A(n2426), .B(n2416), .Z(n4541) );
  XOR U4671 ( .A(n4521), .B(n4549), .Z(n4522) );
  AND U4672 ( .A(g_input[12]), .B(e_input[20]), .Z(n4549) );
  XNOR U4673 ( .A(n4553), .B(n4523), .Z(n4548) );
  NAND U4674 ( .A(e_input[21]), .B(g_input[11]), .Z(n4523) );
  IV U4675 ( .A(n4525), .Z(n4553) );
  XNOR U4676 ( .A(n4531), .B(n4532), .Z(n4527) );
  NAND U4677 ( .A(e_input[23]), .B(g_input[9]), .Z(n4532) );
  XNOR U4678 ( .A(n4529), .B(n4557), .Z(n4531) );
  AND U4679 ( .A(g_input[10]), .B(e_input[22]), .Z(n4557) );
  XNOR U4680 ( .A(n4561), .B(n4558), .Z(n4559) );
  XOR U4681 ( .A(n4562), .B(n4563), .Z(n4536) );
  XNOR U4682 ( .A(n4564), .B(n4547), .Z(n4562) );
  XOR U4683 ( .A(n4565), .B(n4566), .Z(n4547) );
  AND U4684 ( .A(n4567), .B(n4568), .Z(n4566) );
  XOR U4685 ( .A(n4569), .B(n4570), .Z(n4568) );
  XOR U4686 ( .A(n4565), .B(n4571), .Z(n4570) );
  XOR U4687 ( .A(n4555), .B(n4572), .Z(n4567) );
  XOR U4688 ( .A(n4565), .B(n4556), .Z(n4572) );
  NAND U4689 ( .A(e_input[23]), .B(g_input[8]), .Z(n4561) );
  XOR U4690 ( .A(n4558), .B(n4573), .Z(n4560) );
  AND U4691 ( .A(g_input[9]), .B(e_input[22]), .Z(n4573) );
  XNOR U4692 ( .A(n4577), .B(n4574), .Z(n4575) );
  XOR U4693 ( .A(n4550), .B(n4579), .Z(n4551) );
  AND U4694 ( .A(g_input[11]), .B(e_input[20]), .Z(n4579) );
  XNOR U4695 ( .A(n4583), .B(n4552), .Z(n4578) );
  NAND U4696 ( .A(e_input[21]), .B(g_input[10]), .Z(n4552) );
  IV U4697 ( .A(n4554), .Z(n4583) );
  XOR U4698 ( .A(n4587), .B(n4588), .Z(n4565) );
  AND U4699 ( .A(n4589), .B(n4590), .Z(n4588) );
  XOR U4700 ( .A(n4591), .B(n4592), .Z(n4590) );
  XOR U4701 ( .A(n4587), .B(n4593), .Z(n4592) );
  XOR U4702 ( .A(n4585), .B(n4594), .Z(n4589) );
  XOR U4703 ( .A(n4587), .B(n4586), .Z(n4594) );
  NAND U4704 ( .A(e_input[23]), .B(g_input[7]), .Z(n4577) );
  XOR U4705 ( .A(n4574), .B(n4595), .Z(n4576) );
  AND U4706 ( .A(g_input[8]), .B(e_input[22]), .Z(n4595) );
  XNOR U4707 ( .A(n4599), .B(n4596), .Z(n4597) );
  XOR U4708 ( .A(n4580), .B(n4601), .Z(n4581) );
  AND U4709 ( .A(g_input[10]), .B(e_input[20]), .Z(n4601) );
  XNOR U4710 ( .A(n4605), .B(n4582), .Z(n4600) );
  NAND U4711 ( .A(e_input[21]), .B(g_input[9]), .Z(n4582) );
  IV U4712 ( .A(n4584), .Z(n4605) );
  XOR U4713 ( .A(n4609), .B(n4610), .Z(n4587) );
  AND U4714 ( .A(n4611), .B(n4612), .Z(n4610) );
  XOR U4715 ( .A(n4613), .B(n4614), .Z(n4612) );
  XOR U4716 ( .A(n4609), .B(n4615), .Z(n4614) );
  XOR U4717 ( .A(n4607), .B(n4616), .Z(n4611) );
  XOR U4718 ( .A(n4609), .B(n4608), .Z(n4616) );
  NAND U4719 ( .A(e_input[23]), .B(g_input[6]), .Z(n4599) );
  XOR U4720 ( .A(n4596), .B(n4617), .Z(n4598) );
  AND U4721 ( .A(g_input[7]), .B(e_input[22]), .Z(n4617) );
  XNOR U4722 ( .A(n4621), .B(n4618), .Z(n4619) );
  XOR U4723 ( .A(n4602), .B(n4623), .Z(n4603) );
  AND U4724 ( .A(g_input[9]), .B(e_input[20]), .Z(n4623) );
  XNOR U4725 ( .A(n4627), .B(n4604), .Z(n4622) );
  NAND U4726 ( .A(e_input[21]), .B(g_input[8]), .Z(n4604) );
  IV U4727 ( .A(n4606), .Z(n4627) );
  XOR U4728 ( .A(n4631), .B(n4632), .Z(n4609) );
  AND U4729 ( .A(n4633), .B(n4634), .Z(n4632) );
  XOR U4730 ( .A(n4635), .B(n4636), .Z(n4634) );
  XOR U4731 ( .A(n4631), .B(n4637), .Z(n4636) );
  XOR U4732 ( .A(n4629), .B(n4638), .Z(n4633) );
  XOR U4733 ( .A(n4631), .B(n4630), .Z(n4638) );
  NAND U4734 ( .A(e_input[23]), .B(g_input[5]), .Z(n4621) );
  XOR U4735 ( .A(n4618), .B(n4639), .Z(n4620) );
  AND U4736 ( .A(g_input[6]), .B(e_input[22]), .Z(n4639) );
  XNOR U4737 ( .A(n4643), .B(n4640), .Z(n4641) );
  XOR U4738 ( .A(n4624), .B(n4645), .Z(n4625) );
  AND U4739 ( .A(g_input[8]), .B(e_input[20]), .Z(n4645) );
  XNOR U4740 ( .A(n4649), .B(n4626), .Z(n4644) );
  NAND U4741 ( .A(e_input[21]), .B(g_input[7]), .Z(n4626) );
  IV U4742 ( .A(n4628), .Z(n4649) );
  XOR U4743 ( .A(n4653), .B(n4654), .Z(n4631) );
  AND U4744 ( .A(n4655), .B(n4656), .Z(n4654) );
  XOR U4745 ( .A(n4657), .B(n4658), .Z(n4656) );
  XOR U4746 ( .A(n4653), .B(n4659), .Z(n4658) );
  XOR U4747 ( .A(n4651), .B(n4660), .Z(n4655) );
  XOR U4748 ( .A(n4653), .B(n4652), .Z(n4660) );
  NAND U4749 ( .A(e_input[23]), .B(g_input[4]), .Z(n4643) );
  XOR U4750 ( .A(n4640), .B(n4661), .Z(n4642) );
  AND U4751 ( .A(g_input[5]), .B(e_input[22]), .Z(n4661) );
  XNOR U4752 ( .A(n4665), .B(n4662), .Z(n4663) );
  XOR U4753 ( .A(n4646), .B(n4667), .Z(n4647) );
  AND U4754 ( .A(g_input[7]), .B(e_input[20]), .Z(n4667) );
  XNOR U4755 ( .A(n4671), .B(n4648), .Z(n4666) );
  NAND U4756 ( .A(e_input[21]), .B(g_input[6]), .Z(n4648) );
  IV U4757 ( .A(n4650), .Z(n4671) );
  XOR U4758 ( .A(n4675), .B(n4676), .Z(n4653) );
  AND U4759 ( .A(n4677), .B(n4678), .Z(n4676) );
  XOR U4760 ( .A(n4679), .B(n4680), .Z(n4678) );
  XOR U4761 ( .A(n4675), .B(n4681), .Z(n4680) );
  XOR U4762 ( .A(n4673), .B(n4682), .Z(n4677) );
  XOR U4763 ( .A(n4675), .B(n4674), .Z(n4682) );
  NAND U4764 ( .A(e_input[23]), .B(g_input[3]), .Z(n4665) );
  XOR U4765 ( .A(n4662), .B(n4683), .Z(n4664) );
  AND U4766 ( .A(g_input[4]), .B(e_input[22]), .Z(n4683) );
  XNOR U4767 ( .A(n4687), .B(n4684), .Z(n4685) );
  XOR U4768 ( .A(n4668), .B(n4689), .Z(n4669) );
  AND U4769 ( .A(g_input[6]), .B(e_input[20]), .Z(n4689) );
  XNOR U4770 ( .A(n4693), .B(n4670), .Z(n4688) );
  NAND U4771 ( .A(e_input[21]), .B(g_input[5]), .Z(n4670) );
  IV U4772 ( .A(n4672), .Z(n4693) );
  XOR U4773 ( .A(n4697), .B(n4698), .Z(n4675) );
  AND U4774 ( .A(n4699), .B(n4700), .Z(n4698) );
  XOR U4775 ( .A(n4701), .B(n4702), .Z(n4700) );
  XOR U4776 ( .A(n4697), .B(n4703), .Z(n4702) );
  XOR U4777 ( .A(n4695), .B(n4704), .Z(n4699) );
  XOR U4778 ( .A(n4697), .B(n4696), .Z(n4704) );
  NAND U4779 ( .A(e_input[23]), .B(g_input[2]), .Z(n4687) );
  XOR U4780 ( .A(n4684), .B(n4705), .Z(n4686) );
  AND U4781 ( .A(g_input[3]), .B(e_input[22]), .Z(n4705) );
  XNOR U4782 ( .A(n4709), .B(n4706), .Z(n4707) );
  XOR U4783 ( .A(n4690), .B(n4711), .Z(n4691) );
  AND U4784 ( .A(g_input[5]), .B(e_input[20]), .Z(n4711) );
  XNOR U4785 ( .A(n4715), .B(n4692), .Z(n4710) );
  NAND U4786 ( .A(e_input[21]), .B(g_input[4]), .Z(n4692) );
  IV U4787 ( .A(n4694), .Z(n4715) );
  XOR U4788 ( .A(n4720), .B(n4721), .Z(n4540) );
  XNOR U4789 ( .A(n4722), .B(n4719), .Z(n4720) );
  XOR U4790 ( .A(n4712), .B(n4724), .Z(n4713) );
  AND U4791 ( .A(g_input[4]), .B(e_input[20]), .Z(n4724) );
  XOR U4792 ( .A(n4727), .B(n4725), .Z(n4726) );
  AND U4793 ( .A(g_input[3]), .B(e_input[20]), .Z(n4727) );
  AND U4794 ( .A(g_input[2]), .B(e_input[21]), .Z(n4728) );
  XNOR U4795 ( .A(n4732), .B(n4729), .Z(n4730) );
  XNOR U4796 ( .A(n4733), .B(n4714), .Z(n4723) );
  NAND U4797 ( .A(e_input[21]), .B(g_input[3]), .Z(n4714) );
  IV U4798 ( .A(n4716), .Z(n4733) );
  NAND U4799 ( .A(e_input[21]), .B(g_input[1]), .Z(n4732) );
  XOR U4800 ( .A(n4729), .B(n4734), .Z(n4731) );
  AND U4801 ( .A(g_input[2]), .B(e_input[20]), .Z(n4734) );
  AND U4802 ( .A(n4735), .B(g_input[0]), .Z(n4729) );
  NANDN U4803 ( .B(e_input[21]), .A(n4736), .Z(n4735) );
  NAND U4804 ( .A(g_input[1]), .B(e_input[20]), .Z(n4736) );
  XNOR U4805 ( .A(n4708), .B(n4709), .Z(n4718) );
  NAND U4806 ( .A(e_input[23]), .B(g_input[1]), .Z(n4709) );
  XNOR U4807 ( .A(n4706), .B(n4737), .Z(n4708) );
  AND U4808 ( .A(g_input[2]), .B(e_input[22]), .Z(n4737) );
  AND U4809 ( .A(n4738), .B(g_input[0]), .Z(n4706) );
  NANDN U4810 ( .B(e_input[23]), .A(n4739), .Z(n4738) );
  NAND U4811 ( .A(g_input[1]), .B(e_input[22]), .Z(n4739) );
  XOR U4812 ( .A(n4740), .B(n4741), .Z(n4719) );
  XOR U4813 ( .A(n2421), .B(n4743), .Z(n2422) );
  AND U4814 ( .A(g_input[17]), .B(e_input[16]), .Z(n4743) );
  XNOR U4815 ( .A(n4747), .B(n2423), .Z(n4742) );
  NAND U4816 ( .A(e_input[17]), .B(g_input[16]), .Z(n2423) );
  IV U4817 ( .A(n2425), .Z(n4747) );
  XNOR U4818 ( .A(n4545), .B(n4546), .Z(n4563) );
  NAND U4819 ( .A(e_input[19]), .B(g_input[13]), .Z(n4546) );
  XNOR U4820 ( .A(n4543), .B(n4749), .Z(n4545) );
  AND U4821 ( .A(g_input[14]), .B(e_input[18]), .Z(n4749) );
  XNOR U4822 ( .A(n4753), .B(n4750), .Z(n4751) );
  XOR U4823 ( .A(n4744), .B(n4755), .Z(n4745) );
  AND U4824 ( .A(g_input[16]), .B(e_input[16]), .Z(n4755) );
  XNOR U4825 ( .A(n4759), .B(n4746), .Z(n4754) );
  NAND U4826 ( .A(e_input[17]), .B(g_input[15]), .Z(n4746) );
  IV U4827 ( .A(n4748), .Z(n4759) );
  NAND U4828 ( .A(e_input[19]), .B(g_input[12]), .Z(n4753) );
  XOR U4829 ( .A(n4750), .B(n4761), .Z(n4752) );
  AND U4830 ( .A(g_input[13]), .B(e_input[18]), .Z(n4761) );
  XNOR U4831 ( .A(n4765), .B(n4762), .Z(n4763) );
  XOR U4832 ( .A(n4756), .B(n4767), .Z(n4757) );
  AND U4833 ( .A(g_input[15]), .B(e_input[16]), .Z(n4767) );
  XNOR U4834 ( .A(n4771), .B(n4758), .Z(n4766) );
  NAND U4835 ( .A(e_input[17]), .B(g_input[14]), .Z(n4758) );
  IV U4836 ( .A(n4760), .Z(n4771) );
  NAND U4837 ( .A(e_input[19]), .B(g_input[11]), .Z(n4765) );
  XOR U4838 ( .A(n4762), .B(n4773), .Z(n4764) );
  AND U4839 ( .A(g_input[12]), .B(e_input[18]), .Z(n4773) );
  XNOR U4840 ( .A(n4777), .B(n4774), .Z(n4775) );
  XOR U4841 ( .A(n4768), .B(n4779), .Z(n4769) );
  AND U4842 ( .A(g_input[14]), .B(e_input[16]), .Z(n4779) );
  XNOR U4843 ( .A(n4783), .B(n4770), .Z(n4778) );
  NAND U4844 ( .A(e_input[17]), .B(g_input[13]), .Z(n4770) );
  IV U4845 ( .A(n4772), .Z(n4783) );
  NAND U4846 ( .A(e_input[19]), .B(g_input[10]), .Z(n4777) );
  XOR U4847 ( .A(n4774), .B(n4785), .Z(n4776) );
  AND U4848 ( .A(g_input[11]), .B(e_input[18]), .Z(n4785) );
  XNOR U4849 ( .A(n4789), .B(n4786), .Z(n4787) );
  XOR U4850 ( .A(n4780), .B(n4791), .Z(n4781) );
  AND U4851 ( .A(g_input[13]), .B(e_input[16]), .Z(n4791) );
  XNOR U4852 ( .A(n4795), .B(n4782), .Z(n4790) );
  NAND U4853 ( .A(e_input[17]), .B(g_input[12]), .Z(n4782) );
  IV U4854 ( .A(n4784), .Z(n4795) );
  NAND U4855 ( .A(e_input[19]), .B(g_input[9]), .Z(n4789) );
  XOR U4856 ( .A(n4786), .B(n4797), .Z(n4788) );
  AND U4857 ( .A(g_input[10]), .B(e_input[18]), .Z(n4797) );
  XNOR U4858 ( .A(n4801), .B(n4798), .Z(n4799) );
  XOR U4859 ( .A(n4792), .B(n4803), .Z(n4793) );
  AND U4860 ( .A(g_input[12]), .B(e_input[16]), .Z(n4803) );
  XNOR U4861 ( .A(n4807), .B(n4794), .Z(n4802) );
  NAND U4862 ( .A(e_input[17]), .B(g_input[11]), .Z(n4794) );
  IV U4863 ( .A(n4796), .Z(n4807) );
  NAND U4864 ( .A(e_input[19]), .B(g_input[8]), .Z(n4801) );
  XOR U4865 ( .A(n4798), .B(n4809), .Z(n4800) );
  AND U4866 ( .A(g_input[9]), .B(e_input[18]), .Z(n4809) );
  XNOR U4867 ( .A(n4813), .B(n4810), .Z(n4811) );
  XOR U4868 ( .A(n4804), .B(n4815), .Z(n4805) );
  AND U4869 ( .A(g_input[11]), .B(e_input[16]), .Z(n4815) );
  XNOR U4870 ( .A(n4819), .B(n4806), .Z(n4814) );
  NAND U4871 ( .A(e_input[17]), .B(g_input[10]), .Z(n4806) );
  IV U4872 ( .A(n4808), .Z(n4819) );
  NAND U4873 ( .A(e_input[19]), .B(g_input[7]), .Z(n4813) );
  XOR U4874 ( .A(n4810), .B(n4821), .Z(n4812) );
  AND U4875 ( .A(g_input[8]), .B(e_input[18]), .Z(n4821) );
  XNOR U4876 ( .A(n4825), .B(n4822), .Z(n4823) );
  XOR U4877 ( .A(n4816), .B(n4827), .Z(n4817) );
  AND U4878 ( .A(g_input[10]), .B(e_input[16]), .Z(n4827) );
  XNOR U4879 ( .A(n4831), .B(n4818), .Z(n4826) );
  NAND U4880 ( .A(e_input[17]), .B(g_input[9]), .Z(n4818) );
  IV U4881 ( .A(n4820), .Z(n4831) );
  NAND U4882 ( .A(e_input[19]), .B(g_input[6]), .Z(n4825) );
  XOR U4883 ( .A(n4822), .B(n4833), .Z(n4824) );
  AND U4884 ( .A(g_input[7]), .B(e_input[18]), .Z(n4833) );
  XNOR U4885 ( .A(n4837), .B(n4834), .Z(n4835) );
  XOR U4886 ( .A(n4828), .B(n4839), .Z(n4829) );
  AND U4887 ( .A(g_input[9]), .B(e_input[16]), .Z(n4839) );
  XNOR U4888 ( .A(n4843), .B(n4830), .Z(n4838) );
  NAND U4889 ( .A(e_input[17]), .B(g_input[8]), .Z(n4830) );
  IV U4890 ( .A(n4832), .Z(n4843) );
  NAND U4891 ( .A(e_input[19]), .B(g_input[5]), .Z(n4837) );
  XOR U4892 ( .A(n4834), .B(n4845), .Z(n4836) );
  AND U4893 ( .A(g_input[6]), .B(e_input[18]), .Z(n4845) );
  XNOR U4894 ( .A(n4849), .B(n4846), .Z(n4848) );
  XOR U4895 ( .A(n4840), .B(n4851), .Z(n4841) );
  AND U4896 ( .A(g_input[8]), .B(e_input[16]), .Z(n4851) );
  XNOR U4897 ( .A(n4855), .B(n4852), .Z(n4854) );
  XNOR U4898 ( .A(n4856), .B(n4842), .Z(n4850) );
  NAND U4899 ( .A(e_input[17]), .B(g_input[7]), .Z(n4842) );
  IV U4900 ( .A(n4844), .Z(n4856) );
  XOR U4901 ( .A(n4857), .B(n4858), .Z(n4844) );
  AND U4902 ( .A(n4859), .B(n4860), .Z(n4858) );
  XOR U4903 ( .A(n4853), .B(n4861), .Z(n4860) );
  XNOR U4904 ( .A(n4855), .B(n4857), .Z(n4861) );
  NAND U4905 ( .A(e_input[17]), .B(g_input[6]), .Z(n4855) );
  XOR U4906 ( .A(n4852), .B(n4862), .Z(n4853) );
  AND U4907 ( .A(g_input[7]), .B(e_input[16]), .Z(n4862) );
  XNOR U4908 ( .A(n4866), .B(n4863), .Z(n4865) );
  XOR U4909 ( .A(n4847), .B(n4867), .Z(n4859) );
  XNOR U4910 ( .A(n4849), .B(n4857), .Z(n4867) );
  NAND U4911 ( .A(e_input[19]), .B(g_input[4]), .Z(n4849) );
  XOR U4912 ( .A(n4846), .B(n4868), .Z(n4847) );
  AND U4913 ( .A(g_input[5]), .B(e_input[18]), .Z(n4868) );
  XNOR U4914 ( .A(n4872), .B(n4869), .Z(n4871) );
  XOR U4915 ( .A(n4873), .B(n4874), .Z(n4857) );
  AND U4916 ( .A(n4875), .B(n4876), .Z(n4874) );
  XOR U4917 ( .A(n4864), .B(n4877), .Z(n4876) );
  XNOR U4918 ( .A(n4866), .B(n4873), .Z(n4877) );
  NAND U4919 ( .A(e_input[17]), .B(g_input[5]), .Z(n4866) );
  XOR U4920 ( .A(n4863), .B(n4878), .Z(n4864) );
  AND U4921 ( .A(g_input[6]), .B(e_input[16]), .Z(n4878) );
  XNOR U4922 ( .A(n4882), .B(n4879), .Z(n4881) );
  XOR U4923 ( .A(n4870), .B(n4883), .Z(n4875) );
  XNOR U4924 ( .A(n4872), .B(n4873), .Z(n4883) );
  NAND U4925 ( .A(e_input[19]), .B(g_input[3]), .Z(n4872) );
  XOR U4926 ( .A(n4869), .B(n4884), .Z(n4870) );
  AND U4927 ( .A(g_input[4]), .B(e_input[18]), .Z(n4884) );
  XNOR U4928 ( .A(n4888), .B(n4885), .Z(n4887) );
  XOR U4929 ( .A(n4889), .B(n4890), .Z(n4873) );
  AND U4930 ( .A(n4891), .B(n4892), .Z(n4890) );
  XOR U4931 ( .A(n4880), .B(n4893), .Z(n4892) );
  XNOR U4932 ( .A(n4882), .B(n4889), .Z(n4893) );
  NAND U4933 ( .A(e_input[17]), .B(g_input[4]), .Z(n4882) );
  XOR U4934 ( .A(n4879), .B(n4894), .Z(n4880) );
  AND U4935 ( .A(g_input[5]), .B(e_input[16]), .Z(n4894) );
  XOR U4936 ( .A(n4886), .B(n4898), .Z(n4891) );
  XNOR U4937 ( .A(n4888), .B(n4889), .Z(n4898) );
  NAND U4938 ( .A(e_input[19]), .B(g_input[2]), .Z(n4888) );
  XOR U4939 ( .A(n4885), .B(n4899), .Z(n4886) );
  AND U4940 ( .A(g_input[3]), .B(e_input[18]), .Z(n4899) );
  XNOR U4941 ( .A(n4903), .B(n4900), .Z(n4901) );
  NAND U4942 ( .A(e_input[19]), .B(g_input[1]), .Z(n4903) );
  XOR U4943 ( .A(n4900), .B(n4905), .Z(n4902) );
  AND U4944 ( .A(g_input[2]), .B(e_input[18]), .Z(n4905) );
  AND U4945 ( .A(n4906), .B(g_input[0]), .Z(n4900) );
  NANDN U4946 ( .B(e_input[19]), .A(n4907), .Z(n4906) );
  NAND U4947 ( .A(g_input[1]), .B(e_input[18]), .Z(n4907) );
  XOR U4948 ( .A(n4895), .B(n4909), .Z(n4896) );
  AND U4949 ( .A(g_input[4]), .B(e_input[16]), .Z(n4909) );
  XOR U4950 ( .A(n4912), .B(n4910), .Z(n4911) );
  AND U4951 ( .A(g_input[3]), .B(e_input[16]), .Z(n4912) );
  AND U4952 ( .A(g_input[2]), .B(e_input[17]), .Z(n4913) );
  XNOR U4953 ( .A(n4917), .B(n4914), .Z(n4915) );
  XNOR U4954 ( .A(n4918), .B(n4897), .Z(n4908) );
  NAND U4955 ( .A(e_input[17]), .B(g_input[3]), .Z(n4897) );
  IV U4956 ( .A(n4904), .Z(n4918) );
  NAND U4957 ( .A(e_input[17]), .B(g_input[1]), .Z(n4917) );
  XOR U4958 ( .A(n4914), .B(n4919), .Z(n4916) );
  AND U4959 ( .A(g_input[2]), .B(e_input[16]), .Z(n4919) );
  AND U4960 ( .A(n4920), .B(g_input[0]), .Z(n4914) );
  NANDN U4961 ( .B(e_input[17]), .A(n4921), .Z(n4920) );
  NAND U4962 ( .A(g_input[1]), .B(e_input[16]), .Z(n4921) );
  XOR U4963 ( .A(n4922), .B(n2445), .Z(n2435) );
  XNOR U4964 ( .A(n2432), .B(n2433), .Z(n2445) );
  NAND U4965 ( .A(e_input[27]), .B(g_input[6]), .Z(n2433) );
  XNOR U4966 ( .A(n2430), .B(n4923), .Z(n2432) );
  AND U4967 ( .A(g_input[7]), .B(e_input[26]), .Z(n4923) );
  XNOR U4968 ( .A(n4927), .B(n4924), .Z(n4925) );
  XNOR U4969 ( .A(n2444), .B(n2434), .Z(n4922) );
  XOR U4970 ( .A(n4929), .B(n4930), .Z(n4538) );
  XNOR U4971 ( .A(n4931), .B(n4928), .Z(n4929) );
  XOR U4972 ( .A(n4934), .B(n4935), .Z(n4928) );
  XOR U4973 ( .A(n2439), .B(n4937), .Z(n2440) );
  AND U4974 ( .A(g_input[9]), .B(e_input[24]), .Z(n4937) );
  XNOR U4975 ( .A(n4941), .B(n2441), .Z(n4936) );
  NAND U4976 ( .A(e_input[25]), .B(g_input[8]), .Z(n2441) );
  IV U4977 ( .A(n2443), .Z(n4941) );
  XNOR U4978 ( .A(n4926), .B(n4927), .Z(n4930) );
  NAND U4979 ( .A(e_input[27]), .B(g_input[5]), .Z(n4927) );
  XNOR U4980 ( .A(n4924), .B(n4943), .Z(n4926) );
  AND U4981 ( .A(g_input[6]), .B(e_input[26]), .Z(n4943) );
  XNOR U4982 ( .A(n4947), .B(n4944), .Z(n4946) );
  XOR U4983 ( .A(n4938), .B(n4949), .Z(n4939) );
  AND U4984 ( .A(g_input[8]), .B(e_input[24]), .Z(n4949) );
  XNOR U4985 ( .A(n4953), .B(n4950), .Z(n4952) );
  XNOR U4986 ( .A(n4954), .B(n4940), .Z(n4948) );
  NAND U4987 ( .A(e_input[25]), .B(g_input[7]), .Z(n4940) );
  IV U4988 ( .A(n4942), .Z(n4954) );
  XOR U4989 ( .A(n4955), .B(n4956), .Z(n4942) );
  AND U4990 ( .A(n4957), .B(n4958), .Z(n4956) );
  XOR U4991 ( .A(n4951), .B(n4959), .Z(n4958) );
  XNOR U4992 ( .A(n4953), .B(n4955), .Z(n4959) );
  NAND U4993 ( .A(e_input[25]), .B(g_input[6]), .Z(n4953) );
  XOR U4994 ( .A(n4950), .B(n4960), .Z(n4951) );
  AND U4995 ( .A(g_input[7]), .B(e_input[24]), .Z(n4960) );
  XNOR U4996 ( .A(n4964), .B(n4961), .Z(n4963) );
  XOR U4997 ( .A(n4945), .B(n4965), .Z(n4957) );
  XNOR U4998 ( .A(n4947), .B(n4955), .Z(n4965) );
  NAND U4999 ( .A(e_input[27]), .B(g_input[4]), .Z(n4947) );
  XOR U5000 ( .A(n4944), .B(n4966), .Z(n4945) );
  AND U5001 ( .A(g_input[5]), .B(e_input[26]), .Z(n4966) );
  XNOR U5002 ( .A(n4970), .B(n4967), .Z(n4969) );
  XOR U5003 ( .A(n4971), .B(n4972), .Z(n4955) );
  AND U5004 ( .A(n4973), .B(n4974), .Z(n4972) );
  XOR U5005 ( .A(n4962), .B(n4975), .Z(n4974) );
  XNOR U5006 ( .A(n4964), .B(n4971), .Z(n4975) );
  NAND U5007 ( .A(e_input[25]), .B(g_input[5]), .Z(n4964) );
  XOR U5008 ( .A(n4961), .B(n4976), .Z(n4962) );
  AND U5009 ( .A(g_input[6]), .B(e_input[24]), .Z(n4976) );
  XNOR U5010 ( .A(n4980), .B(n4977), .Z(n4979) );
  XOR U5011 ( .A(n4968), .B(n4981), .Z(n4973) );
  XNOR U5012 ( .A(n4970), .B(n4971), .Z(n4981) );
  NAND U5013 ( .A(e_input[27]), .B(g_input[3]), .Z(n4970) );
  XOR U5014 ( .A(n4967), .B(n4982), .Z(n4968) );
  AND U5015 ( .A(g_input[4]), .B(e_input[26]), .Z(n4982) );
  XNOR U5016 ( .A(n4986), .B(n4983), .Z(n4985) );
  XOR U5017 ( .A(n4987), .B(n4988), .Z(n4971) );
  AND U5018 ( .A(n4989), .B(n4990), .Z(n4988) );
  XOR U5019 ( .A(n4978), .B(n4991), .Z(n4990) );
  XNOR U5020 ( .A(n4980), .B(n4987), .Z(n4991) );
  NAND U5021 ( .A(e_input[25]), .B(g_input[4]), .Z(n4980) );
  XOR U5022 ( .A(n4977), .B(n4992), .Z(n4978) );
  AND U5023 ( .A(g_input[5]), .B(e_input[24]), .Z(n4992) );
  XOR U5024 ( .A(n4984), .B(n4996), .Z(n4989) );
  XNOR U5025 ( .A(n4986), .B(n4987), .Z(n4996) );
  NAND U5026 ( .A(e_input[27]), .B(g_input[2]), .Z(n4986) );
  XOR U5027 ( .A(n4983), .B(n4997), .Z(n4984) );
  AND U5028 ( .A(g_input[3]), .B(e_input[26]), .Z(n4997) );
  XNOR U5029 ( .A(n5001), .B(n4998), .Z(n4999) );
  NAND U5030 ( .A(e_input[27]), .B(g_input[1]), .Z(n5001) );
  XOR U5031 ( .A(n4998), .B(n5003), .Z(n5000) );
  AND U5032 ( .A(g_input[2]), .B(e_input[26]), .Z(n5003) );
  AND U5033 ( .A(n5004), .B(g_input[0]), .Z(n4998) );
  NANDN U5034 ( .B(e_input[27]), .A(n5005), .Z(n5004) );
  NAND U5035 ( .A(g_input[1]), .B(e_input[26]), .Z(n5005) );
  XOR U5036 ( .A(n4993), .B(n5007), .Z(n4994) );
  AND U5037 ( .A(g_input[4]), .B(e_input[24]), .Z(n5007) );
  XOR U5038 ( .A(n5010), .B(n5008), .Z(n5009) );
  AND U5039 ( .A(g_input[3]), .B(e_input[24]), .Z(n5010) );
  AND U5040 ( .A(g_input[2]), .B(e_input[25]), .Z(n5011) );
  XNOR U5041 ( .A(n5015), .B(n5012), .Z(n5013) );
  XNOR U5042 ( .A(n5016), .B(n4995), .Z(n5006) );
  NAND U5043 ( .A(e_input[25]), .B(g_input[3]), .Z(n4995) );
  IV U5044 ( .A(n5002), .Z(n5016) );
  NAND U5045 ( .A(e_input[25]), .B(g_input[1]), .Z(n5015) );
  XOR U5046 ( .A(n5012), .B(n5017), .Z(n5014) );
  AND U5047 ( .A(g_input[2]), .B(e_input[24]), .Z(n5017) );
  AND U5048 ( .A(n5018), .B(g_input[0]), .Z(n5012) );
  NANDN U5049 ( .B(e_input[25]), .A(n5019), .Z(n5018) );
  NAND U5050 ( .A(g_input[1]), .B(e_input[24]), .Z(n5019) );
  XOR U5051 ( .A(n2448), .B(n5021), .Z(n2449) );
  AND U5052 ( .A(g_input[5]), .B(e_input[28]), .Z(n5021) );
  XNOR U5053 ( .A(n5025), .B(n2450), .Z(n5020) );
  NAND U5054 ( .A(e_input[29]), .B(g_input[4]), .Z(n2450) );
  IV U5055 ( .A(n2452), .Z(n5025) );
  XOR U5056 ( .A(n5022), .B(n5028), .Z(n5023) );
  AND U5057 ( .A(g_input[4]), .B(e_input[28]), .Z(n5028) );
  XOR U5058 ( .A(n5031), .B(n5029), .Z(n5030) );
  AND U5059 ( .A(g_input[3]), .B(e_input[28]), .Z(n5031) );
  AND U5060 ( .A(g_input[2]), .B(e_input[29]), .Z(n5032) );
  XNOR U5061 ( .A(n5036), .B(n5033), .Z(n5034) );
  XNOR U5062 ( .A(n5037), .B(n5024), .Z(n5027) );
  NAND U5063 ( .A(e_input[29]), .B(g_input[3]), .Z(n5024) );
  IV U5064 ( .A(n5026), .Z(n5037) );
  XNOR U5065 ( .A(n5038), .B(n5039), .Z(n4932) );
  NAND U5066 ( .A(e_input[29]), .B(g_input[1]), .Z(n5036) );
  XOR U5067 ( .A(n5033), .B(n5040), .Z(n5035) );
  AND U5068 ( .A(g_input[2]), .B(e_input[28]), .Z(n5040) );
  AND U5069 ( .A(n5041), .B(g_input[0]), .Z(n5033) );
  NANDN U5070 ( .B(e_input[29]), .A(n5042), .Z(n5041) );
  NAND U5071 ( .A(g_input[1]), .B(e_input[28]), .Z(n5042) );
  XNOR U5072 ( .A(n2458), .B(n2459), .Z(n2454) );
  NAND U5073 ( .A(e_input[31]), .B(g_input[2]), .Z(n2459) );
  XNOR U5074 ( .A(n2456), .B(n5043), .Z(n2458) );
  AND U5075 ( .A(g_input[3]), .B(e_input[30]), .Z(n5043) );
  XNOR U5076 ( .A(n5044), .B(n5045), .Z(n5038) );
  AND U5077 ( .A(g_input[2]), .B(e_input[30]), .Z(n5045) );
  NAND U5078 ( .A(e_input[31]), .B(g_input[1]), .Z(n5039) );
  AND U5079 ( .A(n5046), .B(g_input[0]), .Z(n5044) );
  NANDN U5080 ( .B(e_input[31]), .A(n5047), .Z(n5046) );
  NAND U5081 ( .A(g_input[1]), .B(e_input[30]), .Z(n5047) );
endmodule

