
module MxM_W16_N1000 ( clk, rst, A, X, Y );
  input [15:0] A;
  input [15:0] X;
  output [15:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, \add_25/carry[9] , \add_25/carry[8] ,
         \add_25/carry[7] , \add_25/carry[6] , \add_25/carry[5] ,
         \add_25/carry[4] , \add_25/carry[3] , \add_25/carry[2] , n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736;
  wire   [15:0] Y0;
  wire   [9:0] n;

  DFF \n_reg[0]  ( .D(n244), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n243), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n242), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n241), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n240), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n239), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n238), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \n_reg[7]  ( .D(n237), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[7]) );
  DFF \n_reg[8]  ( .D(n236), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[8]) );
  DFF \n_reg[9]  ( .D(n235), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[9]) );
  DFF \Y0_reg[0]  ( .D(n234), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n233), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n232), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n231), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n230), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n229), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n228), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n227), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y0_reg[8]  ( .D(n226), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[8]) );
  DFF \Y0_reg[9]  ( .D(n225), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[9]) );
  DFF \Y0_reg[10]  ( .D(n224), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[10]) );
  DFF \Y0_reg[11]  ( .D(n223), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[11]) );
  DFF \Y0_reg[12]  ( .D(n222), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[12]) );
  DFF \Y0_reg[13]  ( .D(n221), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[13]) );
  DFF \Y0_reg[14]  ( .D(n220), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[14]) );
  DFF \Y0_reg[15]  ( .D(n219), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[15]) );
  DFF \Y_reg[15]  ( .D(n218), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[15]) );
  DFF \Y_reg[14]  ( .D(n217), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[14]) );
  DFF \Y_reg[13]  ( .D(n216), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[13]) );
  DFF \Y_reg[12]  ( .D(n215), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[12]) );
  DFF \Y_reg[11]  ( .D(n214), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[11]) );
  DFF \Y_reg[10]  ( .D(n213), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[10]) );
  DFF \Y_reg[9]  ( .D(n212), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[9]) );
  DFF \Y_reg[8]  ( .D(n211), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[8]) );
  DFF \Y_reg[7]  ( .D(n210), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n209), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n208), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n207), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n206), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n205), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n204), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n203), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  HADDER \add_25/U1_1_6  ( .IN0(n[6]), .IN1(\add_25/carry[6] ), .COUT(
        \add_25/carry[7] ), .SUM(N13) );
  HADDER \add_25/U1_1_7  ( .IN0(n[7]), .IN1(\add_25/carry[7] ), .COUT(
        \add_25/carry[8] ), .SUM(N14) );
  HADDER \add_25/U1_1_8  ( .IN0(n[8]), .IN1(\add_25/carry[8] ), .COUT(
        \add_25/carry[9] ), .SUM(N15) );
  MUX U247 ( .IN0(n245), .IN1(n1561), .SEL(n1562), .F(n1545) );
  IV U248 ( .A(n1563), .Z(n245) );
  MUX U249 ( .IN0(n246), .IN1(n1228), .SEL(n1229), .F(n1205) );
  IV U250 ( .A(n1230), .Z(n246) );
  MUX U251 ( .IN0(n1636), .IN1(n1654), .SEL(n1638), .F(n1617) );
  XOR U252 ( .A(n1419), .B(n1409), .Z(n1225) );
  XOR U253 ( .A(n1231), .B(n1213), .Z(n1217) );
  MUX U254 ( .IN0(n247), .IN1(n978), .SEL(n979), .F(n908) );
  IV U255 ( .A(n980), .Z(n247) );
  MUX U256 ( .IN0(n248), .IN1(n1139), .SEL(n1140), .F(n1064) );
  IV U257 ( .A(n1141), .Z(n248) );
  MUX U258 ( .IN0(n249), .IN1(n1205), .SEL(n1206), .F(n1182) );
  IV U259 ( .A(n1207), .Z(n249) );
  MUX U260 ( .IN0(n250), .IN1(n1401), .SEL(n1402), .F(n1391) );
  IV U261 ( .A(n1403), .Z(n250) );
  XOR U262 ( .A(n1404), .B(n1396), .Z(n1202) );
  MUX U263 ( .IN0(n1356), .IN1(n1359), .SEL(n1357), .F(n1341) );
  MUX U264 ( .IN0(n251), .IN1(n703), .SEL(n704), .F(n652) );
  IV U265 ( .A(n705), .Z(n251) );
  MUX U266 ( .IN0(n252), .IN1(n1055), .SEL(n1056), .F(n978) );
  IV U267 ( .A(n1057), .Z(n252) );
  XNOR U268 ( .A(n1699), .B(n1700), .Z(n1143) );
  XOR U269 ( .A(n1206), .B(n1207), .Z(n1218) );
  MUX U270 ( .IN0(n253), .IN1(n1155), .SEL(n1156), .F(n1093) );
  IV U271 ( .A(n1157), .Z(n253) );
  XOR U272 ( .A(n1392), .B(n1393), .Z(n1200) );
  MUX U273 ( .IN0(n254), .IN1(n832), .SEL(n833), .F(n767) );
  IV U274 ( .A(n834), .Z(n254) );
  MUX U275 ( .IN0(X[8]), .IN1(n1684), .SEL(X[15]), .F(n715) );
  MUX U276 ( .IN0(n1397), .IN1(n255), .SEL(n1396), .F(n1388) );
  IV U277 ( .A(n1395), .Z(n255) );
  MUX U278 ( .IN0(X[13]), .IN1(n1710), .SEL(X[15]), .F(n497) );
  MUX U279 ( .IN0(n1572), .IN1(n1575), .SEL(n1573), .F(n1556) );
  MUX U280 ( .IN0(n256), .IN1(n1182), .SEL(n1183), .F(n1163) );
  IV U281 ( .A(n1184), .Z(n256) );
  MUX U282 ( .IN0(n257), .IN1(n1391), .SEL(n1392), .F(n1170) );
  IV U283 ( .A(n1393), .Z(n257) );
  XOR U284 ( .A(n1208), .B(n1190), .Z(n1194) );
  MUX U285 ( .IN0(X[9]), .IN1(n1685), .SEL(X[15]), .F(n661) );
  MUX U286 ( .IN0(n538), .IN1(n258), .SEL(n537), .F(n499) );
  IV U287 ( .A(n536), .Z(n258) );
  MUX U288 ( .IN0(X[11]), .IN1(n1665), .SEL(X[15]), .F(n567) );
  MUX U289 ( .IN0(n628), .IN1(n626), .SEL(n627), .F(n581) );
  MUX U290 ( .IN0(n259), .IN1(n421), .SEL(n420), .F(n429) );
  IV U291 ( .A(n432), .Z(n259) );
  MUX U292 ( .IN0(n260), .IN1(n1576), .SEL(n1577), .F(n1572) );
  IV U293 ( .A(n1578), .Z(n260) );
  XOR U294 ( .A(n1402), .B(n1403), .Z(n1223) );
  MUX U295 ( .IN0(n261), .IN1(n959), .SEL(n960), .F(n890) );
  IV U296 ( .A(n961), .Z(n261) );
  MUX U297 ( .IN0(n262), .IN1(n1018), .SEL(n1019), .F(n955) );
  IV U298 ( .A(n1020), .Z(n262) );
  MUX U299 ( .IN0(X[10]), .IN1(n1664), .SEL(X[15]), .F(n608) );
  MUX U300 ( .IN0(n718), .IN1(n263), .SEL(n717), .F(n663) );
  IV U301 ( .A(n716), .Z(n263) );
  MUX U302 ( .IN0(n794), .IN1(n792), .SEL(n793), .F(n727) );
  XNOR U303 ( .A(n1686), .B(n1140), .Z(n1144) );
  XOR U304 ( .A(n430), .B(n451), .Z(n449) );
  MUX U305 ( .IN0(n1617), .IN1(n1635), .SEL(n1619), .F(n1586) );
  MUX U306 ( .IN0(n1505), .IN1(n1527), .SEL(n1507), .F(n1487) );
  MUX U307 ( .IN0(n264), .IN1(n1163), .SEL(n1164), .F(n1101) );
  IV U308 ( .A(n1165), .Z(n264) );
  MUX U309 ( .IN0(n265), .IN1(n1408), .SEL(n1409), .F(n1395) );
  IV U310 ( .A(n1410), .Z(n265) );
  MUX U311 ( .IN0(n266), .IN1(n1130), .SEL(n1131), .F(n1055) );
  IV U312 ( .A(n1132), .Z(n266) );
  MUX U313 ( .IN0(A[11]), .IN1(n1439), .SEL(A[15]), .F(n584) );
  MUX U314 ( .IN0(n666), .IN1(n271), .SEL(n665), .F(n615) );
  MUX U315 ( .IN0(n927), .IN1(n925), .SEL(n926), .F(n857) );
  MUX U316 ( .IN0(n957), .IN1(n267), .SEL(n956), .F(n885) );
  IV U317 ( .A(n955), .Z(n267) );
  NAND U318 ( .A(n499), .B(n534), .Z(n533) );
  XOR U319 ( .A(n477), .B(n485), .Z(n483) );
  MUX U320 ( .IN0(n268), .IN1(n1423), .SEL(n1424), .F(n1408) );
  IV U321 ( .A(n1425), .Z(n268) );
  MUX U322 ( .IN0(n269), .IN1(n970), .SEL(n971), .F(n900) );
  IV U323 ( .A(n972), .Z(n269) );
  MUX U324 ( .IN0(n270), .IN1(n1026), .SEL(n1027), .F(n959) );
  IV U325 ( .A(n1028), .Z(n270) );
  MUX U326 ( .IN0(X[4]), .IN1(n1370), .SEL(X[15]), .F(n954) );
  XOR U327 ( .A(n1666), .B(n1651), .Z(n1591) );
  MUX U328 ( .IN0(n710), .IN1(n712), .SEL(n711), .F(n271) );
  IV U329 ( .A(n271), .Z(n664) );
  MUX U330 ( .IN0(n888), .IN1(n272), .SEL(n887), .F(n815) );
  IV U331 ( .A(n886), .Z(n272) );
  MUX U332 ( .IN0(n995), .IN1(n993), .SEL(n994), .F(n925) );
  MUX U333 ( .IN0(n1113), .IN1(n273), .SEL(n1112), .F(n1036) );
  IV U334 ( .A(n1111), .Z(n273) );
  XNOR U335 ( .A(n618), .B(n578), .Z(n582) );
  XOR U336 ( .A(n508), .B(n516), .Z(n514) );
  XOR U337 ( .A(n1183), .B(n1184), .Z(n1195) );
  MUX U338 ( .IN0(n1511), .IN1(n1521), .SEL(n1513), .F(n1497) );
  MUX U339 ( .IN0(n1586), .IN1(n1616), .SEL(n1588), .F(n1122) );
  XNOR U340 ( .A(n1363), .B(n1364), .Z(n1347) );
  MUX U341 ( .IN0(A[9]), .IN1(n1477), .SEL(A[15]), .F(n678) );
  MUX U342 ( .IN0(A[12]), .IN1(n1421), .SEL(A[15]), .F(n539) );
  XOR U343 ( .A(n587), .B(n630), .Z(n588) );
  MUX U344 ( .IN0(n982), .IN1(n984), .SEL(n983), .F(n914) );
  MUX U345 ( .IN0(n1024), .IN1(n1022), .SEL(n1023), .F(n949) );
  XOR U346 ( .A(n1112), .B(n1113), .Z(n1119) );
  XNOR U347 ( .A(n615), .B(n658), .Z(n616) );
  XNOR U348 ( .A(n719), .B(n672), .Z(n676) );
  MUX U349 ( .IN0(n274), .IN1(n903), .SEL(n904), .F(n835) );
  IV U350 ( .A(n905), .Z(n274) );
  MUX U351 ( .IN0(n762), .IN1(n764), .SEL(n763), .F(n275) );
  IV U352 ( .A(n275), .Z(n698) );
  XOR U353 ( .A(n545), .B(n553), .Z(n551) );
  MUX U354 ( .IN0(n1503), .IN1(n276), .SEL(n1353), .F(n1484) );
  IV U355 ( .A(n1352), .Z(n276) );
  MUX U356 ( .IN0(n1349), .IN1(n1347), .SEL(n1348), .F(n1320) );
  XOR U357 ( .A(n1394), .B(n1388), .Z(n1179) );
  MUX U358 ( .IN0(n277), .IN1(n1122), .SEL(n1123), .F(n1047) );
  IV U359 ( .A(n1124), .Z(n277) );
  MUX U360 ( .IN0(n278), .IN1(n1170), .SEL(n1171), .F(n1111) );
  IV U361 ( .A(n1172), .Z(n278) );
  XOR U362 ( .A(n1185), .B(n1156), .Z(n1160) );
  MUX U363 ( .IN0(n846), .IN1(n848), .SEL(n847), .F(n781) );
  MUX U364 ( .IN0(n1072), .IN1(n1070), .SEL(n1071), .F(n993) );
  XOR U365 ( .A(n1592), .B(n1131), .Z(n1135) );
  XNOR U366 ( .A(n667), .B(n623), .Z(n627) );
  MUX U367 ( .IN0(n279), .IN1(n706), .SEL(n707), .F(n655) );
  IV U368 ( .A(n708), .Z(n279) );
  MUX U369 ( .IN0(n280), .IN1(n821), .SEL(n822), .F(n761) );
  IV U370 ( .A(n823), .Z(n280) );
  NAND U371 ( .A(n885), .B(n953), .Z(n952) );
  MUX U372 ( .IN0(n827), .IN1(n829), .SEL(n828), .F(n762) );
  MUX U373 ( .IN0(n281), .IN1(n801), .SEL(n802), .F(n736) );
  IV U374 ( .A(Y0[5]), .Z(n281) );
  XOR U375 ( .A(n590), .B(n598), .Z(n596) );
  MUX U376 ( .IN0(n282), .IN1(n1556), .SEL(n1557), .F(n1539) );
  IV U377 ( .A(n1558), .Z(n282) );
  MUX U378 ( .IN0(A[1]), .IN1(n1712), .SEL(A[15]), .F(n1366) );
  MUX U379 ( .IN0(n283), .IN1(n767), .SEL(n768), .F(n703) );
  IV U380 ( .A(n769), .Z(n283) );
  MUX U381 ( .IN0(A[6]), .IN1(n1608), .SEL(A[15]), .F(n860) );
  MUX U382 ( .IN0(A[7]), .IN1(n1595), .SEL(A[15]), .F(n795) );
  MUX U383 ( .IN0(A[5]), .IN1(n1628), .SEL(A[15]), .F(n928) );
  MUX U384 ( .IN0(n284), .IN1(n1101), .SEL(n1102), .F(n1026) );
  IV U385 ( .A(n1103), .Z(n284) );
  XOR U386 ( .A(n1171), .B(n1172), .Z(n1177) );
  MUX U387 ( .IN0(n914), .IN1(n916), .SEL(n915), .F(n846) );
  XNOR U388 ( .A(n1153), .B(n1094), .Z(n1098) );
  XOR U389 ( .A(n505), .B(n540), .Z(n506) );
  MUX U390 ( .IN0(n285), .IN1(n570), .SEL(n571), .F(n523) );
  IV U391 ( .A(n572), .Z(n285) );
  NAND U392 ( .A(n663), .B(n714), .Z(n713) );
  MUX U393 ( .IN0(n817), .IN1(n815), .SEL(n816), .F(n759) );
  XNOR U394 ( .A(n849), .B(n789), .Z(n793) );
  MUX U395 ( .IN0(n286), .IN1(n1050), .SEL(n1051), .F(n973) );
  IV U396 ( .A(n1052), .Z(n286) );
  MUX U397 ( .IN0(n287), .IN1(n897), .SEL(n896), .F(n827) );
  IV U398 ( .A(n895), .Z(n287) );
  MUX U399 ( .IN0(n288), .IN1(n866), .SEL(n867), .F(n801) );
  IV U400 ( .A(Y0[4]), .Z(n288) );
  XOR U401 ( .A(n635), .B(n643), .Z(n641) );
  MUX U402 ( .IN0(n1320), .IN1(n289), .SEL(n1321), .F(n1293) );
  IV U403 ( .A(n1322), .Z(n289) );
  MUX U404 ( .IN0(n1412), .IN1(n290), .SEL(n1225), .F(n1399) );
  IV U405 ( .A(n1223), .Z(n290) );
  XNOR U406 ( .A(n1577), .B(n1578), .Z(n1564) );
  MUX U407 ( .IN0(n291), .IN1(n900), .SEL(n901), .F(n832) );
  IV U408 ( .A(n902), .Z(n291) );
  MUX U409 ( .IN0(A[3]), .IN1(n1689), .SEL(A[15]), .F(n292) );
  IV U410 ( .A(n292), .Z(n1073) );
  MUX U411 ( .IN0(A[4]), .IN1(n1646), .SEL(A[15]), .F(n293) );
  IV U412 ( .A(n293), .Z(n996) );
  MUX U413 ( .IN0(n1159), .IN1(n294), .SEL(n1160), .F(n1097) );
  IV U414 ( .A(n1161), .Z(n294) );
  XOR U415 ( .A(n1490), .B(n1491), .Z(n1352) );
  MUX U416 ( .IN0(n583), .IN1(n581), .SEL(n582), .F(n528) );
  MUX U417 ( .IN0(n295), .IN1(n890), .SEL(n891), .F(n821) );
  IV U418 ( .A(n892), .Z(n295) );
  XOR U419 ( .A(n798), .B(n861), .Z(n799) );
  MUX U420 ( .IN0(n1059), .IN1(n1061), .SEL(n1060), .F(n982) );
  MUX U421 ( .IN0(n1145), .IN1(n1143), .SEL(n1144), .F(n1070) );
  MUX U422 ( .IN0(n296), .IN1(n612), .SEL(n613), .F(n570) );
  IV U423 ( .A(n614), .Z(n296) );
  XOR U424 ( .A(n773), .B(n717), .Z(n711) );
  XNOR U425 ( .A(n784), .B(n724), .Z(n728) );
  MUX U426 ( .IN0(n297), .IN1(n835), .SEL(n836), .F(n770) );
  IV U427 ( .A(n837), .Z(n297) );
  XOR U428 ( .A(n948), .B(n886), .Z(n887) );
  MUX U429 ( .IN0(n1044), .IN1(n298), .SEL(n1043), .F(n965) );
  IV U430 ( .A(n1042), .Z(n298) );
  MUX U431 ( .IN0(n962), .IN1(n299), .SEL(n963), .F(n895) );
  IV U432 ( .A(n964), .Z(n299) );
  MUX U433 ( .IN0(n300), .IN1(n934), .SEL(n935), .F(n866) );
  IV U434 ( .A(Y0[3]), .Z(n300) );
  XOR U435 ( .A(n690), .B(n696), .Z(n685) );
  MUX U436 ( .IN0(n301), .IN1(n1350), .SEL(n1167), .F(n1323) );
  IV U437 ( .A(n1166), .Z(n301) );
  MUX U438 ( .IN0(n1266), .IN1(n302), .SEL(n1267), .F(n1239) );
  IV U439 ( .A(n1268), .Z(n302) );
  MUX U440 ( .IN0(X[1]), .IN1(n303), .SEL(X[15]), .F(n1383) );
  IV U441 ( .A(n1583), .Z(n303) );
  MUX U442 ( .IN0(X[6]), .IN1(n1375), .SEL(X[15]), .F(n820) );
  MUX U443 ( .IN0(X[3]), .IN1(n1569), .SEL(X[15]), .F(n1039) );
  MUX U444 ( .IN0(n1134), .IN1(n1136), .SEL(n1135), .F(n1059) );
  MUX U445 ( .IN0(X[14]), .IN1(n1715), .SEL(X[15]), .F(n466) );
  NAND U446 ( .A(n564), .B(n607), .Z(n606) );
  XOR U447 ( .A(n838), .B(n778), .Z(n782) );
  XNOR U448 ( .A(n917), .B(n854), .Z(n858) );
  MUX U449 ( .IN0(n304), .IN1(n973), .SEL(n974), .F(n903) );
  IV U450 ( .A(n975), .Z(n304) );
  XNOR U451 ( .A(n1016), .B(n956), .Z(n950) );
  MUX U452 ( .IN0(n1029), .IN1(n305), .SEL(n1030), .F(n962) );
  IV U453 ( .A(n1031), .Z(n305) );
  MUX U454 ( .IN0(n306), .IN1(n508), .SEL(n509), .F(n477) );
  IV U455 ( .A(Y0[11]), .Z(n306) );
  XOR U456 ( .A(n736), .B(n744), .Z(n742) );
  MUX U457 ( .IN0(n1484), .IN1(n307), .SEL(n1329), .F(n1465) );
  IV U458 ( .A(n1327), .Z(n307) );
  MUX U459 ( .IN0(n1539), .IN1(n1555), .SEL(n1541), .F(n1522) );
  MUX U460 ( .IN0(n1216), .IN1(n308), .SEL(n1217), .F(n1193) );
  IV U461 ( .A(n1218), .Z(n308) );
  XOR U462 ( .A(n1164), .B(n1165), .Z(n1161) );
  XOR U463 ( .A(n1562), .B(n1563), .Z(n1377) );
  MUX U464 ( .IN0(n309), .IN1(n1047), .SEL(n1048), .F(n970) );
  IV U465 ( .A(n1049), .Z(n309) );
  MUX U466 ( .IN0(A[10]), .IN1(n1457), .SEL(A[15]), .F(n629) );
  XNOR U467 ( .A(n1354), .B(n1344), .Z(n1348) );
  XOR U468 ( .A(n681), .B(n731), .Z(n682) );
  MUX U469 ( .IN0(n729), .IN1(n727), .SEL(n728), .F(n675) );
  MUX U470 ( .IN0(n951), .IN1(n949), .SEL(n950), .F(n886) );
  MUX U471 ( .IN0(A[13]), .IN1(n1407), .SEL(A[15]), .F(n502) );
  MUX U472 ( .IN0(n310), .IN1(n770), .SEL(n771), .F(n706) );
  IV U473 ( .A(n772), .Z(n310) );
  XOR U474 ( .A(n906), .B(n843), .Z(n847) );
  XNOR U475 ( .A(n1062), .B(n990), .Z(n994) );
  MUX U476 ( .IN0(n311), .IN1(n1125), .SEL(n1126), .F(n1050) );
  IV U477 ( .A(n1127), .Z(n311) );
  MUX U478 ( .IN0(n312), .IN1(n1114), .SEL(n1115), .F(n1042) );
  IV U479 ( .A(n1116), .Z(n312) );
  MUX U480 ( .IN0(A[14]), .IN1(n1384), .SEL(A[15]), .F(n467) );
  MUX U481 ( .IN0(n525), .IN1(n313), .SEL(n524), .F(n493) );
  IV U482 ( .A(n523), .Z(n313) );
  XNOR U483 ( .A(n827), .B(n826), .Z(n879) );
  MUX U484 ( .IN0(Y0[13]), .IN1(n314), .SEL(n431), .F(n423) );
  IV U485 ( .A(n430), .Z(n314) );
  MUX U486 ( .IN0(n315), .IN1(n590), .SEL(n591), .F(n545) );
  IV U487 ( .A(Y0[9]), .Z(n315) );
  MUX U488 ( .IN0(n316), .IN1(n1079), .SEL(n1080), .F(n1002) );
  IV U489 ( .A(Y0[1]), .Z(n316) );
  XOR U490 ( .A(n801), .B(n809), .Z(n807) );
  MUX U491 ( .IN0(n1465), .IN1(n317), .SEL(n1302), .F(n1446) );
  IV U492 ( .A(n1300), .Z(n317) );
  MUX U493 ( .IN0(n1239), .IN1(n318), .SEL(n1240), .F(n1216) );
  IV U494 ( .A(n1241), .Z(n318) );
  MUX U495 ( .IN0(n1522), .IN1(n1538), .SEL(n1524), .F(n1511) );
  MUX U496 ( .IN0(n1399), .IN1(n319), .SEL(n1202), .F(n1389) );
  IV U497 ( .A(n1200), .Z(n319) );
  MUX U498 ( .IN0(A[8]), .IN1(n1495), .SEL(A[15]), .F(n730) );
  MUX U499 ( .IN0(A[2]), .IN1(n1702), .SEL(A[15]), .F(n1146) );
  MUX U500 ( .IN0(n320), .IN1(n1093), .SEL(n1094), .F(n1018) );
  IV U501 ( .A(n1095), .Z(n320) );
  MUX U502 ( .IN0(n321), .IN1(n652), .SEL(n653), .F(n609) );
  IV U503 ( .A(n654), .Z(n321) );
  MUX U504 ( .IN0(n781), .IN1(n783), .SEL(n782), .F(n710) );
  MUX U505 ( .IN0(n859), .IN1(n857), .SEL(n858), .F(n792) );
  XOR U506 ( .A(n1076), .B(n1147), .Z(n1077) );
  MUX U507 ( .IN0(n1099), .IN1(n1097), .SEL(n1098), .F(n1022) );
  XNOR U508 ( .A(n528), .B(n529), .Z(n527) );
  MUX U509 ( .IN0(n322), .IN1(n655), .SEL(n656), .F(n612) );
  IV U510 ( .A(n657), .Z(n322) );
  XOR U511 ( .A(n822), .B(n823), .Z(n817) );
  XOR U512 ( .A(n1053), .B(n979), .Z(n983) );
  XNOR U513 ( .A(n1137), .B(n1067), .Z(n1071) );
  NAND U514 ( .A(n1036), .B(n1109), .Z(n1108) );
  XNOR U515 ( .A(n532), .B(n531), .Z(n525) );
  XNOR U516 ( .A(n927), .B(n926), .Z(n905) );
  MUX U517 ( .IN0(n967), .IN1(n965), .SEL(n966), .F(n323) );
  IV U518 ( .A(n323), .Z(n894) );
  MUX U519 ( .IN0(n1104), .IN1(n324), .SEL(n1105), .F(n1029) );
  IV U520 ( .A(n1106), .Z(n324) );
  MUX U521 ( .IN0(n698), .IN1(n325), .SEL(n699), .F(n649) );
  IV U522 ( .A(n700), .Z(n325) );
  MUX U523 ( .IN0(n326), .IN1(n477), .SEL(n478), .F(n430) );
  IV U524 ( .A(Y0[12]), .Z(n326) );
  MUX U525 ( .IN0(n327), .IN1(n635), .SEL(n636), .F(n590) );
  IV U526 ( .A(Y0[8]), .Z(n327) );
  XOR U527 ( .A(n866), .B(n874), .Z(n872) );
  MUX U528 ( .IN0(n1446), .IN1(n328), .SEL(n1275), .F(n1427) );
  IV U529 ( .A(n1273), .Z(n328) );
  MUX U530 ( .IN0(n329), .IN1(n1590), .SEL(n1591), .F(n1640) );
  IV U531 ( .A(n1660), .Z(n329) );
  NOR U532 ( .A(A[0]), .B(n1712), .Z(n1703) );
  XOR U533 ( .A(n1570), .B(n1557), .Z(n1378) );
  MUX U534 ( .IN0(n1389), .IN1(n330), .SEL(n1179), .F(n1117) );
  IV U535 ( .A(n1177), .Z(n330) );
  MUX U536 ( .IN0(n677), .IN1(n675), .SEL(n676), .F(n626) );
  XOR U537 ( .A(n931), .B(n997), .Z(n932) );
  MUX U538 ( .IN0(n611), .IN1(n331), .SEL(n610), .F(n564) );
  IV U539 ( .A(n609), .Z(n331) );
  MUX U540 ( .IN0(X[7]), .IN1(n1376), .SEL(X[15]), .F(n753) );
  XNOR U541 ( .A(n985), .B(n922), .Z(n926) );
  XOR U542 ( .A(n976), .B(n911), .Z(n915) );
  XNOR U543 ( .A(n1091), .B(n1019), .Z(n1023) );
  XNOR U544 ( .A(n1145), .B(n1144), .Z(n1127) );
  MUX U545 ( .IN0(n501), .IN1(n527), .SEL(n500), .F(n472) );
  XNOR U546 ( .A(n583), .B(n582), .Z(n572) );
  XNOR U547 ( .A(n794), .B(n793), .Z(n772) );
  XNOR U548 ( .A(n859), .B(n858), .Z(n837) );
  XNOR U549 ( .A(n965), .B(n1032), .Z(n966) );
  XNOR U550 ( .A(n708), .B(n707), .Z(n700) );
  XOR U551 ( .A(n814), .B(n755), .Z(n763) );
  XNOR U552 ( .A(n975), .B(n974), .Z(n964) );
  XNOR U553 ( .A(n1052), .B(n1051), .Z(n1031) );
  XNOR U554 ( .A(n491), .B(n490), .Z(n515) );
  MUX U555 ( .IN0(n332), .IN1(n684), .SEL(n685), .F(n635) );
  IV U556 ( .A(Y0[7]), .Z(n332) );
  MUX U557 ( .IN0(Y0[14]), .IN1(n423), .SEL(n424), .F(n413) );
  XOR U558 ( .A(n934), .B(n942), .Z(n940) );
  MUX U559 ( .IN0(n1293), .IN1(n333), .SEL(n1294), .F(n1266) );
  IV U560 ( .A(n1295), .Z(n333) );
  MUX U561 ( .IN0(n334), .IN1(n1377), .SEL(n1378), .F(n1550) );
  IV U562 ( .A(n1564), .Z(n334) );
  MUX U563 ( .IN0(n1427), .IN1(n335), .SEL(n1248), .F(n1412) );
  IV U564 ( .A(n1246), .Z(n335) );
  XOR U565 ( .A(n1688), .B(A[3]), .Z(n1689) );
  MUX U566 ( .IN0(n1193), .IN1(n336), .SEL(n1194), .F(n1159) );
  IV U567 ( .A(n1195), .Z(n336) );
  XOR U568 ( .A(n1658), .B(n1659), .Z(n1590) );
  XOR U569 ( .A(n1509), .B(n1500), .Z(n1353) );
  MUX U570 ( .IN0(X[5]), .IN1(n1371), .SEL(X[15]), .F(n883) );
  MUX U571 ( .IN0(X[2]), .IN1(n1568), .SEL(X[15]), .F(n1110) );
  XNOR U572 ( .A(n1349), .B(n1348), .Z(n1166) );
  XNOR U573 ( .A(n573), .B(n537), .Z(n531) );
  MUX U574 ( .IN0(n617), .IN1(n615), .SEL(n616), .F(n337) );
  IV U575 ( .A(n337), .Z(n569) );
  XOR U576 ( .A(n891), .B(n892), .Z(n888) );
  XOR U577 ( .A(n1128), .B(n1056), .Z(n1060) );
  MUX U578 ( .IN0(n1119), .IN1(n1379), .SEL(n1118), .F(n1041) );
  XNOR U579 ( .A(n1099), .B(n1098), .Z(n1116) );
  AND U580 ( .A(n461), .B(n438), .Z(n460) );
  XNOR U581 ( .A(n628), .B(n627), .Z(n614) );
  XNOR U582 ( .A(n677), .B(n676), .Z(n657) );
  XNOR U583 ( .A(n729), .B(n728), .Z(n708) );
  XNOR U584 ( .A(n951), .B(n950), .Z(n967) );
  XNOR U585 ( .A(n995), .B(n994), .Z(n975) );
  XNOR U586 ( .A(n1072), .B(n1071), .Z(n1052) );
  XNOR U587 ( .A(n1024), .B(n1023), .Z(n1044) );
  XNOR U588 ( .A(n1127), .B(n1126), .Z(n1106) );
  XNOR U589 ( .A(n492), .B(n493), .Z(n491) );
  XNOR U590 ( .A(n772), .B(n771), .Z(n764) );
  XNOR U591 ( .A(n837), .B(n836), .Z(n829) );
  XNOR U592 ( .A(n905), .B(n904), .Z(n897) );
  MUX U593 ( .IN0(n338), .IN1(n545), .SEL(n546), .F(n508) );
  IV U594 ( .A(Y0[10]), .Z(n338) );
  MUX U595 ( .IN0(n339), .IN1(n736), .SEL(n737), .F(n684) );
  IV U596 ( .A(Y0[6]), .Z(n339) );
  MUX U597 ( .IN0(n340), .IN1(n1002), .SEL(n1003), .F(n934) );
  IV U598 ( .A(Y0[2]), .Z(n340) );
  MUX U599 ( .IN0(Y0[15]), .IN1(n413), .SEL(n414), .F(n341) );
  IV U600 ( .A(n341), .Z(n410) );
  XOR U601 ( .A(n1080), .B(Y0[1]), .Z(n355) );
  ANDN U602 ( .A(n342), .B(n[0]), .Z(n244) );
  AND U603 ( .A(N8), .B(n342), .Z(n243) );
  AND U604 ( .A(N9), .B(n342), .Z(n242) );
  AND U605 ( .A(N10), .B(n342), .Z(n241) );
  AND U606 ( .A(N11), .B(n342), .Z(n240) );
  AND U607 ( .A(N12), .B(n342), .Z(n239) );
  AND U608 ( .A(N13), .B(n342), .Z(n238) );
  AND U609 ( .A(N14), .B(n342), .Z(n237) );
  AND U610 ( .A(N15), .B(n342), .Z(n236) );
  AND U611 ( .A(n342), .B(n343), .Z(n235) );
  XOR U612 ( .A(n[9]), .B(\add_25/carry[9] ), .Z(n343) );
  ANDN U613 ( .A(n344), .B(rst), .Z(n342) );
  NAND U614 ( .A(n345), .B(n346), .Z(n344) );
  AND U615 ( .A(n347), .B(n348), .Z(n346) );
  AND U616 ( .A(n[1]), .B(n349), .Z(n348) );
  ANDN U617 ( .A(n[0]), .B(n350), .Z(n349) );
  AND U618 ( .A(n[5]), .B(n[2]), .Z(n347) );
  AND U619 ( .A(n351), .B(n352), .Z(n345) );
  AND U620 ( .A(n[7]), .B(n[6]), .Z(n352) );
  AND U621 ( .A(n[8]), .B(n[9]), .Z(n351) );
  NAND U622 ( .A(n353), .B(n354), .Z(n234) );
  OR U623 ( .A(n355), .B(n356), .Z(n354) );
  NANDN U624 ( .B(n357), .A(Y0[0]), .Z(n353) );
  NAND U625 ( .A(n358), .B(n359), .Z(n233) );
  NANDN U626 ( .B(n356), .A(n360), .Z(n359) );
  NANDN U627 ( .B(n361), .A(rst), .Z(n358) );
  NAND U628 ( .A(n362), .B(n363), .Z(n232) );
  NANDN U629 ( .B(n356), .A(n364), .Z(n363) );
  NANDN U630 ( .B(n357), .A(Y0[2]), .Z(n362) );
  NAND U631 ( .A(n365), .B(n366), .Z(n231) );
  NANDN U632 ( .B(n356), .A(n367), .Z(n366) );
  NANDN U633 ( .B(n357), .A(Y0[3]), .Z(n365) );
  NAND U634 ( .A(n368), .B(n369), .Z(n230) );
  NANDN U635 ( .B(n356), .A(n370), .Z(n369) );
  NANDN U636 ( .B(n357), .A(Y0[4]), .Z(n368) );
  NAND U637 ( .A(n371), .B(n372), .Z(n229) );
  NANDN U638 ( .B(n356), .A(n373), .Z(n372) );
  NANDN U639 ( .B(n357), .A(Y0[5]), .Z(n371) );
  NAND U640 ( .A(n374), .B(n375), .Z(n228) );
  NANDN U641 ( .B(n356), .A(n376), .Z(n375) );
  NANDN U642 ( .B(n357), .A(Y0[6]), .Z(n374) );
  NAND U643 ( .A(n377), .B(n378), .Z(n227) );
  NANDN U644 ( .B(n356), .A(n379), .Z(n378) );
  NANDN U645 ( .B(n357), .A(Y0[7]), .Z(n377) );
  NAND U646 ( .A(n380), .B(n381), .Z(n226) );
  NANDN U647 ( .B(n356), .A(n382), .Z(n381) );
  NANDN U648 ( .B(n357), .A(Y0[8]), .Z(n380) );
  NAND U649 ( .A(n383), .B(n384), .Z(n225) );
  NANDN U650 ( .B(n356), .A(n385), .Z(n384) );
  NANDN U651 ( .B(n357), .A(Y0[9]), .Z(n383) );
  NAND U652 ( .A(n386), .B(n387), .Z(n224) );
  NANDN U653 ( .B(n356), .A(n388), .Z(n387) );
  NANDN U654 ( .B(n357), .A(Y0[10]), .Z(n386) );
  NAND U655 ( .A(n389), .B(n390), .Z(n223) );
  NANDN U656 ( .B(n356), .A(n391), .Z(n390) );
  NANDN U657 ( .B(n357), .A(Y0[11]), .Z(n389) );
  NAND U658 ( .A(n392), .B(n393), .Z(n222) );
  NANDN U659 ( .B(n356), .A(n394), .Z(n393) );
  NANDN U660 ( .B(n357), .A(Y0[12]), .Z(n392) );
  NAND U661 ( .A(n395), .B(n396), .Z(n221) );
  NANDN U662 ( .B(n356), .A(n397), .Z(n396) );
  NANDN U663 ( .B(n357), .A(Y0[13]), .Z(n395) );
  NAND U664 ( .A(n398), .B(n399), .Z(n220) );
  OR U665 ( .A(n400), .B(n356), .Z(n399) );
  NANDN U666 ( .B(n357), .A(Y0[14]), .Z(n398) );
  NAND U667 ( .A(n401), .B(n402), .Z(n219) );
  OR U668 ( .A(n356), .B(n403), .Z(n402) );
  NANDN U669 ( .B(n404), .A(n357), .Z(n356) );
  NANDN U670 ( .B(n357), .A(Y0[15]), .Z(n401) );
  NAND U671 ( .A(n405), .B(n406), .Z(n218) );
  NANDN U672 ( .B(n357), .A(Y[15]), .Z(n406) );
  AND U673 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U674 ( .B(n404), .A(Y[15]), .Z(n408) );
  OR U675 ( .A(n403), .B(n409), .Z(n407) );
  XOR U676 ( .A(n410), .B(n411), .Z(n403) );
  XNOR U677 ( .A(Y0[15]), .B(n412), .Z(n411) );
  NAND U678 ( .A(n415), .B(n416), .Z(n217) );
  NANDN U679 ( .B(n357), .A(Y[14]), .Z(n416) );
  AND U680 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U681 ( .B(n404), .A(Y[14]), .Z(n418) );
  OR U682 ( .A(n400), .B(n409), .Z(n417) );
  XOR U683 ( .A(n414), .B(Y0[15]), .Z(n400) );
  XOR U684 ( .A(n413), .B(n412), .Z(n414) );
  NAND U685 ( .A(n419), .B(n420), .Z(n412) );
  OR U686 ( .A(n421), .B(n422), .Z(n419) );
  NAND U687 ( .A(n425), .B(n426), .Z(n216) );
  NANDN U688 ( .B(n357), .A(Y[13]), .Z(n426) );
  AND U689 ( .A(n427), .B(n428), .Z(n425) );
  NANDN U690 ( .B(n404), .A(Y[13]), .Z(n428) );
  NANDN U691 ( .B(n409), .A(n397), .Z(n427) );
  XNOR U692 ( .A(n424), .B(Y0[14]), .Z(n397) );
  XNOR U693 ( .A(n429), .B(n423), .Z(n424) );
  XNOR U694 ( .A(n422), .B(n432), .Z(n421) );
  OR U695 ( .A(n433), .B(n434), .Z(n422) );
  AND U696 ( .A(n435), .B(n436), .Z(n432) );
  OR U697 ( .A(n437), .B(n438), .Z(n436) );
  AND U698 ( .A(n439), .B(n440), .Z(n435) );
  OR U699 ( .A(n441), .B(n442), .Z(n440) );
  OR U700 ( .A(n443), .B(n444), .Z(n439) );
  NAND U701 ( .A(n445), .B(n446), .Z(n215) );
  NANDN U702 ( .B(n357), .A(Y[12]), .Z(n446) );
  AND U703 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U704 ( .B(n404), .A(Y[12]), .Z(n448) );
  NANDN U705 ( .B(n409), .A(n394), .Z(n447) );
  XNOR U706 ( .A(n431), .B(Y0[13]), .Z(n394) );
  XNOR U707 ( .A(n449), .B(n450), .Z(n431) );
  AND U708 ( .A(n420), .B(n452), .Z(n451) );
  XOR U709 ( .A(n433), .B(n453), .Z(n452) );
  XOR U710 ( .A(n453), .B(n434), .Z(n433) );
  OR U711 ( .A(n454), .B(n455), .Z(n434) );
  IV U712 ( .A(n450), .Z(n453) );
  XNOR U713 ( .A(n444), .B(n443), .Z(n450) );
  OR U714 ( .A(n456), .B(n457), .Z(n443) );
  AND U715 ( .A(n458), .B(n459), .Z(n444) );
  XNOR U716 ( .A(n437), .B(n460), .Z(n459) );
  NAND U717 ( .A(n462), .B(n463), .Z(n438) );
  NANDN U718 ( .B(n464), .A(n465), .Z(n462) );
  NANDN U719 ( .B(n441), .A(n466), .Z(n461) );
  NANDN U720 ( .B(n442), .A(n467), .Z(n437) );
  AND U721 ( .A(n468), .B(n469), .Z(n458) );
  OR U722 ( .A(n470), .B(n471), .Z(n469) );
  XNOR U723 ( .A(n472), .B(n473), .Z(n468) );
  ANDN U724 ( .A(n474), .B(n475), .Z(n473) );
  XOR U725 ( .A(n472), .B(n476), .Z(n474) );
  NAND U726 ( .A(n479), .B(n480), .Z(n214) );
  NANDN U727 ( .B(n357), .A(Y[11]), .Z(n480) );
  AND U728 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U729 ( .B(n404), .A(Y[11]), .Z(n482) );
  NANDN U730 ( .B(n409), .A(n391), .Z(n481) );
  XNOR U731 ( .A(n478), .B(Y0[12]), .Z(n391) );
  XNOR U732 ( .A(n483), .B(n484), .Z(n478) );
  AND U733 ( .A(n420), .B(n486), .Z(n485) );
  XOR U734 ( .A(n454), .B(n487), .Z(n486) );
  XOR U735 ( .A(n487), .B(n455), .Z(n454) );
  OR U736 ( .A(n488), .B(n489), .Z(n455) );
  IV U737 ( .A(n484), .Z(n487) );
  XNOR U738 ( .A(n457), .B(n456), .Z(n484) );
  OR U739 ( .A(n490), .B(n491), .Z(n456) );
  XNOR U740 ( .A(n471), .B(n470), .Z(n457) );
  OR U741 ( .A(n492), .B(n493), .Z(n470) );
  XOR U742 ( .A(n476), .B(n475), .Z(n471) );
  XOR U743 ( .A(n472), .B(n494), .Z(n475) );
  AND U744 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U745 ( .B(n441), .A(n497), .Z(n496) );
  OR U746 ( .A(n498), .B(n499), .Z(n495) );
  XOR U747 ( .A(n464), .B(n465), .Z(n476) );
  NANDN U748 ( .B(n442), .A(n502), .Z(n465) );
  XNOR U749 ( .A(n463), .B(n503), .Z(n464) );
  AND U750 ( .A(n467), .B(n466), .Z(n503) );
  ANDN U751 ( .A(n504), .B(n505), .Z(n463) );
  NANDN U752 ( .B(n506), .A(n507), .Z(n504) );
  NAND U753 ( .A(n510), .B(n511), .Z(n213) );
  NANDN U754 ( .B(n357), .A(Y[10]), .Z(n511) );
  AND U755 ( .A(n512), .B(n513), .Z(n510) );
  NANDN U756 ( .B(n404), .A(Y[10]), .Z(n513) );
  NANDN U757 ( .B(n409), .A(n388), .Z(n512) );
  XNOR U758 ( .A(n509), .B(Y0[11]), .Z(n388) );
  XNOR U759 ( .A(n514), .B(n515), .Z(n509) );
  AND U760 ( .A(n420), .B(n517), .Z(n516) );
  XOR U761 ( .A(n488), .B(n518), .Z(n517) );
  XOR U762 ( .A(n518), .B(n489), .Z(n488) );
  OR U763 ( .A(n519), .B(n520), .Z(n489) );
  IV U764 ( .A(n515), .Z(n518) );
  OR U765 ( .A(n521), .B(n522), .Z(n490) );
  XOR U766 ( .A(n501), .B(n500), .Z(n492) );
  XNOR U767 ( .A(n526), .B(n527), .Z(n500) );
  ANDN U768 ( .A(n530), .B(n531), .Z(n529) );
  XOR U769 ( .A(n528), .B(n532), .Z(n530) );
  XNOR U770 ( .A(n533), .B(n498), .Z(n526) );
  NAND U771 ( .A(n497), .B(n467), .Z(n498) );
  NANDN U772 ( .B(n441), .A(n535), .Z(n534) );
  XOR U773 ( .A(n506), .B(n507), .Z(n501) );
  NANDN U774 ( .B(n442), .A(n539), .Z(n507) );
  AND U775 ( .A(n502), .B(n466), .Z(n540) );
  NAND U776 ( .A(n541), .B(n542), .Z(n505) );
  NANDN U777 ( .B(n543), .A(n544), .Z(n541) );
  NAND U778 ( .A(n547), .B(n548), .Z(n212) );
  NANDN U779 ( .B(n357), .A(Y[9]), .Z(n548) );
  AND U780 ( .A(n549), .B(n550), .Z(n547) );
  NANDN U781 ( .B(n404), .A(Y[9]), .Z(n550) );
  NANDN U782 ( .B(n409), .A(n385), .Z(n549) );
  XNOR U783 ( .A(n546), .B(Y0[10]), .Z(n385) );
  XNOR U784 ( .A(n551), .B(n552), .Z(n546) );
  AND U785 ( .A(n420), .B(n554), .Z(n553) );
  XOR U786 ( .A(n519), .B(n555), .Z(n554) );
  XOR U787 ( .A(n555), .B(n520), .Z(n519) );
  OR U788 ( .A(n556), .B(n557), .Z(n520) );
  IV U789 ( .A(n552), .Z(n555) );
  XNOR U790 ( .A(n522), .B(n521), .Z(n552) );
  OR U791 ( .A(n558), .B(n559), .Z(n521) );
  XNOR U792 ( .A(n525), .B(n524), .Z(n522) );
  XOR U793 ( .A(n523), .B(n560), .Z(n524) );
  AND U794 ( .A(n561), .B(n562), .Z(n560) );
  OR U795 ( .A(n563), .B(n564), .Z(n562) );
  AND U796 ( .A(n565), .B(n566), .Z(n561) );
  NANDN U797 ( .B(n441), .A(n567), .Z(n566) );
  NAND U798 ( .A(n568), .B(n569), .Z(n565) );
  XNOR U799 ( .A(n536), .B(n574), .Z(n537) );
  AND U800 ( .A(n467), .B(n535), .Z(n574) );
  XOR U801 ( .A(n575), .B(n576), .Z(n536) );
  ANDN U802 ( .A(n577), .B(n578), .Z(n576) );
  XNOR U803 ( .A(n579), .B(n575), .Z(n577) );
  XOR U804 ( .A(n580), .B(n538), .Z(n573) );
  NAND U805 ( .A(n497), .B(n502), .Z(n538) );
  IV U806 ( .A(n528), .Z(n580) );
  XNOR U807 ( .A(n543), .B(n544), .Z(n532) );
  NANDN U808 ( .B(n442), .A(n584), .Z(n544) );
  XNOR U809 ( .A(n542), .B(n585), .Z(n543) );
  AND U810 ( .A(n539), .B(n466), .Z(n585) );
  ANDN U811 ( .A(n586), .B(n587), .Z(n542) );
  NANDN U812 ( .B(n588), .A(n589), .Z(n586) );
  NAND U813 ( .A(n592), .B(n593), .Z(n211) );
  NANDN U814 ( .B(n357), .A(Y[8]), .Z(n593) );
  AND U815 ( .A(n594), .B(n595), .Z(n592) );
  NANDN U816 ( .B(n404), .A(Y[8]), .Z(n595) );
  NANDN U817 ( .B(n409), .A(n382), .Z(n594) );
  XNOR U818 ( .A(n591), .B(Y0[9]), .Z(n382) );
  XNOR U819 ( .A(n596), .B(n597), .Z(n591) );
  AND U820 ( .A(n420), .B(n599), .Z(n598) );
  XOR U821 ( .A(n556), .B(n600), .Z(n599) );
  XOR U822 ( .A(n600), .B(n557), .Z(n556) );
  OR U823 ( .A(n601), .B(n602), .Z(n557) );
  IV U824 ( .A(n597), .Z(n600) );
  XNOR U825 ( .A(n559), .B(n558), .Z(n597) );
  OR U826 ( .A(n603), .B(n604), .Z(n558) );
  XNOR U827 ( .A(n572), .B(n571), .Z(n559) );
  XOR U828 ( .A(n605), .B(n568), .Z(n571) );
  XNOR U829 ( .A(n606), .B(n563), .Z(n568) );
  NAND U830 ( .A(n567), .B(n467), .Z(n563) );
  NANDN U831 ( .B(n441), .A(n608), .Z(n607) );
  XNOR U832 ( .A(n569), .B(n570), .Z(n605) );
  XNOR U833 ( .A(n575), .B(n619), .Z(n578) );
  AND U834 ( .A(n502), .B(n535), .Z(n619) );
  XOR U835 ( .A(n620), .B(n621), .Z(n575) );
  ANDN U836 ( .A(n622), .B(n623), .Z(n621) );
  XNOR U837 ( .A(n624), .B(n620), .Z(n622) );
  XOR U838 ( .A(n625), .B(n579), .Z(n618) );
  NAND U839 ( .A(n497), .B(n539), .Z(n579) );
  IV U840 ( .A(n581), .Z(n625) );
  XNOR U841 ( .A(n588), .B(n589), .Z(n583) );
  NANDN U842 ( .B(n442), .A(n629), .Z(n589) );
  AND U843 ( .A(n584), .B(n466), .Z(n630) );
  NAND U844 ( .A(n631), .B(n632), .Z(n587) );
  NANDN U845 ( .B(n633), .A(n634), .Z(n631) );
  NAND U846 ( .A(n637), .B(n638), .Z(n210) );
  NANDN U847 ( .B(n357), .A(Y[7]), .Z(n638) );
  AND U848 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U849 ( .B(n404), .A(Y[7]), .Z(n640) );
  NANDN U850 ( .B(n409), .A(n379), .Z(n639) );
  XNOR U851 ( .A(n636), .B(Y0[8]), .Z(n379) );
  XNOR U852 ( .A(n641), .B(n642), .Z(n636) );
  AND U853 ( .A(n420), .B(n644), .Z(n643) );
  XOR U854 ( .A(n601), .B(n645), .Z(n644) );
  XOR U855 ( .A(n645), .B(n602), .Z(n601) );
  OR U856 ( .A(n646), .B(n647), .Z(n602) );
  IV U857 ( .A(n642), .Z(n645) );
  XNOR U858 ( .A(n604), .B(n603), .Z(n642) );
  NANDN U859 ( .B(n648), .A(n649), .Z(n603) );
  XNOR U860 ( .A(n614), .B(n613), .Z(n604) );
  XOR U861 ( .A(n650), .B(n617), .Z(n613) );
  XNOR U862 ( .A(n610), .B(n611), .Z(n617) );
  NAND U863 ( .A(n567), .B(n502), .Z(n611) );
  XNOR U864 ( .A(n609), .B(n651), .Z(n610) );
  AND U865 ( .A(n467), .B(n608), .Z(n651) );
  XNOR U866 ( .A(n616), .B(n612), .Z(n650) );
  AND U867 ( .A(n659), .B(n660), .Z(n658) );
  NANDN U868 ( .B(n441), .A(n661), .Z(n660) );
  OR U869 ( .A(n662), .B(n663), .Z(n659) );
  XNOR U870 ( .A(n620), .B(n668), .Z(n623) );
  AND U871 ( .A(n539), .B(n535), .Z(n668) );
  XOR U872 ( .A(n669), .B(n670), .Z(n620) );
  ANDN U873 ( .A(n671), .B(n672), .Z(n670) );
  XNOR U874 ( .A(n673), .B(n669), .Z(n671) );
  XOR U875 ( .A(n674), .B(n624), .Z(n667) );
  NAND U876 ( .A(n497), .B(n584), .Z(n624) );
  IV U877 ( .A(n626), .Z(n674) );
  XNOR U878 ( .A(n633), .B(n634), .Z(n628) );
  NANDN U879 ( .B(n442), .A(n678), .Z(n634) );
  XNOR U880 ( .A(n632), .B(n679), .Z(n633) );
  AND U881 ( .A(n629), .B(n466), .Z(n679) );
  ANDN U882 ( .A(n680), .B(n681), .Z(n632) );
  NANDN U883 ( .B(n682), .A(n683), .Z(n680) );
  NAND U884 ( .A(n686), .B(n687), .Z(n209) );
  NANDN U885 ( .B(n357), .A(Y[6]), .Z(n687) );
  AND U886 ( .A(n688), .B(n689), .Z(n686) );
  NANDN U887 ( .B(n404), .A(Y[6]), .Z(n689) );
  NANDN U888 ( .B(n409), .A(n376), .Z(n688) );
  XNOR U889 ( .A(n685), .B(Y0[7]), .Z(n376) );
  XNOR U890 ( .A(n691), .B(n692), .Z(n690) );
  AND U891 ( .A(n420), .B(n693), .Z(n692) );
  XOR U892 ( .A(n646), .B(n696), .Z(n693) );
  XOR U893 ( .A(n696), .B(n647), .Z(n646) );
  OR U894 ( .A(n694), .B(n695), .Z(n647) );
  XNOR U895 ( .A(n648), .B(n649), .Z(n696) );
  XNOR U896 ( .A(n657), .B(n656), .Z(n648) );
  XOR U897 ( .A(n701), .B(n666), .Z(n656) );
  XNOR U898 ( .A(n653), .B(n654), .Z(n666) );
  NAND U899 ( .A(n567), .B(n539), .Z(n654) );
  XNOR U900 ( .A(n652), .B(n702), .Z(n653) );
  AND U901 ( .A(n502), .B(n608), .Z(n702) );
  XNOR U902 ( .A(n665), .B(n655), .Z(n701) );
  XNOR U903 ( .A(n709), .B(n664), .Z(n665) );
  XNOR U904 ( .A(n713), .B(n662), .Z(n709) );
  NAND U905 ( .A(n661), .B(n467), .Z(n662) );
  NANDN U906 ( .B(n441), .A(n715), .Z(n714) );
  XNOR U907 ( .A(n669), .B(n720), .Z(n672) );
  AND U908 ( .A(n584), .B(n535), .Z(n720) );
  XOR U909 ( .A(n721), .B(n722), .Z(n669) );
  ANDN U910 ( .A(n723), .B(n724), .Z(n722) );
  XNOR U911 ( .A(n725), .B(n721), .Z(n723) );
  XOR U912 ( .A(n726), .B(n673), .Z(n719) );
  NAND U913 ( .A(n497), .B(n629), .Z(n673) );
  IV U914 ( .A(n675), .Z(n726) );
  XNOR U915 ( .A(n682), .B(n683), .Z(n677) );
  NANDN U916 ( .B(n442), .A(n730), .Z(n683) );
  AND U917 ( .A(n678), .B(n466), .Z(n731) );
  NAND U918 ( .A(n732), .B(n733), .Z(n681) );
  NANDN U919 ( .B(n734), .A(n735), .Z(n732) );
  IV U920 ( .A(n684), .Z(n691) );
  NAND U921 ( .A(n738), .B(n739), .Z(n208) );
  NANDN U922 ( .B(n357), .A(Y[5]), .Z(n739) );
  AND U923 ( .A(n740), .B(n741), .Z(n738) );
  NANDN U924 ( .B(n404), .A(Y[5]), .Z(n741) );
  NANDN U925 ( .B(n409), .A(n373), .Z(n740) );
  XNOR U926 ( .A(n737), .B(Y0[6]), .Z(n373) );
  XNOR U927 ( .A(n742), .B(n743), .Z(n737) );
  AND U928 ( .A(n420), .B(n745), .Z(n744) );
  XOR U929 ( .A(n694), .B(n746), .Z(n745) );
  XOR U930 ( .A(n746), .B(n695), .Z(n694) );
  OR U931 ( .A(n747), .B(n748), .Z(n695) );
  IV U932 ( .A(n743), .Z(n746) );
  XOR U933 ( .A(n700), .B(n699), .Z(n743) );
  XNOR U934 ( .A(n698), .B(n749), .Z(n699) );
  AND U935 ( .A(n697), .B(n750), .Z(n749) );
  AND U936 ( .A(n751), .B(n752), .Z(n750) );
  NANDN U937 ( .B(n441), .A(n753), .Z(n752) );
  OR U938 ( .A(n754), .B(n755), .Z(n751) );
  AND U939 ( .A(n756), .B(n757), .Z(n697) );
  NANDN U940 ( .B(n758), .A(n759), .Z(n757) );
  NANDN U941 ( .B(n760), .A(n761), .Z(n756) );
  XNOR U942 ( .A(n765), .B(n712), .Z(n707) );
  XNOR U943 ( .A(n704), .B(n705), .Z(n712) );
  NAND U944 ( .A(n567), .B(n584), .Z(n705) );
  XNOR U945 ( .A(n703), .B(n766), .Z(n704) );
  AND U946 ( .A(n539), .B(n608), .Z(n766) );
  XNOR U947 ( .A(n711), .B(n706), .Z(n765) );
  XNOR U948 ( .A(n716), .B(n774), .Z(n717) );
  AND U949 ( .A(n467), .B(n715), .Z(n774) );
  XOR U950 ( .A(n775), .B(n776), .Z(n716) );
  ANDN U951 ( .A(n777), .B(n778), .Z(n776) );
  XNOR U952 ( .A(n779), .B(n775), .Z(n777) );
  XOR U953 ( .A(n780), .B(n718), .Z(n773) );
  NAND U954 ( .A(n661), .B(n502), .Z(n718) );
  IV U955 ( .A(n710), .Z(n780) );
  XNOR U956 ( .A(n721), .B(n785), .Z(n724) );
  AND U957 ( .A(n629), .B(n535), .Z(n785) );
  XOR U958 ( .A(n786), .B(n787), .Z(n721) );
  ANDN U959 ( .A(n788), .B(n789), .Z(n787) );
  XNOR U960 ( .A(n790), .B(n786), .Z(n788) );
  XOR U961 ( .A(n791), .B(n725), .Z(n784) );
  NAND U962 ( .A(n497), .B(n678), .Z(n725) );
  IV U963 ( .A(n727), .Z(n791) );
  XNOR U964 ( .A(n734), .B(n735), .Z(n729) );
  NANDN U965 ( .B(n442), .A(n795), .Z(n735) );
  XNOR U966 ( .A(n733), .B(n796), .Z(n734) );
  AND U967 ( .A(n730), .B(n466), .Z(n796) );
  ANDN U968 ( .A(n797), .B(n798), .Z(n733) );
  NANDN U969 ( .B(n799), .A(n800), .Z(n797) );
  NAND U970 ( .A(n803), .B(n804), .Z(n207) );
  NANDN U971 ( .B(n357), .A(Y[4]), .Z(n804) );
  AND U972 ( .A(n805), .B(n806), .Z(n803) );
  NANDN U973 ( .B(n404), .A(Y[4]), .Z(n806) );
  NANDN U974 ( .B(n409), .A(n370), .Z(n805) );
  XNOR U975 ( .A(n802), .B(Y0[5]), .Z(n370) );
  XNOR U976 ( .A(n807), .B(n808), .Z(n802) );
  AND U977 ( .A(n420), .B(n810), .Z(n809) );
  XOR U978 ( .A(n747), .B(n811), .Z(n810) );
  XOR U979 ( .A(n811), .B(n748), .Z(n747) );
  OR U980 ( .A(n812), .B(n813), .Z(n748) );
  IV U981 ( .A(n808), .Z(n811) );
  XOR U982 ( .A(n764), .B(n763), .Z(n808) );
  XOR U983 ( .A(n758), .B(n759), .Z(n755) );
  XOR U984 ( .A(n818), .B(n760), .Z(n758) );
  NAND U985 ( .A(n467), .B(n753), .Z(n760) );
  NANDN U986 ( .B(n761), .A(n819), .Z(n818) );
  NANDN U987 ( .B(n441), .A(n820), .Z(n819) );
  XOR U988 ( .A(n824), .B(n754), .Z(n814) );
  OR U989 ( .A(n825), .B(n826), .Z(n754) );
  IV U990 ( .A(n762), .Z(n824) );
  XNOR U991 ( .A(n830), .B(n783), .Z(n771) );
  XNOR U992 ( .A(n768), .B(n769), .Z(n783) );
  NAND U993 ( .A(n567), .B(n629), .Z(n769) );
  XNOR U994 ( .A(n767), .B(n831), .Z(n768) );
  AND U995 ( .A(n584), .B(n608), .Z(n831) );
  XNOR U996 ( .A(n782), .B(n770), .Z(n830) );
  XNOR U997 ( .A(n775), .B(n839), .Z(n778) );
  AND U998 ( .A(n502), .B(n715), .Z(n839) );
  XOR U999 ( .A(n840), .B(n841), .Z(n775) );
  ANDN U1000 ( .A(n842), .B(n843), .Z(n841) );
  XNOR U1001 ( .A(n844), .B(n840), .Z(n842) );
  XOR U1002 ( .A(n845), .B(n779), .Z(n838) );
  NAND U1003 ( .A(n661), .B(n539), .Z(n779) );
  IV U1004 ( .A(n781), .Z(n845) );
  XNOR U1005 ( .A(n786), .B(n850), .Z(n789) );
  AND U1006 ( .A(n678), .B(n535), .Z(n850) );
  XOR U1007 ( .A(n851), .B(n852), .Z(n786) );
  ANDN U1008 ( .A(n853), .B(n854), .Z(n852) );
  XNOR U1009 ( .A(n855), .B(n851), .Z(n853) );
  XOR U1010 ( .A(n856), .B(n790), .Z(n849) );
  NAND U1011 ( .A(n497), .B(n730), .Z(n790) );
  IV U1012 ( .A(n792), .Z(n856) );
  XNOR U1013 ( .A(n799), .B(n800), .Z(n794) );
  NANDN U1014 ( .B(n442), .A(n860), .Z(n800) );
  AND U1015 ( .A(n795), .B(n466), .Z(n861) );
  NAND U1016 ( .A(n862), .B(n863), .Z(n798) );
  NANDN U1017 ( .B(n864), .A(n865), .Z(n862) );
  NAND U1018 ( .A(n868), .B(n869), .Z(n206) );
  NANDN U1019 ( .B(n357), .A(Y[3]), .Z(n869) );
  AND U1020 ( .A(n870), .B(n871), .Z(n868) );
  NANDN U1021 ( .B(n404), .A(Y[3]), .Z(n871) );
  NANDN U1022 ( .B(n409), .A(n367), .Z(n870) );
  XNOR U1023 ( .A(n867), .B(Y0[4]), .Z(n367) );
  XNOR U1024 ( .A(n872), .B(n873), .Z(n867) );
  AND U1025 ( .A(n420), .B(n875), .Z(n874) );
  XOR U1026 ( .A(n812), .B(n876), .Z(n875) );
  XOR U1027 ( .A(n876), .B(n813), .Z(n812) );
  OR U1028 ( .A(n877), .B(n878), .Z(n813) );
  IV U1029 ( .A(n873), .Z(n876) );
  XOR U1030 ( .A(n829), .B(n828), .Z(n873) );
  XOR U1031 ( .A(n879), .B(n825), .Z(n828) );
  XOR U1032 ( .A(n817), .B(n816), .Z(n825) );
  XOR U1033 ( .A(n815), .B(n880), .Z(n816) );
  AND U1034 ( .A(n881), .B(n882), .Z(n880) );
  NANDN U1035 ( .B(n441), .A(n883), .Z(n882) );
  OR U1036 ( .A(n884), .B(n885), .Z(n881) );
  NAND U1037 ( .A(n502), .B(n753), .Z(n823) );
  XNOR U1038 ( .A(n821), .B(n889), .Z(n822) );
  AND U1039 ( .A(n820), .B(n467), .Z(n889) );
  NANDN U1040 ( .B(n893), .A(n894), .Z(n826) );
  XNOR U1041 ( .A(n898), .B(n848), .Z(n836) );
  XNOR U1042 ( .A(n833), .B(n834), .Z(n848) );
  NAND U1043 ( .A(n567), .B(n678), .Z(n834) );
  XNOR U1044 ( .A(n832), .B(n899), .Z(n833) );
  AND U1045 ( .A(n629), .B(n608), .Z(n899) );
  XNOR U1046 ( .A(n847), .B(n835), .Z(n898) );
  XNOR U1047 ( .A(n840), .B(n907), .Z(n843) );
  AND U1048 ( .A(n539), .B(n715), .Z(n907) );
  XOR U1049 ( .A(n908), .B(n909), .Z(n840) );
  ANDN U1050 ( .A(n910), .B(n911), .Z(n909) );
  XNOR U1051 ( .A(n912), .B(n908), .Z(n910) );
  XOR U1052 ( .A(n913), .B(n844), .Z(n906) );
  NAND U1053 ( .A(n661), .B(n584), .Z(n844) );
  IV U1054 ( .A(n846), .Z(n913) );
  XNOR U1055 ( .A(n851), .B(n918), .Z(n854) );
  AND U1056 ( .A(n730), .B(n535), .Z(n918) );
  XOR U1057 ( .A(n919), .B(n920), .Z(n851) );
  ANDN U1058 ( .A(n921), .B(n922), .Z(n920) );
  XNOR U1059 ( .A(n923), .B(n919), .Z(n921) );
  XOR U1060 ( .A(n924), .B(n855), .Z(n917) );
  NAND U1061 ( .A(n497), .B(n795), .Z(n855) );
  IV U1062 ( .A(n857), .Z(n924) );
  XNOR U1063 ( .A(n864), .B(n865), .Z(n859) );
  NANDN U1064 ( .B(n442), .A(n928), .Z(n865) );
  XNOR U1065 ( .A(n863), .B(n929), .Z(n864) );
  AND U1066 ( .A(n860), .B(n466), .Z(n929) );
  ANDN U1067 ( .A(n930), .B(n931), .Z(n863) );
  NANDN U1068 ( .B(n932), .A(n933), .Z(n930) );
  NAND U1069 ( .A(n936), .B(n937), .Z(n205) );
  NANDN U1070 ( .B(n357), .A(Y[2]), .Z(n937) );
  AND U1071 ( .A(n938), .B(n939), .Z(n936) );
  NANDN U1072 ( .B(n404), .A(Y[2]), .Z(n939) );
  NANDN U1073 ( .B(n409), .A(n364), .Z(n938) );
  XNOR U1074 ( .A(n935), .B(Y0[3]), .Z(n364) );
  XNOR U1075 ( .A(n940), .B(n941), .Z(n935) );
  AND U1076 ( .A(n420), .B(n943), .Z(n942) );
  XOR U1077 ( .A(n877), .B(n944), .Z(n943) );
  XOR U1078 ( .A(n944), .B(n878), .Z(n877) );
  OR U1079 ( .A(n945), .B(n946), .Z(n878) );
  IV U1080 ( .A(n941), .Z(n944) );
  XOR U1081 ( .A(n897), .B(n896), .Z(n941) );
  XOR U1082 ( .A(n947), .B(n893), .Z(n896) );
  XOR U1083 ( .A(n888), .B(n887), .Z(n893) );
  XNOR U1084 ( .A(n952), .B(n884), .Z(n948) );
  NAND U1085 ( .A(n467), .B(n883), .Z(n884) );
  NANDN U1086 ( .B(n441), .A(n954), .Z(n953) );
  NAND U1087 ( .A(n539), .B(n753), .Z(n892) );
  XNOR U1088 ( .A(n890), .B(n958), .Z(n891) );
  AND U1089 ( .A(n820), .B(n502), .Z(n958) );
  XNOR U1090 ( .A(n894), .B(n895), .Z(n947) );
  XNOR U1091 ( .A(n968), .B(n916), .Z(n904) );
  XNOR U1092 ( .A(n901), .B(n902), .Z(n916) );
  NAND U1093 ( .A(n567), .B(n730), .Z(n902) );
  XNOR U1094 ( .A(n900), .B(n969), .Z(n901) );
  AND U1095 ( .A(n678), .B(n608), .Z(n969) );
  XNOR U1096 ( .A(n915), .B(n903), .Z(n968) );
  XNOR U1097 ( .A(n908), .B(n977), .Z(n911) );
  AND U1098 ( .A(n584), .B(n715), .Z(n977) );
  XOR U1099 ( .A(n981), .B(n912), .Z(n976) );
  NAND U1100 ( .A(n661), .B(n629), .Z(n912) );
  IV U1101 ( .A(n914), .Z(n981) );
  XNOR U1102 ( .A(n919), .B(n986), .Z(n922) );
  AND U1103 ( .A(n795), .B(n535), .Z(n986) );
  XOR U1104 ( .A(n987), .B(n988), .Z(n919) );
  ANDN U1105 ( .A(n989), .B(n990), .Z(n988) );
  XNOR U1106 ( .A(n991), .B(n987), .Z(n989) );
  XOR U1107 ( .A(n992), .B(n923), .Z(n985) );
  NAND U1108 ( .A(n497), .B(n860), .Z(n923) );
  IV U1109 ( .A(n925), .Z(n992) );
  XNOR U1110 ( .A(n932), .B(n933), .Z(n927) );
  OR U1111 ( .A(n996), .B(n442), .Z(n933) );
  AND U1112 ( .A(n928), .B(n466), .Z(n997) );
  NAND U1113 ( .A(n998), .B(n999), .Z(n931) );
  NANDN U1114 ( .B(n1000), .A(n1001), .Z(n998) );
  NAND U1115 ( .A(n1004), .B(n1005), .Z(n204) );
  NANDN U1116 ( .B(n357), .A(Y[1]), .Z(n1005) );
  AND U1117 ( .A(n1006), .B(n1007), .Z(n1004) );
  NANDN U1118 ( .B(n404), .A(Y[1]), .Z(n1007) );
  NANDN U1119 ( .B(n409), .A(n360), .Z(n1006) );
  XNOR U1120 ( .A(n1003), .B(Y0[2]), .Z(n360) );
  XNOR U1121 ( .A(n1008), .B(n1009), .Z(n1003) );
  XOR U1122 ( .A(n1002), .B(n1010), .Z(n1008) );
  AND U1123 ( .A(n420), .B(n1011), .Z(n1010) );
  XOR U1124 ( .A(n945), .B(n1012), .Z(n1011) );
  XOR U1125 ( .A(n1012), .B(n946), .Z(n945) );
  NANDN U1126 ( .B(n1013), .A(n1014), .Z(n946) );
  IV U1127 ( .A(n1009), .Z(n1012) );
  XOR U1128 ( .A(n964), .B(n963), .Z(n1009) );
  XNOR U1129 ( .A(n1015), .B(n967), .Z(n963) );
  XNOR U1130 ( .A(n955), .B(n1017), .Z(n956) );
  AND U1131 ( .A(n954), .B(n467), .Z(n1017) );
  XOR U1132 ( .A(n1021), .B(n957), .Z(n1016) );
  NAND U1133 ( .A(n502), .B(n883), .Z(n957) );
  IV U1134 ( .A(n949), .Z(n1021) );
  XNOR U1135 ( .A(n960), .B(n961), .Z(n951) );
  NAND U1136 ( .A(n584), .B(n753), .Z(n961) );
  XNOR U1137 ( .A(n959), .B(n1025), .Z(n960) );
  AND U1138 ( .A(n820), .B(n539), .Z(n1025) );
  XNOR U1139 ( .A(n966), .B(n962), .Z(n1015) );
  AND U1140 ( .A(n1033), .B(n1034), .Z(n1032) );
  OR U1141 ( .A(n1035), .B(n1036), .Z(n1034) );
  AND U1142 ( .A(n1037), .B(n1038), .Z(n1033) );
  NANDN U1143 ( .B(n441), .A(n1039), .Z(n1038) );
  NANDN U1144 ( .B(n1040), .A(n1041), .Z(n1037) );
  XNOR U1145 ( .A(n1045), .B(n984), .Z(n974) );
  XNOR U1146 ( .A(n971), .B(n972), .Z(n984) );
  NAND U1147 ( .A(n567), .B(n795), .Z(n972) );
  XNOR U1148 ( .A(n970), .B(n1046), .Z(n971) );
  AND U1149 ( .A(n730), .B(n608), .Z(n1046) );
  XNOR U1150 ( .A(n983), .B(n973), .Z(n1045) );
  XNOR U1151 ( .A(n978), .B(n1054), .Z(n979) );
  AND U1152 ( .A(n629), .B(n715), .Z(n1054) );
  XOR U1153 ( .A(n1058), .B(n980), .Z(n1053) );
  NAND U1154 ( .A(n661), .B(n678), .Z(n980) );
  IV U1155 ( .A(n982), .Z(n1058) );
  XNOR U1156 ( .A(n987), .B(n1063), .Z(n990) );
  AND U1157 ( .A(n860), .B(n535), .Z(n1063) );
  XOR U1158 ( .A(n1064), .B(n1065), .Z(n987) );
  ANDN U1159 ( .A(n1066), .B(n1067), .Z(n1065) );
  XNOR U1160 ( .A(n1068), .B(n1064), .Z(n1066) );
  XOR U1161 ( .A(n1069), .B(n991), .Z(n1062) );
  NAND U1162 ( .A(n497), .B(n928), .Z(n991) );
  IV U1163 ( .A(n993), .Z(n1069) );
  XNOR U1164 ( .A(n1000), .B(n1001), .Z(n995) );
  OR U1165 ( .A(n1073), .B(n442), .Z(n1001) );
  XNOR U1166 ( .A(n999), .B(n1074), .Z(n1000) );
  ANDN U1167 ( .A(n466), .B(n996), .Z(n1074) );
  ANDN U1168 ( .A(n1075), .B(n1076), .Z(n999) );
  NANDN U1169 ( .B(n1077), .A(n1078), .Z(n1075) );
  NAND U1170 ( .A(n1081), .B(n1082), .Z(n203) );
  NANDN U1171 ( .B(n357), .A(Y[0]), .Z(n1082) );
  AND U1172 ( .A(n1083), .B(n1084), .Z(n1081) );
  NANDN U1173 ( .B(n404), .A(Y[0]), .Z(n1084) );
  IV U1174 ( .A(n1085), .Z(n404) );
  OR U1175 ( .A(n409), .B(n355), .Z(n1083) );
  IV U1176 ( .A(Y0[1]), .Z(n361) );
  XOR U1177 ( .A(n1086), .B(n1087), .Z(n1080) );
  XNOR U1178 ( .A(n1088), .B(n1079), .Z(n1086) );
  NAND U1179 ( .A(Y0[0]), .B(n1013), .Z(n1079) );
  NAND U1180 ( .A(n1089), .B(n420), .Z(n1088) );
  XOR U1181 ( .A(A[15]), .B(X[15]), .Z(n420) );
  XNOR U1182 ( .A(n1014), .B(n1087), .Z(n1089) );
  XNOR U1183 ( .A(n1013), .B(n1087), .Z(n1014) );
  XNOR U1184 ( .A(n1031), .B(n1030), .Z(n1087) );
  XNOR U1185 ( .A(n1090), .B(n1044), .Z(n1030) );
  XNOR U1186 ( .A(n1018), .B(n1092), .Z(n1019) );
  AND U1187 ( .A(n954), .B(n502), .Z(n1092) );
  XOR U1188 ( .A(n1096), .B(n1020), .Z(n1091) );
  NAND U1189 ( .A(n539), .B(n883), .Z(n1020) );
  IV U1190 ( .A(n1022), .Z(n1096) );
  XNOR U1191 ( .A(n1027), .B(n1028), .Z(n1024) );
  NAND U1192 ( .A(n629), .B(n753), .Z(n1028) );
  XNOR U1193 ( .A(n1026), .B(n1100), .Z(n1027) );
  AND U1194 ( .A(n820), .B(n584), .Z(n1100) );
  XNOR U1195 ( .A(n1043), .B(n1029), .Z(n1090) );
  XNOR U1196 ( .A(n1107), .B(n1040), .Z(n1043) );
  XOR U1197 ( .A(n1108), .B(n1035), .Z(n1040) );
  NAND U1198 ( .A(n467), .B(n1039), .Z(n1035) );
  NANDN U1199 ( .B(n441), .A(n1110), .Z(n1109) );
  XNOR U1200 ( .A(n1041), .B(n1042), .Z(n1107) );
  XNOR U1201 ( .A(n1120), .B(n1061), .Z(n1051) );
  XNOR U1202 ( .A(n1048), .B(n1049), .Z(n1061) );
  NAND U1203 ( .A(n567), .B(n860), .Z(n1049) );
  XNOR U1204 ( .A(n1047), .B(n1121), .Z(n1048) );
  AND U1205 ( .A(n795), .B(n608), .Z(n1121) );
  XNOR U1206 ( .A(n1060), .B(n1050), .Z(n1120) );
  XNOR U1207 ( .A(n1055), .B(n1129), .Z(n1056) );
  AND U1208 ( .A(n678), .B(n715), .Z(n1129) );
  XOR U1209 ( .A(n1133), .B(n1057), .Z(n1128) );
  NAND U1210 ( .A(n661), .B(n730), .Z(n1057) );
  IV U1211 ( .A(n1059), .Z(n1133) );
  XNOR U1212 ( .A(n1064), .B(n1138), .Z(n1067) );
  AND U1213 ( .A(n928), .B(n535), .Z(n1138) );
  XOR U1214 ( .A(n1142), .B(n1068), .Z(n1137) );
  NANDN U1215 ( .B(n996), .A(n497), .Z(n1068) );
  IV U1216 ( .A(n1070), .Z(n1142) );
  XNOR U1217 ( .A(n1077), .B(n1078), .Z(n1072) );
  NANDN U1218 ( .B(n442), .A(n1146), .Z(n1078) );
  ANDN U1219 ( .A(n466), .B(n1073), .Z(n1147) );
  NAND U1220 ( .A(n1148), .B(n1149), .Z(n1076) );
  NANDN U1221 ( .B(n1150), .A(n1151), .Z(n1148) );
  XNOR U1222 ( .A(n1106), .B(n1105), .Z(n1013) );
  XNOR U1223 ( .A(n1152), .B(n1116), .Z(n1105) );
  XNOR U1224 ( .A(n1093), .B(n1154), .Z(n1094) );
  AND U1225 ( .A(n954), .B(n539), .Z(n1154) );
  XOR U1226 ( .A(n1158), .B(n1095), .Z(n1153) );
  NAND U1227 ( .A(n584), .B(n883), .Z(n1095) );
  IV U1228 ( .A(n1097), .Z(n1158) );
  XNOR U1229 ( .A(n1102), .B(n1103), .Z(n1099) );
  NAND U1230 ( .A(n678), .B(n753), .Z(n1103) );
  XNOR U1231 ( .A(n1101), .B(n1162), .Z(n1102) );
  AND U1232 ( .A(n820), .B(n629), .Z(n1162) );
  XNOR U1233 ( .A(n1115), .B(n1104), .Z(n1152) );
  XOR U1234 ( .A(n1166), .B(n1167), .Z(n1104) );
  XNOR U1235 ( .A(n1168), .B(n1119), .Z(n1115) );
  NAND U1236 ( .A(n502), .B(n1039), .Z(n1113) );
  XNOR U1237 ( .A(n1111), .B(n1169), .Z(n1112) );
  AND U1238 ( .A(n1110), .B(n467), .Z(n1169) );
  XNOR U1239 ( .A(n1118), .B(n1114), .Z(n1168) );
  XOR U1240 ( .A(n1173), .B(n1174), .Z(n1114) );
  AND U1241 ( .A(n1175), .B(n1176), .Z(n1174) );
  XOR U1242 ( .A(n1177), .B(n1178), .Z(n1176) );
  XOR U1243 ( .A(n1173), .B(n1179), .Z(n1178) );
  XOR U1244 ( .A(n1160), .B(n1180), .Z(n1175) );
  XOR U1245 ( .A(n1173), .B(n1161), .Z(n1180) );
  NAND U1246 ( .A(n753), .B(n730), .Z(n1165) );
  XNOR U1247 ( .A(n1163), .B(n1181), .Z(n1164) );
  AND U1248 ( .A(n820), .B(n678), .Z(n1181) );
  XNOR U1249 ( .A(n1155), .B(n1186), .Z(n1156) );
  AND U1250 ( .A(n954), .B(n584), .Z(n1186) );
  XOR U1251 ( .A(n1187), .B(n1188), .Z(n1155) );
  ANDN U1252 ( .A(n1189), .B(n1190), .Z(n1188) );
  XNOR U1253 ( .A(n1191), .B(n1187), .Z(n1189) );
  XOR U1254 ( .A(n1192), .B(n1157), .Z(n1185) );
  NAND U1255 ( .A(n629), .B(n883), .Z(n1157) );
  IV U1256 ( .A(n1159), .Z(n1192) );
  XOR U1257 ( .A(n1196), .B(n1197), .Z(n1173) );
  AND U1258 ( .A(n1198), .B(n1199), .Z(n1197) );
  XOR U1259 ( .A(n1200), .B(n1201), .Z(n1199) );
  XOR U1260 ( .A(n1196), .B(n1202), .Z(n1201) );
  XOR U1261 ( .A(n1194), .B(n1203), .Z(n1198) );
  XOR U1262 ( .A(n1196), .B(n1195), .Z(n1203) );
  NAND U1263 ( .A(n753), .B(n795), .Z(n1184) );
  XNOR U1264 ( .A(n1182), .B(n1204), .Z(n1183) );
  AND U1265 ( .A(n730), .B(n820), .Z(n1204) );
  XNOR U1266 ( .A(n1187), .B(n1209), .Z(n1190) );
  AND U1267 ( .A(n954), .B(n629), .Z(n1209) );
  XOR U1268 ( .A(n1210), .B(n1211), .Z(n1187) );
  ANDN U1269 ( .A(n1212), .B(n1213), .Z(n1211) );
  XNOR U1270 ( .A(n1214), .B(n1210), .Z(n1212) );
  XOR U1271 ( .A(n1215), .B(n1191), .Z(n1208) );
  NAND U1272 ( .A(n678), .B(n883), .Z(n1191) );
  IV U1273 ( .A(n1193), .Z(n1215) );
  XOR U1274 ( .A(n1219), .B(n1220), .Z(n1196) );
  AND U1275 ( .A(n1221), .B(n1222), .Z(n1220) );
  XOR U1276 ( .A(n1223), .B(n1224), .Z(n1222) );
  XOR U1277 ( .A(n1219), .B(n1225), .Z(n1224) );
  XOR U1278 ( .A(n1217), .B(n1226), .Z(n1221) );
  XOR U1279 ( .A(n1219), .B(n1218), .Z(n1226) );
  NAND U1280 ( .A(n753), .B(n860), .Z(n1207) );
  XNOR U1281 ( .A(n1205), .B(n1227), .Z(n1206) );
  AND U1282 ( .A(n795), .B(n820), .Z(n1227) );
  XNOR U1283 ( .A(n1210), .B(n1232), .Z(n1213) );
  AND U1284 ( .A(n954), .B(n678), .Z(n1232) );
  XOR U1285 ( .A(n1233), .B(n1234), .Z(n1210) );
  ANDN U1286 ( .A(n1235), .B(n1236), .Z(n1234) );
  XNOR U1287 ( .A(n1237), .B(n1233), .Z(n1235) );
  XOR U1288 ( .A(n1238), .B(n1214), .Z(n1231) );
  NAND U1289 ( .A(n883), .B(n730), .Z(n1214) );
  IV U1290 ( .A(n1216), .Z(n1238) );
  XOR U1291 ( .A(n1242), .B(n1243), .Z(n1219) );
  AND U1292 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U1293 ( .A(n1246), .B(n1247), .Z(n1245) );
  XOR U1294 ( .A(n1242), .B(n1248), .Z(n1247) );
  XOR U1295 ( .A(n1240), .B(n1249), .Z(n1244) );
  XOR U1296 ( .A(n1242), .B(n1241), .Z(n1249) );
  XNOR U1297 ( .A(n1250), .B(n1230), .Z(n1241) );
  NAND U1298 ( .A(n753), .B(n928), .Z(n1230) );
  IV U1299 ( .A(n1229), .Z(n1250) );
  XNOR U1300 ( .A(n1228), .B(n1251), .Z(n1229) );
  AND U1301 ( .A(n860), .B(n820), .Z(n1251) );
  XOR U1302 ( .A(n1252), .B(n1253), .Z(n1228) );
  ANDN U1303 ( .A(n1254), .B(n1255), .Z(n1253) );
  XNOR U1304 ( .A(n1256), .B(n1252), .Z(n1254) );
  XNOR U1305 ( .A(n1257), .B(n1258), .Z(n1240) );
  IV U1306 ( .A(n1236), .Z(n1258) );
  XNOR U1307 ( .A(n1233), .B(n1259), .Z(n1236) );
  AND U1308 ( .A(n730), .B(n954), .Z(n1259) );
  XOR U1309 ( .A(n1260), .B(n1261), .Z(n1233) );
  ANDN U1310 ( .A(n1262), .B(n1263), .Z(n1261) );
  XNOR U1311 ( .A(n1264), .B(n1260), .Z(n1262) );
  XOR U1312 ( .A(n1265), .B(n1237), .Z(n1257) );
  NAND U1313 ( .A(n883), .B(n795), .Z(n1237) );
  IV U1314 ( .A(n1239), .Z(n1265) );
  XOR U1315 ( .A(n1269), .B(n1270), .Z(n1242) );
  AND U1316 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U1317 ( .A(n1273), .B(n1274), .Z(n1272) );
  XOR U1318 ( .A(n1269), .B(n1275), .Z(n1274) );
  XOR U1319 ( .A(n1267), .B(n1276), .Z(n1271) );
  XOR U1320 ( .A(n1269), .B(n1268), .Z(n1276) );
  XNOR U1321 ( .A(n1277), .B(n1256), .Z(n1268) );
  NANDN U1322 ( .B(n996), .A(n753), .Z(n1256) );
  IV U1323 ( .A(n1255), .Z(n1277) );
  XNOR U1324 ( .A(n1252), .B(n1278), .Z(n1255) );
  AND U1325 ( .A(n928), .B(n820), .Z(n1278) );
  XOR U1326 ( .A(n1279), .B(n1280), .Z(n1252) );
  ANDN U1327 ( .A(n1281), .B(n1282), .Z(n1280) );
  XNOR U1328 ( .A(n1283), .B(n1279), .Z(n1281) );
  XNOR U1329 ( .A(n1284), .B(n1285), .Z(n1267) );
  IV U1330 ( .A(n1263), .Z(n1285) );
  XNOR U1331 ( .A(n1260), .B(n1286), .Z(n1263) );
  AND U1332 ( .A(n795), .B(n954), .Z(n1286) );
  XOR U1333 ( .A(n1287), .B(n1288), .Z(n1260) );
  ANDN U1334 ( .A(n1289), .B(n1290), .Z(n1288) );
  XNOR U1335 ( .A(n1291), .B(n1287), .Z(n1289) );
  XOR U1336 ( .A(n1292), .B(n1264), .Z(n1284) );
  NAND U1337 ( .A(n883), .B(n860), .Z(n1264) );
  IV U1338 ( .A(n1266), .Z(n1292) );
  XOR U1339 ( .A(n1296), .B(n1297), .Z(n1269) );
  AND U1340 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U1341 ( .A(n1300), .B(n1301), .Z(n1299) );
  XOR U1342 ( .A(n1296), .B(n1302), .Z(n1301) );
  XOR U1343 ( .A(n1294), .B(n1303), .Z(n1298) );
  XOR U1344 ( .A(n1296), .B(n1295), .Z(n1303) );
  XNOR U1345 ( .A(n1304), .B(n1283), .Z(n1295) );
  NANDN U1346 ( .B(n1073), .A(n753), .Z(n1283) );
  IV U1347 ( .A(n1282), .Z(n1304) );
  XNOR U1348 ( .A(n1279), .B(n1305), .Z(n1282) );
  ANDN U1349 ( .A(n820), .B(n996), .Z(n1305) );
  XOR U1350 ( .A(n1306), .B(n1307), .Z(n1279) );
  ANDN U1351 ( .A(n1308), .B(n1309), .Z(n1307) );
  XNOR U1352 ( .A(n1310), .B(n1306), .Z(n1308) );
  XNOR U1353 ( .A(n1311), .B(n1312), .Z(n1294) );
  IV U1354 ( .A(n1290), .Z(n1312) );
  XNOR U1355 ( .A(n1287), .B(n1313), .Z(n1290) );
  AND U1356 ( .A(n860), .B(n954), .Z(n1313) );
  XOR U1357 ( .A(n1314), .B(n1315), .Z(n1287) );
  ANDN U1358 ( .A(n1316), .B(n1317), .Z(n1315) );
  XNOR U1359 ( .A(n1318), .B(n1314), .Z(n1316) );
  XOR U1360 ( .A(n1319), .B(n1291), .Z(n1311) );
  NAND U1361 ( .A(n883), .B(n928), .Z(n1291) );
  IV U1362 ( .A(n1293), .Z(n1319) );
  XOR U1363 ( .A(n1323), .B(n1324), .Z(n1296) );
  AND U1364 ( .A(n1325), .B(n1326), .Z(n1324) );
  XOR U1365 ( .A(n1327), .B(n1328), .Z(n1326) );
  XOR U1366 ( .A(n1323), .B(n1329), .Z(n1328) );
  XOR U1367 ( .A(n1321), .B(n1330), .Z(n1325) );
  XOR U1368 ( .A(n1323), .B(n1322), .Z(n1330) );
  XNOR U1369 ( .A(n1331), .B(n1310), .Z(n1322) );
  NAND U1370 ( .A(n753), .B(n1146), .Z(n1310) );
  IV U1371 ( .A(n1309), .Z(n1331) );
  XNOR U1372 ( .A(n1306), .B(n1332), .Z(n1309) );
  ANDN U1373 ( .A(n820), .B(n1073), .Z(n1332) );
  XOR U1374 ( .A(n1333), .B(n1334), .Z(n1306) );
  ANDN U1375 ( .A(n1335), .B(n1336), .Z(n1334) );
  XNOR U1376 ( .A(n1337), .B(n1333), .Z(n1335) );
  XNOR U1377 ( .A(n1338), .B(n1339), .Z(n1321) );
  IV U1378 ( .A(n1317), .Z(n1339) );
  XNOR U1379 ( .A(n1314), .B(n1340), .Z(n1317) );
  AND U1380 ( .A(n928), .B(n954), .Z(n1340) );
  XOR U1381 ( .A(n1341), .B(n1342), .Z(n1314) );
  ANDN U1382 ( .A(n1343), .B(n1344), .Z(n1342) );
  XNOR U1383 ( .A(n1345), .B(n1341), .Z(n1343) );
  XOR U1384 ( .A(n1346), .B(n1318), .Z(n1338) );
  NANDN U1385 ( .B(n996), .A(n883), .Z(n1318) );
  IV U1386 ( .A(n1320), .Z(n1346) );
  XOR U1387 ( .A(n1351), .B(n1352), .Z(n1167) );
  XNOR U1388 ( .A(n1353), .B(n1350), .Z(n1351) );
  XNOR U1389 ( .A(n1341), .B(n1355), .Z(n1344) );
  ANDN U1390 ( .A(n954), .B(n996), .Z(n1355) );
  XOR U1391 ( .A(n1358), .B(n1356), .Z(n1357) );
  ANDN U1392 ( .A(n954), .B(n1073), .Z(n1358) );
  AND U1393 ( .A(n1146), .B(n883), .Z(n1359) );
  XOR U1394 ( .A(n1360), .B(n1361), .Z(n1356) );
  ANDN U1395 ( .A(n1362), .B(n1363), .Z(n1361) );
  XNOR U1396 ( .A(n1364), .B(n1360), .Z(n1362) );
  XOR U1397 ( .A(n1365), .B(n1345), .Z(n1354) );
  NANDN U1398 ( .B(n1073), .A(n883), .Z(n1345) );
  IV U1399 ( .A(n1347), .Z(n1365) );
  NAND U1400 ( .A(n883), .B(n1366), .Z(n1364) );
  XNOR U1401 ( .A(n1360), .B(n1367), .Z(n1363) );
  AND U1402 ( .A(n1146), .B(n954), .Z(n1367) );
  AND U1403 ( .A(n1368), .B(A[0]), .Z(n1360) );
  NANDN U1404 ( .B(n883), .A(n1369), .Z(n1368) );
  NAND U1405 ( .A(n1366), .B(n954), .Z(n1369) );
  XNOR U1406 ( .A(n1336), .B(n1337), .Z(n1349) );
  NAND U1407 ( .A(n753), .B(n1366), .Z(n1337) );
  XNOR U1408 ( .A(n1333), .B(n1372), .Z(n1336) );
  AND U1409 ( .A(n1146), .B(n820), .Z(n1372) );
  AND U1410 ( .A(n1373), .B(A[0]), .Z(n1333) );
  NANDN U1411 ( .B(n753), .A(n1374), .Z(n1373) );
  NAND U1412 ( .A(n1366), .B(n820), .Z(n1374) );
  XOR U1413 ( .A(n1377), .B(n1378), .Z(n1350) );
  XOR U1414 ( .A(n1379), .B(n1380), .Z(n1118) );
  AND U1415 ( .A(n1381), .B(n1382), .Z(n1380) );
  NANDN U1416 ( .B(n441), .A(n1383), .Z(n1382) );
  NANDN U1417 ( .B(n1384), .A(n1385), .Z(n441) );
  AND U1418 ( .A(n1386), .B(A[15]), .Z(n1385) );
  OR U1419 ( .A(n1387), .B(n1388), .Z(n1381) );
  IV U1420 ( .A(n1117), .Z(n1379) );
  NAND U1421 ( .A(n539), .B(n1039), .Z(n1172) );
  XNOR U1422 ( .A(n1170), .B(n1390), .Z(n1171) );
  AND U1423 ( .A(n1110), .B(n502), .Z(n1390) );
  XOR U1424 ( .A(n1398), .B(n1387), .Z(n1394) );
  NAND U1425 ( .A(n467), .B(n1383), .Z(n1387) );
  IV U1426 ( .A(n1389), .Z(n1398) );
  NAND U1427 ( .A(n584), .B(n1039), .Z(n1393) );
  XNOR U1428 ( .A(n1391), .B(n1400), .Z(n1392) );
  AND U1429 ( .A(n1110), .B(n539), .Z(n1400) );
  XNOR U1430 ( .A(n1395), .B(n1405), .Z(n1396) );
  AND U1431 ( .A(n467), .B(X[0]), .Z(n1405) );
  XNOR U1432 ( .A(n1386), .B(A[14]), .Z(n1384) );
  NOR U1433 ( .A(n1406), .B(n1407), .Z(n1386) );
  XOR U1434 ( .A(n1411), .B(n1397), .Z(n1404) );
  NAND U1435 ( .A(n502), .B(n1383), .Z(n1397) );
  IV U1436 ( .A(n1399), .Z(n1411) );
  NAND U1437 ( .A(n629), .B(n1039), .Z(n1403) );
  XNOR U1438 ( .A(n1401), .B(n1413), .Z(n1402) );
  AND U1439 ( .A(n1110), .B(n584), .Z(n1413) );
  XOR U1440 ( .A(n1414), .B(n1415), .Z(n1401) );
  ANDN U1441 ( .A(n1416), .B(n1417), .Z(n1415) );
  XNOR U1442 ( .A(n1418), .B(n1414), .Z(n1416) );
  XNOR U1443 ( .A(n1408), .B(n1420), .Z(n1409) );
  AND U1444 ( .A(n502), .B(X[0]), .Z(n1420) );
  XOR U1445 ( .A(n1406), .B(A[13]), .Z(n1407) );
  NANDN U1446 ( .B(n1421), .A(n1422), .Z(n1406) );
  XOR U1447 ( .A(n1426), .B(n1410), .Z(n1419) );
  NAND U1448 ( .A(n539), .B(n1383), .Z(n1410) );
  IV U1449 ( .A(n1412), .Z(n1426) );
  XNOR U1450 ( .A(n1428), .B(n1418), .Z(n1246) );
  NAND U1451 ( .A(n678), .B(n1039), .Z(n1418) );
  IV U1452 ( .A(n1417), .Z(n1428) );
  XNOR U1453 ( .A(n1414), .B(n1429), .Z(n1417) );
  AND U1454 ( .A(n1110), .B(n629), .Z(n1429) );
  XOR U1455 ( .A(n1430), .B(n1431), .Z(n1414) );
  ANDN U1456 ( .A(n1432), .B(n1433), .Z(n1431) );
  XNOR U1457 ( .A(n1434), .B(n1430), .Z(n1432) );
  XNOR U1458 ( .A(n1435), .B(n1436), .Z(n1248) );
  IV U1459 ( .A(n1424), .Z(n1436) );
  XNOR U1460 ( .A(n1423), .B(n1437), .Z(n1424) );
  AND U1461 ( .A(n539), .B(X[0]), .Z(n1437) );
  XNOR U1462 ( .A(n1422), .B(A[12]), .Z(n1421) );
  NOR U1463 ( .A(n1438), .B(n1439), .Z(n1422) );
  XOR U1464 ( .A(n1440), .B(n1441), .Z(n1423) );
  ANDN U1465 ( .A(n1442), .B(n1443), .Z(n1441) );
  XNOR U1466 ( .A(n1444), .B(n1440), .Z(n1442) );
  XOR U1467 ( .A(n1445), .B(n1425), .Z(n1435) );
  NAND U1468 ( .A(n584), .B(n1383), .Z(n1425) );
  IV U1469 ( .A(n1427), .Z(n1445) );
  XNOR U1470 ( .A(n1447), .B(n1434), .Z(n1273) );
  NAND U1471 ( .A(n730), .B(n1039), .Z(n1434) );
  IV U1472 ( .A(n1433), .Z(n1447) );
  XNOR U1473 ( .A(n1430), .B(n1448), .Z(n1433) );
  AND U1474 ( .A(n1110), .B(n678), .Z(n1448) );
  XOR U1475 ( .A(n1449), .B(n1450), .Z(n1430) );
  ANDN U1476 ( .A(n1451), .B(n1452), .Z(n1450) );
  XNOR U1477 ( .A(n1453), .B(n1449), .Z(n1451) );
  XNOR U1478 ( .A(n1454), .B(n1455), .Z(n1275) );
  IV U1479 ( .A(n1443), .Z(n1455) );
  XNOR U1480 ( .A(n1440), .B(n1456), .Z(n1443) );
  AND U1481 ( .A(n584), .B(X[0]), .Z(n1456) );
  XOR U1482 ( .A(n1438), .B(A[11]), .Z(n1439) );
  NANDN U1483 ( .B(n1457), .A(n1458), .Z(n1438) );
  XOR U1484 ( .A(n1459), .B(n1460), .Z(n1440) );
  ANDN U1485 ( .A(n1461), .B(n1462), .Z(n1460) );
  XNOR U1486 ( .A(n1463), .B(n1459), .Z(n1461) );
  XOR U1487 ( .A(n1464), .B(n1444), .Z(n1454) );
  NAND U1488 ( .A(n629), .B(n1383), .Z(n1444) );
  IV U1489 ( .A(n1446), .Z(n1464) );
  XNOR U1490 ( .A(n1466), .B(n1453), .Z(n1300) );
  NAND U1491 ( .A(n795), .B(n1039), .Z(n1453) );
  IV U1492 ( .A(n1452), .Z(n1466) );
  XNOR U1493 ( .A(n1449), .B(n1467), .Z(n1452) );
  AND U1494 ( .A(n1110), .B(n730), .Z(n1467) );
  XOR U1495 ( .A(n1468), .B(n1469), .Z(n1449) );
  ANDN U1496 ( .A(n1470), .B(n1471), .Z(n1469) );
  XNOR U1497 ( .A(n1472), .B(n1468), .Z(n1470) );
  XNOR U1498 ( .A(n1473), .B(n1474), .Z(n1302) );
  IV U1499 ( .A(n1462), .Z(n1474) );
  XNOR U1500 ( .A(n1459), .B(n1475), .Z(n1462) );
  AND U1501 ( .A(n629), .B(X[0]), .Z(n1475) );
  XNOR U1502 ( .A(n1458), .B(A[10]), .Z(n1457) );
  NOR U1503 ( .A(n1476), .B(n1477), .Z(n1458) );
  XOR U1504 ( .A(n1478), .B(n1479), .Z(n1459) );
  ANDN U1505 ( .A(n1480), .B(n1481), .Z(n1479) );
  XNOR U1506 ( .A(n1482), .B(n1478), .Z(n1480) );
  XOR U1507 ( .A(n1483), .B(n1463), .Z(n1473) );
  NAND U1508 ( .A(n678), .B(n1383), .Z(n1463) );
  IV U1509 ( .A(n1465), .Z(n1483) );
  XNOR U1510 ( .A(n1485), .B(n1472), .Z(n1327) );
  NAND U1511 ( .A(n860), .B(n1039), .Z(n1472) );
  IV U1512 ( .A(n1471), .Z(n1485) );
  XNOR U1513 ( .A(n1468), .B(n1486), .Z(n1471) );
  AND U1514 ( .A(n1110), .B(n795), .Z(n1486) );
  XOR U1515 ( .A(n1487), .B(n1488), .Z(n1468) );
  ANDN U1516 ( .A(n1489), .B(n1490), .Z(n1488) );
  XNOR U1517 ( .A(n1491), .B(n1487), .Z(n1489) );
  XNOR U1518 ( .A(n1492), .B(n1493), .Z(n1329) );
  IV U1519 ( .A(n1481), .Z(n1493) );
  XNOR U1520 ( .A(n1478), .B(n1494), .Z(n1481) );
  AND U1521 ( .A(n678), .B(X[0]), .Z(n1494) );
  XOR U1522 ( .A(n1476), .B(A[9]), .Z(n1477) );
  NANDN U1523 ( .B(n1495), .A(n1496), .Z(n1476) );
  XOR U1524 ( .A(n1497), .B(n1498), .Z(n1478) );
  ANDN U1525 ( .A(n1499), .B(n1500), .Z(n1498) );
  XNOR U1526 ( .A(n1501), .B(n1497), .Z(n1499) );
  XOR U1527 ( .A(n1502), .B(n1482), .Z(n1492) );
  NAND U1528 ( .A(n730), .B(n1383), .Z(n1482) );
  IV U1529 ( .A(n1484), .Z(n1502) );
  NAND U1530 ( .A(n928), .B(n1039), .Z(n1491) );
  XNOR U1531 ( .A(n1487), .B(n1504), .Z(n1490) );
  AND U1532 ( .A(n1110), .B(n860), .Z(n1504) );
  XNOR U1533 ( .A(n1508), .B(n1505), .Z(n1507) );
  XNOR U1534 ( .A(n1497), .B(n1510), .Z(n1500) );
  AND U1535 ( .A(n730), .B(X[0]), .Z(n1510) );
  XNOR U1536 ( .A(n1514), .B(n1511), .Z(n1513) );
  XOR U1537 ( .A(n1515), .B(n1501), .Z(n1509) );
  NAND U1538 ( .A(n795), .B(n1383), .Z(n1501) );
  IV U1539 ( .A(n1503), .Z(n1515) );
  XNOR U1540 ( .A(n1516), .B(n1517), .Z(n1503) );
  AND U1541 ( .A(n1518), .B(n1519), .Z(n1517) );
  XOR U1542 ( .A(n1512), .B(n1520), .Z(n1519) );
  XNOR U1543 ( .A(n1514), .B(n1516), .Z(n1520) );
  NAND U1544 ( .A(n860), .B(n1383), .Z(n1514) );
  XOR U1545 ( .A(n1511), .B(n1521), .Z(n1512) );
  AND U1546 ( .A(n795), .B(X[0]), .Z(n1521) );
  XNOR U1547 ( .A(n1525), .B(n1522), .Z(n1524) );
  XOR U1548 ( .A(n1506), .B(n1526), .Z(n1518) );
  XNOR U1549 ( .A(n1508), .B(n1516), .Z(n1526) );
  NANDN U1550 ( .B(n996), .A(n1039), .Z(n1508) );
  XOR U1551 ( .A(n1505), .B(n1527), .Z(n1506) );
  AND U1552 ( .A(n1110), .B(n928), .Z(n1527) );
  XOR U1553 ( .A(n1528), .B(n1529), .Z(n1505) );
  AND U1554 ( .A(n1530), .B(n1531), .Z(n1529) );
  XNOR U1555 ( .A(n1532), .B(n1528), .Z(n1531) );
  XOR U1556 ( .A(n1533), .B(n1534), .Z(n1516) );
  AND U1557 ( .A(n1535), .B(n1536), .Z(n1534) );
  XOR U1558 ( .A(n1523), .B(n1537), .Z(n1536) );
  XNOR U1559 ( .A(n1525), .B(n1533), .Z(n1537) );
  NAND U1560 ( .A(n928), .B(n1383), .Z(n1525) );
  XOR U1561 ( .A(n1522), .B(n1538), .Z(n1523) );
  AND U1562 ( .A(n860), .B(X[0]), .Z(n1538) );
  XNOR U1563 ( .A(n1542), .B(n1539), .Z(n1541) );
  XOR U1564 ( .A(n1530), .B(n1543), .Z(n1535) );
  XNOR U1565 ( .A(n1532), .B(n1533), .Z(n1543) );
  NANDN U1566 ( .B(n1073), .A(n1039), .Z(n1532) );
  XOR U1567 ( .A(n1528), .B(n1544), .Z(n1530) );
  ANDN U1568 ( .A(n1110), .B(n996), .Z(n1544) );
  XOR U1569 ( .A(n1545), .B(n1546), .Z(n1528) );
  AND U1570 ( .A(n1547), .B(n1548), .Z(n1546) );
  XNOR U1571 ( .A(n1549), .B(n1545), .Z(n1548) );
  XOR U1572 ( .A(n1550), .B(n1551), .Z(n1533) );
  AND U1573 ( .A(n1552), .B(n1553), .Z(n1551) );
  XOR U1574 ( .A(n1540), .B(n1554), .Z(n1553) );
  XNOR U1575 ( .A(n1542), .B(n1550), .Z(n1554) );
  NANDN U1576 ( .B(n996), .A(n1383), .Z(n1542) );
  XOR U1577 ( .A(n1539), .B(n1555), .Z(n1540) );
  AND U1578 ( .A(n928), .B(X[0]), .Z(n1555) );
  XOR U1579 ( .A(n1547), .B(n1559), .Z(n1552) );
  XNOR U1580 ( .A(n1549), .B(n1550), .Z(n1559) );
  NAND U1581 ( .A(n1039), .B(n1146), .Z(n1549) );
  XOR U1582 ( .A(n1545), .B(n1560), .Z(n1547) );
  ANDN U1583 ( .A(n1110), .B(n1073), .Z(n1560) );
  NAND U1584 ( .A(n1039), .B(n1366), .Z(n1563) );
  XNOR U1585 ( .A(n1561), .B(n1565), .Z(n1562) );
  AND U1586 ( .A(n1146), .B(n1110), .Z(n1565) );
  AND U1587 ( .A(n1566), .B(A[0]), .Z(n1561) );
  NANDN U1588 ( .B(n1039), .A(n1567), .Z(n1566) );
  NAND U1589 ( .A(n1366), .B(n1110), .Z(n1567) );
  XNOR U1590 ( .A(n1556), .B(n1571), .Z(n1557) );
  ANDN U1591 ( .A(X[0]), .B(n996), .Z(n1571) );
  XOR U1592 ( .A(n1574), .B(n1572), .Z(n1573) );
  ANDN U1593 ( .A(X[0]), .B(n1073), .Z(n1574) );
  AND U1594 ( .A(n1383), .B(n1146), .Z(n1575) );
  XOR U1595 ( .A(n1579), .B(n1558), .Z(n1570) );
  NANDN U1596 ( .B(n1073), .A(n1383), .Z(n1558) );
  IV U1597 ( .A(n1564), .Z(n1579) );
  NAND U1598 ( .A(n1383), .B(n1366), .Z(n1578) );
  XNOR U1599 ( .A(n1576), .B(n1580), .Z(n1577) );
  AND U1600 ( .A(n1146), .B(X[0]), .Z(n1580) );
  AND U1601 ( .A(n1581), .B(A[0]), .Z(n1576) );
  NANDN U1602 ( .B(n1383), .A(n1582), .Z(n1581) );
  NAND U1603 ( .A(n1366), .B(X[0]), .Z(n1582) );
  XNOR U1604 ( .A(n1584), .B(n1136), .Z(n1126) );
  XNOR U1605 ( .A(n1123), .B(n1124), .Z(n1136) );
  NAND U1606 ( .A(n567), .B(n928), .Z(n1124) );
  XNOR U1607 ( .A(n1122), .B(n1585), .Z(n1123) );
  AND U1608 ( .A(n860), .B(n608), .Z(n1585) );
  XNOR U1609 ( .A(n1589), .B(n1586), .Z(n1588) );
  XNOR U1610 ( .A(n1135), .B(n1125), .Z(n1584) );
  XOR U1611 ( .A(n1590), .B(n1591), .Z(n1125) );
  XNOR U1612 ( .A(n1130), .B(n1593), .Z(n1131) );
  AND U1613 ( .A(n730), .B(n715), .Z(n1593) );
  XNOR U1614 ( .A(n1496), .B(A[8]), .Z(n1495) );
  NOR U1615 ( .A(n1594), .B(n1595), .Z(n1496) );
  XOR U1616 ( .A(n1596), .B(n1597), .Z(n1130) );
  AND U1617 ( .A(n1598), .B(n1599), .Z(n1597) );
  XNOR U1618 ( .A(n1600), .B(n1596), .Z(n1599) );
  XOR U1619 ( .A(n1601), .B(n1132), .Z(n1592) );
  NAND U1620 ( .A(n661), .B(n795), .Z(n1132) );
  IV U1621 ( .A(n1134), .Z(n1601) );
  XNOR U1622 ( .A(n1602), .B(n1603), .Z(n1134) );
  AND U1623 ( .A(n1604), .B(n1605), .Z(n1603) );
  XOR U1624 ( .A(n1598), .B(n1606), .Z(n1605) );
  XNOR U1625 ( .A(n1600), .B(n1602), .Z(n1606) );
  NAND U1626 ( .A(n661), .B(n860), .Z(n1600) );
  XOR U1627 ( .A(n1596), .B(n1607), .Z(n1598) );
  AND U1628 ( .A(n795), .B(n715), .Z(n1607) );
  XOR U1629 ( .A(n1594), .B(A[7]), .Z(n1595) );
  NANDN U1630 ( .B(n1608), .A(n1609), .Z(n1594) );
  XOR U1631 ( .A(n1610), .B(n1611), .Z(n1596) );
  AND U1632 ( .A(n1612), .B(n1613), .Z(n1611) );
  XNOR U1633 ( .A(n1614), .B(n1610), .Z(n1613) );
  XOR U1634 ( .A(n1587), .B(n1615), .Z(n1604) );
  XNOR U1635 ( .A(n1589), .B(n1602), .Z(n1615) );
  NANDN U1636 ( .B(n996), .A(n567), .Z(n1589) );
  XOR U1637 ( .A(n1586), .B(n1616), .Z(n1587) );
  AND U1638 ( .A(n928), .B(n608), .Z(n1616) );
  XNOR U1639 ( .A(n1620), .B(n1617), .Z(n1619) );
  XOR U1640 ( .A(n1621), .B(n1622), .Z(n1602) );
  AND U1641 ( .A(n1623), .B(n1624), .Z(n1622) );
  XOR U1642 ( .A(n1612), .B(n1625), .Z(n1624) );
  XNOR U1643 ( .A(n1614), .B(n1621), .Z(n1625) );
  NAND U1644 ( .A(n661), .B(n928), .Z(n1614) );
  XOR U1645 ( .A(n1610), .B(n1626), .Z(n1612) );
  AND U1646 ( .A(n860), .B(n715), .Z(n1626) );
  XNOR U1647 ( .A(n1609), .B(A[6]), .Z(n1608) );
  NOR U1648 ( .A(n1627), .B(n1628), .Z(n1609) );
  XOR U1649 ( .A(n1629), .B(n1630), .Z(n1610) );
  AND U1650 ( .A(n1631), .B(n1632), .Z(n1630) );
  XNOR U1651 ( .A(n1633), .B(n1629), .Z(n1632) );
  XOR U1652 ( .A(n1618), .B(n1634), .Z(n1623) );
  XNOR U1653 ( .A(n1620), .B(n1621), .Z(n1634) );
  NANDN U1654 ( .B(n1073), .A(n567), .Z(n1620) );
  XOR U1655 ( .A(n1617), .B(n1635), .Z(n1618) );
  ANDN U1656 ( .A(n608), .B(n996), .Z(n1635) );
  XNOR U1657 ( .A(n1639), .B(n1636), .Z(n1638) );
  XOR U1658 ( .A(n1640), .B(n1641), .Z(n1621) );
  AND U1659 ( .A(n1642), .B(n1643), .Z(n1641) );
  XOR U1660 ( .A(n1631), .B(n1644), .Z(n1643) );
  XNOR U1661 ( .A(n1633), .B(n1640), .Z(n1644) );
  NANDN U1662 ( .B(n996), .A(n661), .Z(n1633) );
  XOR U1663 ( .A(n1629), .B(n1645), .Z(n1631) );
  AND U1664 ( .A(n928), .B(n715), .Z(n1645) );
  XOR U1665 ( .A(n1627), .B(A[5]), .Z(n1628) );
  NANDN U1666 ( .B(n1646), .A(n1647), .Z(n1627) );
  XOR U1667 ( .A(n1648), .B(n1649), .Z(n1629) );
  ANDN U1668 ( .A(n1650), .B(n1651), .Z(n1649) );
  XNOR U1669 ( .A(n1652), .B(n1648), .Z(n1650) );
  XOR U1670 ( .A(n1637), .B(n1653), .Z(n1642) );
  XNOR U1671 ( .A(n1639), .B(n1640), .Z(n1653) );
  NAND U1672 ( .A(n567), .B(n1146), .Z(n1639) );
  XOR U1673 ( .A(n1636), .B(n1654), .Z(n1637) );
  ANDN U1674 ( .A(n608), .B(n1073), .Z(n1654) );
  XOR U1675 ( .A(n1655), .B(n1656), .Z(n1636) );
  ANDN U1676 ( .A(n1657), .B(n1658), .Z(n1656) );
  XNOR U1677 ( .A(n1659), .B(n1655), .Z(n1657) );
  NAND U1678 ( .A(n567), .B(n1366), .Z(n1659) );
  XNOR U1679 ( .A(n1655), .B(n1661), .Z(n1658) );
  AND U1680 ( .A(n1146), .B(n608), .Z(n1661) );
  AND U1681 ( .A(n1662), .B(A[0]), .Z(n1655) );
  NANDN U1682 ( .B(n567), .A(n1663), .Z(n1662) );
  NAND U1683 ( .A(n1366), .B(n608), .Z(n1663) );
  XNOR U1684 ( .A(n1648), .B(n1667), .Z(n1651) );
  ANDN U1685 ( .A(n715), .B(n996), .Z(n1667) );
  XOR U1686 ( .A(n1668), .B(n1669), .Z(n1648) );
  AND U1687 ( .A(n1670), .B(n1671), .Z(n1669) );
  XOR U1688 ( .A(n1672), .B(n1668), .Z(n1671) );
  ANDN U1689 ( .A(n715), .B(n1073), .Z(n1672) );
  XOR U1690 ( .A(n1673), .B(n1668), .Z(n1670) );
  AND U1691 ( .A(n1146), .B(n661), .Z(n1673) );
  XOR U1692 ( .A(n1674), .B(n1675), .Z(n1668) );
  ANDN U1693 ( .A(n1676), .B(n1677), .Z(n1675) );
  XNOR U1694 ( .A(n1678), .B(n1674), .Z(n1676) );
  XOR U1695 ( .A(n1679), .B(n1652), .Z(n1666) );
  NANDN U1696 ( .B(n1073), .A(n661), .Z(n1652) );
  IV U1697 ( .A(n1660), .Z(n1679) );
  XOR U1698 ( .A(n1680), .B(n1678), .Z(n1660) );
  NAND U1699 ( .A(n661), .B(n1366), .Z(n1678) );
  IV U1700 ( .A(n1677), .Z(n1680) );
  XNOR U1701 ( .A(n1674), .B(n1681), .Z(n1677) );
  AND U1702 ( .A(n1146), .B(n715), .Z(n1681) );
  AND U1703 ( .A(n1682), .B(A[0]), .Z(n1674) );
  NANDN U1704 ( .B(n661), .A(n1683), .Z(n1682) );
  NAND U1705 ( .A(n1366), .B(n715), .Z(n1683) );
  XNOR U1706 ( .A(n1139), .B(n1687), .Z(n1140) );
  ANDN U1707 ( .A(n535), .B(n996), .Z(n1687) );
  XNOR U1708 ( .A(n1647), .B(A[4]), .Z(n1646) );
  NOR U1709 ( .A(n1688), .B(n1689), .Z(n1647) );
  XOR U1710 ( .A(n1690), .B(n1691), .Z(n1139) );
  AND U1711 ( .A(n1692), .B(n1693), .Z(n1691) );
  XOR U1712 ( .A(n1694), .B(n1690), .Z(n1693) );
  ANDN U1713 ( .A(n535), .B(n1073), .Z(n1694) );
  XOR U1714 ( .A(n1695), .B(n1690), .Z(n1692) );
  AND U1715 ( .A(n1146), .B(n497), .Z(n1695) );
  XOR U1716 ( .A(n1696), .B(n1697), .Z(n1690) );
  ANDN U1717 ( .A(n1698), .B(n1699), .Z(n1697) );
  XNOR U1718 ( .A(n1700), .B(n1696), .Z(n1698) );
  XOR U1719 ( .A(n1701), .B(n1141), .Z(n1686) );
  NANDN U1720 ( .B(n1073), .A(n497), .Z(n1141) );
  NANDN U1721 ( .B(n1702), .A(n1703), .Z(n1688) );
  IV U1722 ( .A(n1143), .Z(n1701) );
  NAND U1723 ( .A(n497), .B(n1366), .Z(n1700) );
  XNOR U1724 ( .A(n1696), .B(n1704), .Z(n1699) );
  AND U1725 ( .A(n1146), .B(n535), .Z(n1704) );
  AND U1726 ( .A(n1705), .B(A[0]), .Z(n1696) );
  NANDN U1727 ( .B(n497), .A(n1706), .Z(n1705) );
  NAND U1728 ( .A(n1366), .B(n535), .Z(n1706) );
  XNOR U1729 ( .A(n1707), .B(X[12]), .Z(n535) );
  NAND U1730 ( .A(n1708), .B(X[15]), .Z(n1707) );
  XOR U1731 ( .A(n1709), .B(X[12]), .Z(n1708) );
  XNOR U1732 ( .A(n1150), .B(n1151), .Z(n1145) );
  NANDN U1733 ( .B(n442), .A(n1366), .Z(n1151) );
  XNOR U1734 ( .A(n1149), .B(n1711), .Z(n1150) );
  AND U1735 ( .A(n1146), .B(n466), .Z(n1711) );
  XNOR U1736 ( .A(n1703), .B(A[2]), .Z(n1702) );
  AND U1737 ( .A(n1713), .B(A[0]), .Z(n1149) );
  NAND U1738 ( .A(n1714), .B(n442), .Z(n1713) );
  NANDN U1739 ( .B(n1715), .A(n1716), .Z(n442) );
  ANDN U1740 ( .A(X[15]), .B(n1717), .Z(n1716) );
  NAND U1741 ( .A(n1366), .B(n466), .Z(n1714) );
  XOR U1742 ( .A(n1717), .B(X[14]), .Z(n1715) );
  OR U1743 ( .A(n1710), .B(n1718), .Z(n1717) );
  XOR U1744 ( .A(n1718), .B(X[13]), .Z(n1710) );
  OR U1745 ( .A(n1709), .B(n1719), .Z(n1718) );
  XOR U1746 ( .A(n1719), .B(X[12]), .Z(n1709) );
  OR U1747 ( .A(n1665), .B(n1720), .Z(n1719) );
  XOR U1748 ( .A(n1720), .B(X[11]), .Z(n1665) );
  OR U1749 ( .A(n1664), .B(n1721), .Z(n1720) );
  XOR U1750 ( .A(n1721), .B(X[10]), .Z(n1664) );
  OR U1751 ( .A(n1685), .B(n1722), .Z(n1721) );
  XOR U1752 ( .A(n1722), .B(X[9]), .Z(n1685) );
  OR U1753 ( .A(n1684), .B(n1723), .Z(n1722) );
  XOR U1754 ( .A(n1723), .B(X[8]), .Z(n1684) );
  OR U1755 ( .A(n1376), .B(n1724), .Z(n1723) );
  XOR U1756 ( .A(n1724), .B(X[7]), .Z(n1376) );
  OR U1757 ( .A(n1375), .B(n1725), .Z(n1724) );
  XOR U1758 ( .A(n1725), .B(X[6]), .Z(n1375) );
  OR U1759 ( .A(n1371), .B(n1726), .Z(n1725) );
  XOR U1760 ( .A(n1726), .B(X[5]), .Z(n1371) );
  OR U1761 ( .A(n1370), .B(n1727), .Z(n1726) );
  XOR U1762 ( .A(n1727), .B(X[4]), .Z(n1370) );
  OR U1763 ( .A(n1569), .B(n1728), .Z(n1727) );
  XOR U1764 ( .A(n1728), .B(X[3]), .Z(n1569) );
  OR U1765 ( .A(n1568), .B(n1729), .Z(n1728) );
  XOR U1766 ( .A(n1729), .B(X[2]), .Z(n1568) );
  NANDN U1767 ( .B(X[0]), .A(n1583), .Z(n1729) );
  XNOR U1768 ( .A(X[0]), .B(X[1]), .Z(n1583) );
  XOR U1769 ( .A(A[0]), .B(A[1]), .Z(n1712) );
  NANDN U1770 ( .B(n1085), .A(n357), .Z(n409) );
  IV U1771 ( .A(rst), .Z(n357) );
  NAND U1772 ( .A(n1730), .B(n1731), .Z(n1085) );
  AND U1773 ( .A(n1732), .B(n1733), .Z(n1731) );
  ANDN U1774 ( .A(n1734), .B(n[7]), .Z(n1733) );
  NOR U1775 ( .A(n[9]), .B(n[8]), .Z(n1734) );
  NOR U1776 ( .A(n[5]), .B(n[6]), .Z(n1732) );
  AND U1777 ( .A(n1735), .B(n1736), .Z(n1730) );
  NOR U1778 ( .A(n[1]), .B(n[2]), .Z(n1736) );
  NOR U1779 ( .A(n[0]), .B(n350), .Z(n1735) );
  OR U1780 ( .A(n[3]), .B(n[4]), .Z(n350) );
endmodule

