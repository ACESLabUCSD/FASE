
module MxM_TG_W16_N1000 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MxM/n97 , \_MxM/n94 , \_MxM/n91 , \_MxM/n88 , \_MxM/n85 ,
         \_MxM/n82 , \_MxM/n79 , \_MxM/n76 , \_MxM/n73 , \_MxM/n70 ,
         \_MxM/n67 , \_MxM/n64 , \_MxM/n61 , \_MxM/n58 , \_MxM/n55 ,
         \_MxM/n52 , \_MxM/N23 , \_MxM/N22 , \_MxM/N21 , \_MxM/N20 ,
         \_MxM/N19 , \_MxM/N18 , \_MxM/N17 , \_MxM/N16 , \_MxM/N15 ,
         \_MxM/N14 , \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 ,
         \_MxM/N7 , \_MxM/N6 , \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/Y1[0] , \_MxM/Y1[1] ,
         \_MxM/Y1[2] , \_MxM/Y1[3] , \_MxM/Y1[4] , \_MxM/Y1[5] , \_MxM/Y1[6] ,
         \_MxM/Y1[7] , \_MxM/Y1[8] , \_MxM/Y1[9] , \_MxM/Y1[10] ,
         \_MxM/Y1[11] , \_MxM/Y1[12] , \_MxM/Y1[13] , \_MxM/Y1[14] ,
         \_MxM/Y1[15] , \_MxM/Y0[15] , \_MxM/Y0[14] , \_MxM/Y0[13] ,
         \_MxM/Y0[12] , \_MxM/Y0[11] , \_MxM/Y0[10] , \_MxM/Y0[9] ,
         \_MxM/Y0[8] , \_MxM/Y0[7] , \_MxM/Y0[6] , \_MxM/Y0[5] , \_MxM/Y0[4] ,
         \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] , \_MxM/Y0[0] ,
         \_MxM/add_43/carry[9] , \_MxM/add_43/carry[8] ,
         \_MxM/add_43/carry[7] , \_MxM/add_43/carry[6] ,
         \_MxM/add_43/carry[5] , \_MxM/add_43/carry[4] ,
         \_MxM/add_43/carry[3] , \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380;

  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n52 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/Y1[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n55 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/Y1[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n58 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/Y1[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n61 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/Y1[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n64 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/Y1[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n67 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/Y1[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n70 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/Y1[9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n73 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/Y1[8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n76 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n79 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n82 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n85 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n88 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n91 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n94 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n97 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N14 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_43/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_43/carry[6] ), .COUT(\_MxM/add_43/carry[7] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_43/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_43/carry[7] ), .COUT(\_MxM/add_43/carry[8] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_43/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_43/carry[8] ), .COUT(\_MxM/add_43/carry[9] ), .SUM(\_MxM/N12 ) );
  MUX U1 ( .IN0(n1), .IN1(n1299), .SEL(n1300), .F(n1280) );
  IV U2 ( .A(n1301), .Z(n1) );
  MUX U3 ( .IN0(n2), .IN1(n844), .SEL(n845), .F(n823) );
  IV U4 ( .A(n846), .Z(n2) );
  XOR U5 ( .A(n1064), .B(n1054), .Z(n864) );
  MUX U6 ( .IN0(n998), .IN1(n1001), .SEL(n999), .F(n983) );
  XOR U7 ( .A(n1036), .B(n1037), .Z(n839) );
  MUX U8 ( .IN0(n3), .IN1(n559), .SEL(n560), .F(n498) );
  IV U9 ( .A(n561), .Z(n3) );
  MUX U10 ( .IN0(e_input[12]), .IN1(n1351), .SEL(e_input[15]), .F(n226) );
  MUX U11 ( .IN0(n1280), .IN1(n1298), .SEL(n1282), .F(n1260) );
  XOR U12 ( .A(n1046), .B(n1047), .Z(n862) );
  MUX U13 ( .IN0(n4), .IN1(n804), .SEL(n805), .F(n737) );
  IV U14 ( .A(n806), .Z(n4) );
  XOR U15 ( .A(n847), .B(n829), .Z(n833) );
  MUX U16 ( .IN0(n1041), .IN1(n5), .SEL(n1040), .F(n1030) );
  IV U17 ( .A(n1039), .Z(n5) );
  MUX U18 ( .IN0(e_input[8]), .IN1(n1327), .SEL(e_input[15]), .F(n385) );
  XNOR U19 ( .A(n1329), .B(n779), .Z(n783) );
  MUX U20 ( .IN0(n6), .IN1(n1085), .SEL(n1086), .F(n1068) );
  IV U21 ( .A(n1087), .Z(n6) );
  MUX U22 ( .IN0(n1229), .IN1(n1259), .SEL(n1231), .F(n757) );
  XOR U23 ( .A(n805), .B(n806), .Z(n802) );
  MUX U24 ( .IN0(n7), .IN1(n1035), .SEL(n1036), .F(n811) );
  IV U25 ( .A(n1037), .Z(n7) );
  MUX U26 ( .IN0(n8), .IN1(n440), .SEL(n441), .F(n386) );
  IV U27 ( .A(n442), .Z(n8) );
  MUX U28 ( .IN0(n601), .IN1(n9), .SEL(n600), .F(n536) );
  IV U29 ( .A(n599), .Z(n9) );
  MUX U30 ( .IN0(e_input[13]), .IN1(n1352), .SEL(e_input[15]), .F(n191) );
  MUX U31 ( .IN0(n10), .IN1(n1045), .SEL(n1046), .F(n1035) );
  IV U32 ( .A(n1047), .Z(n10) );
  MUX U33 ( .IN0(n11), .IN1(n1053), .SEL(n1054), .F(n1039) );
  IV U34 ( .A(n1055), .Z(n11) );
  MUX U35 ( .IN0(n12), .IN1(n737), .SEL(n738), .F(n667) );
  IV U36 ( .A(n739), .Z(n12) );
  MUX U37 ( .IN0(n13), .IN1(n729), .SEL(n730), .F(n659) );
  IV U38 ( .A(n731), .Z(n13) );
  MUX U39 ( .IN0(n14), .IN1(n551), .SEL(n552), .F(n490) );
  IV U40 ( .A(n553), .Z(n14) );
  MUX U41 ( .IN0(e_input[9]), .IN1(n1328), .SEL(e_input[15]), .F(n338) );
  MUX U42 ( .IN0(n576), .IN1(n574), .SEL(n575), .F(n513) );
  MUX U43 ( .IN0(n229), .IN1(n15), .SEL(n228), .F(n193) );
  IV U44 ( .A(n227), .Z(n15) );
  MUX U45 ( .IN0(n16), .IN1(n1197), .SEL(n1198), .F(n1180) );
  IV U46 ( .A(n1199), .Z(n16) );
  XOR U47 ( .A(n824), .B(n825), .Z(n834) );
  MUX U48 ( .IN0(n17), .IN1(n757), .SEL(n758), .F(n688) );
  IV U49 ( .A(n759), .Z(n17) );
  MUX U50 ( .IN0(n18), .IN1(n696), .SEL(n697), .F(n622) );
  IV U51 ( .A(n698), .Z(n18) );
  MUX U52 ( .IN0(n19), .IN1(n659), .SEL(n660), .F(n599) );
  IV U53 ( .A(n661), .Z(n19) );
  MUX U54 ( .IN0(g_input[11]), .IN1(n1084), .SEL(g_input[15]), .F(n270) );
  XOR U55 ( .A(n748), .B(n749), .Z(n754) );
  MUX U56 ( .IN0(n502), .IN1(n504), .SEL(n503), .F(n444) );
  MUX U57 ( .IN0(n539), .IN1(n20), .SEL(n538), .F(n473) );
  IV U58 ( .A(n537), .Z(n20) );
  XNOR U59 ( .A(n774), .B(n708), .Z(n712) );
  XOR U60 ( .A(n845), .B(n846), .Z(n857) );
  MUX U61 ( .IN0(g_input[1]), .IN1(n1354), .SEL(g_input[15]), .F(n1008) );
  XOR U62 ( .A(n1038), .B(n1030), .Z(n820) );
  MUX U63 ( .IN0(g_input[2]), .IN1(n1345), .SEL(g_input[15]), .F(n785) );
  MUX U64 ( .IN0(n21), .IN1(n614), .SEL(n615), .F(n551) );
  IV U65 ( .A(n616), .Z(n21) );
  MUX U66 ( .IN0(n22), .IN1(n498), .SEL(n499), .F(n440) );
  IV U67 ( .A(n500), .Z(n22) );
  MUX U68 ( .IN0(g_input[10]), .IN1(n1100), .SEL(g_input[15]), .F(n310) );
  MUX U69 ( .IN0(n749), .IN1(n23), .SEL(n748), .F(n677) );
  IV U70 ( .A(n747), .Z(n23) );
  MUX U71 ( .IN0(n457), .IN1(n455), .SEL(n456), .F(n397) );
  MUX U72 ( .IN0(n380), .IN1(n382), .SEL(n381), .F(n24) );
  IV U73 ( .A(n24), .Z(n341) );
  XNOR U74 ( .A(n727), .B(n660), .Z(n664) );
  XNOR U75 ( .A(n703), .B(n636), .Z(n640) );
  MUX U76 ( .IN0(n1215), .IN1(n1218), .SEL(n1216), .F(n1197) );
  XOR U77 ( .A(n1300), .B(n1301), .Z(n1233) );
  XOR U78 ( .A(n812), .B(n813), .Z(n818) );
  MUX U79 ( .IN0(n25), .IN1(n667), .SEL(n668), .F(n603) );
  IV U80 ( .A(n669), .Z(n25) );
  MUX U81 ( .IN0(g_input[9]), .IN1(n1120), .SEL(g_input[15]), .F(n353) );
  XNOR U82 ( .A(n792), .B(n730), .Z(n734) );
  MUX U83 ( .IN0(n444), .IN1(n446), .SEL(n445), .F(n380) );
  MUX U84 ( .IN0(n399), .IN1(n397), .SEL(n398), .F(n350) );
  MUX U85 ( .IN0(n388), .IN1(n26), .SEL(n387), .F(n340) );
  IV U86 ( .A(n386), .Z(n26) );
  XNOR U87 ( .A(n631), .B(n571), .Z(n575) );
  NAND U88 ( .A(n536), .B(n597), .Z(n596) );
  MUX U89 ( .IN0(n27), .IN1(n992), .SEL(n808), .F(n965) );
  IV U90 ( .A(n807), .Z(n27) );
  MUX U91 ( .IN0(n1163), .IN1(n1179), .SEL(n1165), .F(n1152) );
  MUX U92 ( .IN0(n28), .IN1(n811), .SEL(n812), .F(n747) );
  IV U93 ( .A(n813), .Z(n28) );
  MUX U94 ( .IN0(n29), .IN1(n603), .SEL(n604), .F(n541) );
  IV U95 ( .A(n605), .Z(n29) );
  XOR U96 ( .A(n717), .B(n786), .Z(n718) );
  MUX U97 ( .IN0(n352), .IN1(n350), .SEL(n351), .F(n307) );
  MUX U98 ( .IN0(e_input[10]), .IN1(n1306), .SEL(e_input[15]), .F(n289) );
  XOR U99 ( .A(n592), .B(n537), .Z(n538) );
  XNOR U100 ( .A(n566), .B(n510), .Z(n514) );
  XOR U101 ( .A(n438), .B(n387), .Z(n381) );
  MUX U102 ( .IN0(n427), .IN1(n429), .SEL(n428), .F(n30) );
  IV U103 ( .A(n30), .Z(n368) );
  XOR U104 ( .A(n583), .B(n586), .Z(n584) );
  MUX U105 ( .IN0(n935), .IN1(n31), .SEL(n936), .F(n908) );
  IV U106 ( .A(n937), .Z(n31) );
  MUX U107 ( .IN0(n32), .IN1(n1068), .SEL(n1069), .F(n1053) );
  IV U108 ( .A(n1070), .Z(n32) );
  XOR U109 ( .A(n1131), .B(n1132), .Z(n994) );
  MUX U110 ( .IN0(n628), .IN1(n630), .SEL(n629), .F(n563) );
  XOR U111 ( .A(n461), .B(n517), .Z(n462) );
  MUX U112 ( .IN0(e_input[6]), .IN1(n1017), .SEL(e_input[15]), .F(n478) );
  MUX U113 ( .IN0(n33), .IN1(n329), .SEL(n330), .F(n290) );
  IV U114 ( .A(n331), .Z(n33) );
  XNOR U115 ( .A(n657), .B(n600), .Z(n594) );
  MUX U116 ( .IN0(n34), .IN1(n554), .SEL(n555), .F(n493) );
  IV U117 ( .A(n556), .Z(n34) );
  XNOR U118 ( .A(n505), .B(n452), .Z(n456) );
  NAND U119 ( .A(n340), .B(n384), .Z(n383) );
  XOR U120 ( .A(n522), .B(n525), .Z(n523) );
  MUX U121 ( .IN0(n35), .IN1(n1121), .SEL(n1122), .F(n1102) );
  IV U122 ( .A(n1123), .Z(n35) );
  MUX U123 ( .IN0(n36), .IN1(n1019), .SEL(n1020), .F(n1191) );
  IV U124 ( .A(n1207), .Z(n36) );
  MUX U125 ( .IN0(n1146), .IN1(n1168), .SEL(n1148), .F(n1128) );
  XOR U126 ( .A(n826), .B(n797), .Z(n801) );
  MUX U127 ( .IN0(g_input[3]), .IN1(n1332), .SEL(g_input[15]), .F(n37) );
  IV U128 ( .A(n37), .Z(n714) );
  MUX U129 ( .IN0(n38), .IN1(n688), .SEL(n689), .F(n614) );
  IV U130 ( .A(n690), .Z(n38) );
  MUX U131 ( .IN0(n784), .IN1(n782), .SEL(n783), .F(n711) );
  XOR U132 ( .A(n580), .B(n643), .Z(n581) );
  MUX U133 ( .IN0(n563), .IN1(n565), .SEL(n564), .F(n502) );
  MUX U134 ( .IN0(n269), .IN1(n267), .SEL(n268), .F(n219) );
  MUX U135 ( .IN0(g_input[12]), .IN1(n1066), .SEL(g_input[15]), .F(n230) );
  XOR U136 ( .A(n480), .B(n481), .Z(n475) );
  MUX U137 ( .IN0(n39), .IN1(n435), .SEL(n436), .F(n376) );
  IV U138 ( .A(n437), .Z(n39) );
  XNOR U139 ( .A(n447), .B(n394), .Z(n398) );
  XNOR U140 ( .A(n296), .B(n335), .Z(n297) );
  MUX U141 ( .IN0(n670), .IN1(n40), .SEL(n671), .F(n606) );
  IV U142 ( .A(n672), .Z(n40) );
  MUX U143 ( .IN0(n41), .IN1(n316), .SEL(n110), .F(n276) );
  IV U144 ( .A(\_MxM/Y0[8] ), .Z(n41) );
  XOR U145 ( .A(n464), .B(n467), .Z(n465) );
  MUX U146 ( .IN0(n1089), .IN1(n42), .SEL(n917), .F(n1072) );
  IV U147 ( .A(n915), .Z(n42) );
  MUX U148 ( .IN0(e_input[1]), .IN1(n43), .SEL(e_input[15]), .F(n1025) );
  IV U149 ( .A(n1226), .Z(n43) );
  MUX U150 ( .IN0(n832), .IN1(n44), .SEL(n833), .F(n800) );
  IV U151 ( .A(n834), .Z(n44) );
  XNOR U152 ( .A(n1005), .B(n1006), .Z(n989) );
  MUX U153 ( .IN0(n771), .IN1(n773), .SEL(n772), .F(n700) );
  MUX U154 ( .IN0(e_input[2]), .IN1(n1211), .SEL(e_input[15]), .F(n746) );
  MUX U155 ( .IN0(n515), .IN1(n513), .SEL(n514), .F(n455) );
  XOR U156 ( .A(n356), .B(n401), .Z(n357) );
  MUX U157 ( .IN0(n45), .IN1(n750), .SEL(n751), .F(n683) );
  IV U158 ( .A(n752), .Z(n45) );
  MUX U159 ( .IN0(n46), .IN1(n691), .SEL(n692), .F(n617) );
  IV U160 ( .A(n693), .Z(n46) );
  XOR U161 ( .A(n557), .B(n499), .Z(n503) );
  MUX U162 ( .IN0(n47), .IN1(n479), .SEL(n480), .F(n426) );
  IV U163 ( .A(n481), .Z(n47) );
  MUX U164 ( .IN0(n48), .IN1(n376), .SEL(n377), .F(n332) );
  IV U165 ( .A(n378), .Z(n48) );
  NAND U166 ( .A(n250), .B(n288), .Z(n287) );
  XNOR U167 ( .A(n299), .B(n264), .Z(n268) );
  MUX U168 ( .IN0(n49), .IN1(n548), .SEL(n547), .F(n485) );
  IV U169 ( .A(n546), .Z(n49) );
  MUX U170 ( .IN0(n50), .IN1(n202), .SEL(n203), .F(n172) );
  IV U171 ( .A(\_MxM/Y0[11] ), .Z(n50) );
  XOR U172 ( .A(n406), .B(n409), .Z(n407) );
  MUX U173 ( .IN0(n962), .IN1(n51), .SEL(n963), .F(n935) );
  IV U174 ( .A(n964), .Z(n51) );
  MUX U175 ( .IN0(n1125), .IN1(n52), .SEL(n971), .F(n1108) );
  IV U176 ( .A(n969), .Z(n52) );
  MUX U177 ( .IN0(n855), .IN1(n53), .SEL(n856), .F(n832) );
  IV U178 ( .A(n857), .Z(n53) );
  MUX U179 ( .IN0(n1057), .IN1(n54), .SEL(n864), .F(n1043) );
  IV U180 ( .A(n862), .Z(n54) );
  XOR U181 ( .A(n1213), .B(n1198), .Z(n1020) );
  MUX U182 ( .IN0(e_input[4]), .IN1(n1012), .SEL(e_input[15]), .F(n598) );
  XOR U183 ( .A(n1235), .B(n768), .Z(n772) );
  MUX U184 ( .IN0(n665), .IN1(n663), .SEL(n664), .F(n593) );
  MUX U185 ( .IN0(n55), .IN1(n541), .SEL(n542), .F(n479) );
  IV U186 ( .A(n543), .Z(n55) );
  MUX U187 ( .IN0(e_input[11]), .IN1(n1307), .SEL(e_input[15]), .F(n253) );
  MUX U188 ( .IN0(n56), .IN1(n617), .SEL(n618), .F(n554) );
  IV U189 ( .A(n619), .Z(n56) );
  XNOR U190 ( .A(n259), .B(n228), .Z(n222) );
  MUX U191 ( .IN0(n57), .IN1(n256), .SEL(n257), .F(n214) );
  IV U192 ( .A(n258), .Z(n57) );
  MUX U193 ( .IN0(e_input[14]), .IN1(n1357), .SEL(e_input[15]), .F(n161) );
  XNOR U194 ( .A(n609), .B(n673), .Z(n610) );
  MUX U195 ( .IN0(n485), .IN1(n487), .SEL(n486), .F(n427) );
  MUX U196 ( .IN0(n58), .IN1(n648), .SEL(n116), .F(n583) );
  IV U197 ( .A(\_MxM/Y0[2] ), .Z(n58) );
  XNOR U198 ( .A(n172), .B(n173), .Z(n130) );
  XOR U199 ( .A(n360), .B(n366), .Z(n111) );
  MUX U200 ( .IN0(n1108), .IN1(n59), .SEL(n944), .F(n1089) );
  IV U201 ( .A(n942), .Z(n59) );
  MUX U202 ( .IN0(n60), .IN1(n1219), .SEL(n1220), .F(n1215) );
  IV U203 ( .A(n1221), .Z(n60) );
  MUX U204 ( .IN0(n1043), .IN1(n61), .SEL(n841), .F(n1031) );
  IV U205 ( .A(n839), .Z(n61) );
  MUX U206 ( .IN0(n800), .IN1(n62), .SEL(n801), .F(n733) );
  IV U207 ( .A(n802), .Z(n62) );
  XNOR U208 ( .A(n996), .B(n986), .Z(n990) );
  MUX U209 ( .IN0(g_input[5]), .IN1(n1272), .SEL(g_input[15]), .F(n577) );
  MUX U210 ( .IN0(n713), .IN1(n711), .SEL(n712), .F(n639) );
  MUX U211 ( .IN0(n343), .IN1(n63), .SEL(n342), .F(n296) );
  IV U212 ( .A(n341), .Z(n63) );
  XOR U213 ( .A(n273), .B(n311), .Z(n274) );
  MUX U214 ( .IN0(n64), .IN1(n760), .SEL(n761), .F(n691) );
  IV U215 ( .A(n762), .Z(n64) );
  NAND U216 ( .A(n677), .B(n745), .Z(n744) );
  XOR U217 ( .A(n694), .B(n625), .Z(n629) );
  XOR U218 ( .A(n542), .B(n543), .Z(n539) );
  MUX U219 ( .IN0(n65), .IN1(n493), .SEL(n494), .F(n435) );
  IV U220 ( .A(n495), .Z(n65) );
  XNOR U221 ( .A(n389), .B(n347), .Z(n351) );
  MUX U222 ( .IN0(n66), .IN1(n293), .SEL(n294), .F(n256) );
  IV U223 ( .A(n295), .Z(n66) );
  MUX U224 ( .IN0(n292), .IN1(n67), .SEL(n291), .F(n250) );
  IV U225 ( .A(n290), .Z(n67) );
  XNOR U226 ( .A(n219), .B(n220), .Z(n218) );
  XNOR U227 ( .A(n595), .B(n594), .Z(n611) );
  XNOR U228 ( .A(n223), .B(n222), .Z(n216) );
  XOR U229 ( .A(n472), .B(n420), .Z(n428) );
  MUX U230 ( .IN0(n68), .IN1(n522), .SEL(n114), .F(n464) );
  IV U231 ( .A(\_MxM/Y0[4] ), .Z(n68) );
  MUX U232 ( .IN0(\_MxM/Y0[13] ), .IN1(n130), .SEL(n129), .F(n126) );
  XOR U233 ( .A(n276), .B(n279), .Z(n277) );
  XOR U234 ( .A(n1150), .B(n1141), .Z(n995) );
  MUX U235 ( .IN0(n69), .IN1(n432), .SEL(n433), .F(n373) );
  IV U236 ( .A(n434), .Z(n69) );
  MUX U237 ( .IN0(e_input[3]), .IN1(n1212), .SEL(e_input[15]), .F(n680) );
  MUX U238 ( .IN0(n641), .IN1(n639), .SEL(n640), .F(n574) );
  MUX U239 ( .IN0(e_input[5]), .IN1(n1013), .SEL(e_input[15]), .F(n534) );
  MUX U240 ( .IN0(n309), .IN1(n307), .SEL(n308), .F(n267) );
  XOR U241 ( .A(n763), .B(n697), .Z(n701) );
  XNOR U242 ( .A(n784), .B(n783), .Z(n762) );
  MUX U243 ( .IN0(n685), .IN1(n70), .SEL(n684), .F(n609) );
  IV U244 ( .A(n683), .Z(n70) );
  MUX U245 ( .IN0(e_input[7]), .IN1(n1018), .SEL(e_input[15]), .F(n418) );
  MUX U246 ( .IN0(n298), .IN1(n296), .SEL(n297), .F(n71) );
  IV U247 ( .A(n71), .Z(n255) );
  NAND U248 ( .A(n193), .B(n225), .Z(n224) );
  XOR U249 ( .A(n199), .B(n231), .Z(n200) );
  MUX U250 ( .IN0(n606), .IN1(n72), .SEL(n607), .F(n546) );
  IV U251 ( .A(n608), .Z(n72) );
  XNOR U252 ( .A(n399), .B(n398), .Z(n378) );
  MUX U253 ( .IN0(n216), .IN1(n73), .SEL(n215), .F(n187) );
  IV U254 ( .A(n214), .Z(n73) );
  XNOR U255 ( .A(n495), .B(n494), .Z(n487) );
  MUX U256 ( .IN0(n74), .IN1(n464), .SEL(n113), .F(n406) );
  IV U257 ( .A(\_MxM/Y0[5] ), .Z(n74) );
  MUX U258 ( .IN0(n75), .IN1(n276), .SEL(n109), .F(n236) );
  IV U259 ( .A(\_MxM/Y0[9] ), .Z(n75) );
  MUX U260 ( .IN0(n76), .IN1(n124), .SEL(n123), .F(n128) );
  IV U261 ( .A(n131), .Z(n76) );
  MUX U262 ( .IN0(n908), .IN1(n77), .SEL(n909), .F(n881) );
  IV U263 ( .A(n910), .Z(n77) );
  MUX U264 ( .IN0(n1187), .IN1(n1201), .SEL(n1189), .F(n1169) );
  XNOR U265 ( .A(n1220), .B(n1221), .Z(n1207) );
  XOR U266 ( .A(n1331), .B(g_input[3]), .Z(n1332) );
  MUX U267 ( .IN0(g_input[6]), .IN1(n1251), .SEL(g_input[15]), .F(n516) );
  MUX U268 ( .IN0(n78), .IN1(n490), .SEL(n491), .F(n432) );
  IV U269 ( .A(n492), .Z(n78) );
  MUX U270 ( .IN0(g_input[7]), .IN1(n1238), .SEL(g_input[15]), .F(n458) );
  MUX U271 ( .IN0(g_input[8]), .IN1(n1136), .SEL(g_input[15]), .F(n400) );
  XNOR U272 ( .A(n1031), .B(n1032), .Z(n1021) );
  XNOR U273 ( .A(n991), .B(n990), .Z(n807) );
  MUX U274 ( .IN0(n595), .IN1(n593), .SEL(n594), .F(n537) );
  XNOR U275 ( .A(n735), .B(n734), .Z(n752) );
  XOR U276 ( .A(n620), .B(n560), .Z(n564) );
  MUX U277 ( .IN0(n79), .IN1(n332), .SEL(n333), .F(n293) );
  IV U278 ( .A(n334), .Z(n79) );
  XNOR U279 ( .A(n344), .B(n304), .Z(n308) );
  MUX U280 ( .IN0(g_input[13]), .IN1(n1052), .SEL(g_input[15]), .F(n196) );
  XNOR U281 ( .A(n665), .B(n664), .Z(n685) );
  XNOR U282 ( .A(n762), .B(n761), .Z(n742) );
  XNOR U283 ( .A(n641), .B(n640), .Z(n619) );
  XNOR U284 ( .A(n576), .B(n575), .Z(n556) );
  AND U285 ( .A(n156), .B(n137), .Z(n155) );
  XNOR U286 ( .A(n693), .B(n692), .Z(n672) );
  XNOR U287 ( .A(n485), .B(n484), .Z(n530) );
  MUX U288 ( .IN0(n80), .IN1(n583), .SEL(n115), .F(n522) );
  IV U289 ( .A(\_MxM/Y0[3] ), .Z(n80) );
  XNOR U290 ( .A(n437), .B(n436), .Z(n429) );
  XNOR U291 ( .A(n378), .B(n377), .Z(n370) );
  MUX U292 ( .IN0(n81), .IN1(n359), .SEL(n111), .F(n316) );
  IV U293 ( .A(\_MxM/Y0[7] ), .Z(n81) );
  XNOR U294 ( .A(n186), .B(n187), .Z(n185) );
  XOR U295 ( .A(n236), .B(n239), .Z(n237) );
  MUX U296 ( .IN0(\_MxM/Y0[14] ), .IN1(n126), .SEL(n127), .F(n120) );
  MUX U297 ( .IN0(n991), .IN1(n989), .SEL(n990), .F(n962) );
  MUX U298 ( .IN0(n1144), .IN1(n82), .SEL(n995), .F(n1125) );
  IV U299 ( .A(n994), .Z(n82) );
  MUX U300 ( .IN0(n83), .IN1(n1233), .SEL(n1234), .F(n1284) );
  IV U301 ( .A(n1302), .Z(n83) );
  MUX U302 ( .IN0(n881), .IN1(n84), .SEL(n882), .F(n855) );
  IV U303 ( .A(n883), .Z(n84) );
  NOR U304 ( .A(g_input[0]), .B(n1354), .Z(n1346) );
  MUX U305 ( .IN0(n1072), .IN1(n85), .SEL(n890), .F(n1057) );
  IV U306 ( .A(n888), .Z(n85) );
  MUX U307 ( .IN0(n86), .IN1(n823), .SEL(n824), .F(n804) );
  IV U308 ( .A(n825), .Z(n86) );
  MUX U309 ( .IN0(n87), .IN1(n828), .SEL(n829), .F(n794) );
  IV U310 ( .A(n830), .Z(n87) );
  MUX U311 ( .IN0(n1152), .IN1(n1162), .SEL(n1154), .F(n1138) );
  XOR U312 ( .A(n1205), .B(n1206), .Z(n1019) );
  MUX U313 ( .IN0(g_input[4]), .IN1(n1290), .SEL(g_input[15]), .F(n88) );
  IV U314 ( .A(n88), .Z(n642) );
  MUX U315 ( .IN0(n89), .IN1(n346), .SEL(n347), .F(n301) );
  IV U316 ( .A(n348), .Z(n89) );
  MUX U317 ( .IN0(n90), .IN1(n373), .SEL(n374), .F(n329) );
  IV U318 ( .A(n375), .Z(n90) );
  MUX U319 ( .IN0(n735), .IN1(n733), .SEL(n734), .F(n663) );
  MUX U320 ( .IN0(n700), .IN1(n702), .SEL(n701), .F(n628) );
  MUX U321 ( .IN0(n754), .IN1(n1021), .SEL(n753), .F(n682) );
  XOR U322 ( .A(n496), .B(n441), .Z(n445) );
  MUX U323 ( .IN0(n475), .IN1(n473), .SEL(n474), .F(n424) );
  XNOR U324 ( .A(n713), .B(n712), .Z(n693) );
  MUX U325 ( .IN0(n740), .IN1(n91), .SEL(n741), .F(n670) );
  IV U326 ( .A(n742), .Z(n91) );
  MUX U327 ( .IN0(n611), .IN1(n609), .SEL(n610), .F(n92) );
  IV U328 ( .A(n92), .Z(n545) );
  XNOR U329 ( .A(n515), .B(n514), .Z(n495) );
  XNOR U330 ( .A(n457), .B(n456), .Z(n437) );
  XNOR U331 ( .A(n352), .B(n351), .Z(n334) );
  XNOR U332 ( .A(n309), .B(n308), .Z(n295) );
  XNOR U333 ( .A(n269), .B(n268), .Z(n258) );
  MUX U334 ( .IN0(n195), .IN1(n218), .SEL(n194), .F(n167) );
  MUX U335 ( .IN0(g_input[14]), .IN1(n1026), .SEL(g_input[15]), .F(n162) );
  XNOR U336 ( .A(n619), .B(n618), .Z(n608) );
  XNOR U337 ( .A(n556), .B(n555), .Z(n548) );
  MUX U338 ( .IN0(n368), .IN1(n93), .SEL(n369), .F(n326) );
  IV U339 ( .A(n370), .Z(n93) );
  MUX U340 ( .IN0(n94), .IN1(n406), .SEL(n112), .F(n359) );
  IV U341 ( .A(\_MxM/Y0[6] ), .Z(n94) );
  MUX U342 ( .IN0(n95), .IN1(n236), .SEL(n108), .F(n202) );
  IV U343 ( .A(\_MxM/Y0[10] ), .Z(n95) );
  MUX U344 ( .IN0(n96), .IN1(n720), .SEL(n721), .F(n648) );
  IV U345 ( .A(\_MxM/Y0[1] ), .Z(n96) );
  XNOR U346 ( .A(n185), .B(n184), .Z(n206) );
  MUX U347 ( .IN0(\_MxM/Y0[15] ), .IN1(n120), .SEL(n121), .F(n97) );
  IV U348 ( .A(n97), .Z(n117) );
  MUX U349 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n98), .F(\_MxM/n97 ) );
  MUX U350 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n98), .F(\_MxM/n94 ) );
  MUX U351 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n98), .F(\_MxM/n91 ) );
  MUX U352 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n98), .F(\_MxM/n88 ) );
  MUX U353 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n98), .F(\_MxM/n85 ) );
  MUX U354 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n98), .F(\_MxM/n82 ) );
  MUX U355 ( .IN0(\_MxM/Y1[6] ), .IN1(o[6]), .SEL(n98), .F(\_MxM/n79 ) );
  MUX U356 ( .IN0(\_MxM/Y1[7] ), .IN1(o[7]), .SEL(n98), .F(\_MxM/n76 ) );
  MUX U357 ( .IN0(\_MxM/Y1[8] ), .IN1(o[8]), .SEL(n98), .F(\_MxM/n73 ) );
  MUX U358 ( .IN0(\_MxM/Y1[9] ), .IN1(o[9]), .SEL(n98), .F(\_MxM/n70 ) );
  MUX U359 ( .IN0(\_MxM/Y1[10] ), .IN1(o[10]), .SEL(n98), .F(\_MxM/n67 ) );
  MUX U360 ( .IN0(\_MxM/Y1[11] ), .IN1(o[11]), .SEL(n98), .F(\_MxM/n64 ) );
  MUX U361 ( .IN0(\_MxM/Y1[12] ), .IN1(o[12]), .SEL(n98), .F(\_MxM/n61 ) );
  MUX U362 ( .IN0(\_MxM/Y1[13] ), .IN1(o[13]), .SEL(n98), .F(\_MxM/n58 ) );
  IV U363 ( .A(n99), .Z(n98) );
  MUX U364 ( .IN0(o[14]), .IN1(\_MxM/Y1[14] ), .SEL(n99), .F(\_MxM/n55 ) );
  MUX U365 ( .IN0(o[15]), .IN1(\_MxM/Y1[15] ), .SEL(n99), .F(\_MxM/n52 ) );
  AND U366 ( .A(n100), .B(n101), .Z(n99) );
  AND U367 ( .A(n102), .B(n103), .Z(n101) );
  ANDN U368 ( .A(n104), .B(\_MxM/n[7] ), .Z(n103) );
  NOR U369 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n104) );
  NOR U370 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n102) );
  AND U371 ( .A(n105), .B(n106), .Z(n100) );
  NOR U372 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n106) );
  NOR U373 ( .A(\_MxM/n[0] ), .B(n107), .Z(n105) );
  XNOR U374 ( .A(n108), .B(\_MxM/Y0[10] ), .Z(\_MxM/Y1[9] ) );
  XNOR U375 ( .A(n109), .B(\_MxM/Y0[9] ), .Z(\_MxM/Y1[8] ) );
  XNOR U376 ( .A(n110), .B(\_MxM/Y0[8] ), .Z(\_MxM/Y1[7] ) );
  XNOR U377 ( .A(n111), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XNOR U378 ( .A(n112), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XNOR U379 ( .A(n113), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U380 ( .A(n114), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U381 ( .A(n115), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U382 ( .A(n116), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U383 ( .A(n117), .B(n118), .Z(\_MxM/Y1[15] ) );
  XNOR U384 ( .A(\_MxM/Y0[15] ), .B(n119), .Z(n118) );
  XNOR U385 ( .A(n121), .B(\_MxM/Y0[15] ), .Z(\_MxM/Y1[14] ) );
  XOR U386 ( .A(n120), .B(n119), .Z(n121) );
  NAND U387 ( .A(n122), .B(n123), .Z(n119) );
  OR U388 ( .A(n124), .B(n125), .Z(n122) );
  XNOR U389 ( .A(n127), .B(\_MxM/Y0[14] ), .Z(\_MxM/Y1[13] ) );
  XNOR U390 ( .A(n128), .B(n126), .Z(n127) );
  XNOR U391 ( .A(n125), .B(n131), .Z(n124) );
  OR U392 ( .A(n132), .B(n133), .Z(n125) );
  AND U393 ( .A(n134), .B(n135), .Z(n131) );
  OR U394 ( .A(n136), .B(n137), .Z(n135) );
  AND U395 ( .A(n138), .B(n139), .Z(n134) );
  OR U396 ( .A(n140), .B(n141), .Z(n139) );
  OR U397 ( .A(n142), .B(n143), .Z(n138) );
  XNOR U398 ( .A(n129), .B(\_MxM/Y0[13] ), .Z(\_MxM/Y1[12] ) );
  XNOR U399 ( .A(n144), .B(n145), .Z(n129) );
  XNOR U400 ( .A(n130), .B(n146), .Z(n144) );
  AND U401 ( .A(n123), .B(n147), .Z(n146) );
  XOR U402 ( .A(n132), .B(n148), .Z(n147) );
  XOR U403 ( .A(n148), .B(n133), .Z(n132) );
  OR U404 ( .A(n149), .B(n150), .Z(n133) );
  IV U405 ( .A(n145), .Z(n148) );
  XNOR U406 ( .A(n143), .B(n142), .Z(n145) );
  OR U407 ( .A(n151), .B(n152), .Z(n142) );
  AND U408 ( .A(n153), .B(n154), .Z(n143) );
  XNOR U409 ( .A(n136), .B(n155), .Z(n154) );
  NAND U410 ( .A(n157), .B(n158), .Z(n137) );
  NANDN U411 ( .B(n159), .A(n160), .Z(n157) );
  NANDN U412 ( .B(n140), .A(n161), .Z(n156) );
  NANDN U413 ( .B(n141), .A(n162), .Z(n136) );
  AND U414 ( .A(n163), .B(n164), .Z(n153) );
  OR U415 ( .A(n165), .B(n166), .Z(n164) );
  XNOR U416 ( .A(n167), .B(n168), .Z(n163) );
  ANDN U417 ( .A(n169), .B(n170), .Z(n168) );
  XOR U418 ( .A(n167), .B(n171), .Z(n169) );
  ANDN U419 ( .A(n174), .B(n175), .Z(n173) );
  XOR U420 ( .A(\_MxM/Y0[12] ), .B(n176), .Z(n174) );
  XNOR U421 ( .A(n175), .B(\_MxM/Y0[12] ), .Z(\_MxM/Y1[11] ) );
  XNOR U422 ( .A(n177), .B(n178), .Z(n175) );
  XNOR U423 ( .A(n176), .B(n179), .Z(n177) );
  AND U424 ( .A(n123), .B(n180), .Z(n179) );
  XOR U425 ( .A(n149), .B(n181), .Z(n180) );
  XOR U426 ( .A(n181), .B(n150), .Z(n149) );
  OR U427 ( .A(n182), .B(n183), .Z(n150) );
  IV U428 ( .A(n178), .Z(n181) );
  XNOR U429 ( .A(n152), .B(n151), .Z(n178) );
  OR U430 ( .A(n184), .B(n185), .Z(n151) );
  XNOR U431 ( .A(n166), .B(n165), .Z(n152) );
  OR U432 ( .A(n186), .B(n187), .Z(n165) );
  XOR U433 ( .A(n171), .B(n170), .Z(n166) );
  XOR U434 ( .A(n167), .B(n188), .Z(n170) );
  AND U435 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U436 ( .B(n140), .A(n191), .Z(n190) );
  OR U437 ( .A(n192), .B(n193), .Z(n189) );
  XOR U438 ( .A(n159), .B(n160), .Z(n171) );
  NANDN U439 ( .B(n141), .A(n196), .Z(n160) );
  XNOR U440 ( .A(n158), .B(n197), .Z(n159) );
  AND U441 ( .A(n162), .B(n161), .Z(n197) );
  ANDN U442 ( .A(n198), .B(n199), .Z(n158) );
  NANDN U443 ( .B(n200), .A(n201), .Z(n198) );
  IV U444 ( .A(n172), .Z(n176) );
  XNOR U445 ( .A(n203), .B(\_MxM/Y0[11] ), .Z(\_MxM/Y1[10] ) );
  XNOR U446 ( .A(n205), .B(n206), .Z(n203) );
  XNOR U447 ( .A(n204), .B(n207), .Z(n205) );
  AND U448 ( .A(n123), .B(n208), .Z(n207) );
  XOR U449 ( .A(n182), .B(n209), .Z(n208) );
  XOR U450 ( .A(n209), .B(n183), .Z(n182) );
  OR U451 ( .A(n210), .B(n211), .Z(n183) );
  IV U452 ( .A(n206), .Z(n209) );
  OR U453 ( .A(n212), .B(n213), .Z(n184) );
  XOR U454 ( .A(n195), .B(n194), .Z(n186) );
  XNOR U455 ( .A(n217), .B(n218), .Z(n194) );
  ANDN U456 ( .A(n221), .B(n222), .Z(n220) );
  XOR U457 ( .A(n219), .B(n223), .Z(n221) );
  XNOR U458 ( .A(n224), .B(n192), .Z(n217) );
  NAND U459 ( .A(n191), .B(n162), .Z(n192) );
  NANDN U460 ( .B(n140), .A(n226), .Z(n225) );
  XOR U461 ( .A(n200), .B(n201), .Z(n195) );
  NANDN U462 ( .B(n141), .A(n230), .Z(n201) );
  AND U463 ( .A(n196), .B(n161), .Z(n231) );
  NAND U464 ( .A(n232), .B(n233), .Z(n199) );
  NANDN U465 ( .B(n234), .A(n235), .Z(n232) );
  IV U466 ( .A(n202), .Z(n204) );
  XNOR U467 ( .A(n237), .B(n238), .Z(n108) );
  AND U468 ( .A(n123), .B(n240), .Z(n239) );
  XOR U469 ( .A(n210), .B(n241), .Z(n240) );
  XOR U470 ( .A(n241), .B(n211), .Z(n210) );
  OR U471 ( .A(n242), .B(n243), .Z(n211) );
  IV U472 ( .A(n238), .Z(n241) );
  XNOR U473 ( .A(n213), .B(n212), .Z(n238) );
  OR U474 ( .A(n244), .B(n245), .Z(n212) );
  XNOR U475 ( .A(n216), .B(n215), .Z(n213) );
  XOR U476 ( .A(n214), .B(n246), .Z(n215) );
  AND U477 ( .A(n247), .B(n248), .Z(n246) );
  OR U478 ( .A(n249), .B(n250), .Z(n248) );
  AND U479 ( .A(n251), .B(n252), .Z(n247) );
  NANDN U480 ( .B(n140), .A(n253), .Z(n252) );
  NAND U481 ( .A(n254), .B(n255), .Z(n251) );
  XNOR U482 ( .A(n227), .B(n260), .Z(n228) );
  AND U483 ( .A(n162), .B(n226), .Z(n260) );
  XOR U484 ( .A(n261), .B(n262), .Z(n227) );
  ANDN U485 ( .A(n263), .B(n264), .Z(n262) );
  XNOR U486 ( .A(n265), .B(n261), .Z(n263) );
  XOR U487 ( .A(n266), .B(n229), .Z(n259) );
  NAND U488 ( .A(n191), .B(n196), .Z(n229) );
  IV U489 ( .A(n219), .Z(n266) );
  XNOR U490 ( .A(n234), .B(n235), .Z(n223) );
  NANDN U491 ( .B(n141), .A(n270), .Z(n235) );
  XNOR U492 ( .A(n233), .B(n271), .Z(n234) );
  AND U493 ( .A(n230), .B(n161), .Z(n271) );
  ANDN U494 ( .A(n272), .B(n273), .Z(n233) );
  NANDN U495 ( .B(n274), .A(n275), .Z(n272) );
  XNOR U496 ( .A(n277), .B(n278), .Z(n109) );
  AND U497 ( .A(n123), .B(n280), .Z(n279) );
  XOR U498 ( .A(n242), .B(n281), .Z(n280) );
  XOR U499 ( .A(n281), .B(n243), .Z(n242) );
  OR U500 ( .A(n282), .B(n283), .Z(n243) );
  IV U501 ( .A(n278), .Z(n281) );
  XNOR U502 ( .A(n245), .B(n244), .Z(n278) );
  OR U503 ( .A(n284), .B(n285), .Z(n244) );
  XNOR U504 ( .A(n258), .B(n257), .Z(n245) );
  XOR U505 ( .A(n286), .B(n254), .Z(n257) );
  XNOR U506 ( .A(n287), .B(n249), .Z(n254) );
  NAND U507 ( .A(n253), .B(n162), .Z(n249) );
  NANDN U508 ( .B(n140), .A(n289), .Z(n288) );
  XNOR U509 ( .A(n255), .B(n256), .Z(n286) );
  XNOR U510 ( .A(n261), .B(n300), .Z(n264) );
  AND U511 ( .A(n196), .B(n226), .Z(n300) );
  XOR U512 ( .A(n301), .B(n302), .Z(n261) );
  ANDN U513 ( .A(n303), .B(n304), .Z(n302) );
  XNOR U514 ( .A(n305), .B(n301), .Z(n303) );
  XOR U515 ( .A(n306), .B(n265), .Z(n299) );
  NAND U516 ( .A(n191), .B(n230), .Z(n265) );
  IV U517 ( .A(n267), .Z(n306) );
  XNOR U518 ( .A(n274), .B(n275), .Z(n269) );
  NANDN U519 ( .B(n141), .A(n310), .Z(n275) );
  AND U520 ( .A(n270), .B(n161), .Z(n311) );
  NAND U521 ( .A(n312), .B(n313), .Z(n273) );
  NANDN U522 ( .B(n314), .A(n315), .Z(n312) );
  XNOR U523 ( .A(n317), .B(n318), .Z(n110) );
  XNOR U524 ( .A(n319), .B(n320), .Z(n317) );
  AND U525 ( .A(n123), .B(n321), .Z(n320) );
  XOR U526 ( .A(n282), .B(n322), .Z(n321) );
  XOR U527 ( .A(n322), .B(n283), .Z(n282) );
  OR U528 ( .A(n323), .B(n324), .Z(n283) );
  IV U529 ( .A(n318), .Z(n322) );
  XNOR U530 ( .A(n285), .B(n284), .Z(n318) );
  NANDN U531 ( .B(n325), .A(n326), .Z(n284) );
  XNOR U532 ( .A(n295), .B(n294), .Z(n285) );
  XOR U533 ( .A(n327), .B(n298), .Z(n294) );
  XNOR U534 ( .A(n291), .B(n292), .Z(n298) );
  NAND U535 ( .A(n253), .B(n196), .Z(n292) );
  XNOR U536 ( .A(n290), .B(n328), .Z(n291) );
  AND U537 ( .A(n162), .B(n289), .Z(n328) );
  XNOR U538 ( .A(n297), .B(n293), .Z(n327) );
  AND U539 ( .A(n336), .B(n337), .Z(n335) );
  NANDN U540 ( .B(n140), .A(n338), .Z(n337) );
  OR U541 ( .A(n339), .B(n340), .Z(n336) );
  XNOR U542 ( .A(n301), .B(n345), .Z(n304) );
  AND U543 ( .A(n230), .B(n226), .Z(n345) );
  XOR U544 ( .A(n349), .B(n305), .Z(n344) );
  NAND U545 ( .A(n191), .B(n270), .Z(n305) );
  IV U546 ( .A(n307), .Z(n349) );
  XNOR U547 ( .A(n314), .B(n315), .Z(n309) );
  NANDN U548 ( .B(n141), .A(n353), .Z(n315) );
  XNOR U549 ( .A(n313), .B(n354), .Z(n314) );
  AND U550 ( .A(n310), .B(n161), .Z(n354) );
  ANDN U551 ( .A(n355), .B(n356), .Z(n313) );
  NANDN U552 ( .B(n357), .A(n358), .Z(n355) );
  IV U553 ( .A(n316), .Z(n319) );
  XNOR U554 ( .A(n361), .B(n362), .Z(n360) );
  AND U555 ( .A(n123), .B(n363), .Z(n362) );
  XOR U556 ( .A(n323), .B(n366), .Z(n363) );
  XOR U557 ( .A(n366), .B(n324), .Z(n323) );
  OR U558 ( .A(n364), .B(n365), .Z(n324) );
  XNOR U559 ( .A(n325), .B(n326), .Z(n366) );
  XNOR U560 ( .A(n334), .B(n333), .Z(n325) );
  XOR U561 ( .A(n371), .B(n343), .Z(n333) );
  XNOR U562 ( .A(n330), .B(n331), .Z(n343) );
  NAND U563 ( .A(n253), .B(n230), .Z(n331) );
  XNOR U564 ( .A(n329), .B(n372), .Z(n330) );
  AND U565 ( .A(n196), .B(n289), .Z(n372) );
  XNOR U566 ( .A(n342), .B(n332), .Z(n371) );
  XNOR U567 ( .A(n379), .B(n341), .Z(n342) );
  XNOR U568 ( .A(n383), .B(n339), .Z(n379) );
  NAND U569 ( .A(n338), .B(n162), .Z(n339) );
  NANDN U570 ( .B(n140), .A(n385), .Z(n384) );
  XNOR U571 ( .A(n346), .B(n390), .Z(n347) );
  AND U572 ( .A(n270), .B(n226), .Z(n390) );
  XOR U573 ( .A(n391), .B(n392), .Z(n346) );
  ANDN U574 ( .A(n393), .B(n394), .Z(n392) );
  XNOR U575 ( .A(n395), .B(n391), .Z(n393) );
  XOR U576 ( .A(n396), .B(n348), .Z(n389) );
  NAND U577 ( .A(n191), .B(n310), .Z(n348) );
  IV U578 ( .A(n350), .Z(n396) );
  XNOR U579 ( .A(n357), .B(n358), .Z(n352) );
  NANDN U580 ( .B(n141), .A(n400), .Z(n358) );
  AND U581 ( .A(n353), .B(n161), .Z(n401) );
  NAND U582 ( .A(n402), .B(n403), .Z(n356) );
  NANDN U583 ( .B(n404), .A(n405), .Z(n402) );
  IV U584 ( .A(n359), .Z(n361) );
  XNOR U585 ( .A(n407), .B(n408), .Z(n112) );
  AND U586 ( .A(n123), .B(n410), .Z(n409) );
  XOR U587 ( .A(n364), .B(n411), .Z(n410) );
  XOR U588 ( .A(n411), .B(n365), .Z(n364) );
  OR U589 ( .A(n412), .B(n413), .Z(n365) );
  IV U590 ( .A(n408), .Z(n411) );
  XOR U591 ( .A(n370), .B(n369), .Z(n408) );
  XNOR U592 ( .A(n368), .B(n414), .Z(n369) );
  AND U593 ( .A(n367), .B(n415), .Z(n414) );
  AND U594 ( .A(n416), .B(n417), .Z(n415) );
  NANDN U595 ( .B(n140), .A(n418), .Z(n417) );
  OR U596 ( .A(n419), .B(n420), .Z(n416) );
  AND U597 ( .A(n421), .B(n422), .Z(n367) );
  NANDN U598 ( .B(n423), .A(n424), .Z(n422) );
  NANDN U599 ( .B(n425), .A(n426), .Z(n421) );
  XNOR U600 ( .A(n430), .B(n382), .Z(n377) );
  XNOR U601 ( .A(n374), .B(n375), .Z(n382) );
  NAND U602 ( .A(n253), .B(n270), .Z(n375) );
  XNOR U603 ( .A(n373), .B(n431), .Z(n374) );
  AND U604 ( .A(n230), .B(n289), .Z(n431) );
  XNOR U605 ( .A(n381), .B(n376), .Z(n430) );
  XNOR U606 ( .A(n386), .B(n439), .Z(n387) );
  AND U607 ( .A(n162), .B(n385), .Z(n439) );
  XOR U608 ( .A(n443), .B(n388), .Z(n438) );
  NAND U609 ( .A(n338), .B(n196), .Z(n388) );
  IV U610 ( .A(n380), .Z(n443) );
  XNOR U611 ( .A(n391), .B(n448), .Z(n394) );
  AND U612 ( .A(n310), .B(n226), .Z(n448) );
  XOR U613 ( .A(n449), .B(n450), .Z(n391) );
  ANDN U614 ( .A(n451), .B(n452), .Z(n450) );
  XNOR U615 ( .A(n453), .B(n449), .Z(n451) );
  XOR U616 ( .A(n454), .B(n395), .Z(n447) );
  NAND U617 ( .A(n191), .B(n353), .Z(n395) );
  IV U618 ( .A(n397), .Z(n454) );
  XNOR U619 ( .A(n404), .B(n405), .Z(n399) );
  NANDN U620 ( .B(n141), .A(n458), .Z(n405) );
  XNOR U621 ( .A(n403), .B(n459), .Z(n404) );
  AND U622 ( .A(n400), .B(n161), .Z(n459) );
  ANDN U623 ( .A(n460), .B(n461), .Z(n403) );
  NANDN U624 ( .B(n462), .A(n463), .Z(n460) );
  XNOR U625 ( .A(n465), .B(n466), .Z(n113) );
  AND U626 ( .A(n123), .B(n468), .Z(n467) );
  XOR U627 ( .A(n412), .B(n469), .Z(n468) );
  XOR U628 ( .A(n469), .B(n413), .Z(n412) );
  OR U629 ( .A(n470), .B(n471), .Z(n413) );
  IV U630 ( .A(n466), .Z(n469) );
  XOR U631 ( .A(n429), .B(n428), .Z(n466) );
  XOR U632 ( .A(n423), .B(n424), .Z(n420) );
  XOR U633 ( .A(n476), .B(n425), .Z(n423) );
  NAND U634 ( .A(n162), .B(n418), .Z(n425) );
  NANDN U635 ( .B(n426), .A(n477), .Z(n476) );
  NANDN U636 ( .B(n140), .A(n478), .Z(n477) );
  XOR U637 ( .A(n482), .B(n419), .Z(n472) );
  OR U638 ( .A(n483), .B(n484), .Z(n419) );
  IV U639 ( .A(n427), .Z(n482) );
  XNOR U640 ( .A(n488), .B(n446), .Z(n436) );
  XNOR U641 ( .A(n433), .B(n434), .Z(n446) );
  NAND U642 ( .A(n253), .B(n310), .Z(n434) );
  XNOR U643 ( .A(n432), .B(n489), .Z(n433) );
  AND U644 ( .A(n270), .B(n289), .Z(n489) );
  XNOR U645 ( .A(n445), .B(n435), .Z(n488) );
  XNOR U646 ( .A(n440), .B(n497), .Z(n441) );
  AND U647 ( .A(n196), .B(n385), .Z(n497) );
  XOR U648 ( .A(n501), .B(n442), .Z(n496) );
  NAND U649 ( .A(n338), .B(n230), .Z(n442) );
  IV U650 ( .A(n444), .Z(n501) );
  XNOR U651 ( .A(n449), .B(n506), .Z(n452) );
  AND U652 ( .A(n353), .B(n226), .Z(n506) );
  XOR U653 ( .A(n507), .B(n508), .Z(n449) );
  ANDN U654 ( .A(n509), .B(n510), .Z(n508) );
  XNOR U655 ( .A(n511), .B(n507), .Z(n509) );
  XOR U656 ( .A(n512), .B(n453), .Z(n505) );
  NAND U657 ( .A(n191), .B(n400), .Z(n453) );
  IV U658 ( .A(n455), .Z(n512) );
  XNOR U659 ( .A(n462), .B(n463), .Z(n457) );
  NANDN U660 ( .B(n141), .A(n516), .Z(n463) );
  AND U661 ( .A(n458), .B(n161), .Z(n517) );
  NAND U662 ( .A(n518), .B(n519), .Z(n461) );
  NANDN U663 ( .B(n520), .A(n521), .Z(n518) );
  XNOR U664 ( .A(n523), .B(n524), .Z(n114) );
  AND U665 ( .A(n123), .B(n526), .Z(n525) );
  XOR U666 ( .A(n470), .B(n527), .Z(n526) );
  XOR U667 ( .A(n527), .B(n471), .Z(n470) );
  OR U668 ( .A(n528), .B(n529), .Z(n471) );
  IV U669 ( .A(n524), .Z(n527) );
  XOR U670 ( .A(n487), .B(n486), .Z(n524) );
  XOR U671 ( .A(n530), .B(n483), .Z(n486) );
  XOR U672 ( .A(n475), .B(n474), .Z(n483) );
  XOR U673 ( .A(n473), .B(n531), .Z(n474) );
  AND U674 ( .A(n532), .B(n533), .Z(n531) );
  NANDN U675 ( .B(n140), .A(n534), .Z(n533) );
  OR U676 ( .A(n535), .B(n536), .Z(n532) );
  NAND U677 ( .A(n196), .B(n418), .Z(n481) );
  XNOR U678 ( .A(n479), .B(n540), .Z(n480) );
  AND U679 ( .A(n478), .B(n162), .Z(n540) );
  NANDN U680 ( .B(n544), .A(n545), .Z(n484) );
  XNOR U681 ( .A(n549), .B(n504), .Z(n494) );
  XNOR U682 ( .A(n491), .B(n492), .Z(n504) );
  NAND U683 ( .A(n253), .B(n353), .Z(n492) );
  XNOR U684 ( .A(n490), .B(n550), .Z(n491) );
  AND U685 ( .A(n310), .B(n289), .Z(n550) );
  XNOR U686 ( .A(n503), .B(n493), .Z(n549) );
  XNOR U687 ( .A(n498), .B(n558), .Z(n499) );
  AND U688 ( .A(n230), .B(n385), .Z(n558) );
  XOR U689 ( .A(n562), .B(n500), .Z(n557) );
  NAND U690 ( .A(n338), .B(n270), .Z(n500) );
  IV U691 ( .A(n502), .Z(n562) );
  XNOR U692 ( .A(n507), .B(n567), .Z(n510) );
  AND U693 ( .A(n400), .B(n226), .Z(n567) );
  XOR U694 ( .A(n568), .B(n569), .Z(n507) );
  ANDN U695 ( .A(n570), .B(n571), .Z(n569) );
  XNOR U696 ( .A(n572), .B(n568), .Z(n570) );
  XOR U697 ( .A(n573), .B(n511), .Z(n566) );
  NAND U698 ( .A(n191), .B(n458), .Z(n511) );
  IV U699 ( .A(n513), .Z(n573) );
  XNOR U700 ( .A(n520), .B(n521), .Z(n515) );
  NANDN U701 ( .B(n141), .A(n577), .Z(n521) );
  XNOR U702 ( .A(n519), .B(n578), .Z(n520) );
  AND U703 ( .A(n516), .B(n161), .Z(n578) );
  ANDN U704 ( .A(n579), .B(n580), .Z(n519) );
  NANDN U705 ( .B(n581), .A(n582), .Z(n579) );
  XNOR U706 ( .A(n584), .B(n585), .Z(n115) );
  AND U707 ( .A(n123), .B(n587), .Z(n586) );
  XOR U708 ( .A(n528), .B(n588), .Z(n587) );
  XOR U709 ( .A(n588), .B(n529), .Z(n528) );
  OR U710 ( .A(n589), .B(n590), .Z(n529) );
  IV U711 ( .A(n585), .Z(n588) );
  XOR U712 ( .A(n548), .B(n547), .Z(n585) );
  XOR U713 ( .A(n591), .B(n544), .Z(n547) );
  XOR U714 ( .A(n539), .B(n538), .Z(n544) );
  XNOR U715 ( .A(n596), .B(n535), .Z(n592) );
  NAND U716 ( .A(n162), .B(n534), .Z(n535) );
  NANDN U717 ( .B(n140), .A(n598), .Z(n597) );
  NAND U718 ( .A(n230), .B(n418), .Z(n543) );
  XNOR U719 ( .A(n541), .B(n602), .Z(n542) );
  AND U720 ( .A(n478), .B(n196), .Z(n602) );
  XNOR U721 ( .A(n545), .B(n546), .Z(n591) );
  XNOR U722 ( .A(n612), .B(n565), .Z(n555) );
  XNOR U723 ( .A(n552), .B(n553), .Z(n565) );
  NAND U724 ( .A(n253), .B(n400), .Z(n553) );
  XNOR U725 ( .A(n551), .B(n613), .Z(n552) );
  AND U726 ( .A(n353), .B(n289), .Z(n613) );
  XNOR U727 ( .A(n564), .B(n554), .Z(n612) );
  XNOR U728 ( .A(n559), .B(n621), .Z(n560) );
  AND U729 ( .A(n270), .B(n385), .Z(n621) );
  XOR U730 ( .A(n622), .B(n623), .Z(n559) );
  ANDN U731 ( .A(n624), .B(n625), .Z(n623) );
  XNOR U732 ( .A(n626), .B(n622), .Z(n624) );
  XOR U733 ( .A(n627), .B(n561), .Z(n620) );
  NAND U734 ( .A(n338), .B(n310), .Z(n561) );
  IV U735 ( .A(n563), .Z(n627) );
  XNOR U736 ( .A(n568), .B(n632), .Z(n571) );
  AND U737 ( .A(n458), .B(n226), .Z(n632) );
  XOR U738 ( .A(n633), .B(n634), .Z(n568) );
  ANDN U739 ( .A(n635), .B(n636), .Z(n634) );
  XNOR U740 ( .A(n637), .B(n633), .Z(n635) );
  XOR U741 ( .A(n638), .B(n572), .Z(n631) );
  NAND U742 ( .A(n191), .B(n516), .Z(n572) );
  IV U743 ( .A(n574), .Z(n638) );
  XNOR U744 ( .A(n581), .B(n582), .Z(n576) );
  OR U745 ( .A(n642), .B(n141), .Z(n582) );
  AND U746 ( .A(n577), .B(n161), .Z(n643) );
  NAND U747 ( .A(n644), .B(n645), .Z(n580) );
  NANDN U748 ( .B(n646), .A(n647), .Z(n644) );
  XNOR U749 ( .A(n649), .B(n650), .Z(n116) );
  XOR U750 ( .A(n648), .B(n651), .Z(n649) );
  AND U751 ( .A(n123), .B(n652), .Z(n651) );
  XOR U752 ( .A(n589), .B(n653), .Z(n652) );
  XOR U753 ( .A(n653), .B(n590), .Z(n589) );
  NANDN U754 ( .B(n654), .A(n655), .Z(n590) );
  IV U755 ( .A(n650), .Z(n653) );
  XOR U756 ( .A(n608), .B(n607), .Z(n650) );
  XNOR U757 ( .A(n656), .B(n611), .Z(n607) );
  XNOR U758 ( .A(n599), .B(n658), .Z(n600) );
  AND U759 ( .A(n598), .B(n162), .Z(n658) );
  XOR U760 ( .A(n662), .B(n601), .Z(n657) );
  NAND U761 ( .A(n196), .B(n534), .Z(n601) );
  IV U762 ( .A(n593), .Z(n662) );
  XNOR U763 ( .A(n604), .B(n605), .Z(n595) );
  NAND U764 ( .A(n270), .B(n418), .Z(n605) );
  XNOR U765 ( .A(n603), .B(n666), .Z(n604) );
  AND U766 ( .A(n478), .B(n230), .Z(n666) );
  XNOR U767 ( .A(n610), .B(n606), .Z(n656) );
  AND U768 ( .A(n674), .B(n675), .Z(n673) );
  OR U769 ( .A(n676), .B(n677), .Z(n675) );
  AND U770 ( .A(n678), .B(n679), .Z(n674) );
  NANDN U771 ( .B(n140), .A(n680), .Z(n679) );
  NANDN U772 ( .B(n681), .A(n682), .Z(n678) );
  XNOR U773 ( .A(n686), .B(n630), .Z(n618) );
  XNOR U774 ( .A(n615), .B(n616), .Z(n630) );
  NAND U775 ( .A(n253), .B(n458), .Z(n616) );
  XNOR U776 ( .A(n614), .B(n687), .Z(n615) );
  AND U777 ( .A(n400), .B(n289), .Z(n687) );
  XNOR U778 ( .A(n629), .B(n617), .Z(n686) );
  XNOR U779 ( .A(n622), .B(n695), .Z(n625) );
  AND U780 ( .A(n310), .B(n385), .Z(n695) );
  XOR U781 ( .A(n699), .B(n626), .Z(n694) );
  NAND U782 ( .A(n338), .B(n353), .Z(n626) );
  IV U783 ( .A(n628), .Z(n699) );
  XNOR U784 ( .A(n633), .B(n704), .Z(n636) );
  AND U785 ( .A(n516), .B(n226), .Z(n704) );
  XOR U786 ( .A(n705), .B(n706), .Z(n633) );
  ANDN U787 ( .A(n707), .B(n708), .Z(n706) );
  XNOR U788 ( .A(n709), .B(n705), .Z(n707) );
  XOR U789 ( .A(n710), .B(n637), .Z(n703) );
  NAND U790 ( .A(n191), .B(n577), .Z(n637) );
  IV U791 ( .A(n639), .Z(n710) );
  XNOR U792 ( .A(n646), .B(n647), .Z(n641) );
  OR U793 ( .A(n714), .B(n141), .Z(n647) );
  XNOR U794 ( .A(n645), .B(n715), .Z(n646) );
  ANDN U795 ( .A(n161), .B(n642), .Z(n715) );
  ANDN U796 ( .A(n716), .B(n717), .Z(n645) );
  NANDN U797 ( .B(n718), .A(n719), .Z(n716) );
  XNOR U798 ( .A(n721), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U799 ( .A(n722), .B(n723), .Z(n721) );
  XNOR U800 ( .A(n724), .B(n720), .Z(n722) );
  NAND U801 ( .A(\_MxM/Y0[0] ), .B(n654), .Z(n720) );
  NAND U802 ( .A(n725), .B(n123), .Z(n724) );
  XOR U803 ( .A(e_input[15]), .B(g_input[15]), .Z(n123) );
  XNOR U804 ( .A(n655), .B(n723), .Z(n725) );
  XNOR U805 ( .A(n654), .B(n723), .Z(n655) );
  XNOR U806 ( .A(n672), .B(n671), .Z(n723) );
  XNOR U807 ( .A(n726), .B(n685), .Z(n671) );
  XNOR U808 ( .A(n659), .B(n728), .Z(n660) );
  AND U809 ( .A(n598), .B(n196), .Z(n728) );
  XOR U810 ( .A(n732), .B(n661), .Z(n727) );
  NAND U811 ( .A(n230), .B(n534), .Z(n661) );
  IV U812 ( .A(n663), .Z(n732) );
  XNOR U813 ( .A(n668), .B(n669), .Z(n665) );
  NAND U814 ( .A(n310), .B(n418), .Z(n669) );
  XNOR U815 ( .A(n667), .B(n736), .Z(n668) );
  AND U816 ( .A(n478), .B(n270), .Z(n736) );
  XNOR U817 ( .A(n684), .B(n670), .Z(n726) );
  XNOR U818 ( .A(n743), .B(n681), .Z(n684) );
  XOR U819 ( .A(n744), .B(n676), .Z(n681) );
  NAND U820 ( .A(n162), .B(n680), .Z(n676) );
  NANDN U821 ( .B(n140), .A(n746), .Z(n745) );
  XNOR U822 ( .A(n682), .B(n683), .Z(n743) );
  XNOR U823 ( .A(n755), .B(n702), .Z(n692) );
  XNOR U824 ( .A(n689), .B(n690), .Z(n702) );
  NAND U825 ( .A(n253), .B(n516), .Z(n690) );
  XNOR U826 ( .A(n688), .B(n756), .Z(n689) );
  AND U827 ( .A(n458), .B(n289), .Z(n756) );
  XNOR U828 ( .A(n701), .B(n691), .Z(n755) );
  XNOR U829 ( .A(n696), .B(n764), .Z(n697) );
  AND U830 ( .A(n353), .B(n385), .Z(n764) );
  XOR U831 ( .A(n765), .B(n766), .Z(n696) );
  ANDN U832 ( .A(n767), .B(n768), .Z(n766) );
  XNOR U833 ( .A(n769), .B(n765), .Z(n767) );
  XOR U834 ( .A(n770), .B(n698), .Z(n763) );
  NAND U835 ( .A(n338), .B(n400), .Z(n698) );
  IV U836 ( .A(n700), .Z(n770) );
  XNOR U837 ( .A(n705), .B(n775), .Z(n708) );
  AND U838 ( .A(n577), .B(n226), .Z(n775) );
  XOR U839 ( .A(n776), .B(n777), .Z(n705) );
  ANDN U840 ( .A(n778), .B(n779), .Z(n777) );
  XNOR U841 ( .A(n780), .B(n776), .Z(n778) );
  XOR U842 ( .A(n781), .B(n709), .Z(n774) );
  NANDN U843 ( .B(n642), .A(n191), .Z(n709) );
  IV U844 ( .A(n711), .Z(n781) );
  XNOR U845 ( .A(n718), .B(n719), .Z(n713) );
  NANDN U846 ( .B(n141), .A(n785), .Z(n719) );
  ANDN U847 ( .A(n161), .B(n714), .Z(n786) );
  NAND U848 ( .A(n787), .B(n788), .Z(n717) );
  NANDN U849 ( .B(n789), .A(n790), .Z(n787) );
  XNOR U850 ( .A(n742), .B(n741), .Z(n654) );
  XNOR U851 ( .A(n791), .B(n752), .Z(n741) );
  XNOR U852 ( .A(n729), .B(n793), .Z(n730) );
  AND U853 ( .A(n598), .B(n230), .Z(n793) );
  XOR U854 ( .A(n794), .B(n795), .Z(n729) );
  ANDN U855 ( .A(n796), .B(n797), .Z(n795) );
  XNOR U856 ( .A(n798), .B(n794), .Z(n796) );
  XOR U857 ( .A(n799), .B(n731), .Z(n792) );
  NAND U858 ( .A(n270), .B(n534), .Z(n731) );
  IV U859 ( .A(n733), .Z(n799) );
  XNOR U860 ( .A(n738), .B(n739), .Z(n735) );
  NAND U861 ( .A(n353), .B(n418), .Z(n739) );
  XNOR U862 ( .A(n737), .B(n803), .Z(n738) );
  AND U863 ( .A(n478), .B(n310), .Z(n803) );
  XNOR U864 ( .A(n751), .B(n740), .Z(n791) );
  XOR U865 ( .A(n807), .B(n808), .Z(n740) );
  XNOR U866 ( .A(n809), .B(n754), .Z(n751) );
  NAND U867 ( .A(n196), .B(n680), .Z(n749) );
  XNOR U868 ( .A(n747), .B(n810), .Z(n748) );
  AND U869 ( .A(n746), .B(n162), .Z(n810) );
  XNOR U870 ( .A(n753), .B(n750), .Z(n809) );
  XOR U871 ( .A(n814), .B(n815), .Z(n750) );
  AND U872 ( .A(n816), .B(n817), .Z(n815) );
  XOR U873 ( .A(n818), .B(n819), .Z(n817) );
  XOR U874 ( .A(n814), .B(n820), .Z(n819) );
  XOR U875 ( .A(n801), .B(n821), .Z(n816) );
  XOR U876 ( .A(n814), .B(n802), .Z(n821) );
  NAND U877 ( .A(n418), .B(n400), .Z(n806) );
  XNOR U878 ( .A(n804), .B(n822), .Z(n805) );
  AND U879 ( .A(n478), .B(n353), .Z(n822) );
  XNOR U880 ( .A(n794), .B(n827), .Z(n797) );
  AND U881 ( .A(n598), .B(n270), .Z(n827) );
  XOR U882 ( .A(n831), .B(n798), .Z(n826) );
  NAND U883 ( .A(n310), .B(n534), .Z(n798) );
  IV U884 ( .A(n800), .Z(n831) );
  XOR U885 ( .A(n835), .B(n836), .Z(n814) );
  AND U886 ( .A(n837), .B(n838), .Z(n836) );
  XOR U887 ( .A(n839), .B(n840), .Z(n838) );
  XOR U888 ( .A(n835), .B(n841), .Z(n840) );
  XOR U889 ( .A(n833), .B(n842), .Z(n837) );
  XOR U890 ( .A(n835), .B(n834), .Z(n842) );
  NAND U891 ( .A(n418), .B(n458), .Z(n825) );
  XNOR U892 ( .A(n823), .B(n843), .Z(n824) );
  AND U893 ( .A(n400), .B(n478), .Z(n843) );
  XNOR U894 ( .A(n828), .B(n848), .Z(n829) );
  AND U895 ( .A(n598), .B(n310), .Z(n848) );
  XOR U896 ( .A(n849), .B(n850), .Z(n828) );
  ANDN U897 ( .A(n851), .B(n852), .Z(n850) );
  XNOR U898 ( .A(n853), .B(n849), .Z(n851) );
  XOR U899 ( .A(n854), .B(n830), .Z(n847) );
  NAND U900 ( .A(n353), .B(n534), .Z(n830) );
  IV U901 ( .A(n832), .Z(n854) );
  XOR U902 ( .A(n858), .B(n859), .Z(n835) );
  AND U903 ( .A(n860), .B(n861), .Z(n859) );
  XOR U904 ( .A(n862), .B(n863), .Z(n861) );
  XOR U905 ( .A(n858), .B(n864), .Z(n863) );
  XOR U906 ( .A(n856), .B(n865), .Z(n860) );
  XOR U907 ( .A(n858), .B(n857), .Z(n865) );
  NAND U908 ( .A(n418), .B(n516), .Z(n846) );
  XNOR U909 ( .A(n844), .B(n866), .Z(n845) );
  AND U910 ( .A(n458), .B(n478), .Z(n866) );
  XOR U911 ( .A(n867), .B(n868), .Z(n844) );
  ANDN U912 ( .A(n869), .B(n870), .Z(n868) );
  XNOR U913 ( .A(n871), .B(n867), .Z(n869) );
  XNOR U914 ( .A(n872), .B(n873), .Z(n856) );
  IV U915 ( .A(n852), .Z(n873) );
  XNOR U916 ( .A(n849), .B(n874), .Z(n852) );
  AND U917 ( .A(n598), .B(n353), .Z(n874) );
  XOR U918 ( .A(n875), .B(n876), .Z(n849) );
  ANDN U919 ( .A(n877), .B(n878), .Z(n876) );
  XNOR U920 ( .A(n879), .B(n875), .Z(n877) );
  XOR U921 ( .A(n880), .B(n853), .Z(n872) );
  NAND U922 ( .A(n534), .B(n400), .Z(n853) );
  IV U923 ( .A(n855), .Z(n880) );
  XOR U924 ( .A(n884), .B(n885), .Z(n858) );
  AND U925 ( .A(n886), .B(n887), .Z(n885) );
  XOR U926 ( .A(n888), .B(n889), .Z(n887) );
  XOR U927 ( .A(n884), .B(n890), .Z(n889) );
  XOR U928 ( .A(n882), .B(n891), .Z(n886) );
  XOR U929 ( .A(n884), .B(n883), .Z(n891) );
  XNOR U930 ( .A(n892), .B(n871), .Z(n883) );
  NAND U931 ( .A(n418), .B(n577), .Z(n871) );
  IV U932 ( .A(n870), .Z(n892) );
  XNOR U933 ( .A(n867), .B(n893), .Z(n870) );
  AND U934 ( .A(n516), .B(n478), .Z(n893) );
  XOR U935 ( .A(n894), .B(n895), .Z(n867) );
  ANDN U936 ( .A(n896), .B(n897), .Z(n895) );
  XNOR U937 ( .A(n898), .B(n894), .Z(n896) );
  XNOR U938 ( .A(n899), .B(n900), .Z(n882) );
  IV U939 ( .A(n878), .Z(n900) );
  XNOR U940 ( .A(n875), .B(n901), .Z(n878) );
  AND U941 ( .A(n400), .B(n598), .Z(n901) );
  XOR U942 ( .A(n902), .B(n903), .Z(n875) );
  ANDN U943 ( .A(n904), .B(n905), .Z(n903) );
  XNOR U944 ( .A(n906), .B(n902), .Z(n904) );
  XOR U945 ( .A(n907), .B(n879), .Z(n899) );
  NAND U946 ( .A(n534), .B(n458), .Z(n879) );
  IV U947 ( .A(n881), .Z(n907) );
  XOR U948 ( .A(n911), .B(n912), .Z(n884) );
  AND U949 ( .A(n913), .B(n914), .Z(n912) );
  XOR U950 ( .A(n915), .B(n916), .Z(n914) );
  XOR U951 ( .A(n911), .B(n917), .Z(n916) );
  XOR U952 ( .A(n909), .B(n918), .Z(n913) );
  XOR U953 ( .A(n911), .B(n910), .Z(n918) );
  XNOR U954 ( .A(n919), .B(n898), .Z(n910) );
  NANDN U955 ( .B(n642), .A(n418), .Z(n898) );
  IV U956 ( .A(n897), .Z(n919) );
  XNOR U957 ( .A(n894), .B(n920), .Z(n897) );
  AND U958 ( .A(n577), .B(n478), .Z(n920) );
  XOR U959 ( .A(n921), .B(n922), .Z(n894) );
  ANDN U960 ( .A(n923), .B(n924), .Z(n922) );
  XNOR U961 ( .A(n925), .B(n921), .Z(n923) );
  XNOR U962 ( .A(n926), .B(n927), .Z(n909) );
  IV U963 ( .A(n905), .Z(n927) );
  XNOR U964 ( .A(n902), .B(n928), .Z(n905) );
  AND U965 ( .A(n458), .B(n598), .Z(n928) );
  XOR U966 ( .A(n929), .B(n930), .Z(n902) );
  ANDN U967 ( .A(n931), .B(n932), .Z(n930) );
  XNOR U968 ( .A(n933), .B(n929), .Z(n931) );
  XOR U969 ( .A(n934), .B(n906), .Z(n926) );
  NAND U970 ( .A(n534), .B(n516), .Z(n906) );
  IV U971 ( .A(n908), .Z(n934) );
  XOR U972 ( .A(n938), .B(n939), .Z(n911) );
  AND U973 ( .A(n940), .B(n941), .Z(n939) );
  XOR U974 ( .A(n942), .B(n943), .Z(n941) );
  XOR U975 ( .A(n938), .B(n944), .Z(n943) );
  XOR U976 ( .A(n936), .B(n945), .Z(n940) );
  XOR U977 ( .A(n938), .B(n937), .Z(n945) );
  XNOR U978 ( .A(n946), .B(n925), .Z(n937) );
  NANDN U979 ( .B(n714), .A(n418), .Z(n925) );
  IV U980 ( .A(n924), .Z(n946) );
  XNOR U981 ( .A(n921), .B(n947), .Z(n924) );
  ANDN U982 ( .A(n478), .B(n642), .Z(n947) );
  XOR U983 ( .A(n948), .B(n949), .Z(n921) );
  ANDN U984 ( .A(n950), .B(n951), .Z(n949) );
  XNOR U985 ( .A(n952), .B(n948), .Z(n950) );
  XNOR U986 ( .A(n953), .B(n954), .Z(n936) );
  IV U987 ( .A(n932), .Z(n954) );
  XNOR U988 ( .A(n929), .B(n955), .Z(n932) );
  AND U989 ( .A(n516), .B(n598), .Z(n955) );
  XOR U990 ( .A(n956), .B(n957), .Z(n929) );
  ANDN U991 ( .A(n958), .B(n959), .Z(n957) );
  XNOR U992 ( .A(n960), .B(n956), .Z(n958) );
  XOR U993 ( .A(n961), .B(n933), .Z(n953) );
  NAND U994 ( .A(n534), .B(n577), .Z(n933) );
  IV U995 ( .A(n935), .Z(n961) );
  XOR U996 ( .A(n965), .B(n966), .Z(n938) );
  AND U997 ( .A(n967), .B(n968), .Z(n966) );
  XOR U998 ( .A(n969), .B(n970), .Z(n968) );
  XOR U999 ( .A(n965), .B(n971), .Z(n970) );
  XOR U1000 ( .A(n963), .B(n972), .Z(n967) );
  XOR U1001 ( .A(n965), .B(n964), .Z(n972) );
  XNOR U1002 ( .A(n973), .B(n952), .Z(n964) );
  NAND U1003 ( .A(n418), .B(n785), .Z(n952) );
  IV U1004 ( .A(n951), .Z(n973) );
  XNOR U1005 ( .A(n948), .B(n974), .Z(n951) );
  ANDN U1006 ( .A(n478), .B(n714), .Z(n974) );
  XOR U1007 ( .A(n975), .B(n976), .Z(n948) );
  ANDN U1008 ( .A(n977), .B(n978), .Z(n976) );
  XNOR U1009 ( .A(n979), .B(n975), .Z(n977) );
  XNOR U1010 ( .A(n980), .B(n981), .Z(n963) );
  IV U1011 ( .A(n959), .Z(n981) );
  XNOR U1012 ( .A(n956), .B(n982), .Z(n959) );
  AND U1013 ( .A(n577), .B(n598), .Z(n982) );
  XOR U1014 ( .A(n983), .B(n984), .Z(n956) );
  ANDN U1015 ( .A(n985), .B(n986), .Z(n984) );
  XNOR U1016 ( .A(n987), .B(n983), .Z(n985) );
  XOR U1017 ( .A(n988), .B(n960), .Z(n980) );
  NANDN U1018 ( .B(n642), .A(n534), .Z(n960) );
  IV U1019 ( .A(n962), .Z(n988) );
  XOR U1020 ( .A(n993), .B(n994), .Z(n808) );
  XNOR U1021 ( .A(n995), .B(n992), .Z(n993) );
  XNOR U1022 ( .A(n983), .B(n997), .Z(n986) );
  ANDN U1023 ( .A(n598), .B(n642), .Z(n997) );
  XOR U1024 ( .A(n1000), .B(n998), .Z(n999) );
  ANDN U1025 ( .A(n598), .B(n714), .Z(n1000) );
  AND U1026 ( .A(n785), .B(n534), .Z(n1001) );
  XOR U1027 ( .A(n1002), .B(n1003), .Z(n998) );
  ANDN U1028 ( .A(n1004), .B(n1005), .Z(n1003) );
  XNOR U1029 ( .A(n1006), .B(n1002), .Z(n1004) );
  XOR U1030 ( .A(n1007), .B(n987), .Z(n996) );
  NANDN U1031 ( .B(n714), .A(n534), .Z(n987) );
  IV U1032 ( .A(n989), .Z(n1007) );
  NAND U1033 ( .A(n534), .B(n1008), .Z(n1006) );
  XNOR U1034 ( .A(n1002), .B(n1009), .Z(n1005) );
  AND U1035 ( .A(n785), .B(n598), .Z(n1009) );
  AND U1036 ( .A(n1010), .B(g_input[0]), .Z(n1002) );
  NANDN U1037 ( .B(n534), .A(n1011), .Z(n1010) );
  NAND U1038 ( .A(n1008), .B(n598), .Z(n1011) );
  XNOR U1039 ( .A(n978), .B(n979), .Z(n991) );
  NAND U1040 ( .A(n418), .B(n1008), .Z(n979) );
  XNOR U1041 ( .A(n975), .B(n1014), .Z(n978) );
  AND U1042 ( .A(n785), .B(n478), .Z(n1014) );
  AND U1043 ( .A(n1015), .B(g_input[0]), .Z(n975) );
  NANDN U1044 ( .B(n418), .A(n1016), .Z(n1015) );
  NAND U1045 ( .A(n1008), .B(n478), .Z(n1016) );
  XOR U1046 ( .A(n1019), .B(n1020), .Z(n992) );
  XOR U1047 ( .A(n1021), .B(n1022), .Z(n753) );
  AND U1048 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U1049 ( .B(n140), .A(n1025), .Z(n1024) );
  NANDN U1050 ( .B(n1026), .A(n1027), .Z(n140) );
  AND U1051 ( .A(n1028), .B(g_input[15]), .Z(n1027) );
  OR U1052 ( .A(n1029), .B(n1030), .Z(n1023) );
  AND U1053 ( .A(n820), .B(n1033), .Z(n1032) );
  XNOR U1054 ( .A(n1031), .B(n818), .Z(n1033) );
  NAND U1055 ( .A(n230), .B(n680), .Z(n813) );
  XNOR U1056 ( .A(n811), .B(n1034), .Z(n812) );
  AND U1057 ( .A(n746), .B(n196), .Z(n1034) );
  XOR U1058 ( .A(n1042), .B(n1029), .Z(n1038) );
  NAND U1059 ( .A(n162), .B(n1025), .Z(n1029) );
  IV U1060 ( .A(n1031), .Z(n1042) );
  NAND U1061 ( .A(n270), .B(n680), .Z(n1037) );
  XNOR U1062 ( .A(n1035), .B(n1044), .Z(n1036) );
  AND U1063 ( .A(n746), .B(n230), .Z(n1044) );
  XNOR U1064 ( .A(n1048), .B(n1049), .Z(n841) );
  IV U1065 ( .A(n1040), .Z(n1049) );
  XNOR U1066 ( .A(n1039), .B(n1050), .Z(n1040) );
  AND U1067 ( .A(n162), .B(e_input[0]), .Z(n1050) );
  XNOR U1068 ( .A(n1028), .B(g_input[14]), .Z(n1026) );
  NOR U1069 ( .A(n1051), .B(n1052), .Z(n1028) );
  XOR U1070 ( .A(n1056), .B(n1041), .Z(n1048) );
  NAND U1071 ( .A(n196), .B(n1025), .Z(n1041) );
  IV U1072 ( .A(n1043), .Z(n1056) );
  NAND U1073 ( .A(n310), .B(n680), .Z(n1047) );
  XNOR U1074 ( .A(n1045), .B(n1058), .Z(n1046) );
  AND U1075 ( .A(n746), .B(n270), .Z(n1058) );
  XOR U1076 ( .A(n1059), .B(n1060), .Z(n1045) );
  ANDN U1077 ( .A(n1061), .B(n1062), .Z(n1060) );
  XNOR U1078 ( .A(n1063), .B(n1059), .Z(n1061) );
  XNOR U1079 ( .A(n1053), .B(n1065), .Z(n1054) );
  AND U1080 ( .A(n196), .B(e_input[0]), .Z(n1065) );
  XOR U1081 ( .A(n1051), .B(g_input[13]), .Z(n1052) );
  NANDN U1082 ( .B(n1066), .A(n1067), .Z(n1051) );
  XOR U1083 ( .A(n1071), .B(n1055), .Z(n1064) );
  NAND U1084 ( .A(n230), .B(n1025), .Z(n1055) );
  IV U1085 ( .A(n1057), .Z(n1071) );
  XNOR U1086 ( .A(n1073), .B(n1063), .Z(n888) );
  NAND U1087 ( .A(n353), .B(n680), .Z(n1063) );
  IV U1088 ( .A(n1062), .Z(n1073) );
  XNOR U1089 ( .A(n1059), .B(n1074), .Z(n1062) );
  AND U1090 ( .A(n746), .B(n310), .Z(n1074) );
  XOR U1091 ( .A(n1075), .B(n1076), .Z(n1059) );
  ANDN U1092 ( .A(n1077), .B(n1078), .Z(n1076) );
  XNOR U1093 ( .A(n1079), .B(n1075), .Z(n1077) );
  XNOR U1094 ( .A(n1080), .B(n1081), .Z(n890) );
  IV U1095 ( .A(n1069), .Z(n1081) );
  XNOR U1096 ( .A(n1068), .B(n1082), .Z(n1069) );
  AND U1097 ( .A(n230), .B(e_input[0]), .Z(n1082) );
  XNOR U1098 ( .A(n1067), .B(g_input[12]), .Z(n1066) );
  NOR U1099 ( .A(n1083), .B(n1084), .Z(n1067) );
  XOR U1100 ( .A(n1088), .B(n1070), .Z(n1080) );
  NAND U1101 ( .A(n270), .B(n1025), .Z(n1070) );
  IV U1102 ( .A(n1072), .Z(n1088) );
  XNOR U1103 ( .A(n1090), .B(n1079), .Z(n915) );
  NAND U1104 ( .A(n400), .B(n680), .Z(n1079) );
  IV U1105 ( .A(n1078), .Z(n1090) );
  XNOR U1106 ( .A(n1075), .B(n1091), .Z(n1078) );
  AND U1107 ( .A(n746), .B(n353), .Z(n1091) );
  XOR U1108 ( .A(n1092), .B(n1093), .Z(n1075) );
  ANDN U1109 ( .A(n1094), .B(n1095), .Z(n1093) );
  XNOR U1110 ( .A(n1096), .B(n1092), .Z(n1094) );
  XNOR U1111 ( .A(n1097), .B(n1098), .Z(n917) );
  IV U1112 ( .A(n1086), .Z(n1098) );
  XNOR U1113 ( .A(n1085), .B(n1099), .Z(n1086) );
  AND U1114 ( .A(n270), .B(e_input[0]), .Z(n1099) );
  XOR U1115 ( .A(n1083), .B(g_input[11]), .Z(n1084) );
  NANDN U1116 ( .B(n1100), .A(n1101), .Z(n1083) );
  XOR U1117 ( .A(n1102), .B(n1103), .Z(n1085) );
  ANDN U1118 ( .A(n1104), .B(n1105), .Z(n1103) );
  XNOR U1119 ( .A(n1106), .B(n1102), .Z(n1104) );
  XOR U1120 ( .A(n1107), .B(n1087), .Z(n1097) );
  NAND U1121 ( .A(n310), .B(n1025), .Z(n1087) );
  IV U1122 ( .A(n1089), .Z(n1107) );
  XNOR U1123 ( .A(n1109), .B(n1096), .Z(n942) );
  NAND U1124 ( .A(n458), .B(n680), .Z(n1096) );
  IV U1125 ( .A(n1095), .Z(n1109) );
  XNOR U1126 ( .A(n1092), .B(n1110), .Z(n1095) );
  AND U1127 ( .A(n746), .B(n400), .Z(n1110) );
  XOR U1128 ( .A(n1111), .B(n1112), .Z(n1092) );
  ANDN U1129 ( .A(n1113), .B(n1114), .Z(n1112) );
  XNOR U1130 ( .A(n1115), .B(n1111), .Z(n1113) );
  XNOR U1131 ( .A(n1116), .B(n1117), .Z(n944) );
  IV U1132 ( .A(n1105), .Z(n1117) );
  XNOR U1133 ( .A(n1102), .B(n1118), .Z(n1105) );
  AND U1134 ( .A(n310), .B(e_input[0]), .Z(n1118) );
  XNOR U1135 ( .A(n1101), .B(g_input[10]), .Z(n1100) );
  NOR U1136 ( .A(n1119), .B(n1120), .Z(n1101) );
  XOR U1137 ( .A(n1124), .B(n1106), .Z(n1116) );
  NAND U1138 ( .A(n353), .B(n1025), .Z(n1106) );
  IV U1139 ( .A(n1108), .Z(n1124) );
  XNOR U1140 ( .A(n1126), .B(n1115), .Z(n969) );
  NAND U1141 ( .A(n516), .B(n680), .Z(n1115) );
  IV U1142 ( .A(n1114), .Z(n1126) );
  XNOR U1143 ( .A(n1111), .B(n1127), .Z(n1114) );
  AND U1144 ( .A(n746), .B(n458), .Z(n1127) );
  XOR U1145 ( .A(n1128), .B(n1129), .Z(n1111) );
  ANDN U1146 ( .A(n1130), .B(n1131), .Z(n1129) );
  XNOR U1147 ( .A(n1132), .B(n1128), .Z(n1130) );
  XNOR U1148 ( .A(n1133), .B(n1134), .Z(n971) );
  IV U1149 ( .A(n1122), .Z(n1134) );
  XNOR U1150 ( .A(n1121), .B(n1135), .Z(n1122) );
  AND U1151 ( .A(n353), .B(e_input[0]), .Z(n1135) );
  XOR U1152 ( .A(n1119), .B(g_input[9]), .Z(n1120) );
  NANDN U1153 ( .B(n1136), .A(n1137), .Z(n1119) );
  XOR U1154 ( .A(n1138), .B(n1139), .Z(n1121) );
  ANDN U1155 ( .A(n1140), .B(n1141), .Z(n1139) );
  XNOR U1156 ( .A(n1142), .B(n1138), .Z(n1140) );
  XOR U1157 ( .A(n1143), .B(n1123), .Z(n1133) );
  NAND U1158 ( .A(n400), .B(n1025), .Z(n1123) );
  IV U1159 ( .A(n1125), .Z(n1143) );
  NAND U1160 ( .A(n577), .B(n680), .Z(n1132) );
  XNOR U1161 ( .A(n1128), .B(n1145), .Z(n1131) );
  AND U1162 ( .A(n746), .B(n516), .Z(n1145) );
  XNOR U1163 ( .A(n1149), .B(n1146), .Z(n1148) );
  XNOR U1164 ( .A(n1138), .B(n1151), .Z(n1141) );
  AND U1165 ( .A(n400), .B(e_input[0]), .Z(n1151) );
  XNOR U1166 ( .A(n1155), .B(n1152), .Z(n1154) );
  XOR U1167 ( .A(n1156), .B(n1142), .Z(n1150) );
  NAND U1168 ( .A(n458), .B(n1025), .Z(n1142) );
  IV U1169 ( .A(n1144), .Z(n1156) );
  XNOR U1170 ( .A(n1157), .B(n1158), .Z(n1144) );
  AND U1171 ( .A(n1159), .B(n1160), .Z(n1158) );
  XOR U1172 ( .A(n1153), .B(n1161), .Z(n1160) );
  XNOR U1173 ( .A(n1155), .B(n1157), .Z(n1161) );
  NAND U1174 ( .A(n516), .B(n1025), .Z(n1155) );
  XOR U1175 ( .A(n1152), .B(n1162), .Z(n1153) );
  AND U1176 ( .A(n458), .B(e_input[0]), .Z(n1162) );
  XNOR U1177 ( .A(n1166), .B(n1163), .Z(n1165) );
  XOR U1178 ( .A(n1147), .B(n1167), .Z(n1159) );
  XNOR U1179 ( .A(n1149), .B(n1157), .Z(n1167) );
  NANDN U1180 ( .B(n642), .A(n680), .Z(n1149) );
  XOR U1181 ( .A(n1146), .B(n1168), .Z(n1147) );
  AND U1182 ( .A(n746), .B(n577), .Z(n1168) );
  XOR U1183 ( .A(n1169), .B(n1170), .Z(n1146) );
  AND U1184 ( .A(n1171), .B(n1172), .Z(n1170) );
  XNOR U1185 ( .A(n1173), .B(n1169), .Z(n1172) );
  XOR U1186 ( .A(n1174), .B(n1175), .Z(n1157) );
  AND U1187 ( .A(n1176), .B(n1177), .Z(n1175) );
  XOR U1188 ( .A(n1164), .B(n1178), .Z(n1177) );
  XNOR U1189 ( .A(n1166), .B(n1174), .Z(n1178) );
  NAND U1190 ( .A(n577), .B(n1025), .Z(n1166) );
  XOR U1191 ( .A(n1163), .B(n1179), .Z(n1164) );
  AND U1192 ( .A(n516), .B(e_input[0]), .Z(n1179) );
  XOR U1193 ( .A(n1180), .B(n1181), .Z(n1163) );
  AND U1194 ( .A(n1182), .B(n1183), .Z(n1181) );
  XNOR U1195 ( .A(n1184), .B(n1180), .Z(n1183) );
  XOR U1196 ( .A(n1171), .B(n1185), .Z(n1176) );
  XNOR U1197 ( .A(n1173), .B(n1174), .Z(n1185) );
  NANDN U1198 ( .B(n714), .A(n680), .Z(n1173) );
  XOR U1199 ( .A(n1169), .B(n1186), .Z(n1171) );
  ANDN U1200 ( .A(n746), .B(n642), .Z(n1186) );
  XNOR U1201 ( .A(n1190), .B(n1187), .Z(n1189) );
  XOR U1202 ( .A(n1191), .B(n1192), .Z(n1174) );
  AND U1203 ( .A(n1193), .B(n1194), .Z(n1192) );
  XOR U1204 ( .A(n1182), .B(n1195), .Z(n1194) );
  XNOR U1205 ( .A(n1184), .B(n1191), .Z(n1195) );
  NANDN U1206 ( .B(n642), .A(n1025), .Z(n1184) );
  XOR U1207 ( .A(n1180), .B(n1196), .Z(n1182) );
  AND U1208 ( .A(n577), .B(e_input[0]), .Z(n1196) );
  XOR U1209 ( .A(n1188), .B(n1200), .Z(n1193) );
  XNOR U1210 ( .A(n1190), .B(n1191), .Z(n1200) );
  NAND U1211 ( .A(n680), .B(n785), .Z(n1190) );
  XOR U1212 ( .A(n1187), .B(n1201), .Z(n1188) );
  ANDN U1213 ( .A(n746), .B(n714), .Z(n1201) );
  XOR U1214 ( .A(n1202), .B(n1203), .Z(n1187) );
  ANDN U1215 ( .A(n1204), .B(n1205), .Z(n1203) );
  XNOR U1216 ( .A(n1206), .B(n1202), .Z(n1204) );
  NAND U1217 ( .A(n680), .B(n1008), .Z(n1206) );
  XNOR U1218 ( .A(n1202), .B(n1208), .Z(n1205) );
  AND U1219 ( .A(n785), .B(n746), .Z(n1208) );
  AND U1220 ( .A(n1209), .B(g_input[0]), .Z(n1202) );
  NANDN U1221 ( .B(n680), .A(n1210), .Z(n1209) );
  NAND U1222 ( .A(n1008), .B(n746), .Z(n1210) );
  XNOR U1223 ( .A(n1197), .B(n1214), .Z(n1198) );
  ANDN U1224 ( .A(e_input[0]), .B(n642), .Z(n1214) );
  XOR U1225 ( .A(n1217), .B(n1215), .Z(n1216) );
  ANDN U1226 ( .A(e_input[0]), .B(n714), .Z(n1217) );
  AND U1227 ( .A(n1025), .B(n785), .Z(n1218) );
  XOR U1228 ( .A(n1222), .B(n1199), .Z(n1213) );
  NANDN U1229 ( .B(n714), .A(n1025), .Z(n1199) );
  IV U1230 ( .A(n1207), .Z(n1222) );
  NAND U1231 ( .A(n1025), .B(n1008), .Z(n1221) );
  XNOR U1232 ( .A(n1219), .B(n1223), .Z(n1220) );
  AND U1233 ( .A(n785), .B(e_input[0]), .Z(n1223) );
  AND U1234 ( .A(n1224), .B(g_input[0]), .Z(n1219) );
  NANDN U1235 ( .B(n1025), .A(n1225), .Z(n1224) );
  NAND U1236 ( .A(n1008), .B(e_input[0]), .Z(n1225) );
  XNOR U1237 ( .A(n1227), .B(n773), .Z(n761) );
  XNOR U1238 ( .A(n758), .B(n759), .Z(n773) );
  NAND U1239 ( .A(n253), .B(n577), .Z(n759) );
  XNOR U1240 ( .A(n757), .B(n1228), .Z(n758) );
  AND U1241 ( .A(n516), .B(n289), .Z(n1228) );
  XNOR U1242 ( .A(n1232), .B(n1229), .Z(n1231) );
  XNOR U1243 ( .A(n772), .B(n760), .Z(n1227) );
  XOR U1244 ( .A(n1233), .B(n1234), .Z(n760) );
  XNOR U1245 ( .A(n765), .B(n1236), .Z(n768) );
  AND U1246 ( .A(n400), .B(n385), .Z(n1236) );
  XNOR U1247 ( .A(n1137), .B(g_input[8]), .Z(n1136) );
  NOR U1248 ( .A(n1237), .B(n1238), .Z(n1137) );
  XOR U1249 ( .A(n1239), .B(n1240), .Z(n765) );
  AND U1250 ( .A(n1241), .B(n1242), .Z(n1240) );
  XNOR U1251 ( .A(n1243), .B(n1239), .Z(n1242) );
  XOR U1252 ( .A(n1244), .B(n769), .Z(n1235) );
  NAND U1253 ( .A(n338), .B(n458), .Z(n769) );
  IV U1254 ( .A(n771), .Z(n1244) );
  XNOR U1255 ( .A(n1245), .B(n1246), .Z(n771) );
  AND U1256 ( .A(n1247), .B(n1248), .Z(n1246) );
  XOR U1257 ( .A(n1241), .B(n1249), .Z(n1248) );
  XNOR U1258 ( .A(n1243), .B(n1245), .Z(n1249) );
  NAND U1259 ( .A(n338), .B(n516), .Z(n1243) );
  XOR U1260 ( .A(n1239), .B(n1250), .Z(n1241) );
  AND U1261 ( .A(n458), .B(n385), .Z(n1250) );
  XOR U1262 ( .A(n1237), .B(g_input[7]), .Z(n1238) );
  NANDN U1263 ( .B(n1251), .A(n1252), .Z(n1237) );
  XOR U1264 ( .A(n1253), .B(n1254), .Z(n1239) );
  AND U1265 ( .A(n1255), .B(n1256), .Z(n1254) );
  XNOR U1266 ( .A(n1257), .B(n1253), .Z(n1256) );
  XOR U1267 ( .A(n1230), .B(n1258), .Z(n1247) );
  XNOR U1268 ( .A(n1232), .B(n1245), .Z(n1258) );
  NANDN U1269 ( .B(n642), .A(n253), .Z(n1232) );
  XOR U1270 ( .A(n1229), .B(n1259), .Z(n1230) );
  AND U1271 ( .A(n577), .B(n289), .Z(n1259) );
  XOR U1272 ( .A(n1260), .B(n1261), .Z(n1229) );
  AND U1273 ( .A(n1262), .B(n1263), .Z(n1261) );
  XNOR U1274 ( .A(n1264), .B(n1260), .Z(n1263) );
  XOR U1275 ( .A(n1265), .B(n1266), .Z(n1245) );
  AND U1276 ( .A(n1267), .B(n1268), .Z(n1266) );
  XOR U1277 ( .A(n1255), .B(n1269), .Z(n1268) );
  XNOR U1278 ( .A(n1257), .B(n1265), .Z(n1269) );
  NAND U1279 ( .A(n338), .B(n577), .Z(n1257) );
  XOR U1280 ( .A(n1253), .B(n1270), .Z(n1255) );
  AND U1281 ( .A(n516), .B(n385), .Z(n1270) );
  XNOR U1282 ( .A(n1252), .B(g_input[6]), .Z(n1251) );
  NOR U1283 ( .A(n1271), .B(n1272), .Z(n1252) );
  XOR U1284 ( .A(n1273), .B(n1274), .Z(n1253) );
  AND U1285 ( .A(n1275), .B(n1276), .Z(n1274) );
  XNOR U1286 ( .A(n1277), .B(n1273), .Z(n1276) );
  XOR U1287 ( .A(n1262), .B(n1278), .Z(n1267) );
  XNOR U1288 ( .A(n1264), .B(n1265), .Z(n1278) );
  NANDN U1289 ( .B(n714), .A(n253), .Z(n1264) );
  XOR U1290 ( .A(n1260), .B(n1279), .Z(n1262) );
  ANDN U1291 ( .A(n289), .B(n642), .Z(n1279) );
  XNOR U1292 ( .A(n1283), .B(n1280), .Z(n1282) );
  XOR U1293 ( .A(n1284), .B(n1285), .Z(n1265) );
  AND U1294 ( .A(n1286), .B(n1287), .Z(n1285) );
  XOR U1295 ( .A(n1275), .B(n1288), .Z(n1287) );
  XNOR U1296 ( .A(n1277), .B(n1284), .Z(n1288) );
  NANDN U1297 ( .B(n642), .A(n338), .Z(n1277) );
  XOR U1298 ( .A(n1273), .B(n1289), .Z(n1275) );
  AND U1299 ( .A(n577), .B(n385), .Z(n1289) );
  XOR U1300 ( .A(n1271), .B(g_input[5]), .Z(n1272) );
  NANDN U1301 ( .B(n1290), .A(n1291), .Z(n1271) );
  XOR U1302 ( .A(n1292), .B(n1293), .Z(n1273) );
  ANDN U1303 ( .A(n1294), .B(n1295), .Z(n1293) );
  XNOR U1304 ( .A(n1296), .B(n1292), .Z(n1294) );
  XOR U1305 ( .A(n1281), .B(n1297), .Z(n1286) );
  XNOR U1306 ( .A(n1283), .B(n1284), .Z(n1297) );
  NAND U1307 ( .A(n253), .B(n785), .Z(n1283) );
  XOR U1308 ( .A(n1280), .B(n1298), .Z(n1281) );
  ANDN U1309 ( .A(n289), .B(n714), .Z(n1298) );
  NAND U1310 ( .A(n253), .B(n1008), .Z(n1301) );
  XNOR U1311 ( .A(n1299), .B(n1303), .Z(n1300) );
  AND U1312 ( .A(n785), .B(n289), .Z(n1303) );
  AND U1313 ( .A(n1304), .B(g_input[0]), .Z(n1299) );
  NANDN U1314 ( .B(n253), .A(n1305), .Z(n1304) );
  NAND U1315 ( .A(n1008), .B(n289), .Z(n1305) );
  XNOR U1316 ( .A(n1308), .B(n1309), .Z(n1234) );
  IV U1317 ( .A(n1295), .Z(n1309) );
  XNOR U1318 ( .A(n1292), .B(n1310), .Z(n1295) );
  ANDN U1319 ( .A(n385), .B(n642), .Z(n1310) );
  XOR U1320 ( .A(n1311), .B(n1312), .Z(n1292) );
  AND U1321 ( .A(n1313), .B(n1314), .Z(n1312) );
  XOR U1322 ( .A(n1315), .B(n1311), .Z(n1314) );
  ANDN U1323 ( .A(n385), .B(n714), .Z(n1315) );
  XOR U1324 ( .A(n1316), .B(n1311), .Z(n1313) );
  AND U1325 ( .A(n785), .B(n338), .Z(n1316) );
  XOR U1326 ( .A(n1317), .B(n1318), .Z(n1311) );
  ANDN U1327 ( .A(n1319), .B(n1320), .Z(n1318) );
  XNOR U1328 ( .A(n1321), .B(n1317), .Z(n1319) );
  XOR U1329 ( .A(n1322), .B(n1296), .Z(n1308) );
  NANDN U1330 ( .B(n714), .A(n338), .Z(n1296) );
  IV U1331 ( .A(n1302), .Z(n1322) );
  XOR U1332 ( .A(n1323), .B(n1321), .Z(n1302) );
  NAND U1333 ( .A(n338), .B(n1008), .Z(n1321) );
  IV U1334 ( .A(n1320), .Z(n1323) );
  XNOR U1335 ( .A(n1317), .B(n1324), .Z(n1320) );
  AND U1336 ( .A(n785), .B(n385), .Z(n1324) );
  AND U1337 ( .A(n1325), .B(g_input[0]), .Z(n1317) );
  NANDN U1338 ( .B(n338), .A(n1326), .Z(n1325) );
  NAND U1339 ( .A(n1008), .B(n385), .Z(n1326) );
  XNOR U1340 ( .A(n776), .B(n1330), .Z(n779) );
  ANDN U1341 ( .A(n226), .B(n642), .Z(n1330) );
  XNOR U1342 ( .A(n1291), .B(g_input[4]), .Z(n1290) );
  NOR U1343 ( .A(n1331), .B(n1332), .Z(n1291) );
  XOR U1344 ( .A(n1333), .B(n1334), .Z(n776) );
  AND U1345 ( .A(n1335), .B(n1336), .Z(n1334) );
  XOR U1346 ( .A(n1337), .B(n1333), .Z(n1336) );
  ANDN U1347 ( .A(n226), .B(n714), .Z(n1337) );
  XOR U1348 ( .A(n1338), .B(n1333), .Z(n1335) );
  AND U1349 ( .A(n785), .B(n191), .Z(n1338) );
  XOR U1350 ( .A(n1339), .B(n1340), .Z(n1333) );
  ANDN U1351 ( .A(n1341), .B(n1342), .Z(n1340) );
  XNOR U1352 ( .A(n1343), .B(n1339), .Z(n1341) );
  XOR U1353 ( .A(n1344), .B(n780), .Z(n1329) );
  NANDN U1354 ( .B(n714), .A(n191), .Z(n780) );
  NANDN U1355 ( .B(n1345), .A(n1346), .Z(n1331) );
  IV U1356 ( .A(n782), .Z(n1344) );
  XOR U1357 ( .A(n1347), .B(n1343), .Z(n782) );
  NAND U1358 ( .A(n191), .B(n1008), .Z(n1343) );
  IV U1359 ( .A(n1342), .Z(n1347) );
  XNOR U1360 ( .A(n1339), .B(n1348), .Z(n1342) );
  AND U1361 ( .A(n785), .B(n226), .Z(n1348) );
  AND U1362 ( .A(n1349), .B(g_input[0]), .Z(n1339) );
  NANDN U1363 ( .B(n191), .A(n1350), .Z(n1349) );
  NAND U1364 ( .A(n1008), .B(n226), .Z(n1350) );
  XNOR U1365 ( .A(n789), .B(n790), .Z(n784) );
  NANDN U1366 ( .B(n141), .A(n1008), .Z(n790) );
  XNOR U1367 ( .A(n788), .B(n1353), .Z(n789) );
  AND U1368 ( .A(n785), .B(n161), .Z(n1353) );
  XNOR U1369 ( .A(n1346), .B(g_input[2]), .Z(n1345) );
  AND U1370 ( .A(n1355), .B(g_input[0]), .Z(n788) );
  NAND U1371 ( .A(n1356), .B(n141), .Z(n1355) );
  NANDN U1372 ( .B(n1357), .A(n1358), .Z(n141) );
  ANDN U1373 ( .A(e_input[15]), .B(n1359), .Z(n1358) );
  NAND U1374 ( .A(n1008), .B(n161), .Z(n1356) );
  XOR U1375 ( .A(n1359), .B(e_input[14]), .Z(n1357) );
  OR U1376 ( .A(n1352), .B(n1360), .Z(n1359) );
  XOR U1377 ( .A(n1360), .B(e_input[13]), .Z(n1352) );
  OR U1378 ( .A(n1351), .B(n1361), .Z(n1360) );
  XOR U1379 ( .A(n1361), .B(e_input[12]), .Z(n1351) );
  OR U1380 ( .A(n1307), .B(n1362), .Z(n1361) );
  XOR U1381 ( .A(n1362), .B(e_input[11]), .Z(n1307) );
  OR U1382 ( .A(n1306), .B(n1363), .Z(n1362) );
  XOR U1383 ( .A(n1363), .B(e_input[10]), .Z(n1306) );
  OR U1384 ( .A(n1328), .B(n1364), .Z(n1363) );
  XOR U1385 ( .A(n1364), .B(e_input[9]), .Z(n1328) );
  OR U1386 ( .A(n1327), .B(n1365), .Z(n1364) );
  XOR U1387 ( .A(n1365), .B(e_input[8]), .Z(n1327) );
  OR U1388 ( .A(n1018), .B(n1366), .Z(n1365) );
  XOR U1389 ( .A(n1366), .B(e_input[7]), .Z(n1018) );
  OR U1390 ( .A(n1017), .B(n1367), .Z(n1366) );
  XOR U1391 ( .A(n1367), .B(e_input[6]), .Z(n1017) );
  OR U1392 ( .A(n1013), .B(n1368), .Z(n1367) );
  XOR U1393 ( .A(n1368), .B(e_input[5]), .Z(n1013) );
  OR U1394 ( .A(n1012), .B(n1369), .Z(n1368) );
  XOR U1395 ( .A(n1369), .B(e_input[4]), .Z(n1012) );
  OR U1396 ( .A(n1212), .B(n1370), .Z(n1369) );
  XOR U1397 ( .A(n1370), .B(e_input[3]), .Z(n1212) );
  OR U1398 ( .A(n1211), .B(n1371), .Z(n1370) );
  XOR U1399 ( .A(n1371), .B(e_input[2]), .Z(n1211) );
  NANDN U1400 ( .B(e_input[0]), .A(n1226), .Z(n1371) );
  XNOR U1401 ( .A(e_input[0]), .B(e_input[1]), .Z(n1226) );
  XOR U1402 ( .A(g_input[0]), .B(g_input[1]), .Z(n1354) );
  AND U1403 ( .A(n1372), .B(n1373), .Z(\_MxM/N23 ) );
  XOR U1404 ( .A(\_MxM/n[9] ), .B(\_MxM/add_43/carry[9] ), .Z(n1373) );
  AND U1405 ( .A(\_MxM/N12 ), .B(n1372), .Z(\_MxM/N22 ) );
  AND U1406 ( .A(\_MxM/N11 ), .B(n1372), .Z(\_MxM/N21 ) );
  AND U1407 ( .A(\_MxM/N10 ), .B(n1372), .Z(\_MxM/N20 ) );
  AND U1408 ( .A(\_MxM/N9 ), .B(n1372), .Z(\_MxM/N19 ) );
  AND U1409 ( .A(\_MxM/N8 ), .B(n1372), .Z(\_MxM/N18 ) );
  AND U1410 ( .A(\_MxM/N7 ), .B(n1372), .Z(\_MxM/N17 ) );
  AND U1411 ( .A(\_MxM/N6 ), .B(n1372), .Z(\_MxM/N16 ) );
  AND U1412 ( .A(\_MxM/N5 ), .B(n1372), .Z(\_MxM/N15 ) );
  NAND U1413 ( .A(n1374), .B(n1375), .Z(n1372) );
  AND U1414 ( .A(n1376), .B(n1377), .Z(n1375) );
  AND U1415 ( .A(\_MxM/n[1] ), .B(n1378), .Z(n1377) );
  NOR U1416 ( .A(\_MxM/N14 ), .B(n107), .Z(n1378) );
  OR U1417 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n107) );
  AND U1418 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n1376) );
  AND U1419 ( .A(n1379), .B(n1380), .Z(n1374) );
  AND U1420 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n1380) );
  AND U1421 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n1379) );
  IV U1422 ( .A(\_MxM/n[0] ), .Z(\_MxM/N14 ) );
endmodule

