
module MxM_TG_W32_N1000 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MxM/n372 , \_MxM/n371 , \_MxM/n370 , \_MxM/n369 , \_MxM/n368 ,
         \_MxM/n367 , \_MxM/n366 , \_MxM/n365 , \_MxM/n364 , \_MxM/n363 ,
         \_MxM/n362 , \_MxM/n361 , \_MxM/n360 , \_MxM/n359 , \_MxM/n358 ,
         \_MxM/n357 , \_MxM/n356 , \_MxM/n355 , \_MxM/n354 , \_MxM/n353 ,
         \_MxM/n352 , \_MxM/n351 , \_MxM/n350 , \_MxM/n349 , \_MxM/n348 ,
         \_MxM/n347 , \_MxM/n346 , \_MxM/n345 , \_MxM/n344 , \_MxM/n343 ,
         \_MxM/n342 , \_MxM/n341 , \_MxM/n340 , \_MxM/n339 , \_MxM/n338 ,
         \_MxM/n337 , \_MxM/n336 , \_MxM/n335 , \_MxM/n334 , \_MxM/n333 ,
         \_MxM/n332 , \_MxM/n331 , \_MxM/n330 , \_MxM/n329 , \_MxM/n328 ,
         \_MxM/n327 , \_MxM/n326 , \_MxM/n325 , \_MxM/n324 , \_MxM/n323 ,
         \_MxM/n322 , \_MxM/n321 , \_MxM/n320 , \_MxM/n319 , \_MxM/n318 ,
         \_MxM/n317 , \_MxM/n316 , \_MxM/n315 , \_MxM/n314 , \_MxM/n313 ,
         \_MxM/n312 , \_MxM/n311 , \_MxM/n310 , \_MxM/n309 , \_MxM/n308 ,
         \_MxM/n307 , \_MxM/n306 , \_MxM/n305 , \_MxM/n304 , \_MxM/n303 ,
         \_MxM/n302 , \_MxM/n301 , \_MxM/n300 , \_MxM/n299 , \_MxM/N15 ,
         \_MxM/N14 , \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 ,
         \_MxM/N8 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] ,
         \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] ,
         \_MxM/n[9] , \_MxM/Y0[0] , \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] ,
         \_MxM/Y0[4] , \_MxM/Y0[5] , \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/Y0[8] ,
         \_MxM/Y0[9] , \_MxM/Y0[10] , \_MxM/Y0[11] , \_MxM/Y0[12] ,
         \_MxM/Y0[13] , \_MxM/Y0[14] , \_MxM/Y0[15] , \_MxM/Y0[16] ,
         \_MxM/Y0[17] , \_MxM/Y0[18] , \_MxM/Y0[19] , \_MxM/Y0[20] ,
         \_MxM/Y0[21] , \_MxM/Y0[22] , \_MxM/Y0[23] , \_MxM/Y0[24] ,
         \_MxM/Y0[25] , \_MxM/Y0[26] , \_MxM/Y0[27] , \_MxM/Y0[28] ,
         \_MxM/Y0[29] , \_MxM/Y0[30] , \_MxM/Y0[31] , \_MxM/add_39/carry[9] ,
         \_MxM/add_39/carry[8] , \_MxM/add_39/carry[7] ,
         \_MxM/add_39/carry[6] , \_MxM/add_39/carry[5] ,
         \_MxM/add_39/carry[4] , \_MxM/add_39/carry[3] ,
         \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n299 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n300 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n301 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n302 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n303 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n304 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n305 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n306 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n307 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n308 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n309 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n310 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n311 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n312 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n313 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n314 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y_reg[16]  ( .D(\_MxM/n315 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[16]) );
  DFF \_MxM/Y_reg[17]  ( .D(\_MxM/n316 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[17]) );
  DFF \_MxM/Y_reg[18]  ( .D(\_MxM/n317 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[18]) );
  DFF \_MxM/Y_reg[19]  ( .D(\_MxM/n318 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[19]) );
  DFF \_MxM/Y_reg[20]  ( .D(\_MxM/n319 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[20]) );
  DFF \_MxM/Y_reg[21]  ( .D(\_MxM/n320 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[21]) );
  DFF \_MxM/Y_reg[22]  ( .D(\_MxM/n321 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[22]) );
  DFF \_MxM/Y_reg[23]  ( .D(\_MxM/n322 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[23]) );
  DFF \_MxM/Y_reg[24]  ( .D(\_MxM/n323 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[24]) );
  DFF \_MxM/Y_reg[25]  ( .D(\_MxM/n324 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[25]) );
  DFF \_MxM/Y_reg[26]  ( .D(\_MxM/n325 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[26]) );
  DFF \_MxM/Y_reg[27]  ( .D(\_MxM/n326 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[27]) );
  DFF \_MxM/Y_reg[28]  ( .D(\_MxM/n327 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[28]) );
  DFF \_MxM/Y_reg[29]  ( .D(\_MxM/n328 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[29]) );
  DFF \_MxM/Y_reg[30]  ( .D(\_MxM/n329 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[30]) );
  DFF \_MxM/Y_reg[31]  ( .D(\_MxM/n330 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[31]) );
  DFF \_MxM/Y0_reg[31]  ( .D(\_MxM/n331 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[31] ) );
  DFF \_MxM/Y0_reg[30]  ( .D(\_MxM/n332 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[30] ) );
  DFF \_MxM/Y0_reg[29]  ( .D(\_MxM/n333 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[29] ) );
  DFF \_MxM/Y0_reg[28]  ( .D(\_MxM/n334 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[28] ) );
  DFF \_MxM/Y0_reg[27]  ( .D(\_MxM/n335 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[27] ) );
  DFF \_MxM/Y0_reg[26]  ( .D(\_MxM/n336 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[26] ) );
  DFF \_MxM/Y0_reg[25]  ( .D(\_MxM/n337 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[25] ) );
  DFF \_MxM/Y0_reg[24]  ( .D(\_MxM/n338 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[24] ) );
  DFF \_MxM/Y0_reg[23]  ( .D(\_MxM/n339 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[23] ) );
  DFF \_MxM/Y0_reg[22]  ( .D(\_MxM/n340 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[22] ) );
  DFF \_MxM/Y0_reg[21]  ( .D(\_MxM/n341 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[21] ) );
  DFF \_MxM/Y0_reg[20]  ( .D(\_MxM/n342 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[20] ) );
  DFF \_MxM/Y0_reg[19]  ( .D(\_MxM/n343 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[19] ) );
  DFF \_MxM/Y0_reg[18]  ( .D(\_MxM/n344 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[18] ) );
  DFF \_MxM/Y0_reg[17]  ( .D(\_MxM/n345 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[17] ) );
  DFF \_MxM/Y0_reg[16]  ( .D(\_MxM/n346 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[16] ) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/n347 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/n348 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/n349 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/n350 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/n351 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/n352 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/n353 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/n354 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n355 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n356 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n357 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n358 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n359 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n360 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n361 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n362 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/n363 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/n364 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/n365 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n366 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n367 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n368 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n369 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n370 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n371 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n372 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N14 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N15 ) );
  MUX U1 ( .IN0(n3708), .IN1(n1), .SEL(n3709), .F(n3662) );
  IV U2 ( .A(n3710), .Z(n1) );
  MUX U3 ( .IN0(n3536), .IN1(n3538), .SEL(n3537), .F(n3490) );
  MUX U4 ( .IN0(n4309), .IN1(n4311), .SEL(n4310), .F(n4285) );
  MUX U5 ( .IN0(n3361), .IN1(n3363), .SEL(n3362), .F(n3315) );
  XNOR U6 ( .A(n4297), .B(n4296), .Z(n4312) );
  XNOR U7 ( .A(n4680), .B(n4678), .Z(n4685) );
  MUX U8 ( .IN0(n3265), .IN1(n3267), .SEL(n3266), .F(n3222) );
  MUX U9 ( .IN0(n5013), .IN1(n5015), .SEL(n5014), .F(n5001) );
  MUX U10 ( .IN0(n4871), .IN1(n2), .SEL(n4872), .F(n4851) );
  IV U11 ( .A(n4873), .Z(n2) );
  MUX U12 ( .IN0(n5020), .IN1(n3), .SEL(n5021), .F(n5008) );
  IV U13 ( .A(n5022), .Z(n3) );
  MUX U14 ( .IN0(n4230), .IN1(n4), .SEL(n4231), .F(n4210) );
  IV U15 ( .A(n4232), .Z(n4) );
  XNOR U16 ( .A(n3218), .B(n3217), .Z(n3254) );
  MUX U17 ( .IN0(n4635), .IN1(n5), .SEL(n4636), .F(n4625) );
  IV U18 ( .A(n4637), .Z(n5) );
  XNOR U19 ( .A(n3243), .B(n3241), .Z(n3278) );
  XNOR U20 ( .A(n4406), .B(n4404), .Z(n4413) );
  NANDN U21 ( .B(n1294), .A(n3019), .Z(n18) );
  MUX U22 ( .IN0(n3095), .IN1(n3097), .SEL(n3096), .F(n3056) );
  MUX U23 ( .IN0(n3088), .IN1(n6), .SEL(n3089), .F(n3049) );
  IV U24 ( .A(n3090), .Z(n6) );
  MUX U25 ( .IN0(n3100), .IN1(n3102), .SEL(n3101), .F(n3029) );
  MUX U26 ( .IN0(n1005), .IN1(n7), .SEL(n1006), .F(n936) );
  IV U27 ( .A(n1007), .Z(n7) );
  MUX U28 ( .IN0(n1302), .IN1(n1304), .SEL(n1303), .F(n1218) );
  MUX U29 ( .IN0(n1357), .IN1(n8), .SEL(n1358), .F(n1266) );
  IV U30 ( .A(n1359), .Z(n8) );
  MUX U31 ( .IN0(n1405), .IN1(n9), .SEL(n1406), .F(n1310) );
  IV U32 ( .A(n1407), .Z(n9) );
  MUX U33 ( .IN0(n1510), .IN1(n10), .SEL(n1511), .F(n1413) );
  IV U34 ( .A(n1512), .Z(n10) );
  MUX U35 ( .IN0(n1769), .IN1(n1771), .SEL(n1770), .F(n1668) );
  MUX U36 ( .IN0(n1885), .IN1(n11), .SEL(n1886), .F(n1777) );
  IV U37 ( .A(n1887), .Z(n11) );
  MUX U38 ( .IN0(n2058), .IN1(n12), .SEL(n2059), .F(n1949) );
  IV U39 ( .A(n2060), .Z(n12) );
  MUX U40 ( .IN0(g_input[29]), .IN1(n4381), .SEL(g_input[31]), .F(n13) );
  IV U41 ( .A(n13), .Z(n629) );
  MUX U42 ( .IN0(n14), .IN1(n4370), .SEL(g_input[31]), .F(n585) );
  IV U43 ( .A(g_input[30]), .Z(n14) );
  MUX U44 ( .IN0(n4932), .IN1(n4934), .SEL(n4933), .F(n4908) );
  MUX U45 ( .IN0(n4682), .IN1(n4684), .SEL(n4683), .F(n4667) );
  XNOR U46 ( .A(n5054), .B(n5052), .Z(n5059) );
  MUX U47 ( .IN0(n4265), .IN1(n4267), .SEL(n4266), .F(n4245) );
  MUX U48 ( .IN0(n4270), .IN1(n15), .SEL(n4271), .F(n4250) );
  IV U49 ( .A(n4272), .Z(n15) );
  XNOR U50 ( .A(n4920), .B(n4919), .Z(n4935) );
  MUX U51 ( .IN0(n5001), .IN1(n5003), .SEL(n5002), .F(n4989) );
  MUX U52 ( .IN0(n4851), .IN1(n16), .SEL(n4852), .F(n4831) );
  IV U53 ( .A(n4853), .Z(n16) );
  MUX U54 ( .IN0(n5008), .IN1(n17), .SEL(n5009), .F(n4996) );
  IV U55 ( .A(n5010), .Z(n17) );
  MUX U56 ( .IN0(n3180), .IN1(n3182), .SEL(n3181), .F(n3135) );
  XNOR U57 ( .A(n4638), .B(n4637), .Z(n4643) );
  MUX U58 ( .IN0(n4630), .IN1(n4632), .SEL(n4631), .F(n4620) );
  MUX U59 ( .IN0(n5125), .IN1(n18), .SEL(n5126), .F(n5114) );
  XNOR U60 ( .A(n3131), .B(n3130), .Z(n3169) );
  MUX U61 ( .IN0(n4615), .IN1(n19), .SEL(n4616), .F(n4602) );
  IV U62 ( .A(n4617), .Z(n19) );
  MUX U63 ( .IN0(n3049), .IN1(n20), .SEL(n3050), .F(n2919) );
  IV U64 ( .A(n3051), .Z(n20) );
  MUX U65 ( .IN0(n1157), .IN1(n21), .SEL(n1158), .F(n1077) );
  IV U66 ( .A(n1159), .Z(n21) );
  MUX U67 ( .IN0(n1218), .IN1(n1220), .SEL(n1219), .F(n1137) );
  MUX U68 ( .IN0(n1275), .IN1(n1277), .SEL(n1276), .F(n1193) );
  MUX U69 ( .IN0(n1590), .IN1(n1592), .SEL(n1591), .F(n1494) );
  MUX U70 ( .IN0(n1598), .IN1(n22), .SEL(n1599), .F(n1502) );
  IV U71 ( .A(n1600), .Z(n22) );
  MUX U72 ( .IN0(n1606), .IN1(n23), .SEL(n1607), .F(n1510) );
  IV U73 ( .A(n1608), .Z(n23) );
  MUX U74 ( .IN0(n1653), .IN1(n24), .SEL(n1654), .F(n1553) );
  IV U75 ( .A(n1655), .Z(n24) );
  MUX U76 ( .IN0(n1850), .IN1(n1852), .SEL(n1851), .F(n1742) );
  MUX U77 ( .IN0(n1992), .IN1(n25), .SEL(n1993), .F(n1885) );
  IV U78 ( .A(n1994), .Z(n25) );
  MUX U79 ( .IN0(n2172), .IN1(n26), .SEL(n2173), .F(n2058) );
  IV U80 ( .A(n2174), .Z(n26) );
  MUX U81 ( .IN0(n2798), .IN1(n27), .SEL(n2799), .F(n2673) );
  IV U82 ( .A(n2800), .Z(n27) );
  MUX U83 ( .IN0(n705), .IN1(n28), .SEL(n706), .F(n659) );
  IV U84 ( .A(n707), .Z(n28) );
  MUX U85 ( .IN0(n2952), .IN1(n2954), .SEL(n2953), .F(n2814) );
  MUX U86 ( .IN0(n29), .IN1(n740), .SEL(n739), .F(n702) );
  IV U87 ( .A(n738), .Z(n29) );
  MUX U88 ( .IN0(n3716), .IN1(n3718), .SEL(n3717), .F(n3672) );
  MUX U89 ( .IN0(n4694), .IN1(n4696), .SEL(n4695), .F(n4682) );
  XNOR U90 ( .A(n4692), .B(n4691), .Z(n4697) );
  MUX U91 ( .IN0(n4886), .IN1(n4888), .SEL(n4887), .F(n4866) );
  MUX U92 ( .IN0(n5034), .IN1(n30), .SEL(n5035), .F(n5020) );
  IV U93 ( .A(n5036), .Z(n30) );
  MUX U94 ( .IN0(n4245), .IN1(n4247), .SEL(n4246), .F(n4225) );
  MUX U95 ( .IN0(n4250), .IN1(n31), .SEL(n4251), .F(n4230) );
  IV U96 ( .A(n4252), .Z(n31) );
  MUX U97 ( .IN0(n3229), .IN1(n3231), .SEL(n3230), .F(n3185) );
  XNOR U98 ( .A(n4854), .B(n4853), .Z(n4869) );
  MUX U99 ( .IN0(n4989), .IN1(n4991), .SEL(n4990), .F(n4977) );
  XNOR U100 ( .A(n4999), .B(n4998), .Z(n5004) );
  NANDN U101 ( .B(n2050), .A(n3019), .Z(n44) );
  MUX U102 ( .IN0(n4625), .IN1(n32), .SEL(n4626), .F(n4615) );
  IV U103 ( .A(n4627), .Z(n32) );
  MUX U104 ( .IN0(n4620), .IN1(n4622), .SEL(n4621), .F(n4610) );
  XNOR U105 ( .A(n3091), .B(n3090), .Z(n3124) );
  MUX U106 ( .IN0(n1397), .IN1(n1399), .SEL(n1398), .F(n1302) );
  MUX U107 ( .IN0(n1694), .IN1(n33), .SEL(n1695), .F(n1598) );
  IV U108 ( .A(n1696), .Z(n33) );
  MUX U109 ( .IN0(n1702), .IN1(n34), .SEL(n1703), .F(n1606) );
  IV U110 ( .A(n1704), .Z(n34) );
  MUX U111 ( .IN0(n1660), .IN1(n1662), .SEL(n1661), .F(n1562) );
  MUX U112 ( .IN0(n1668), .IN1(n1670), .SEL(n1669), .F(n1570) );
  MUX U113 ( .IN0(n1754), .IN1(n35), .SEL(n1755), .F(n1653) );
  IV U114 ( .A(n1756), .Z(n35) );
  MUX U115 ( .IN0(n1787), .IN1(n1789), .SEL(n1788), .F(n1686) );
  MUX U116 ( .IN0(n1958), .IN1(n1960), .SEL(n1959), .F(n1850) );
  MUX U117 ( .IN0(n2100), .IN1(n36), .SEL(n2101), .F(n1992) );
  IV U118 ( .A(n2102), .Z(n36) );
  MUX U119 ( .IN0(n2268), .IN1(n2270), .SEL(n2269), .F(n2149) );
  MUX U120 ( .IN0(n2406), .IN1(n37), .SEL(n2407), .F(n2286) );
  IV U121 ( .A(n2408), .Z(n37) );
  MUX U122 ( .IN0(n2935), .IN1(n38), .SEL(n2936), .F(n2798) );
  IV U123 ( .A(n2937), .Z(n38) );
  MUX U124 ( .IN0(n731), .IN1(n733), .SEL(n732), .F(n689) );
  MUX U125 ( .IN0(n621), .IN1(n39), .SEL(n622), .F(n575) );
  IV U126 ( .A(n623), .Z(n39) );
  MUX U127 ( .IN0(n40), .IN1(n967), .SEL(n966), .F(n902) );
  IV U128 ( .A(n965), .Z(n40) );
  MUX U129 ( .IN0(n5056), .IN1(n5058), .SEL(n5057), .F(n5039) );
  MUX U130 ( .IN0(n4937), .IN1(n41), .SEL(n4938), .F(n4915) );
  IV U131 ( .A(n4939), .Z(n41) );
  MUX U132 ( .IN0(n4755), .IN1(n4757), .SEL(n4756), .F(n4739) );
  MUX U133 ( .IN0(n4866), .IN1(n4868), .SEL(n4867), .F(n4846) );
  MUX U134 ( .IN0(n4640), .IN1(n4642), .SEL(n4641), .F(n4630) );
  XNOR U135 ( .A(n4422), .B(n4421), .Z(n4429) );
  MUX U136 ( .IN0(n4205), .IN1(n4207), .SEL(n4206), .F(n4185) );
  XNOR U137 ( .A(n4233), .B(n4232), .Z(n4248) );
  MUX U138 ( .IN0(n4831), .IN1(n42), .SEL(n4832), .F(n4811) );
  IV U139 ( .A(n4833), .Z(n42) );
  MUX U140 ( .IN0(n4996), .IN1(n43), .SEL(n4997), .F(n4984) );
  IV U141 ( .A(n4998), .Z(n43) );
  MUX U142 ( .IN0(n3801), .IN1(n44), .SEL(n3802), .F(n3790) );
  MUX U143 ( .IN0(n4977), .IN1(n4979), .SEL(n4978), .F(n4794) );
  MUX U144 ( .IN0(n4166), .IN1(n45), .SEL(n4167), .F(n4145) );
  IV U145 ( .A(n4168), .Z(n45) );
  XNOR U146 ( .A(n4618), .B(n4617), .Z(n4623) );
  MUX U147 ( .IN0(n3056), .IN1(n3058), .SEL(n3057), .F(n2926) );
  MUX U148 ( .IN0(n1466), .IN1(n1468), .SEL(n1467), .F(n1364) );
  MUX U149 ( .IN0(n1502), .IN1(n46), .SEL(n1503), .F(n1405) );
  IV U150 ( .A(n1504), .Z(n46) );
  MUX U151 ( .IN0(n1494), .IN1(n1496), .SEL(n1495), .F(n1397) );
  MUX U152 ( .IN0(n1803), .IN1(n47), .SEL(n1804), .F(n1702) );
  IV U153 ( .A(n1805), .Z(n47) );
  MUX U154 ( .IN0(n1976), .IN1(n1978), .SEL(n1977), .F(n1869) );
  MUX U155 ( .IN0(n1969), .IN1(n48), .SEL(n1970), .F(n1862) );
  IV U156 ( .A(n1971), .Z(n48) );
  MUX U157 ( .IN0(n2008), .IN1(n49), .SEL(n2009), .F(n1901) );
  IV U158 ( .A(n2010), .Z(n49) );
  MUX U159 ( .IN0(n2065), .IN1(n2067), .SEL(n2066), .F(n1958) );
  MUX U160 ( .IN0(n2219), .IN1(n50), .SEL(n2220), .F(n2100) );
  IV U161 ( .A(n2221), .Z(n50) );
  MUX U162 ( .IN0(n2636), .IN1(n2638), .SEL(n2637), .F(n2512) );
  MUX U163 ( .IN0(n2644), .IN1(n51), .SEL(n2645), .F(n2520) );
  IV U164 ( .A(n2646), .Z(n51) );
  MUX U165 ( .IN0(g_input[28]), .IN1(n4399), .SEL(g_input[31]), .F(n52) );
  IV U166 ( .A(n52), .Z(n669) );
  MUX U167 ( .IN0(n689), .IN1(n691), .SEL(n690), .F(n648) );
  XNOR U168 ( .A(n970), .B(n967), .Z(n1030) );
  MUX U169 ( .IN0(n5119), .IN1(n5121), .SEL(n5120), .F(n5103) );
  MUX U170 ( .IN0(n53), .IN1(n4734), .SEL(n4735), .F(n4720) );
  IV U171 ( .A(n4736), .Z(n53) );
  XNOR U172 ( .A(n4253), .B(n4252), .Z(n4268) );
  MUX U173 ( .IN0(n5197), .IN1(n54), .SEL(n5198), .F(n5179) );
  IV U174 ( .A(n5199), .Z(n54) );
  MUX U175 ( .IN0(n4846), .IN1(n4848), .SEL(n4847), .F(n4826) );
  MUX U176 ( .IN0(n4185), .IN1(n4187), .SEL(n4186), .F(n4173) );
  NANDN U177 ( .B(n2545), .A(n3019), .Z(n67) );
  MUX U178 ( .IN0(n4190), .IN1(n55), .SEL(n4191), .F(n4166) );
  IV U179 ( .A(n4192), .Z(n55) );
  XNOR U180 ( .A(n3900), .B(n3898), .Z(n3913) );
  XNOR U181 ( .A(n4834), .B(n4833), .Z(n4849) );
  MUX U182 ( .IN0(n4984), .IN1(n56), .SEL(n4985), .F(n4972) );
  IV U183 ( .A(n4986), .Z(n56) );
  MUX U184 ( .IN0(n4610), .IN1(n4612), .SEL(n4611), .F(n4593) );
  MUX U185 ( .IN0(n4780), .IN1(n57), .SEL(n4781), .F(n2966) );
  IV U186 ( .A(n4782), .Z(n57) );
  MUX U187 ( .IN0(n1413), .IN1(n58), .SEL(n1414), .F(n1320) );
  IV U188 ( .A(n1415), .Z(n58) );
  MUX U189 ( .IN0(n1562), .IN1(n1564), .SEL(n1563), .F(n1466) );
  MUX U190 ( .IN0(n1686), .IN1(n1688), .SEL(n1687), .F(n1590) );
  MUX U191 ( .IN0(n1862), .IN1(n59), .SEL(n1863), .F(n1754) );
  IV U192 ( .A(n1864), .Z(n59) );
  MUX U193 ( .IN0(n2016), .IN1(n60), .SEL(n2017), .F(n1909) );
  IV U194 ( .A(n2018), .Z(n60) );
  MUX U195 ( .IN0(n2116), .IN1(n61), .SEL(n2117), .F(n2008) );
  IV U196 ( .A(n2118), .Z(n61) );
  MUX U197 ( .IN0(n2211), .IN1(n2213), .SEL(n2212), .F(n2092) );
  MUX U198 ( .IN0(n2203), .IN1(n2205), .SEL(n2204), .F(n2084) );
  MUX U199 ( .IN0(n2293), .IN1(n2295), .SEL(n2294), .F(n2179) );
  MUX U200 ( .IN0(n2586), .IN1(n62), .SEL(n2587), .F(n2461) );
  IV U201 ( .A(n2588), .Z(n62) );
  MUX U202 ( .IN0(n670), .IN1(n672), .SEL(n671), .F(n630) );
  MUX U203 ( .IN0(n1042), .IN1(n1044), .SEL(n1043), .F(n974) );
  MUX U204 ( .IN0(g_input[25]), .IN1(n4448), .SEL(g_input[31]), .F(n63) );
  IV U205 ( .A(n63), .Z(n814) );
  MUX U206 ( .IN0(n2041), .IN1(n2043), .SEL(n2042), .F(n1936) );
  XNOR U207 ( .A(n801), .B(n800), .Z(n856) );
  XNOR U208 ( .A(n290), .B(n1291), .Z(n1214) );
  AND U209 ( .A(n570), .B(n572), .Z(n541) );
  MUX U210 ( .IN0(n4750), .IN1(n64), .SEL(n4751), .F(n4734) );
  IV U211 ( .A(n4752), .Z(n64) );
  XNOR U212 ( .A(n4896), .B(n4895), .Z(n4913) );
  MUX U213 ( .IN0(n3795), .IN1(n3797), .SEL(n3796), .F(n3781) );
  MUX U214 ( .IN0(n4210), .IN1(n65), .SEL(n4211), .F(n4190) );
  IV U215 ( .A(n4212), .Z(n65) );
  XNOR U216 ( .A(n3176), .B(n3175), .Z(n3211) );
  MUX U217 ( .IN0(n66), .IN1(n5179), .SEL(n5180), .F(n5163) );
  IV U218 ( .A(n5181), .Z(n66) );
  MUX U219 ( .IN0(n4826), .IN1(n4828), .SEL(n4827), .F(n4806) );
  MUX U220 ( .IN0(n4328), .IN1(n67), .SEL(n4329), .F(n4314) );
  XNOR U221 ( .A(n4628), .B(n4627), .Z(n4633) );
  MUX U222 ( .IN0(n4811), .IN1(n68), .SEL(n4812), .F(n4780) );
  IV U223 ( .A(n4813), .Z(n68) );
  XNOR U224 ( .A(n3158), .B(n3156), .Z(n3193) );
  MUX U225 ( .IN0(n4972), .IN1(n69), .SEL(n4973), .F(n2989) );
  IV U226 ( .A(n4974), .Z(n69) );
  MUX U227 ( .IN0(n1909), .IN1(n70), .SEL(n1910), .F(n1803) );
  IV U228 ( .A(n1911), .Z(n70) );
  MUX U229 ( .IN0(n2347), .IN1(n2349), .SEL(n2348), .F(n2227) );
  MUX U230 ( .IN0(n2477), .IN1(n71), .SEL(n2478), .F(n2355) );
  IV U231 ( .A(n2479), .Z(n71) );
  MUX U232 ( .IN0(n2485), .IN1(n72), .SEL(n2486), .F(n2363) );
  IV U233 ( .A(n2487), .Z(n72) );
  MUX U234 ( .IN0(g_input[22]), .IN1(n4499), .SEL(g_input[31]), .F(n73) );
  IV U235 ( .A(n73), .Z(n1013) );
  MUX U236 ( .IN0(g_input[24]), .IN1(n4465), .SEL(g_input[31]), .F(n74) );
  IV U237 ( .A(n74), .Z(n878) );
  MUX U238 ( .IN0(g_input[17]), .IN1(n4584), .SEL(g_input[31]), .F(n75) );
  IV U239 ( .A(n75), .Z(n1421) );
  MUX U240 ( .IN0(g_input[19]), .IN1(n4550), .SEL(g_input[31]), .F(n76) );
  IV U241 ( .A(n76), .Z(n1246) );
  MUX U242 ( .IN0(g_input[26]), .IN1(n4432), .SEL(g_input[31]), .F(n77) );
  IV U243 ( .A(n77), .Z(n755) );
  MUX U244 ( .IN0(g_input[27]), .IN1(n4416), .SEL(g_input[31]), .F(n78) );
  IV U245 ( .A(n78), .Z(n713) );
  MUX U246 ( .IN0(n875), .IN1(n873), .SEL(n874), .F(n809) );
  MUX U247 ( .IN0(n2552), .IN1(n2554), .SEL(n2553), .F(n2426) );
  XNOR U248 ( .A(n1038), .B(n1037), .Z(n1104) );
  XOR U249 ( .A(n1382), .B(n1297), .Z(n1298) );
  ANDN U250 ( .A(n592), .B(n572), .Z(n561) );
  XNOR U251 ( .A(n5023), .B(n5022), .Z(n5030) );
  MUX U252 ( .IN0(n3790), .IN1(n79), .SEL(n3791), .F(n3776) );
  IV U253 ( .A(n3792), .Z(n79) );
  MUX U254 ( .IN0(n4765), .IN1(n4767), .SEL(n4766), .F(n4761) );
  MUX U255 ( .IN0(n80), .IN1(n5098), .SEL(n5099), .F(n5084) );
  IV U256 ( .A(n5100), .Z(n80) );
  MUX U257 ( .IN0(n81), .IN1(n4720), .SEL(n4721), .F(n4711) );
  IV U258 ( .A(n4722), .Z(n81) );
  XNOR U259 ( .A(n4213), .B(n4212), .Z(n4228) );
  NANDN U260 ( .B(n5211), .A(n3019), .Z(n97) );
  MUX U261 ( .IN0(n4806), .IN1(n4808), .SEL(n4807), .F(n4787) );
  XNOR U262 ( .A(n4987), .B(n4986), .Z(n4992) );
  XNOR U263 ( .A(n4814), .B(n4813), .Z(n4829) );
  XNOR U264 ( .A(n3052), .B(n3051), .Z(n3086) );
  MUX U265 ( .IN0(n1901), .IN1(n82), .SEL(n1902), .F(n1795) );
  IV U266 ( .A(n1903), .Z(n82) );
  MUX U267 ( .IN0(n2196), .IN1(n83), .SEL(n2197), .F(n2077) );
  IV U268 ( .A(n2198), .Z(n83) );
  MUX U269 ( .IN0(n2388), .IN1(n2390), .SEL(n2389), .F(n2268) );
  MUX U270 ( .IN0(n2610), .IN1(n84), .SEL(n2611), .F(n2485) );
  IV U271 ( .A(n2612), .Z(n84) );
  MUX U272 ( .IN0(g_input[12]), .IN1(n5007), .SEL(g_input[31]), .F(n85) );
  IV U273 ( .A(n85), .Z(n1917) );
  MUX U274 ( .IN0(n2805), .IN1(n2807), .SEL(n2806), .F(n2680) );
  MUX U275 ( .IN0(g_input[20]), .IN1(n4533), .SEL(g_input[31]), .F(n86) );
  IV U276 ( .A(n86), .Z(n1165) );
  MUX U277 ( .IN0(n2774), .IN1(n87), .SEL(n2775), .F(n2644) );
  IV U278 ( .A(n2776), .Z(n87) );
  MUX U279 ( .IN0(g_input[15]), .IN1(n4971), .SEL(g_input[31]), .F(n88) );
  IV U280 ( .A(n88), .Z(n1614) );
  MUX U281 ( .IN0(g_input[23]), .IN1(n4482), .SEL(g_input[31]), .F(n89) );
  IV U282 ( .A(n89), .Z(n946) );
  MUX U283 ( .IN0(g_input[21]), .IN1(n4516), .SEL(g_input[31]), .F(n90) );
  IV U284 ( .A(n90), .Z(n1087) );
  MUX U285 ( .IN0(n787), .IN1(n789), .SEL(n788), .F(n731) );
  MUX U286 ( .IN0(n943), .IN1(n941), .SEL(n942), .F(n873) );
  MUX U287 ( .IN0(n1002), .IN1(n1000), .SEL(n1001), .F(n931) );
  MUX U288 ( .IN0(n1191), .IN1(n1189), .SEL(n1190), .F(n1111) );
  MUX U289 ( .IN0(n91), .IN1(n1325), .SEL(n1326), .F(n1241) );
  IV U290 ( .A(n1327), .Z(n91) );
  MUX U291 ( .IN0(n1956), .IN1(n1954), .SEL(n1955), .F(n1846) );
  MUX U292 ( .IN0(n92), .IN1(n2246), .SEL(n2247), .F(n2127) );
  IV U293 ( .A(n2248), .Z(n92) );
  MUX U294 ( .IN0(n666), .IN1(n664), .SEL(n665), .F(n624) );
  MUX U295 ( .IN0(n974), .IN1(n976), .SEL(n975), .F(n905) );
  MUX U296 ( .IN0(n93), .IN1(n1142), .SEL(n1143), .F(n1062) );
  IV U297 ( .A(n1144), .Z(n93) );
  XOR U298 ( .A(n348), .B(n1631), .Z(n1535) );
  MUX U299 ( .IN0(n1936), .IN1(n1938), .SEL(n1937), .F(n1829) );
  ANDN U300 ( .A(n561), .B(n543), .Z(n532) );
  AND U301 ( .A(n601), .B(n603), .Z(n570) );
  MUX U302 ( .IN0(n1353), .IN1(n1351), .SEL(n1352), .F(n1260) );
  MUX U303 ( .IN0(n5114), .IN1(n94), .SEL(n5115), .F(n5098) );
  IV U304 ( .A(n5116), .Z(n94) );
  MUX U305 ( .IN0(n4225), .IN1(n4227), .SEL(n4226), .F(n4205) );
  MUX U306 ( .IN0(n5202), .IN1(n5204), .SEL(n5203), .F(n5184) );
  XNOR U307 ( .A(n5011), .B(n5010), .Z(n5016) );
  MUX U308 ( .IN0(n95), .IN1(n3776), .SEL(n3777), .F(n3762) );
  IV U309 ( .A(n3778), .Z(n95) );
  MUX U310 ( .IN0(n96), .IN1(n4711), .SEL(n4712), .F(n4699) );
  IV U311 ( .A(n4713), .Z(n96) );
  MUX U312 ( .IN0(n5208), .IN1(n97), .SEL(n5209), .F(n5197) );
  MUX U313 ( .IN0(n4787), .IN1(n4789), .SEL(n4788), .F(n2973) );
  MUX U314 ( .IN0(n2124), .IN1(n98), .SEL(n2125), .F(n2016) );
  IV U315 ( .A(n2126), .Z(n98) );
  MUX U316 ( .IN0(n2092), .IN1(n2094), .SEL(n2093), .F(n1984) );
  MUX U317 ( .IN0(n2286), .IN1(n99), .SEL(n2287), .F(n2172) );
  IV U318 ( .A(n2288), .Z(n99) );
  MUX U319 ( .IN0(n2461), .IN1(n100), .SEL(n2462), .F(n2339) );
  IV U320 ( .A(n2463), .Z(n100) );
  MUX U321 ( .IN0(n2413), .IN1(n2415), .SEL(n2414), .F(n2293) );
  MUX U322 ( .IN0(n2726), .IN1(n2728), .SEL(n2727), .F(n2594) );
  MUX U323 ( .IN0(n2734), .IN1(n101), .SEL(n2735), .F(n2602) );
  IV U324 ( .A(n2736), .Z(n101) );
  MUX U325 ( .IN0(g_input[16]), .IN1(n4601), .SEL(g_input[31]), .F(n102) );
  IV U326 ( .A(n102), .Z(n1518) );
  MUX U327 ( .IN0(g_input[18]), .IN1(n4567), .SEL(g_input[31]), .F(n103) );
  IV U328 ( .A(n103), .Z(n1330) );
  MUX U329 ( .IN0(g_input[14]), .IN1(n4983), .SEL(g_input[31]), .F(n104) );
  IV U330 ( .A(n104), .Z(n1710) );
  MUX U331 ( .IN0(n2766), .IN1(n2768), .SEL(n2767), .F(n2636) );
  MUX U332 ( .IN0(g_input[13]), .IN1(n4995), .SEL(g_input[31]), .F(n105) );
  IV U333 ( .A(n105), .Z(n1811) );
  MUX U334 ( .IN0(n2911), .IN1(n106), .SEL(n2912), .F(n2774) );
  IV U335 ( .A(n2913), .Z(n106) );
  XNOR U336 ( .A(n3069), .B(n3068), .Z(n3848) );
  MUX U337 ( .IN0(n806), .IN1(n107), .SEL(n807), .F(n747) );
  IV U338 ( .A(n808), .Z(n107) );
  MUX U339 ( .IN0(n1040), .IN1(n1038), .SEL(n1039), .F(n970) );
  MUX U340 ( .IN0(n108), .IN1(n1082), .SEL(n1083), .F(n1008) );
  IV U341 ( .A(n1084), .Z(n108) );
  MUX U342 ( .IN0(n1742), .IN1(n1744), .SEL(n1743), .F(n1641) );
  MUX U343 ( .IN0(n1362), .IN1(n1360), .SEL(n1361), .F(n1271) );
  MUX U344 ( .IN0(n1410), .IN1(n1408), .SEL(n1409), .F(n1315) );
  MUX U345 ( .IN0(n1906), .IN1(n1904), .SEL(n1905), .F(n1798) );
  MUX U346 ( .IN0(n1867), .IN1(n1865), .SEL(n1866), .F(n1757) );
  MUX U347 ( .IN0(n1890), .IN1(n1888), .SEL(n1889), .F(n1782) );
  MUX U348 ( .IN0(n2321), .IN1(n2319), .SEL(n2320), .F(n2199) );
  MUX U349 ( .IN0(n2482), .IN1(n2480), .SEL(n2481), .F(n2358) );
  MUX U350 ( .IN0(n109), .IN1(n2488), .SEL(n2489), .F(n2366) );
  IV U351 ( .A(n2490), .Z(n109) );
  MUX U352 ( .IN0(n699), .IN1(n697), .SEL(n698), .F(n654) );
  MUX U353 ( .IN0(n710), .IN1(n708), .SEL(n709), .F(n664) );
  XNOR U354 ( .A(n863), .B(n862), .Z(n924) );
  MUX U355 ( .IN0(n110), .IN1(n1305), .SEL(n1306), .F(n1221) );
  IV U356 ( .A(n1307), .Z(n110) );
  XNOR U357 ( .A(n1383), .B(n1393), .Z(n1482) );
  MUX U358 ( .IN0(n1836), .IN1(n111), .SEL(n1837), .F(n1725) );
  IV U359 ( .A(n1838), .Z(n111) );
  XOR U360 ( .A(n574), .B(n551), .Z(n548) );
  MUX U361 ( .IN0(n648), .IN1(n650), .SEL(n649), .F(n112) );
  IV U362 ( .A(n112), .Z(n614) );
  AND U363 ( .A(n682), .B(n684), .Z(n642) );
  NOR U364 ( .A(n1349), .B(n1350), .Z(n1348) );
  NANDN U365 ( .B(n520), .A(n532), .Z(n500) );
  MUX U366 ( .IN0(n535), .IN1(\_MxM/Y0[29] ), .SEL(n536), .F(n512) );
  MUX U367 ( .IN0(n4132), .IN1(n4130), .SEL(n4131), .F(n4109) );
  MUX U368 ( .IN0(n5068), .IN1(n4945), .SEL(n4946), .F(n5054) );
  MUX U369 ( .IN0(n5128), .IN1(n5130), .SEL(n5129), .F(n5125) );
  MUX U370 ( .IN0(n113), .IN1(n4725), .SEL(n4726), .F(n4706) );
  IV U371 ( .A(n4727), .Z(n113) );
  MUX U372 ( .IN0(n114), .IN1(n5084), .SEL(n5085), .F(n5075) );
  IV U373 ( .A(n5086), .Z(n114) );
  NANDN U374 ( .B(n4952), .A(n3019), .Z(n135) );
  MUX U375 ( .IN0(n4173), .IN1(n4175), .SEL(n4174), .F(n4155) );
  XNOR U376 ( .A(n4193), .B(n4192), .Z(n4208) );
  MUX U377 ( .IN0(n115), .IN1(n5152), .SEL(n5153), .F(n3005) );
  IV U378 ( .A(n5154), .Z(n115) );
  XNOR U379 ( .A(n4975), .B(n4974), .Z(n4980) );
  XNOR U380 ( .A(n4704), .B(n4703), .Z(n4709) );
  MUX U381 ( .IN0(n1869), .IN1(n1871), .SEL(n1870), .F(n1761) );
  MUX U382 ( .IN0(n1984), .IN1(n1986), .SEL(n1985), .F(n1877) );
  MUX U383 ( .IN0(n2227), .IN1(n2229), .SEL(n2228), .F(n2108) );
  MUX U384 ( .IN0(n2235), .IN1(n116), .SEL(n2236), .F(n2116) );
  IV U385 ( .A(n2237), .Z(n116) );
  MUX U386 ( .IN0(n2179), .IN1(n2181), .SEL(n2180), .F(n2065) );
  MUX U387 ( .IN0(n2316), .IN1(n117), .SEL(n2317), .F(n2196) );
  IV U388 ( .A(n2318), .Z(n117) );
  MUX U389 ( .IN0(n2512), .IN1(n2514), .SEL(n2513), .F(n2388) );
  MUX U390 ( .IN0(n2520), .IN1(n118), .SEL(n2521), .F(n2396) );
  IV U391 ( .A(n2522), .Z(n118) );
  MUX U392 ( .IN0(n2659), .IN1(n2661), .SEL(n2660), .F(n2535) );
  MUX U393 ( .IN0(n2710), .IN1(n2712), .SEL(n2711), .F(n2578) );
  MUX U394 ( .IN0(n2718), .IN1(n119), .SEL(n2719), .F(n2586) );
  IV U395 ( .A(n2720), .Z(n119) );
  MUX U396 ( .IN0(n2834), .IN1(n2836), .SEL(n2835), .F(n2702) );
  MUX U397 ( .IN0(n2827), .IN1(n120), .SEL(n2828), .F(n2695) );
  IV U398 ( .A(n2829), .Z(n120) );
  MUX U399 ( .IN0(n2874), .IN1(n121), .SEL(n2875), .F(n2742) );
  IV U400 ( .A(n2876), .Z(n121) );
  MUX U401 ( .IN0(n2782), .IN1(n122), .SEL(n2783), .F(n2652) );
  IV U402 ( .A(n2784), .Z(n122) );
  MUX U403 ( .IN0(n4785), .IN1(n4783), .SEL(n4784), .F(n2969) );
  MUX U404 ( .IN0(n3054), .IN1(n3052), .SEL(n3053), .F(n2922) );
  XNOR U405 ( .A(n3044), .B(n3043), .Z(n3106) );
  MUX U406 ( .IN0(n714), .IN1(n716), .SEL(n715), .F(n670) );
  MUX U407 ( .IN0(n1317), .IN1(n1315), .SEL(n1316), .F(n1231) );
  MUX U408 ( .IN0(n123), .IN1(n1705), .SEL(n1706), .F(n1609) );
  IV U409 ( .A(n1707), .Z(n123) );
  MUX U410 ( .IN0(n1683), .IN1(n1681), .SEL(n1682), .F(n1585) );
  MUX U411 ( .IN0(n1974), .IN1(n1972), .SEL(n1973), .F(n1865) );
  MUX U412 ( .IN0(n2013), .IN1(n2011), .SEL(n2012), .F(n1904) );
  MUX U413 ( .IN0(n2053), .IN1(n2055), .SEL(n2054), .F(n124) );
  IV U414 ( .A(n124), .Z(n1943) );
  MUX U415 ( .IN0(n2224), .IN1(n2222), .SEL(n2223), .F(n2103) );
  MUX U416 ( .IN0(n2411), .IN1(n2409), .SEL(n2410), .F(n2289) );
  MUX U417 ( .IN0(n125), .IN1(n2613), .SEL(n2614), .F(n2488) );
  IV U418 ( .A(n2615), .Z(n125) );
  MUX U419 ( .IN0(n2607), .IN1(n2605), .SEL(n2606), .F(n2480) );
  MUX U420 ( .IN0(n2568), .IN1(n2566), .SEL(n2567), .F(n2441) );
  MUX U421 ( .IN0(n2550), .IN1(n2548), .SEL(n2549), .F(n126) );
  IV U422 ( .A(n126), .Z(n2420) );
  MUX U423 ( .IN0(n2649), .IN1(n2647), .SEL(n2648), .F(n2523) );
  XNOR U424 ( .A(n2938), .B(n2937), .Z(n3062) );
  MUX U425 ( .IN0(n626), .IN1(n624), .SEL(n625), .F(n580) );
  MUX U426 ( .IN0(n811), .IN1(n809), .SEL(n810), .F(n750) );
  MUX U427 ( .IN0(n982), .IN1(n980), .SEL(n981), .F(n911) );
  MUX U428 ( .IN0(n127), .IN1(n990), .SEL(n991), .F(n921) );
  IV U429 ( .A(n992), .Z(n127) );
  XNOR U430 ( .A(n1111), .B(n1110), .Z(n1182) );
  MUX U431 ( .IN0(n128), .IN1(n1400), .SEL(n1401), .F(n1305) );
  IV U432 ( .A(n1402), .Z(n128) );
  XNOR U433 ( .A(n1728), .B(n1637), .Z(n1638) );
  MUX U434 ( .IN0(n1940), .IN1(n129), .SEL(n1941), .F(n1836) );
  IV U435 ( .A(n1942), .Z(n129) );
  MUX U436 ( .IN0(n2426), .IN1(n2428), .SEL(n2427), .F(n2308) );
  ANDN U437 ( .A(n607), .B(n611), .Z(n610) );
  MUX U438 ( .IN0(n130), .IN1(n841), .SEL(n842), .F(n782) );
  IV U439 ( .A(n843), .Z(n130) );
  ANDN U440 ( .A(n1547), .B(n1549), .Z(n1438) );
  MUX U441 ( .IN0(n178), .IN1(n2188), .SEL(n2187), .F(n2071) );
  NANDN U442 ( .B(n593), .A(n594), .Z(n562) );
  AND U443 ( .A(n642), .B(n644), .Z(n601) );
  NANDN U444 ( .B(n762), .A(n763), .Z(n718) );
  AND U445 ( .A(n960), .B(n962), .Z(n892) );
  MUX U446 ( .IN0(n1453), .IN1(n131), .SEL(n1452), .F(n1351) );
  IV U447 ( .A(n1451), .Z(n131) );
  AND U448 ( .A(n508), .B(n509), .Z(n503) );
  MUX U449 ( .IN0(n564), .IN1(\_MxM/Y0[28] ), .SEL(n565), .F(n535) );
  MUX U450 ( .IN0(n3739), .IN1(n3737), .SEL(n3738), .F(n3695) );
  MUX U451 ( .IN0(n3804), .IN1(n3806), .SEL(n3805), .F(n3801) );
  MUX U452 ( .IN0(n132), .IN1(n5089), .SEL(n5090), .F(n5070) );
  IV U453 ( .A(n5091), .Z(n132) );
  MUX U454 ( .IN0(n133), .IN1(n3762), .SEL(n3763), .F(n3753) );
  IV U455 ( .A(n3764), .Z(n133) );
  MUX U456 ( .IN0(n134), .IN1(n4706), .SEL(n4707), .F(n4694) );
  IV U457 ( .A(n4708), .Z(n134) );
  MUX U458 ( .IN0(n4949), .IN1(n135), .SEL(n4950), .F(n4937) );
  MUX U459 ( .IN0(n136), .IN1(n5075), .SEL(n5076), .F(n5063) );
  IV U460 ( .A(n5077), .Z(n136) );
  XNOR U461 ( .A(n4169), .B(n4168), .Z(n4188) );
  MUX U462 ( .IN0(n1761), .IN1(n1763), .SEL(n1762), .F(n1660) );
  MUX U463 ( .IN0(n1795), .IN1(n137), .SEL(n1796), .F(n1694) );
  IV U464 ( .A(n1797), .Z(n137) );
  MUX U465 ( .IN0(n2243), .IN1(n138), .SEL(n2244), .F(n2124) );
  IV U466 ( .A(n2245), .Z(n138) );
  MUX U467 ( .IN0(n2355), .IN1(n139), .SEL(n2356), .F(n2235) );
  IV U468 ( .A(n2357), .Z(n139) );
  MUX U469 ( .IN0(n2331), .IN1(n2333), .SEL(n2332), .F(n2211) );
  MUX U470 ( .IN0(n2445), .IN1(n2447), .SEL(n2446), .F(n2323) );
  MUX U471 ( .IN0(n2438), .IN1(n140), .SEL(n2439), .F(n2316) );
  IV U472 ( .A(n2440), .Z(n140) );
  MUX U473 ( .IN0(n2594), .IN1(n2596), .SEL(n2595), .F(n2469) );
  MUX U474 ( .IN0(n2528), .IN1(n141), .SEL(n2529), .F(n2406) );
  IV U475 ( .A(n2530), .Z(n141) );
  MUX U476 ( .IN0(n2842), .IN1(n2844), .SEL(n2843), .F(n2710) );
  MUX U477 ( .IN0(n2850), .IN1(n142), .SEL(n2851), .F(n2718) );
  IV U478 ( .A(n2852), .Z(n142) );
  MUX U479 ( .IN0(n3005), .IN1(n143), .SEL(n3006), .F(n2866) );
  IV U480 ( .A(n3007), .Z(n143) );
  MUX U481 ( .IN0(n2966), .IN1(n144), .SEL(n2967), .F(n2827) );
  IV U482 ( .A(n2968), .Z(n144) );
  MUX U483 ( .IN0(n2903), .IN1(n2905), .SEL(n2904), .F(n2766) );
  MUX U484 ( .IN0(n4975), .IN1(n4801), .SEL(n4803), .F(n2992) );
  MUX U485 ( .IN0(n756), .IN1(n758), .SEL(n757), .F(n714) );
  MUX U486 ( .IN0(n1560), .IN1(n1558), .SEL(n1559), .F(n1462) );
  MUX U487 ( .IN0(n1603), .IN1(n1601), .SEL(n1602), .F(n1505) );
  MUX U488 ( .IN0(n145), .IN1(n1609), .SEL(n1610), .F(n1513) );
  IV U489 ( .A(n1611), .Z(n145) );
  MUX U490 ( .IN0(n1997), .IN1(n1995), .SEL(n1996), .F(n1888) );
  MUX U491 ( .IN0(n146), .IN1(n2019), .SEL(n2020), .F(n1912) );
  IV U492 ( .A(n2021), .Z(n146) );
  MUX U493 ( .IN0(n2121), .IN1(n2119), .SEL(n2120), .F(n2011) );
  MUX U494 ( .IN0(n2082), .IN1(n2080), .SEL(n2081), .F(n1972) );
  MUX U495 ( .IN0(n2177), .IN1(n2175), .SEL(n2176), .F(n2061) );
  MUX U496 ( .IN0(n2591), .IN1(n2589), .SEL(n2590), .F(n2464) );
  MUX U497 ( .IN0(n2525), .IN1(n2523), .SEL(n2524), .F(n2401) );
  MUX U498 ( .IN0(n2739), .IN1(n2737), .SEL(n2738), .F(n2605) );
  MUX U499 ( .IN0(n147), .IN1(n2745), .SEL(n2746), .F(n2613) );
  IV U500 ( .A(n2747), .Z(n147) );
  MUX U501 ( .IN0(n2700), .IN1(n2698), .SEL(n2699), .F(n2566) );
  MUX U502 ( .IN0(n2787), .IN1(n2785), .SEL(n2786), .F(n2655) );
  XNOR U503 ( .A(n2914), .B(n2913), .Z(n3037) );
  MUX U504 ( .IN0(n744), .IN1(n742), .SEL(n743), .F(n697) );
  XNOR U505 ( .A(n809), .B(n808), .Z(n866) );
  MUX U506 ( .IN0(n1050), .IN1(n1052), .SEL(n1051), .F(n980) );
  XNOR U507 ( .A(n1000), .B(n999), .Z(n1065) );
  XNOR U508 ( .A(n1160), .B(n1159), .Z(n1234) );
  XNOR U509 ( .A(n1189), .B(n1188), .Z(n1264) );
  MUX U510 ( .IN0(n1641), .IN1(n1643), .SEL(n1642), .F(n1540) );
  MUX U511 ( .IN0(n148), .IN1(n1379), .SEL(n1380), .F(n1288) );
  IV U512 ( .A(n1381), .Z(n148) );
  XNOR U513 ( .A(n1729), .B(n1739), .Z(n1839) );
  XOR U514 ( .A(n2157), .B(n2053), .Z(n2054) );
  MUX U515 ( .IN0(n149), .IN1(n2350), .SEL(n2351), .F(n2230) );
  IV U516 ( .A(n2352), .Z(n149) );
  MUX U517 ( .IN0(n2422), .IN1(n150), .SEL(n2421), .F(n2306) );
  IV U518 ( .A(n2420), .Z(n150) );
  MUX U519 ( .IN0(n617), .IN1(n151), .SEL(n616), .F(n589) );
  IV U520 ( .A(n615), .Z(n151) );
  XNOR U521 ( .A(n780), .B(n779), .Z(n833) );
  AND U522 ( .A(n1170), .B(n1172), .Z(n1092) );
  MUX U523 ( .IN0(n152), .IN1(n1278), .SEL(n1279), .F(n1198) );
  IV U524 ( .A(n1280), .Z(n152) );
  MUX U525 ( .IN0(n2432), .IN1(n2434), .SEL(n2433), .F(n2310) );
  NANDN U526 ( .B(n634), .A(n635), .Z(n593) );
  ANDN U527 ( .A(n673), .B(n644), .Z(n633) );
  NANDN U528 ( .B(n821), .A(n822), .Z(n762) );
  NAND U529 ( .A(n1438), .B(n1437), .Z(n1349) );
  MUX U530 ( .IN0(n153), .IN1(n1961), .SEL(n1962), .F(n1853) );
  IV U531 ( .A(n1963), .Z(n153) );
  ANDN U532 ( .A(n1101), .B(n1102), .Z(n1027) );
  MUX U533 ( .IN0(\_MxM/Y0[3] ), .IN1(n2623), .SEL(n2624), .F(n2500) );
  MUX U534 ( .IN0(n500), .IN1(n502), .SEL(n501), .F(n154) );
  IV U535 ( .A(n154), .Z(n499) );
  MUX U536 ( .IN0(n595), .IN1(\_MxM/Y0[27] ), .SEL(n596), .F(n564) );
  MUX U537 ( .IN0(n764), .IN1(\_MxM/Y0[23] ), .SEL(n765), .F(n720) );
  MUX U538 ( .IN0(n1021), .IN1(\_MxM/Y0[19] ), .SEL(n1022), .F(n954) );
  MUX U539 ( .IN0(n1338), .IN1(\_MxM/Y0[15] ), .SEL(n1339), .F(n1254) );
  MUX U540 ( .IN0(n1718), .IN1(\_MxM/Y0[11] ), .SEL(n1719), .F(n1622) );
  MUX U541 ( .IN0(n2140), .IN1(\_MxM/Y0[7] ), .SEL(n2141), .F(n2032) );
  MUX U542 ( .IN0(n4608), .IN1(n4162), .SEL(n4163), .F(n4591) );
  MUX U543 ( .IN0(n155), .IN1(n4139), .SEL(n3704), .F(n4118) );
  IV U544 ( .A(n3702), .Z(n155) );
  MUX U545 ( .IN0(n3578), .IN1(n3576), .SEL(n3577), .F(n3532) );
  MUX U546 ( .IN0(n4299), .IN1(n4297), .SEL(n4298), .F(n4273) );
  XNOR U547 ( .A(n4874), .B(n4873), .Z(n4889) );
  MUX U548 ( .IN0(n4331), .IN1(n4333), .SEL(n4332), .F(n4328) );
  MUX U549 ( .IN0(n156), .IN1(n3767), .SEL(n3768), .F(n3746) );
  IV U550 ( .A(n3769), .Z(n156) );
  NANDN U551 ( .B(n1634), .A(n3019), .Z(n188) );
  MUX U552 ( .IN0(n157), .IN1(n5143), .SEL(n5144), .F(n2997) );
  IV U553 ( .A(n5145), .Z(n157) );
  MUX U554 ( .IN0(n4794), .IN1(n4796), .SEL(n4795), .F(n2981) );
  MUX U555 ( .IN0(n3857), .IN1(n3855), .SEL(n3856), .F(n3069) );
  MUX U556 ( .IN0(n1877), .IN1(n1879), .SEL(n1878), .F(n1769) );
  MUX U557 ( .IN0(n2000), .IN1(n2002), .SEL(n2001), .F(n1893) );
  MUX U558 ( .IN0(n2084), .IN1(n2086), .SEL(n2085), .F(n1976) );
  MUX U559 ( .IN0(n2077), .IN1(n158), .SEL(n2078), .F(n1969) );
  IV U560 ( .A(n2079), .Z(n158) );
  MUX U561 ( .IN0(n2339), .IN1(n159), .SEL(n2340), .F(n2219) );
  IV U562 ( .A(n2341), .Z(n159) );
  MUX U563 ( .IN0(n2453), .IN1(n2455), .SEL(n2454), .F(n2331) );
  MUX U564 ( .IN0(n2469), .IN1(n2471), .SEL(n2470), .F(n2347) );
  MUX U565 ( .IN0(n2602), .IN1(n160), .SEL(n2603), .F(n2477) );
  IV U566 ( .A(n2604), .Z(n160) );
  MUX U567 ( .IN0(n2563), .IN1(n161), .SEL(n2564), .F(n2438) );
  IV U568 ( .A(n2565), .Z(n161) );
  MUX U569 ( .IN0(n2652), .IN1(n162), .SEL(n2653), .F(n2528) );
  IV U570 ( .A(n2654), .Z(n162) );
  MUX U571 ( .IN0(n2742), .IN1(n163), .SEL(n2743), .F(n2610) );
  IV U572 ( .A(n2744), .Z(n163) );
  MUX U573 ( .IN0(n2702), .IN1(n2704), .SEL(n2703), .F(n2570) );
  MUX U574 ( .IN0(g_input[8]), .IN1(n5062), .SEL(g_input[31]), .F(n164) );
  IV U575 ( .A(n164), .Z(n2371) );
  MUX U576 ( .IN0(n2989), .IN1(n165), .SEL(n2990), .F(n2850) );
  IV U577 ( .A(n2991), .Z(n165) );
  MUX U578 ( .IN0(n2942), .IN1(n2944), .SEL(n2943), .F(n2805) );
  MUX U579 ( .IN0(n865), .IN1(n863), .SEL(n864), .F(n801) );
  MUX U580 ( .IN0(n1759), .IN1(n1757), .SEL(n1758), .F(n1656) );
  MUX U581 ( .IN0(n1800), .IN1(n1798), .SEL(n1799), .F(n1697) );
  MUX U582 ( .IN0(n1731), .IN1(n1729), .SEL(n1730), .F(n1637) );
  MUX U583 ( .IN0(n166), .IN1(n1912), .SEL(n1913), .F(n1806) );
  IV U584 ( .A(n1914), .Z(n166) );
  MUX U585 ( .IN0(n2105), .IN1(n2103), .SEL(n2104), .F(n1995) );
  MUX U586 ( .IN0(n2201), .IN1(n2199), .SEL(n2200), .F(n2080) );
  MUX U587 ( .IN0(n2240), .IN1(n2238), .SEL(n2239), .F(n2119) );
  MUX U588 ( .IN0(n2160), .IN1(n2158), .SEL(n2159), .F(n2053) );
  MUX U589 ( .IN0(n2291), .IN1(n2289), .SEL(n2290), .F(n2175) );
  MUX U590 ( .IN0(n167), .IN1(n2366), .SEL(n2367), .F(n2246) );
  IV U591 ( .A(n2368), .Z(n167) );
  MUX U592 ( .IN0(n2669), .IN1(n2667), .SEL(n2668), .F(n2548) );
  MUX U593 ( .IN0(n2723), .IN1(n2721), .SEL(n2722), .F(n2589) );
  MUX U594 ( .IN0(n2832), .IN1(n2830), .SEL(n2831), .F(n2698) );
  MUX U595 ( .IN0(n2871), .IN1(n2869), .SEL(n2870), .F(n2737) );
  MUX U596 ( .IN0(n168), .IN1(n2877), .SEL(n2878), .F(n2745) );
  IV U597 ( .A(n2879), .Z(n168) );
  MUX U598 ( .IN0(n2779), .IN1(n2777), .SEL(n2778), .F(n2647) );
  MUX U599 ( .IN0(n2924), .IN1(n2922), .SEL(n2923), .F(n2785) );
  MUX U600 ( .IN0(n630), .IN1(n632), .SEL(n631), .F(n586) );
  MUX U601 ( .IN0(n752), .IN1(n750), .SEL(n751), .F(n708) );
  XNOR U602 ( .A(n941), .B(n940), .Z(n1003) );
  XNOR U603 ( .A(n1152), .B(n1151), .Z(n1224) );
  XNOR U604 ( .A(n1241), .B(n1240), .Z(n1318) );
  XNOR U605 ( .A(n1271), .B(n1270), .Z(n1355) );
  MUX U606 ( .IN0(n169), .IN1(n1497), .SEL(n1498), .F(n1400) );
  IV U607 ( .A(n1499), .Z(n169) );
  XNOR U608 ( .A(n1489), .B(n1488), .Z(n1578) );
  MUX U609 ( .IN0(n2044), .IN1(n170), .SEL(n2045), .F(n1940) );
  IV U610 ( .A(n2046), .Z(n170) );
  MUX U611 ( .IN0(n171), .IN1(n2111), .SEL(n2112), .F(n2003) );
  IV U612 ( .A(n2113), .Z(n171) );
  MUX U613 ( .IN0(n172), .IN1(n2334), .SEL(n2335), .F(n2214) );
  IV U614 ( .A(n2336), .Z(n172) );
  MUX U615 ( .IN0(n173), .IN1(n2597), .SEL(n2598), .F(n2472) );
  IV U616 ( .A(n2599), .Z(n173) );
  MUX U617 ( .IN0(n174), .IN1(n2515), .SEL(n2516), .F(n2391) );
  IV U618 ( .A(n2517), .Z(n174) );
  MUX U619 ( .IN0(n175), .IN1(n577), .SEL(n576), .F(n551) );
  IV U620 ( .A(n575), .Z(n175) );
  AND U621 ( .A(n613), .B(n614), .Z(n609) );
  MUX U622 ( .IN0(n900), .IN1(n898), .SEL(n899), .F(n838) );
  MUX U623 ( .IN0(n176), .IN1(n1045), .SEL(n1046), .F(n977) );
  IV U624 ( .A(n1047), .Z(n176) );
  AND U625 ( .A(n1251), .B(n1253), .Z(n1170) );
  MUX U626 ( .IN0(n1540), .IN1(n1542), .SEL(n1541), .F(n1449) );
  MUX U627 ( .IN0(n177), .IN1(n1764), .SEL(n1765), .F(n1663) );
  IV U628 ( .A(n1766), .Z(n177) );
  ANDN U629 ( .A(n1748), .B(n1750), .Z(n1647) );
  AND U630 ( .A(n2029), .B(n2031), .Z(n1922) );
  MUX U631 ( .IN0(n2312), .IN1(n2310), .SEL(n2311), .F(n178) );
  IV U632 ( .A(n178), .Z(n2186) );
  NANDN U633 ( .B(n674), .A(n675), .Z(n634) );
  MUX U634 ( .IN0(n761), .IN1(n179), .SEL(n760), .F(n717) );
  IV U635 ( .A(n759), .Z(n179) );
  AND U636 ( .A(n829), .B(n831), .Z(n818) );
  NANDN U637 ( .B(n884), .A(n885), .Z(n821) );
  MUX U638 ( .IN0(n180), .IN1(n1544), .SEL(n1545), .F(n1451) );
  IV U639 ( .A(n1546), .Z(n180) );
  MUX U640 ( .IN0(n181), .IN1(n2068), .SEL(n2069), .F(n1961) );
  IV U641 ( .A(n2070), .Z(n181) );
  MUX U642 ( .IN0(n2540), .IN1(n208), .SEL(n2539), .F(n182) );
  IV U643 ( .A(n182), .Z(n2416) );
  AND U644 ( .A(n541), .B(n543), .Z(n518) );
  ANDN U645 ( .A(n1179), .B(n1180), .Z(n1101) );
  NAND U646 ( .A(n489), .B(n491), .Z(n488) );
  MUX U647 ( .IN0(n636), .IN1(\_MxM/Y0[26] ), .SEL(n637), .F(n595) );
  MUX U648 ( .IN0(n823), .IN1(\_MxM/Y0[22] ), .SEL(n824), .F(n764) );
  MUX U649 ( .IN0(n1095), .IN1(\_MxM/Y0[18] ), .SEL(n1096), .F(n1021) );
  MUX U650 ( .IN0(n1429), .IN1(\_MxM/Y0[14] ), .SEL(n1430), .F(n1338) );
  MUX U651 ( .IN0(n1819), .IN1(\_MxM/Y0[10] ), .SEL(n1820), .F(n1718) );
  MUX U652 ( .IN0(n2259), .IN1(\_MxM/Y0[6] ), .SEL(n2260), .F(n2140) );
  MUX U653 ( .IN0(n4153), .IN1(n4151), .SEL(n4152), .F(n4130) );
  MUX U654 ( .IN0(n3728), .IN1(n3726), .SEL(n3727), .F(n183) );
  IV U655 ( .A(n183), .Z(n3684) );
  MUX U656 ( .IN0(n3651), .IN1(n3649), .SEL(n3650), .F(n3603) );
  MUX U657 ( .IN0(n4574), .IN1(n4120), .SEL(n4121), .F(n4557) );
  MUX U658 ( .IN0(n184), .IN1(n4055), .SEL(n3522), .F(n4034) );
  IV U659 ( .A(n3520), .Z(n184) );
  MUX U660 ( .IN0(n4704), .IN1(n4324), .SEL(n4325), .F(n4692) );
  MUX U661 ( .IN0(n4942), .IN1(n4940), .SEL(n4941), .F(n4920) );
  XNOR U662 ( .A(n4273), .B(n4272), .Z(n4290) );
  MUX U663 ( .IN0(n185), .IN1(n3971), .SEL(n3340), .F(n3950) );
  IV U664 ( .A(n3338), .Z(n185) );
  MUX U665 ( .IN0(n4650), .IN1(n4240), .SEL(n4242), .F(n4638) );
  MUX U666 ( .IN0(n5212), .IN1(n5214), .SEL(n5213), .F(n5208) );
  MUX U667 ( .IN0(n4856), .IN1(n4854), .SEL(n4855), .F(n4834) );
  MUX U668 ( .IN0(n186), .IN1(n5168), .SEL(n5169), .F(n5143) );
  IV U669 ( .A(n5170), .Z(n186) );
  MUX U670 ( .IN0(n187), .IN1(n5070), .SEL(n5071), .F(n5056) );
  IV U671 ( .A(n5072), .Z(n187) );
  MUX U672 ( .IN0(n3822), .IN1(n188), .SEL(n3823), .F(n3708) );
  MUX U673 ( .IN0(n189), .IN1(n3888), .SEL(n3167), .F(n3867) );
  IV U674 ( .A(n3165), .Z(n189) );
  MUX U675 ( .IN0(n1893), .IN1(n1895), .SEL(n1894), .F(n1787) );
  MUX U676 ( .IN0(n2866), .IN1(n190), .SEL(n2867), .F(n2734) );
  IV U677 ( .A(n2868), .Z(n190) );
  MUX U678 ( .IN0(g_input[7]), .IN1(n5151), .SEL(g_input[31]), .F(n191) );
  IV U679 ( .A(n191), .Z(n2493) );
  MUX U680 ( .IN0(g_input[11]), .IN1(n5019), .SEL(g_input[31]), .F(n192) );
  IV U681 ( .A(n192), .Z(n2024) );
  MUX U682 ( .IN0(n2926), .IN1(n2928), .SEL(n2927), .F(n2789) );
  MUX U683 ( .IN0(n2919), .IN1(n193), .SEL(n2920), .F(n2782) );
  IV U684 ( .A(n2921), .Z(n193) );
  MUX U685 ( .IN0(n3046), .IN1(n3044), .SEL(n3045), .F(n2914) );
  MUX U686 ( .IN0(n815), .IN1(n817), .SEL(n816), .F(n756) );
  MUX U687 ( .IN0(n1233), .IN1(n1231), .SEL(n1232), .F(n1152) );
  MUX U688 ( .IN0(n1385), .IN1(n1383), .SEL(n1384), .F(n1297) );
  MUX U689 ( .IN0(n1784), .IN1(n1782), .SEL(n1783), .F(n1681) );
  MUX U690 ( .IN0(n2344), .IN1(n2342), .SEL(n2343), .F(n2222) );
  MUX U691 ( .IN0(n2443), .IN1(n2441), .SEL(n2442), .F(n2319) );
  MUX U692 ( .IN0(n2657), .IN1(n2655), .SEL(n2656), .F(n2531) );
  MUX U693 ( .IN0(n2855), .IN1(n2853), .SEL(n2854), .F(n2721) );
  MUX U694 ( .IN0(n194), .IN1(n3016), .SEL(n3017), .F(n2877) );
  IV U695 ( .A(n3018), .Z(n194) );
  MUX U696 ( .IN0(n3010), .IN1(n3008), .SEL(n3009), .F(n2869) );
  MUX U697 ( .IN0(n2971), .IN1(n2969), .SEL(n2970), .F(n2830) );
  XNOR U698 ( .A(n873), .B(n872), .Z(n934) );
  XNOR U699 ( .A(n931), .B(n930), .Z(n993) );
  XNOR U700 ( .A(n1082), .B(n1081), .Z(n1155) );
  MUX U701 ( .IN0(n1211), .IN1(n195), .SEL(n1212), .F(n1132) );
  IV U702 ( .A(n1213), .Z(n195) );
  XNOR U703 ( .A(n1325), .B(n1324), .Z(n1411) );
  XNOR U704 ( .A(n1360), .B(n1359), .Z(n1455) );
  XNOR U705 ( .A(n1505), .B(n1504), .Z(n1596) );
  MUX U706 ( .IN0(n196), .IN1(n1689), .SEL(n1690), .F(n1593) );
  IV U707 ( .A(n1691), .Z(n196) );
  XNOR U708 ( .A(n1609), .B(n1608), .Z(n1700) );
  XNOR U709 ( .A(n1656), .B(n1655), .Z(n1752) );
  MUX U710 ( .IN0(n197), .IN1(n1880), .SEL(n1881), .F(n1772) );
  IV U711 ( .A(n1882), .Z(n197) );
  XNOR U712 ( .A(n1904), .B(n1903), .Z(n2006) );
  XNOR U713 ( .A(n1912), .B(n1911), .Z(n2014) );
  XNOR U714 ( .A(n2061), .B(n2060), .Z(n2170) );
  XNOR U715 ( .A(n2238), .B(n2237), .Z(n2353) );
  XNOR U716 ( .A(n2246), .B(n2245), .Z(n2361) );
  XNOR U717 ( .A(n2281), .B(n2280), .Z(n2394) );
  MUX U718 ( .IN0(n198), .IN1(n2581), .SEL(n2582), .F(n2456) );
  IV U719 ( .A(n2583), .Z(n198) );
  XNOR U720 ( .A(n2667), .B(n2677), .Z(n2796) );
  MUX U721 ( .IN0(n199), .IN1(n2769), .SEL(n2770), .F(n2639) );
  IV U722 ( .A(n2771), .Z(n199) );
  XNOR U723 ( .A(n580), .B(n577), .Z(n618) );
  MUX U724 ( .IN0(n656), .IN1(n654), .SEL(n655), .F(n607) );
  MUX U725 ( .IN0(n200), .IN1(n692), .SEL(n693), .F(n651) );
  IV U726 ( .A(n694), .Z(n200) );
  AND U727 ( .A(n911), .B(n913), .Z(n844) );
  MUX U728 ( .IN0(n201), .IN1(n1120), .SEL(n1121), .F(n1045) );
  IV U729 ( .A(n1122), .Z(n201) );
  MUX U730 ( .IN0(n1536), .IN1(n348), .SEL(n1535), .F(n1448) );
  AND U731 ( .A(n1619), .B(n1621), .Z(n1523) );
  ANDN U732 ( .A(n1856), .B(n1858), .Z(n1748) );
  MUX U733 ( .IN0(n202), .IN1(n1979), .SEL(n1980), .F(n1872) );
  IV U734 ( .A(n1981), .Z(n202) );
  AND U735 ( .A(n2256), .B(n2258), .Z(n2137) );
  MUX U736 ( .IN0(n203), .IN1(n2448), .SEL(n2449), .F(n2326) );
  IV U737 ( .A(n2450), .Z(n203) );
  MUX U738 ( .IN0(n204), .IN1(n2559), .SEL(n2558), .F(n2432) );
  IV U739 ( .A(n2557), .Z(n204) );
  NANDN U740 ( .B(n562), .A(n563), .Z(n533) );
  ANDN U741 ( .A(n717), .B(n684), .Z(n673) );
  NANDN U742 ( .B(n718), .A(n719), .Z(n674) );
  MUX U743 ( .IN0(n840), .IN1(n838), .SEL(n839), .F(n205) );
  IV U744 ( .A(n205), .Z(n778) );
  OR U745 ( .A(n1019), .B(n1020), .Z(n952) );
  MUX U746 ( .IN0(n206), .IN1(n1644), .SEL(n1645), .F(n1544) );
  IV U747 ( .A(n1646), .Z(n206) );
  MUX U748 ( .IN0(n207), .IN1(n2182), .SEL(n2183), .F(n2068) );
  IV U749 ( .A(n2184), .Z(n207) );
  MUX U750 ( .IN0(n2664), .IN1(n241), .SEL(n2663), .F(n208) );
  IV U751 ( .A(n208), .Z(n2538) );
  AND U752 ( .A(n818), .B(n820), .Z(n726) );
  MUX U753 ( .IN0(n209), .IN1(n1260), .SEL(n1261), .F(n1179) );
  IV U754 ( .A(n1262), .Z(n209) );
  ANDN U755 ( .A(n493), .B(n494), .Z(n485) );
  MUX U756 ( .IN0(n676), .IN1(\_MxM/Y0[25] ), .SEL(n677), .F(n636) );
  MUX U757 ( .IN0(n886), .IN1(\_MxM/Y0[21] ), .SEL(n887), .F(n823) );
  MUX U758 ( .IN0(n1173), .IN1(\_MxM/Y0[17] ), .SEL(n1174), .F(n1095) );
  MUX U759 ( .IN0(n1526), .IN1(\_MxM/Y0[13] ), .SEL(n1527), .F(n1429) );
  MUX U760 ( .IN0(n1925), .IN1(\_MxM/Y0[9] ), .SEL(n1926), .F(n1819) );
  MUX U761 ( .IN0(n2379), .IN1(\_MxM/Y0[5] ), .SEL(n2380), .F(n2259) );
  MUX U762 ( .IN0(n512), .IN1(\_MxM/Y0[30] ), .SEL(n513), .F(n478) );
  MUX U763 ( .IN0(n3059), .IN1(n3740), .SEL(n3060), .F(n210) );
  IV U764 ( .A(n210), .Z(n3698) );
  MUX U765 ( .IN0(n211), .IN1(n3684), .SEL(n3685), .F(n3638) );
  IV U766 ( .A(n3686), .Z(n211) );
  MUX U767 ( .IN0(n4090), .IN1(n4088), .SEL(n4089), .F(n4067) );
  MUX U768 ( .IN0(n3605), .IN1(n3603), .SEL(n3604), .F(n3557) );
  MUX U769 ( .IN0(n212), .IN1(n3502), .SEL(n3503), .F(n3456) );
  IV U770 ( .A(n3504), .Z(n212) );
  MUX U771 ( .IN0(n4506), .IN1(n4036), .SEL(n4037), .F(n4489) );
  MUX U772 ( .IN0(n3396), .IN1(n3394), .SEL(n3395), .F(n3350) );
  MUX U773 ( .IN0(n4006), .IN1(n4004), .SEL(n4005), .F(n3983) );
  MUX U774 ( .IN0(n3423), .IN1(n3421), .SEL(n3422), .F(n3375) );
  MUX U775 ( .IN0(n4790), .IN1(n4943), .SEL(n4791), .F(n213) );
  IV U776 ( .A(n213), .Z(n4923) );
  MUX U777 ( .IN0(n214), .IN1(n3320), .SEL(n3321), .F(n3275) );
  IV U778 ( .A(n3322), .Z(n214) );
  MUX U779 ( .IN0(n4438), .IN1(n3952), .SEL(n3953), .F(n4422) );
  MUX U780 ( .IN0(n5023), .IN1(n4881), .SEL(n4883), .F(n5011) );
  MUX U781 ( .IN0(n3220), .IN1(n3218), .SEL(n3219), .F(n3176) );
  MUX U782 ( .IN0(n4761), .IN1(n215), .SEL(n4762), .F(n4750) );
  IV U783 ( .A(n4764), .Z(n215) );
  MUX U784 ( .IN0(n3922), .IN1(n3920), .SEL(n3921), .F(n3900) );
  MUX U785 ( .IN0(n3245), .IN1(n3243), .SEL(n3244), .F(n3200) );
  MUX U786 ( .IN0(n4953), .IN1(n4955), .SEL(n4954), .F(n4949) );
  MUX U787 ( .IN0(n4215), .IN1(n4213), .SEL(n4214), .F(n4193) );
  NANDN U788 ( .B(n5232), .A(n3019), .Z(n250) );
  MUX U789 ( .IN0(n216), .IN1(n3147), .SEL(n3148), .F(n3103) );
  IV U790 ( .A(n3149), .Z(n216) );
  MUX U791 ( .IN0(n2323), .IN1(n2325), .SEL(n2324), .F(n2203) );
  MUX U792 ( .IN0(n2695), .IN1(n217), .SEL(n2696), .F(n2563) );
  IV U793 ( .A(n2697), .Z(n217) );
  MUX U794 ( .IN0(g_input[10]), .IN1(n5033), .SEL(g_input[31]), .F(n218) );
  IV U795 ( .A(n218), .Z(n2132) );
  MUX U796 ( .IN0(g_input[6]), .IN1(n5162), .SEL(g_input[31]), .F(n219) );
  IV U797 ( .A(n219), .Z(n2618) );
  MUX U798 ( .IN0(g_input[5]), .IN1(n5178), .SEL(g_input[31]), .F(n220) );
  IV U799 ( .A(n220), .Z(n2750) );
  MUX U800 ( .IN0(n4372), .IN1(n3869), .SEL(n3870), .F(n4352) );
  XNOR U801 ( .A(n4608), .B(n4606), .Z(n4613) );
  MUX U802 ( .IN0(n3071), .IN1(n3069), .SEL(n3070), .F(n2938) );
  MUX U803 ( .IN0(n747), .IN1(n221), .SEL(n748), .F(n705) );
  IV U804 ( .A(n749), .Z(n221) );
  MUX U805 ( .IN0(n290), .IN1(n1215), .SEL(n1214), .F(n1126) );
  MUX U806 ( .IN0(n1587), .IN1(n1585), .SEL(n1586), .F(n1489) );
  MUX U807 ( .IN0(n222), .IN1(n1806), .SEL(n1807), .F(n1705) );
  IV U808 ( .A(n1808), .Z(n222) );
  MUX U809 ( .IN0(n2466), .IN1(n2464), .SEL(n2465), .F(n2342) );
  MUX U810 ( .IN0(n2403), .IN1(n2401), .SEL(n2402), .F(n2281) );
  MUX U811 ( .IN0(n2533), .IN1(n2531), .SEL(n2532), .F(n2409) );
  MUX U812 ( .IN0(n2994), .IN1(n2992), .SEL(n2993), .F(n2853) );
  MUX U813 ( .IN0(n2916), .IN1(n2914), .SEL(n2915), .F(n2777) );
  XNOR U814 ( .A(n3008), .B(n3007), .Z(n5148) );
  XNOR U815 ( .A(n2969), .B(n2968), .Z(n4778) );
  XNOR U816 ( .A(n2922), .B(n2921), .Z(n3047) );
  MUX U817 ( .IN0(n972), .IN1(n970), .SEL(n971), .F(n898) );
  MUX U818 ( .IN0(n803), .IN1(n801), .SEL(n802), .F(n742) );
  XNOR U819 ( .A(n1008), .B(n1007), .Z(n1075) );
  MUX U820 ( .IN0(n1134), .IN1(n223), .SEL(n1133), .F(n1050) );
  IV U821 ( .A(n1132), .Z(n223) );
  XNOR U822 ( .A(n1072), .B(n1071), .Z(n1145) );
  XNOR U823 ( .A(n1408), .B(n1407), .Z(n1500) );
  XNOR U824 ( .A(n1416), .B(n1415), .Z(n1508) );
  XNOR U825 ( .A(n1462), .B(n1461), .Z(n1551) );
  MUX U826 ( .IN0(n224), .IN1(n1671), .SEL(n1672), .F(n1575) );
  IV U827 ( .A(n1673), .Z(n224) );
  XNOR U828 ( .A(n1697), .B(n1696), .Z(n1793) );
  MUX U829 ( .IN0(n225), .IN1(n1896), .SEL(n1897), .F(n1790) );
  IV U830 ( .A(n1898), .Z(n225) );
  XNOR U831 ( .A(n1865), .B(n1864), .Z(n1967) );
  XNOR U832 ( .A(n1954), .B(n1953), .Z(n2056) );
  XNOR U833 ( .A(n1995), .B(n1994), .Z(n2098) );
  MUX U834 ( .IN0(n226), .IN1(n2214), .SEL(n2215), .F(n2095) );
  IV U835 ( .A(n2216), .Z(n226) );
  MUX U836 ( .IN0(n227), .IN1(n2271), .SEL(n2272), .F(n2154) );
  IV U837 ( .A(n2273), .Z(n227) );
  XNOR U838 ( .A(n2319), .B(n2318), .Z(n2436) );
  XNOR U839 ( .A(n2358), .B(n2357), .Z(n2475) );
  XNOR U840 ( .A(n2366), .B(n2365), .Z(n2483) );
  XNOR U841 ( .A(n2666), .B(n2548), .Z(n2549) );
  MUX U842 ( .IN0(n228), .IN1(n2845), .SEL(n2846), .F(n2713) );
  IV U843 ( .A(n2847), .Z(n228) );
  MUX U844 ( .IN0(n2863), .IN1(n298), .SEL(n2862), .F(n229) );
  IV U845 ( .A(n229), .Z(n2729) );
  MUX U846 ( .IN0(n230), .IN1(n2821), .SEL(n2822), .F(n2688) );
  IV U847 ( .A(n2823), .Z(n230) );
  MUX U848 ( .IN0(n586), .IN1(n588), .SEL(n587), .F(n556) );
  XNOR U849 ( .A(n624), .B(n623), .Z(n657) );
  MUX U850 ( .IN0(n231), .IN1(n734), .SEL(n735), .F(n692) );
  IV U851 ( .A(n736), .Z(n231) );
  MUX U852 ( .IN0(n232), .IN1(n908), .SEL(n909), .F(n841) );
  IV U853 ( .A(n910), .Z(n232) );
  MUX U854 ( .IN0(n233), .IN1(n1198), .SEL(n1199), .F(n1120) );
  IV U855 ( .A(n1200), .Z(n233) );
  AND U856 ( .A(n1426), .B(n1428), .Z(n1335) );
  MUX U857 ( .IN0(n234), .IN1(n1565), .SEL(n1566), .F(n1469) );
  IV U858 ( .A(n1567), .Z(n234) );
  XNOR U859 ( .A(n1447), .B(n1448), .Z(n1444) );
  AND U860 ( .A(n1647), .B(n1649), .Z(n1547) );
  AND U861 ( .A(n1816), .B(n1818), .Z(n1715) );
  MUX U862 ( .IN0(n235), .IN1(n2087), .SEL(n2088), .F(n1979) );
  IV U863 ( .A(n2089), .Z(n235) );
  AND U864 ( .A(n2376), .B(n2378), .Z(n2256) );
  MUX U865 ( .IN0(n236), .IN1(n2573), .SEL(n2574), .F(n2448) );
  IV U866 ( .A(n2575), .Z(n236) );
  MUX U867 ( .IN0(n237), .IN1(n2685), .SEL(n2686), .F(n2557) );
  IV U868 ( .A(n2687), .Z(n237) );
  NAND U869 ( .A(n551), .B(n550), .Z(n545) );
  XNOR U870 ( .A(n589), .B(n614), .Z(n605) );
  ANDN U871 ( .A(n726), .B(n727), .Z(n682) );
  AND U872 ( .A(n774), .B(n775), .Z(n773) );
  ANDN U873 ( .A(n1027), .B(n1028), .Z(n960) );
  NAND U874 ( .A(n1092), .B(n1094), .Z(n1019) );
  MUX U875 ( .IN0(n238), .IN1(n1853), .SEL(n1854), .F(n1745) );
  IV U876 ( .A(n1855), .Z(n238) );
  MUX U877 ( .IN0(n239), .IN1(n2071), .SEL(n2072), .F(n1964) );
  IV U878 ( .A(n2073), .Z(n239) );
  MUX U879 ( .IN0(n240), .IN1(n2296), .SEL(n2297), .F(n2182) );
  IV U880 ( .A(n2298), .Z(n240) );
  MUX U881 ( .IN0(n2794), .IN1(n272), .SEL(n2793), .F(n241) );
  IV U882 ( .A(n241), .Z(n2662) );
  XNOR U883 ( .A(n562), .B(n567), .Z(n563) );
  XNOR U884 ( .A(n674), .B(n679), .Z(n675) );
  XNOR U885 ( .A(n821), .B(n826), .Z(n822) );
  XOR U886 ( .A(n1260), .B(n1349), .Z(n1344) );
  XNOR U887 ( .A(n2931), .B(n2930), .Z(n2762) );
  MUX U888 ( .IN0(n720), .IN1(\_MxM/Y0[24] ), .SEL(n721), .F(n676) );
  MUX U889 ( .IN0(n954), .IN1(\_MxM/Y0[20] ), .SEL(n955), .F(n886) );
  MUX U890 ( .IN0(n1254), .IN1(\_MxM/Y0[16] ), .SEL(n1255), .F(n1173) );
  MUX U891 ( .IN0(n1622), .IN1(\_MxM/Y0[12] ), .SEL(n1623), .F(n1526) );
  MUX U892 ( .IN0(n2032), .IN1(\_MxM/Y0[8] ), .SEL(n2033), .F(n1925) );
  MUX U893 ( .IN0(\_MxM/Y0[4] ), .IN1(n2500), .SEL(n2501), .F(n2379) );
  XNOR U894 ( .A(n512), .B(n516), .Z(n514) );
  MUX U895 ( .IN0(n3670), .IN1(n3668), .SEL(n3669), .F(n3622) );
  MUX U896 ( .IN0(n4591), .IN1(n4141), .SEL(n4142), .F(n4574) );
  MUX U897 ( .IN0(n242), .IN1(n4118), .SEL(n3658), .F(n4097) );
  IV U898 ( .A(n3656), .Z(n242) );
  MUX U899 ( .IN0(n4069), .IN1(n4067), .SEL(n4068), .F(n4046) );
  MUX U900 ( .IN0(n3559), .IN1(n3557), .SEL(n3558), .F(n3513) );
  MUX U901 ( .IN0(n243), .IN1(n3592), .SEL(n3593), .F(n3546) );
  IV U902 ( .A(n3594), .Z(n243) );
  MUX U903 ( .IN0(n3488), .IN1(n3486), .SEL(n3487), .F(n3440) );
  MUX U904 ( .IN0(n4523), .IN1(n4057), .SEL(n4058), .F(n4506) );
  MUX U905 ( .IN0(n4321), .IN1(n4319), .SEL(n4320), .F(n4297) );
  MUX U906 ( .IN0(n244), .IN1(n4034), .SEL(n3476), .F(n4013) );
  IV U907 ( .A(n3474), .Z(n244) );
  MUX U908 ( .IN0(n4692), .IN1(n4304), .SEL(n4306), .F(n4680) );
  MUX U909 ( .IN0(n3985), .IN1(n3983), .SEL(n3984), .F(n3962) );
  MUX U910 ( .IN0(n3377), .IN1(n3375), .SEL(n3376), .F(n3331) );
  MUX U911 ( .IN0(n245), .IN1(n3410), .SEL(n3411), .F(n3364) );
  IV U912 ( .A(n3412), .Z(n245) );
  MUX U913 ( .IN0(n3306), .IN1(n3304), .SEL(n3305), .F(n3261) );
  MUX U914 ( .IN0(n4455), .IN1(n3973), .SEL(n3974), .F(n4438) );
  MUX U915 ( .IN0(n4758), .IN1(n4344), .SEL(n4345), .F(n246) );
  IV U916 ( .A(n246), .Z(n4744) );
  MUX U917 ( .IN0(n4876), .IN1(n4874), .SEL(n4875), .F(n4854) );
  MUX U918 ( .IN0(n4235), .IN1(n4233), .SEL(n4234), .F(n4213) );
  MUX U919 ( .IN0(n247), .IN1(n3950), .SEL(n3294), .F(n3929) );
  IV U920 ( .A(n3292), .Z(n247) );
  MUX U921 ( .IN0(n5011), .IN1(n4861), .SEL(n4863), .F(n4999) );
  MUX U922 ( .IN0(n3825), .IN1(n3827), .SEL(n3826), .F(n3822) );
  MUX U923 ( .IN0(n4638), .IN1(n4220), .SEL(n4222), .F(n4628) );
  MUX U924 ( .IN0(n3902), .IN1(n3900), .SEL(n3901), .F(n3879) );
  MUX U925 ( .IN0(n3202), .IN1(n3200), .SEL(n3201), .F(n3158) );
  MUX U926 ( .IN0(n248), .IN1(n3232), .SEL(n3233), .F(n3190) );
  IV U927 ( .A(n3234), .Z(n248) );
  MUX U928 ( .IN0(n3133), .IN1(n3131), .SEL(n3132), .F(n3091) );
  MUX U929 ( .IN0(n249), .IN1(n3746), .SEL(n3747), .F(n3721) );
  IV U930 ( .A(n3748), .Z(n249) );
  XNOR U931 ( .A(n5227), .B(g_input[3]), .Z(n5228) );
  XNOR U932 ( .A(n4481), .B(g_input[23]), .Z(n4482) );
  MUX U933 ( .IN0(n4389), .IN1(n3890), .SEL(n3891), .F(n4372) );
  MUX U934 ( .IN0(n5229), .IN1(n250), .SEL(n5230), .F(n3013) );
  MUX U935 ( .IN0(n2108), .IN1(n2110), .SEL(n2109), .F(n2000) );
  MUX U936 ( .IN0(n2363), .IN1(n251), .SEL(n2364), .F(n2243) );
  IV U937 ( .A(n2365), .Z(n251) );
  MUX U938 ( .IN0(n2578), .IN1(n2580), .SEL(n2579), .F(n2453) );
  MUX U939 ( .IN0(n2535), .IN1(n2537), .SEL(n2536), .F(n2413) );
  MUX U940 ( .IN0(n2858), .IN1(n2860), .SEL(n2859), .F(n2726) );
  XNOR U941 ( .A(n5068), .B(n5067), .Z(n5073) );
  XNOR U942 ( .A(n4783), .B(n4782), .Z(n4809) );
  XNOR U943 ( .A(n4151), .B(n4149), .Z(n4164) );
  MUX U944 ( .IN0(n252), .IN1(n3867), .SEL(n3122), .F(n3847) );
  IV U945 ( .A(n3120), .Z(n252) );
  MUX U946 ( .IN0(n933), .IN1(n931), .SEL(n932), .F(n863) );
  MUX U947 ( .IN0(n1010), .IN1(n1008), .SEL(n1009), .F(n941) );
  MUX U948 ( .IN0(n253), .IN1(n5135), .SEL(e_input[31]), .F(n1129) );
  IV U949 ( .A(e_input[19]), .Z(n253) );
  MUX U950 ( .IN0(n254), .IN1(n1416), .SEL(n1417), .F(n1325) );
  IV U951 ( .A(n1418), .Z(n254) );
  MUX U952 ( .IN0(n255), .IN1(n3832), .SEL(e_input[31]), .F(n1634) );
  IV U953 ( .A(e_input[13]), .Z(n255) );
  MUX U954 ( .IN0(n1658), .IN1(n1656), .SEL(n1657), .F(n1558) );
  MUX U955 ( .IN0(n1848), .IN1(n1846), .SEL(n1847), .F(n1729) );
  MUX U956 ( .IN0(n256), .IN1(n2127), .SEL(n2128), .F(n2019) );
  IV U957 ( .A(n2129), .Z(n256) );
  MUX U958 ( .IN0(n2360), .IN1(n2358), .SEL(n2359), .F(n2238) );
  MUX U959 ( .IN0(n2940), .IN1(n2938), .SEL(n2939), .F(n2801) );
  XNOR U960 ( .A(n2992), .B(n2991), .Z(n4968) );
  MUX U961 ( .IN0(n257), .IN1(n3034), .SEL(n3035), .F(n2906) );
  IV U962 ( .A(n3036), .Z(n257) );
  XOR U963 ( .A(n964), .B(n902), .Z(n899) );
  MUX U964 ( .IN0(n258), .IN1(n1062), .SEL(n1063), .F(n990) );
  IV U965 ( .A(n1064), .Z(n258) );
  ANDN U966 ( .A(n1126), .B(n1125), .Z(n1053) );
  XNOR U967 ( .A(n1231), .B(n1230), .Z(n1308) );
  MUX U968 ( .IN0(n1288), .IN1(n259), .SEL(n1289), .F(n1211) );
  IV U969 ( .A(n1290), .Z(n259) );
  XNOR U970 ( .A(n1601), .B(n1600), .Z(n1692) );
  XNOR U971 ( .A(n1585), .B(n1584), .Z(n1674) );
  MUX U972 ( .IN0(n260), .IN1(n1772), .SEL(n1773), .F(n1671) );
  IV U973 ( .A(n1774), .Z(n260) );
  MUX U974 ( .IN0(n261), .IN1(n1790), .SEL(n1791), .F(n1689) );
  IV U975 ( .A(n1792), .Z(n261) );
  XNOR U976 ( .A(n1705), .B(n1704), .Z(n1801) );
  XNOR U977 ( .A(n1888), .B(n1887), .Z(n1990) );
  MUX U978 ( .IN0(n262), .IN1(n2230), .SEL(n2231), .F(n2111) );
  IV U979 ( .A(n2232), .Z(n262) );
  XNOR U980 ( .A(n2158), .B(n2168), .Z(n2274) );
  XNOR U981 ( .A(n2175), .B(n2174), .Z(n2284) );
  XNOR U982 ( .A(n2199), .B(n2198), .Z(n2314) );
  XNOR U983 ( .A(n2222), .B(n2221), .Z(n2337) );
  MUX U984 ( .IN0(n263), .IN1(n2456), .SEL(n2457), .F(n2334) );
  IV U985 ( .A(n2458), .Z(n263) );
  XNOR U986 ( .A(n2531), .B(n2530), .Z(n2650) );
  XNOR U987 ( .A(n2523), .B(n2522), .Z(n2642) );
  XNOR U988 ( .A(n2589), .B(n2588), .Z(n2716) );
  XNOR U989 ( .A(n2698), .B(n2697), .Z(n2825) );
  XNOR U990 ( .A(n2737), .B(n2736), .Z(n2864) );
  XNOR U991 ( .A(n2745), .B(n2744), .Z(n2872) );
  MUX U992 ( .IN0(n591), .IN1(n589), .SEL(n590), .F(n559) );
  NAND U993 ( .A(n702), .B(n701), .Z(n695) );
  XNOR U994 ( .A(n664), .B(n663), .Z(n703) );
  MUX U995 ( .IN0(n264), .IN1(n790), .SEL(n791), .F(n734) );
  IV U996 ( .A(n792), .Z(n264) );
  AND U997 ( .A(n1335), .B(n1337), .Z(n1251) );
  MUX U998 ( .IN0(n265), .IN1(n1369), .SEL(n1370), .F(n1278) );
  IV U999 ( .A(n1371), .Z(n265) );
  MUX U1000 ( .IN0(n266), .IN1(n1872), .SEL(n1873), .F(n1764) );
  IV U1001 ( .A(n1874), .Z(n266) );
  AND U1002 ( .A(n1922), .B(n1924), .Z(n1816) );
  MUX U1003 ( .IN0(n267), .IN1(n2326), .SEL(n2327), .F(n2206) );
  IV U1004 ( .A(n2328), .Z(n267) );
  XNOR U1005 ( .A(n2307), .B(n2306), .Z(n2304) );
  ANDN U1006 ( .A(n2498), .B(n2499), .Z(n2376) );
  MUX U1007 ( .IN0(n2688), .IN1(n2811), .SEL(n2690), .F(n2555) );
  MUX U1008 ( .IN0(n2839), .IN1(n361), .SEL(n2838), .F(n268) );
  IV U1009 ( .A(n268), .Z(n2705) );
  MUX U1010 ( .IN0(n269), .IN1(n2808), .SEL(n2809), .F(n2685) );
  IV U1011 ( .A(n2810), .Z(n269) );
  ANDN U1012 ( .A(n633), .B(n603), .Z(n592) );
  MUX U1013 ( .IN0(n835), .IN1(n837), .SEL(n836), .F(n270) );
  IV U1014 ( .A(n270), .Z(n780) );
  AND U1015 ( .A(n892), .B(n894), .Z(n829) );
  XOR U1016 ( .A(n844), .B(n841), .Z(n895) );
  NANDN U1017 ( .B(n952), .A(n953), .Z(n884) );
  XNOR U1018 ( .A(n1629), .B(n1630), .Z(n1649) );
  MUX U1019 ( .IN0(n271), .IN1(n2416), .SEL(n2417), .F(n2296) );
  IV U1020 ( .A(n2418), .Z(n271) );
  MUX U1021 ( .IN0(n2931), .IN1(n2929), .SEL(n2930), .F(n272) );
  IV U1022 ( .A(n272), .Z(n2792) );
  MUX U1023 ( .IN0(n529), .IN1(n527), .SEL(n528), .F(n273) );
  IV U1024 ( .A(n273), .Z(n506) );
  NANDN U1025 ( .B(n533), .A(n534), .Z(n490) );
  XOR U1026 ( .A(n1122), .B(n1121), .Z(n1102) );
  XOR U1027 ( .A(n1351), .B(n1350), .Z(n1435) );
  XOR U1028 ( .A(n1964), .B(n1961), .Z(n2038) );
  AND U1029 ( .A(n518), .B(n520), .Z(n493) );
  MUX U1030 ( .IN0(n2887), .IN1(\_MxM/Y0[1] ), .SEL(n2888), .F(n2755) );
  XNOR U1031 ( .A(n564), .B(n568), .Z(n566) );
  XNOR U1032 ( .A(n676), .B(n680), .Z(n678) );
  XNOR U1033 ( .A(n823), .B(n827), .Z(n825) );
  XNOR U1034 ( .A(n1021), .B(n1025), .Z(n1023) );
  XNOR U1035 ( .A(n1254), .B(n1258), .Z(n1256) );
  XNOR U1036 ( .A(n1526), .B(n1530), .Z(n1528) );
  XNOR U1037 ( .A(n1819), .B(n1823), .Z(n1821) );
  XNOR U1038 ( .A(n2140), .B(n2144), .Z(n2142) );
  MUX U1039 ( .IN0(n274), .IN1(n4160), .SEL(n3743), .F(n4139) );
  IV U1040 ( .A(n3742), .Z(n274) );
  MUX U1041 ( .IN0(n3624), .IN1(n3622), .SEL(n3623), .F(n3576) );
  MUX U1042 ( .IN0(n4111), .IN1(n4109), .SEL(n4110), .F(n4088) );
  MUX U1043 ( .IN0(n4557), .IN1(n4099), .SEL(n4100), .F(n4540) );
  MUX U1044 ( .IN0(n275), .IN1(n3546), .SEL(n3547), .F(n3502) );
  IV U1045 ( .A(n3548), .Z(n275) );
  MUX U1046 ( .IN0(n276), .IN1(n4076), .SEL(n3566), .F(n4055) );
  IV U1047 ( .A(n3564), .Z(n276) );
  MUX U1048 ( .IN0(n3442), .IN1(n3440), .SEL(n3441), .F(n3394) );
  MUX U1049 ( .IN0(n4027), .IN1(n4025), .SEL(n4026), .F(n4004) );
  MUX U1050 ( .IN0(n3469), .IN1(n3467), .SEL(n3468), .F(n3421) );
  MUX U1051 ( .IN0(n4489), .IN1(n4015), .SEL(n4016), .F(n4472) );
  MUX U1052 ( .IN0(n3838), .IN1(n4322), .SEL(n3839), .F(n277) );
  IV U1053 ( .A(n277), .Z(n4300) );
  MUX U1054 ( .IN0(n4680), .IN1(n4280), .SEL(n4282), .F(n4665) );
  MUX U1055 ( .IN0(n4275), .IN1(n4273), .SEL(n4274), .F(n4253) );
  MUX U1056 ( .IN0(n278), .IN1(n3364), .SEL(n3365), .F(n3320) );
  IV U1057 ( .A(n3366), .Z(n278) );
  MUX U1058 ( .IN0(n279), .IN1(n3992), .SEL(n3384), .F(n3971) );
  IV U1059 ( .A(n3382), .Z(n279) );
  MUX U1060 ( .IN0(n4898), .IN1(n4896), .SEL(n4897), .F(n4874) );
  MUX U1061 ( .IN0(n5037), .IN1(n4903), .SEL(n4905), .F(n5023) );
  MUX U1062 ( .IN0(n3263), .IN1(n3261), .SEL(n3262), .F(n3218) );
  MUX U1063 ( .IN0(n3943), .IN1(n3941), .SEL(n3942), .F(n3920) );
  MUX U1064 ( .IN0(n3287), .IN1(n3285), .SEL(n3286), .F(n3243) );
  MUX U1065 ( .IN0(n4422), .IN1(n3931), .SEL(n3932), .F(n4406) );
  MUX U1066 ( .IN0(g_input[1]), .IN1(n5244), .SEL(g_input[31]), .F(n280) );
  IV U1067 ( .A(n280), .Z(n3812) );
  MUX U1068 ( .IN0(n281), .IN1(n5163), .SEL(n5164), .F(n5152) );
  IV U1069 ( .A(n5165), .Z(n281) );
  MUX U1070 ( .IN0(n4628), .IN1(n4200), .SEL(n4202), .F(n4618) );
  MUX U1071 ( .IN0(n4195), .IN1(n4193), .SEL(n4194), .F(n4169) );
  MUX U1072 ( .IN0(n282), .IN1(n3190), .SEL(n3191), .F(n3147) );
  IV U1073 ( .A(n3192), .Z(n282) );
  MUX U1074 ( .IN0(n283), .IN1(n3909), .SEL(n3209), .F(n3888) );
  IV U1075 ( .A(n3207), .Z(n283) );
  XNOR U1076 ( .A(n5150), .B(g_input[7]), .Z(n5151) );
  XNOR U1077 ( .A(n5018), .B(g_input[11]), .Z(n5019) );
  XNOR U1078 ( .A(n4970), .B(g_input[15]), .Z(n4971) );
  XNOR U1079 ( .A(n4549), .B(g_input[19]), .Z(n4550) );
  MUX U1080 ( .IN0(g_input[2]), .IN1(n5237), .SEL(g_input[31]), .F(n284) );
  IV U1081 ( .A(n284), .Z(n3809) );
  MUX U1082 ( .IN0(n4816), .IN1(n4814), .SEL(n4815), .F(n4783) );
  MUX U1083 ( .IN0(n4987), .IN1(n4821), .SEL(n4823), .F(n4975) );
  MUX U1084 ( .IN0(n3093), .IN1(n3091), .SEL(n3092), .F(n3052) );
  MUX U1085 ( .IN0(n3115), .IN1(n3113), .SEL(n3114), .F(n3044) );
  XNOR U1086 ( .A(n4447), .B(g_input[25]), .Z(n4448) );
  MUX U1087 ( .IN0(n285), .IN1(n3819), .SEL(e_input[31]), .F(n2050) );
  IV U1088 ( .A(e_input[9]), .Z(n285) );
  MUX U1089 ( .IN0(n2570), .IN1(n2572), .SEL(n2571), .F(n2445) );
  MUX U1090 ( .IN0(n2789), .IN1(n2791), .SEL(n2790), .F(n2659) );
  MUX U1091 ( .IN0(g_input[4]), .IN1(n5196), .SEL(g_input[31]), .F(n2748) );
  MUX U1092 ( .IN0(n3013), .IN1(n286), .SEL(n3014), .F(n2874) );
  IV U1093 ( .A(n3015), .Z(n286) );
  MUX U1094 ( .IN0(g_input[9]), .IN1(n5047), .SEL(g_input[31]), .F(n287) );
  IV U1095 ( .A(n287), .Z(n2251) );
  MUX U1096 ( .IN0(n2981), .IN1(n2983), .SEL(n2982), .F(n2842) );
  MUX U1097 ( .IN0(e_input[1]), .IN1(n4776), .SEL(e_input[31]), .F(n288) );
  IV U1098 ( .A(n288), .Z(n4349) );
  XNOR U1099 ( .A(n3737), .B(n3735), .Z(n3751) );
  MUX U1100 ( .IN0(n1074), .IN1(n1072), .SEL(n1073), .F(n1000) );
  MUX U1101 ( .IN0(n289), .IN1(n1241), .SEL(n1242), .F(n1160) );
  IV U1102 ( .A(n1243), .Z(n289) );
  MUX U1103 ( .IN0(n1273), .IN1(n1271), .SEL(n1272), .F(n1189) );
  MUX U1104 ( .IN0(n1297), .IN1(n1299), .SEL(n1298), .F(n290) );
  MUX U1105 ( .IN0(n1699), .IN1(n1697), .SEL(n1698), .F(n1601) );
  MUX U1106 ( .IN0(n2283), .IN1(n2281), .SEL(n2282), .F(n2158) );
  MUX U1107 ( .IN0(n2803), .IN1(n2801), .SEL(n2802), .F(n2667) );
  MUX U1108 ( .IN0(n4352), .IN1(n3865), .SEL(n3866), .F(n291) );
  IV U1109 ( .A(n291), .Z(n2959) );
  XNOR U1110 ( .A(n4946), .B(n4943), .Z(n4944) );
  XNOR U1111 ( .A(n5249), .B(e_input[30]), .Z(n5247) );
  MUX U1112 ( .IN0(n292), .IN1(n853), .SEL(n854), .F(n790) );
  IV U1113 ( .A(n855), .Z(n292) );
  XNOR U1114 ( .A(n1315), .B(n1314), .Z(n1403) );
  MUX U1115 ( .IN0(n293), .IN1(n1479), .SEL(n1480), .F(n1379) );
  IV U1116 ( .A(n1481), .Z(n293) );
  MUX U1117 ( .IN0(n294), .IN1(n1593), .SEL(n1594), .F(n1497) );
  IV U1118 ( .A(n1595), .Z(n294) );
  XNOR U1119 ( .A(n1513), .B(n1512), .Z(n1604) );
  XNOR U1120 ( .A(n1558), .B(n1557), .Z(n1651) );
  XNOR U1121 ( .A(n1681), .B(n1680), .Z(n1775) );
  XNOR U1122 ( .A(n1846), .B(n1845), .Z(n1947) );
  XNOR U1123 ( .A(n2011), .B(n2010), .Z(n2114) );
  XNOR U1124 ( .A(n2019), .B(n2018), .Z(n2122) );
  XNOR U1125 ( .A(n1972), .B(n1971), .Z(n2075) );
  MUX U1126 ( .IN0(n295), .IN1(n2095), .SEL(n2096), .F(n1987) );
  IV U1127 ( .A(n2097), .Z(n295) );
  XNOR U1128 ( .A(n2342), .B(n2341), .Z(n2459) );
  MUX U1129 ( .IN0(n296), .IN1(n2472), .SEL(n2473), .F(n2350) );
  IV U1130 ( .A(n2474), .Z(n296) );
  XNOR U1131 ( .A(n2289), .B(n2288), .Z(n2404) );
  MUX U1132 ( .IN0(n297), .IN1(n2391), .SEL(n2392), .F(n2271) );
  IV U1133 ( .A(n2393), .Z(n297) );
  XNOR U1134 ( .A(n2605), .B(n2604), .Z(n2732) );
  XNOR U1135 ( .A(n2613), .B(n2612), .Z(n2740) );
  XNOR U1136 ( .A(n2566), .B(n2565), .Z(n2693) );
  XNOR U1137 ( .A(n2721), .B(n2720), .Z(n2848) );
  XNOR U1138 ( .A(n2655), .B(n2654), .Z(n2780) );
  XNOR U1139 ( .A(n2647), .B(n2646), .Z(n2772) );
  MUX U1140 ( .IN0(n3002), .IN1(n3000), .SEL(n3001), .F(n298) );
  IV U1141 ( .A(n298), .Z(n2861) );
  MUX U1142 ( .IN0(n299), .IN1(n2984), .SEL(n2985), .F(n2845) );
  IV U1143 ( .A(n2986), .Z(n299) );
  MUX U1144 ( .IN0(n300), .IN1(n2906), .SEL(n2907), .F(n2769) );
  IV U1145 ( .A(n2908), .Z(n300) );
  MUX U1146 ( .IN0(n2956), .IN1(n301), .SEL(n2957), .F(n2821) );
  IV U1147 ( .A(n2958), .Z(n301) );
  MUX U1148 ( .IN0(n582), .IN1(n580), .SEL(n581), .F(n547) );
  MUX U1149 ( .IN0(n302), .IN1(n651), .SEL(n652), .F(n615) );
  IV U1150 ( .A(n653), .Z(n302) );
  XNOR U1151 ( .A(n708), .B(n707), .Z(n745) );
  XNOR U1152 ( .A(n742), .B(n740), .Z(n793) );
  AND U1153 ( .A(n844), .B(n845), .Z(n774) );
  MUX U1154 ( .IN0(n303), .IN1(n977), .SEL(n978), .F(n908) );
  IV U1155 ( .A(n979), .Z(n303) );
  XOR U1156 ( .A(n1050), .B(n1054), .Z(n1123) );
  XNOR U1157 ( .A(n1536), .B(n1535), .Z(n1534) );
  MUX U1158 ( .IN0(n304), .IN1(n1663), .SEL(n1664), .F(n1565) );
  IV U1159 ( .A(n1665), .Z(n304) );
  AND U1160 ( .A(n1715), .B(n1717), .Z(n1619) );
  MUX U1161 ( .IN0(n305), .IN1(n1727), .SEL(n1726), .F(n1630) );
  IV U1162 ( .A(n1725), .Z(n305) );
  AND U1163 ( .A(n2137), .B(n2139), .Z(n2029) );
  MUX U1164 ( .IN0(n306), .IN1(n2206), .SEL(n2207), .F(n2087) );
  IV U1165 ( .A(n2208), .Z(n306) );
  MUX U1166 ( .IN0(n307), .IN1(n2705), .SEL(n2706), .F(n2573) );
  IV U1167 ( .A(n2707), .Z(n307) );
  MUX U1168 ( .IN0(n556), .IN1(n558), .SEL(n557), .F(n524) );
  AND U1169 ( .A(n779), .B(n780), .Z(n776) );
  MUX U1170 ( .IN0(n308), .IN1(n1745), .SEL(n1746), .F(n1644) );
  IV U1171 ( .A(n1747), .Z(n308) );
  XOR U1172 ( .A(n2185), .B(n2071), .Z(n2072) );
  XNOR U1173 ( .A(n2432), .B(n2430), .Z(n2541) );
  NANDN U1174 ( .B(n531), .A(n530), .Z(n502) );
  XNOR U1175 ( .A(n533), .B(n538), .Z(n534) );
  XNOR U1176 ( .A(n634), .B(n639), .Z(n635) );
  XNOR U1177 ( .A(n762), .B(n727), .Z(n763) );
  XNOR U1178 ( .A(n952), .B(n957), .Z(n953) );
  XOR U1179 ( .A(n1200), .B(n1199), .Z(n1180) );
  MUX U1180 ( .IN0(\_MxM/Y0[2] ), .IN1(n2755), .SEL(n2756), .F(n2623) );
  XOR U1181 ( .A(n1353), .B(n1352), .Z(n1432) );
  XOR U1182 ( .A(n1963), .B(n1962), .Z(n2035) );
  XOR U1183 ( .A(n2298), .B(n2297), .Z(n2382) );
  XNOR U1184 ( .A(n2628), .B(n2507), .Z(n2508) );
  XOR U1185 ( .A(n2794), .B(n2793), .Z(n2897) );
  XNOR U1186 ( .A(n595), .B(n599), .Z(n597) );
  XNOR U1187 ( .A(n720), .B(n724), .Z(n722) );
  XNOR U1188 ( .A(n886), .B(n890), .Z(n888) );
  XNOR U1189 ( .A(n1095), .B(n1099), .Z(n1097) );
  XNOR U1190 ( .A(n1338), .B(n1342), .Z(n1340) );
  XNOR U1191 ( .A(n1622), .B(n1626), .Z(n1624) );
  XNOR U1192 ( .A(n1925), .B(n1929), .Z(n1927) );
  XNOR U1193 ( .A(n2259), .B(n2263), .Z(n2261) );
  XOR U1194 ( .A(n478), .B(n479), .Z(n365) );
  MUX U1195 ( .IN0(n3714), .IN1(n3712), .SEL(n3713), .F(n3668) );
  MUX U1196 ( .IN0(n3697), .IN1(n3695), .SEL(n3696), .F(n3649) );
  MUX U1197 ( .IN0(n309), .IN1(n3638), .SEL(n3639), .F(n3592) );
  IV U1198 ( .A(n3640), .Z(n309) );
  MUX U1199 ( .IN0(n3534), .IN1(n3532), .SEL(n3533), .F(n3486) );
  MUX U1200 ( .IN0(n310), .IN1(n4097), .SEL(n3612), .F(n4076) );
  IV U1201 ( .A(n3610), .Z(n310) );
  MUX U1202 ( .IN0(n4540), .IN1(n4078), .SEL(n4079), .F(n4523) );
  MUX U1203 ( .IN0(n4048), .IN1(n4046), .SEL(n4047), .F(n4025) );
  MUX U1204 ( .IN0(n3515), .IN1(n3513), .SEL(n3514), .F(n3467) );
  MUX U1205 ( .IN0(n311), .IN1(n3456), .SEL(n3457), .F(n3410) );
  IV U1206 ( .A(n3458), .Z(n311) );
  MUX U1207 ( .IN0(n3352), .IN1(n3350), .SEL(n3351), .F(n3304) );
  MUX U1208 ( .IN0(n312), .IN1(n4013), .SEL(n3430), .F(n3992) );
  IV U1209 ( .A(n3428), .Z(n312) );
  MUX U1210 ( .IN0(n4472), .IN1(n3994), .SEL(n3995), .F(n4455) );
  MUX U1211 ( .IN0(n4922), .IN1(n4920), .SEL(n4921), .F(n4896) );
  MUX U1212 ( .IN0(n5054), .IN1(n4927), .SEL(n4929), .F(n5037) );
  MUX U1213 ( .IN0(n3964), .IN1(n3962), .SEL(n3963), .F(n3941) );
  MUX U1214 ( .IN0(n3333), .IN1(n3331), .SEL(n3332), .F(n3285) );
  MUX U1215 ( .IN0(n4665), .IN1(n4260), .SEL(n4262), .F(n4650) );
  MUX U1216 ( .IN0(n4255), .IN1(n4253), .SEL(n4254), .F(n4233) );
  MUX U1217 ( .IN0(n5122), .IN1(n4966), .SEL(n4967), .F(n313) );
  IV U1218 ( .A(n313), .Z(n5108) );
  MUX U1219 ( .IN0(n3798), .IN1(n3749), .SEL(n3750), .F(n314) );
  IV U1220 ( .A(n314), .Z(n3784) );
  MUX U1221 ( .IN0(n315), .IN1(n3781), .SEL(n3782), .F(n3767) );
  IV U1222 ( .A(n3783), .Z(n315) );
  MUX U1223 ( .IN0(n316), .IN1(n3275), .SEL(n3276), .F(n3232) );
  IV U1224 ( .A(n3277), .Z(n316) );
  MUX U1225 ( .IN0(n5205), .IN1(n5146), .SEL(n5147), .F(n317) );
  IV U1226 ( .A(n317), .Z(n5189) );
  MUX U1227 ( .IN0(n3178), .IN1(n3176), .SEL(n3177), .F(n3131) );
  MUX U1228 ( .IN0(n318), .IN1(n3929), .SEL(n3252), .F(n3909) );
  IV U1229 ( .A(n3250), .Z(n318) );
  MUX U1230 ( .IN0(n4406), .IN1(n3911), .SEL(n3912), .F(n4389) );
  MUX U1231 ( .IN0(n5233), .IN1(n5235), .SEL(n5234), .F(n5229) );
  MUX U1232 ( .IN0(n4836), .IN1(n4834), .SEL(n4835), .F(n4814) );
  MUX U1233 ( .IN0(n4999), .IN1(n4841), .SEL(n4843), .F(n4987) );
  MUX U1234 ( .IN0(n319), .IN1(n3753), .SEL(n3754), .F(n3731) );
  IV U1235 ( .A(n3755), .Z(n319) );
  MUX U1236 ( .IN0(n3881), .IN1(n3879), .SEL(n3880), .F(n3855) );
  MUX U1237 ( .IN0(n3160), .IN1(n3158), .SEL(n3159), .F(n3113) );
  XNOR U1238 ( .A(n5177), .B(g_input[5]), .Z(n5178) );
  XNOR U1239 ( .A(n5046), .B(g_input[9]), .Z(n5047) );
  MUX U1240 ( .IN0(n320), .IN1(n4960), .SEL(e_input[31]), .F(n4952) );
  IV U1241 ( .A(e_input[21]), .Z(n320) );
  XNOR U1242 ( .A(n4994), .B(g_input[13]), .Z(n4995) );
  XNOR U1243 ( .A(n4583), .B(g_input[17]), .Z(n4584) );
  XNOR U1244 ( .A(n4515), .B(g_input[21]), .Z(n4516) );
  AND U1245 ( .A(n5245), .B(g_input[0]), .Z(n3023) );
  MUX U1246 ( .IN0(n4171), .IN1(n4169), .SEL(n4170), .F(n4151) );
  MUX U1247 ( .IN0(n4618), .IN1(n4180), .SEL(n4182), .F(n4608) );
  MUX U1248 ( .IN0(n321), .IN1(n5224), .SEL(e_input[31]), .F(n5211) );
  IV U1249 ( .A(e_input[25]), .Z(n321) );
  MUX U1250 ( .IN0(n322), .IN1(n5242), .SEL(e_input[31]), .F(n5232) );
  IV U1251 ( .A(e_input[29]), .Z(n322) );
  XNOR U1252 ( .A(n4415), .B(g_input[27]), .Z(n4416) );
  MUX U1253 ( .IN0(g_input[3]), .IN1(n5228), .SEL(g_input[31]), .F(n2880) );
  MUX U1254 ( .IN0(n2997), .IN1(n2999), .SEL(n2998), .F(n2858) );
  MUX U1255 ( .IN0(n2973), .IN1(n2975), .SEL(n2974), .F(n2834) );
  MUX U1256 ( .IN0(e_input[20]), .IN1(n323), .SEL(e_input[31]), .F(n1032) );
  IV U1257 ( .A(n4959), .Z(n323) );
  MUX U1258 ( .IN0(e_input[16]), .IN1(n324), .SEL(e_input[31]), .F(n1394) );
  IV U1259 ( .A(n5139), .Z(n324) );
  MUX U1260 ( .IN0(e_input[8]), .IN1(n325), .SEL(e_input[31]), .F(n2169) );
  IV U1261 ( .A(n3818), .Z(n325) );
  MUX U1262 ( .IN0(e_input[12]), .IN1(n326), .SEL(e_input[31]), .F(n1740) );
  IV U1263 ( .A(n3831), .Z(n326) );
  MUX U1264 ( .IN0(e_input[4]), .IN1(n327), .SEL(e_input[31]), .F(n2678) );
  IV U1265 ( .A(n4337), .Z(n327) );
  XNOR U1266 ( .A(n4325), .B(n4322), .Z(n4323) );
  MUX U1267 ( .IN0(n328), .IN1(n3103), .SEL(n3104), .F(n3034) );
  IV U1268 ( .A(n3105), .Z(n328) );
  MUX U1269 ( .IN0(n329), .IN1(n5218), .SEL(e_input[31]), .F(n647) );
  IV U1270 ( .A(e_input[27]), .Z(n329) );
  MUX U1271 ( .IN0(e_input[26]), .IN1(n330), .SEL(e_input[31]), .F(n688) );
  IV U1272 ( .A(n5219), .Z(n330) );
  MUX U1273 ( .IN0(e_input[24]), .IN1(n331), .SEL(e_input[31]), .F(n795) );
  IV U1274 ( .A(n5223), .Z(n331) );
  MUX U1275 ( .IN0(e_input[28]), .IN1(n332), .SEL(e_input[31]), .F(n620) );
  IV U1276 ( .A(n5241), .Z(n332) );
  MUX U1277 ( .IN0(n1113), .IN1(n1111), .SEL(n1112), .F(n1038) );
  MUX U1278 ( .IN0(n333), .IN1(n1160), .SEL(n1161), .F(n1082) );
  IV U1279 ( .A(n1162), .Z(n333) );
  MUX U1280 ( .IN0(n1154), .IN1(n1152), .SEL(n1153), .F(n1072) );
  MUX U1281 ( .IN0(e_input[18]), .IN1(n334), .SEL(e_input[31]), .F(n1210) );
  IV U1282 ( .A(n5134), .Z(n334) );
  MUX U1283 ( .IN0(n335), .IN1(n5140), .SEL(e_input[31]), .F(n1294) );
  IV U1284 ( .A(e_input[17]), .Z(n335) );
  MUX U1285 ( .IN0(n1491), .IN1(n1489), .SEL(n1490), .F(n1383) );
  MUX U1286 ( .IN0(n1464), .IN1(n1462), .SEL(n1463), .F(n1360) );
  MUX U1287 ( .IN0(n1507), .IN1(n1505), .SEL(n1506), .F(n1408) );
  MUX U1288 ( .IN0(n336), .IN1(n1513), .SEL(n1514), .F(n1416) );
  IV U1289 ( .A(n1515), .Z(n336) );
  MUX U1290 ( .IN0(n337), .IN1(n3814), .SEL(e_input[31]), .F(n1833) );
  IV U1291 ( .A(e_input[11]), .Z(n337) );
  MUX U1292 ( .IN0(e_input[10]), .IN1(n338), .SEL(e_input[31]), .F(n1939) );
  IV U1293 ( .A(n3813), .Z(n338) );
  MUX U1294 ( .IN0(n2063), .IN1(n2061), .SEL(n2062), .F(n1954) );
  MUX U1295 ( .IN0(e_input[6]), .IN1(n339), .SEL(e_input[31]), .F(n2429) );
  IV U1296 ( .A(n4342), .Z(n339) );
  MUX U1297 ( .IN0(n340), .IN1(n4338), .SEL(e_input[31]), .F(n2545) );
  IV U1298 ( .A(e_input[5]), .Z(n340) );
  MUX U1299 ( .IN0(n341), .IN1(n4772), .SEL(e_input[31]), .F(n2818) );
  IV U1300 ( .A(e_input[3]), .Z(n341) );
  MUX U1301 ( .IN0(e_input[2]), .IN1(n342), .SEL(e_input[31]), .F(n2955) );
  IV U1302 ( .A(n4771), .Z(n342) );
  MUX U1303 ( .IN0(n3847), .IN1(n343), .SEL(n3084), .F(n2956) );
  IV U1304 ( .A(n3083), .Z(n343) );
  MUX U1305 ( .IN0(e_input[22]), .IN1(n344), .SEL(e_input[31]), .F(n904) );
  IV U1306 ( .A(n4965), .Z(n344) );
  MUX U1307 ( .IN0(n345), .IN1(n4964), .SEL(e_input[31]), .F(n834) );
  IV U1308 ( .A(e_input[23]), .Z(n345) );
  MUX U1309 ( .IN0(n346), .IN1(n921), .SEL(n922), .F(n853) );
  IV U1310 ( .A(n923), .Z(n346) );
  MUX U1311 ( .IN0(n347), .IN1(n1221), .SEL(n1222), .F(n1142) );
  IV U1312 ( .A(n1223), .Z(n347) );
  MUX U1313 ( .IN0(n1639), .IN1(n1637), .SEL(n1638), .F(n348) );
  MUX U1314 ( .IN0(e_input[14]), .IN1(n349), .SEL(e_input[31]), .F(n1543) );
  IV U1315 ( .A(n3836), .Z(n349) );
  MUX U1316 ( .IN0(n350), .IN1(n1575), .SEL(n1576), .F(n1479) );
  IV U1317 ( .A(n1577), .Z(n350) );
  XNOR U1318 ( .A(n1798), .B(n1797), .Z(n1899) );
  XNOR U1319 ( .A(n1806), .B(n1805), .Z(n1907) );
  XNOR U1320 ( .A(n1757), .B(n1756), .Z(n1860) );
  XNOR U1321 ( .A(n1782), .B(n1781), .Z(n1883) );
  MUX U1322 ( .IN0(n351), .IN1(n1987), .SEL(n1988), .F(n1880) );
  IV U1323 ( .A(n1989), .Z(n351) );
  MUX U1324 ( .IN0(n352), .IN1(n2003), .SEL(n2004), .F(n1896) );
  IV U1325 ( .A(n2005), .Z(n352) );
  MUX U1326 ( .IN0(n1943), .IN1(n2047), .SEL(n1945), .F(n1835) );
  XNOR U1327 ( .A(n2103), .B(n2102), .Z(n2217) );
  XNOR U1328 ( .A(n2080), .B(n2079), .Z(n2194) );
  XNOR U1329 ( .A(n2119), .B(n2118), .Z(n2233) );
  XNOR U1330 ( .A(n2127), .B(n2126), .Z(n2241) );
  MUX U1331 ( .IN0(n353), .IN1(n2154), .SEL(n2155), .F(n2044) );
  IV U1332 ( .A(n2156), .Z(n353) );
  MUX U1333 ( .IN0(n354), .IN1(n4343), .SEL(e_input[31]), .F(n2303) );
  IV U1334 ( .A(e_input[7]), .Z(n354) );
  XNOR U1335 ( .A(n2488), .B(n2487), .Z(n2608) );
  XNOR U1336 ( .A(n2480), .B(n2479), .Z(n2600) );
  XNOR U1337 ( .A(n2441), .B(n2440), .Z(n2561) );
  XNOR U1338 ( .A(n2464), .B(n2463), .Z(n2584) );
  XNOR U1339 ( .A(n2401), .B(n2400), .Z(n2518) );
  XNOR U1340 ( .A(n2409), .B(n2408), .Z(n2526) );
  MUX U1341 ( .IN0(n355), .IN1(n2639), .SEL(n2640), .F(n2515) );
  IV U1342 ( .A(n2641), .Z(n355) );
  MUX U1343 ( .IN0(n356), .IN1(n2729), .SEL(n2730), .F(n2597) );
  IV U1344 ( .A(n2731), .Z(n356) );
  MUX U1345 ( .IN0(n357), .IN1(n2713), .SEL(n2714), .F(n2581) );
  IV U1346 ( .A(n2715), .Z(n357) );
  XNOR U1347 ( .A(n2877), .B(n2876), .Z(n3011) );
  XNOR U1348 ( .A(n2869), .B(n2868), .Z(n3003) );
  XNOR U1349 ( .A(n2830), .B(n2829), .Z(n2964) );
  XNOR U1350 ( .A(n2853), .B(n2852), .Z(n2987) );
  XNOR U1351 ( .A(n2777), .B(n2776), .Z(n2909) );
  XNOR U1352 ( .A(n2785), .B(n2784), .Z(n2917) );
  MUX U1353 ( .IN0(n2959), .IN1(n4346), .SEL(n2961), .F(n2820) );
  XNOR U1354 ( .A(n2801), .B(n2800), .Z(n2933) );
  MUX U1355 ( .IN0(e_input[30]), .IN1(n358), .SEL(e_input[31]), .F(n554) );
  IV U1356 ( .A(n5247), .Z(n358) );
  XNOR U1357 ( .A(n697), .B(n701), .Z(n737) );
  NAND U1358 ( .A(n902), .B(n901), .Z(n896) );
  MUX U1359 ( .IN0(n905), .IN1(n907), .SEL(n906), .F(n835) );
  XNOR U1360 ( .A(n750), .B(n749), .Z(n804) );
  NAND U1361 ( .A(n1053), .B(n1054), .Z(n1048) );
  MUX U1362 ( .IN0(n359), .IN1(n1469), .SEL(n1470), .F(n1369) );
  IV U1363 ( .A(n1471), .Z(n359) );
  MUX U1364 ( .IN0(n360), .IN1(n3837), .SEL(e_input[31]), .F(n1442) );
  IV U1365 ( .A(e_input[15]), .Z(n360) );
  AND U1366 ( .A(n1523), .B(n1525), .Z(n1426) );
  ANDN U1367 ( .A(n1964), .B(n1965), .Z(n1856) );
  MUX U1368 ( .IN0(n2978), .IN1(n2976), .SEL(n2977), .F(n361) );
  IV U1369 ( .A(n361), .Z(n2837) );
  MUX U1370 ( .IN0(n362), .IN1(n2945), .SEL(n2946), .F(n2808) );
  IV U1371 ( .A(n2947), .Z(n362) );
  MUX U1372 ( .IN0(n549), .IN1(n547), .SEL(n548), .F(n527) );
  ANDN U1373 ( .A(n559), .B(n560), .Z(n530) );
  MUX U1374 ( .IN0(n363), .IN1(n782), .SEL(n783), .F(n759) );
  IV U1375 ( .A(n784), .Z(n363) );
  XNOR U1376 ( .A(n1444), .B(n1443), .Z(n1437) );
  XNOR U1377 ( .A(n2310), .B(n2305), .Z(n2419) );
  MUX U1378 ( .IN0(n524), .IN1(n526), .SEL(n525), .F(n364) );
  IV U1379 ( .A(n364), .Z(n509) );
  XNOR U1380 ( .A(n593), .B(n598), .Z(n594) );
  XNOR U1381 ( .A(n718), .B(n723), .Z(n719) );
  XNOR U1382 ( .A(n884), .B(n889), .Z(n885) );
  XOR U1383 ( .A(n1047), .B(n1046), .Z(n1028) );
  XOR U1384 ( .A(n1280), .B(n1279), .Z(n1262) );
  XOR U1385 ( .A(n1546), .B(n1545), .Z(n1625) );
  XOR U1386 ( .A(n1747), .B(n1746), .Z(n1822) );
  XOR U1387 ( .A(n1855), .B(n1854), .Z(n1928) );
  XOR U1388 ( .A(n2070), .B(n2069), .Z(n2143) );
  XOR U1389 ( .A(n2184), .B(n2183), .Z(n2262) );
  XOR U1390 ( .A(n2418), .B(n2417), .Z(n2504) );
  XOR U1391 ( .A(n2540), .B(n2539), .Z(n2628) );
  XOR U1392 ( .A(n2664), .B(n2663), .Z(n2758) );
  AND U1393 ( .A(\_MxM/Y0[0] ), .B(n2762), .Z(n2887) );
  XNOR U1394 ( .A(n535), .B(n539), .Z(n537) );
  XNOR U1395 ( .A(n636), .B(n640), .Z(n638) );
  XNOR U1396 ( .A(n764), .B(n767), .Z(n766) );
  XNOR U1397 ( .A(n954), .B(n958), .Z(n956) );
  XNOR U1398 ( .A(n1173), .B(n1177), .Z(n1175) );
  XNOR U1399 ( .A(n1429), .B(n1433), .Z(n1431) );
  XNOR U1400 ( .A(n1718), .B(n1722), .Z(n1720) );
  XNOR U1401 ( .A(n2032), .B(n2036), .Z(n2034) );
  XNOR U1402 ( .A(n2379), .B(n2383), .Z(n2381) );
  MUX U1403 ( .IN0(n365), .IN1(n470), .SEL(n476), .F(n473) );
  ANDN U1404 ( .A(n366), .B(\_MxM/n[0] ), .Z(\_MxM/n372 ) );
  AND U1405 ( .A(\_MxM/N8 ), .B(n366), .Z(\_MxM/n371 ) );
  AND U1406 ( .A(\_MxM/N9 ), .B(n366), .Z(\_MxM/n370 ) );
  AND U1407 ( .A(\_MxM/N10 ), .B(n366), .Z(\_MxM/n369 ) );
  AND U1408 ( .A(\_MxM/N11 ), .B(n366), .Z(\_MxM/n368 ) );
  AND U1409 ( .A(\_MxM/N12 ), .B(n366), .Z(\_MxM/n367 ) );
  AND U1410 ( .A(\_MxM/N13 ), .B(n366), .Z(\_MxM/n366 ) );
  AND U1411 ( .A(\_MxM/N14 ), .B(n366), .Z(\_MxM/n365 ) );
  AND U1412 ( .A(\_MxM/N15 ), .B(n366), .Z(\_MxM/n364 ) );
  AND U1413 ( .A(n366), .B(n367), .Z(\_MxM/n363 ) );
  XOR U1414 ( .A(\_MxM/n[9] ), .B(\_MxM/add_39/carry[9] ), .Z(n367) );
  ANDN U1415 ( .A(n368), .B(rst), .Z(n366) );
  NAND U1416 ( .A(n369), .B(n370), .Z(n368) );
  AND U1417 ( .A(n371), .B(n372), .Z(n370) );
  AND U1418 ( .A(\_MxM/n[1] ), .B(n373), .Z(n372) );
  AND U1419 ( .A(n374), .B(\_MxM/n[0] ), .Z(n373) );
  AND U1420 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n371) );
  AND U1421 ( .A(n375), .B(n376), .Z(n369) );
  AND U1422 ( .A(\_MxM/n[6] ), .B(\_MxM/n[7] ), .Z(n376) );
  AND U1423 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n375) );
  NAND U1424 ( .A(n377), .B(n378), .Z(\_MxM/n362 ) );
  NAND U1425 ( .A(n379), .B(n380), .Z(n378) );
  NAND U1426 ( .A(\_MxM/Y0[0] ), .B(rst), .Z(n377) );
  NAND U1427 ( .A(n381), .B(n382), .Z(\_MxM/n361 ) );
  NAND U1428 ( .A(n383), .B(n380), .Z(n382) );
  NAND U1429 ( .A(\_MxM/Y0[1] ), .B(rst), .Z(n381) );
  NAND U1430 ( .A(n384), .B(n385), .Z(\_MxM/n360 ) );
  NAND U1431 ( .A(n386), .B(n380), .Z(n385) );
  NAND U1432 ( .A(\_MxM/Y0[2] ), .B(rst), .Z(n384) );
  NAND U1433 ( .A(n387), .B(n388), .Z(\_MxM/n359 ) );
  NAND U1434 ( .A(n389), .B(n380), .Z(n388) );
  NAND U1435 ( .A(\_MxM/Y0[3] ), .B(rst), .Z(n387) );
  NAND U1436 ( .A(n390), .B(n391), .Z(\_MxM/n358 ) );
  NAND U1437 ( .A(n392), .B(n380), .Z(n391) );
  NAND U1438 ( .A(\_MxM/Y0[4] ), .B(rst), .Z(n390) );
  NAND U1439 ( .A(n393), .B(n394), .Z(\_MxM/n357 ) );
  NAND U1440 ( .A(n395), .B(n380), .Z(n394) );
  NAND U1441 ( .A(rst), .B(\_MxM/Y0[5] ), .Z(n393) );
  NAND U1442 ( .A(n396), .B(n397), .Z(\_MxM/n356 ) );
  NAND U1443 ( .A(n398), .B(n380), .Z(n397) );
  NAND U1444 ( .A(rst), .B(\_MxM/Y0[6] ), .Z(n396) );
  NAND U1445 ( .A(n399), .B(n400), .Z(\_MxM/n355 ) );
  NAND U1446 ( .A(n401), .B(n380), .Z(n400) );
  NAND U1447 ( .A(rst), .B(\_MxM/Y0[7] ), .Z(n399) );
  NAND U1448 ( .A(n402), .B(n403), .Z(\_MxM/n354 ) );
  NAND U1449 ( .A(n404), .B(n380), .Z(n403) );
  NAND U1450 ( .A(rst), .B(\_MxM/Y0[8] ), .Z(n402) );
  NAND U1451 ( .A(n405), .B(n406), .Z(\_MxM/n353 ) );
  NAND U1452 ( .A(n407), .B(n380), .Z(n406) );
  NAND U1453 ( .A(rst), .B(\_MxM/Y0[9] ), .Z(n405) );
  NAND U1454 ( .A(n408), .B(n409), .Z(\_MxM/n352 ) );
  NAND U1455 ( .A(n410), .B(n380), .Z(n409) );
  NAND U1456 ( .A(rst), .B(\_MxM/Y0[10] ), .Z(n408) );
  NAND U1457 ( .A(n411), .B(n412), .Z(\_MxM/n351 ) );
  NAND U1458 ( .A(n413), .B(n380), .Z(n412) );
  NAND U1459 ( .A(rst), .B(\_MxM/Y0[11] ), .Z(n411) );
  NAND U1460 ( .A(n414), .B(n415), .Z(\_MxM/n350 ) );
  NAND U1461 ( .A(n416), .B(n380), .Z(n415) );
  NAND U1462 ( .A(rst), .B(\_MxM/Y0[12] ), .Z(n414) );
  NAND U1463 ( .A(n417), .B(n418), .Z(\_MxM/n349 ) );
  NAND U1464 ( .A(n419), .B(n380), .Z(n418) );
  NAND U1465 ( .A(rst), .B(\_MxM/Y0[13] ), .Z(n417) );
  NAND U1466 ( .A(n420), .B(n421), .Z(\_MxM/n348 ) );
  NAND U1467 ( .A(n422), .B(n380), .Z(n421) );
  NAND U1468 ( .A(rst), .B(\_MxM/Y0[14] ), .Z(n420) );
  NAND U1469 ( .A(n423), .B(n424), .Z(\_MxM/n347 ) );
  NAND U1470 ( .A(n425), .B(n380), .Z(n424) );
  NAND U1471 ( .A(rst), .B(\_MxM/Y0[15] ), .Z(n423) );
  NAND U1472 ( .A(n426), .B(n427), .Z(\_MxM/n346 ) );
  NAND U1473 ( .A(n428), .B(n380), .Z(n427) );
  NAND U1474 ( .A(rst), .B(\_MxM/Y0[16] ), .Z(n426) );
  NAND U1475 ( .A(n429), .B(n430), .Z(\_MxM/n345 ) );
  NAND U1476 ( .A(n431), .B(n380), .Z(n430) );
  NAND U1477 ( .A(rst), .B(\_MxM/Y0[17] ), .Z(n429) );
  NAND U1478 ( .A(n432), .B(n433), .Z(\_MxM/n344 ) );
  NAND U1479 ( .A(n434), .B(n380), .Z(n433) );
  NAND U1480 ( .A(rst), .B(\_MxM/Y0[18] ), .Z(n432) );
  NAND U1481 ( .A(n435), .B(n436), .Z(\_MxM/n343 ) );
  NAND U1482 ( .A(n437), .B(n380), .Z(n436) );
  NAND U1483 ( .A(rst), .B(\_MxM/Y0[19] ), .Z(n435) );
  NAND U1484 ( .A(n438), .B(n439), .Z(\_MxM/n342 ) );
  NAND U1485 ( .A(n440), .B(n380), .Z(n439) );
  NAND U1486 ( .A(rst), .B(\_MxM/Y0[20] ), .Z(n438) );
  NAND U1487 ( .A(n441), .B(n442), .Z(\_MxM/n341 ) );
  NAND U1488 ( .A(n443), .B(n380), .Z(n442) );
  NAND U1489 ( .A(rst), .B(\_MxM/Y0[21] ), .Z(n441) );
  NAND U1490 ( .A(n444), .B(n445), .Z(\_MxM/n340 ) );
  NAND U1491 ( .A(n446), .B(n380), .Z(n445) );
  NAND U1492 ( .A(rst), .B(\_MxM/Y0[22] ), .Z(n444) );
  NAND U1493 ( .A(n447), .B(n448), .Z(\_MxM/n339 ) );
  NAND U1494 ( .A(n449), .B(n380), .Z(n448) );
  NAND U1495 ( .A(rst), .B(\_MxM/Y0[23] ), .Z(n447) );
  NAND U1496 ( .A(n450), .B(n451), .Z(\_MxM/n338 ) );
  NAND U1497 ( .A(n452), .B(n380), .Z(n451) );
  NAND U1498 ( .A(rst), .B(\_MxM/Y0[24] ), .Z(n450) );
  NAND U1499 ( .A(n453), .B(n454), .Z(\_MxM/n337 ) );
  NAND U1500 ( .A(n455), .B(n380), .Z(n454) );
  NAND U1501 ( .A(rst), .B(\_MxM/Y0[25] ), .Z(n453) );
  NAND U1502 ( .A(n456), .B(n457), .Z(\_MxM/n336 ) );
  NAND U1503 ( .A(n458), .B(n380), .Z(n457) );
  NAND U1504 ( .A(rst), .B(\_MxM/Y0[26] ), .Z(n456) );
  NAND U1505 ( .A(n459), .B(n460), .Z(\_MxM/n335 ) );
  NAND U1506 ( .A(n461), .B(n380), .Z(n460) );
  NAND U1507 ( .A(rst), .B(\_MxM/Y0[27] ), .Z(n459) );
  NAND U1508 ( .A(n462), .B(n463), .Z(\_MxM/n334 ) );
  NAND U1509 ( .A(n464), .B(n380), .Z(n463) );
  NAND U1510 ( .A(rst), .B(\_MxM/Y0[28] ), .Z(n462) );
  NAND U1511 ( .A(n465), .B(n466), .Z(\_MxM/n333 ) );
  NAND U1512 ( .A(n467), .B(n380), .Z(n466) );
  NAND U1513 ( .A(rst), .B(\_MxM/Y0[29] ), .Z(n465) );
  NAND U1514 ( .A(n468), .B(n469), .Z(\_MxM/n332 ) );
  NAND U1515 ( .A(n470), .B(n380), .Z(n469) );
  NAND U1516 ( .A(rst), .B(\_MxM/Y0[30] ), .Z(n468) );
  NAND U1517 ( .A(n471), .B(n472), .Z(\_MxM/n331 ) );
  NAND U1518 ( .A(n473), .B(n380), .Z(n472) );
  NOR U1519 ( .A(rst), .B(n474), .Z(n380) );
  NAND U1520 ( .A(\_MxM/Y0[31] ), .B(rst), .Z(n471) );
  MUX U1521 ( .IN0(o[31]), .IN1(n473), .SEL(n475), .F(\_MxM/n330 ) );
  XNOR U1522 ( .A(\_MxM/Y0[31] ), .B(n477), .Z(n476) );
  AND U1523 ( .A(n480), .B(n481), .Z(n479) );
  XNOR U1524 ( .A(\_MxM/Y0[31] ), .B(n482), .Z(n481) );
  MUX U1525 ( .IN0(o[30]), .IN1(n470), .SEL(n475), .F(\_MxM/n329 ) );
  XOR U1526 ( .A(n480), .B(\_MxM/Y0[31] ), .Z(n470) );
  XOR U1527 ( .A(n482), .B(n477), .Z(n480) );
  XOR U1528 ( .A(n483), .B(n484), .Z(n477) );
  XOR U1529 ( .A(n485), .B(n486), .Z(n484) );
  AND U1530 ( .A(n487), .B(n488), .Z(n486) );
  XOR U1531 ( .A(n495), .B(n493), .Z(n483) );
  XOR U1532 ( .A(n496), .B(n497), .Z(n495) );
  XOR U1533 ( .A(n498), .B(n499), .Z(n497) );
  XOR U1534 ( .A(n503), .B(n504), .Z(n498) );
  ANDN U1535 ( .A(n505), .B(n506), .Z(n504) );
  XOR U1536 ( .A(n510), .B(n511), .Z(n496) );
  XOR U1537 ( .A(n500), .B(n502), .Z(n511) );
  XOR U1538 ( .A(n509), .B(n506), .Z(n510) );
  IV U1539 ( .A(n478), .Z(n482) );
  MUX U1540 ( .IN0(o[29]), .IN1(n467), .SEL(n475), .F(\_MxM/n328 ) );
  XOR U1541 ( .A(n513), .B(\_MxM/Y0[30] ), .Z(n467) );
  XNOR U1542 ( .A(n514), .B(n515), .Z(n513) );
  AND U1543 ( .A(n487), .B(n517), .Z(n516) );
  XNOR U1544 ( .A(n491), .B(n515), .Z(n517) );
  XOR U1545 ( .A(n489), .B(n515), .Z(n491) );
  XNOR U1546 ( .A(n494), .B(n492), .Z(n515) );
  IV U1547 ( .A(n493), .Z(n492) );
  XNOR U1548 ( .A(n500), .B(n501), .Z(n494) );
  XNOR U1549 ( .A(n502), .B(n505), .Z(n501) );
  XNOR U1550 ( .A(n506), .B(n521), .Z(n505) );
  XOR U1551 ( .A(n507), .B(n508), .Z(n521) );
  NAND U1552 ( .A(n522), .B(n523), .Z(n508) );
  IV U1553 ( .A(n509), .Z(n507) );
  IV U1554 ( .A(n490), .Z(n489) );
  MUX U1555 ( .IN0(o[28]), .IN1(n464), .SEL(n475), .F(\_MxM/n327 ) );
  XOR U1556 ( .A(n536), .B(\_MxM/Y0[29] ), .Z(n464) );
  XNOR U1557 ( .A(n537), .B(n538), .Z(n536) );
  AND U1558 ( .A(n487), .B(n540), .Z(n539) );
  XNOR U1559 ( .A(n534), .B(n538), .Z(n540) );
  XNOR U1560 ( .A(n520), .B(n519), .Z(n538) );
  IV U1561 ( .A(n518), .Z(n519) );
  XOR U1562 ( .A(n532), .B(n531), .Z(n520) );
  XOR U1563 ( .A(n530), .B(n544), .Z(n531) );
  XNOR U1564 ( .A(n529), .B(n528), .Z(n544) );
  XNOR U1565 ( .A(n545), .B(n546), .Z(n528) );
  IV U1566 ( .A(n527), .Z(n546) );
  XNOR U1567 ( .A(n525), .B(n526), .Z(n529) );
  NAND U1568 ( .A(n552), .B(n523), .Z(n526) );
  XNOR U1569 ( .A(n524), .B(n553), .Z(n525) );
  ANDN U1570 ( .A(n554), .B(n555), .Z(n553) );
  MUX U1571 ( .IN0(o[27]), .IN1(n461), .SEL(n475), .F(\_MxM/n326 ) );
  XOR U1572 ( .A(n565), .B(\_MxM/Y0[28] ), .Z(n461) );
  XNOR U1573 ( .A(n566), .B(n567), .Z(n565) );
  AND U1574 ( .A(n487), .B(n569), .Z(n568) );
  XNOR U1575 ( .A(n563), .B(n567), .Z(n569) );
  XNOR U1576 ( .A(n543), .B(n542), .Z(n567) );
  IV U1577 ( .A(n541), .Z(n542) );
  XOR U1578 ( .A(n561), .B(n560), .Z(n543) );
  XOR U1579 ( .A(n559), .B(n573), .Z(n560) );
  XNOR U1580 ( .A(n549), .B(n548), .Z(n573) );
  XOR U1581 ( .A(n578), .B(n550), .Z(n574) );
  AND U1582 ( .A(n579), .B(n522), .Z(n550) );
  IV U1583 ( .A(n547), .Z(n578) );
  XNOR U1584 ( .A(n557), .B(n558), .Z(n549) );
  NAND U1585 ( .A(n583), .B(n523), .Z(n558) );
  XNOR U1586 ( .A(n556), .B(n584), .Z(n557) );
  ANDN U1587 ( .A(n554), .B(n585), .Z(n584) );
  MUX U1588 ( .IN0(o[26]), .IN1(n458), .SEL(n475), .F(\_MxM/n325 ) );
  XOR U1589 ( .A(n596), .B(\_MxM/Y0[27] ), .Z(n458) );
  XNOR U1590 ( .A(n597), .B(n598), .Z(n596) );
  AND U1591 ( .A(n487), .B(n600), .Z(n599) );
  XNOR U1592 ( .A(n594), .B(n598), .Z(n600) );
  XNOR U1593 ( .A(n572), .B(n571), .Z(n598) );
  IV U1594 ( .A(n570), .Z(n571) );
  XNOR U1595 ( .A(n592), .B(n604), .Z(n572) );
  XOR U1596 ( .A(n591), .B(n590), .Z(n604) );
  XOR U1597 ( .A(n605), .B(n606), .Z(n590) );
  XOR U1598 ( .A(n607), .B(n608), .Z(n606) );
  XOR U1599 ( .A(n609), .B(n610), .Z(n608) );
  XNOR U1600 ( .A(n582), .B(n581), .Z(n591) );
  XOR U1601 ( .A(n618), .B(n576), .Z(n581) );
  XNOR U1602 ( .A(n575), .B(n619), .Z(n576) );
  ANDN U1603 ( .A(n620), .B(n555), .Z(n619) );
  AND U1604 ( .A(n552), .B(n579), .Z(n577) );
  XNOR U1605 ( .A(n587), .B(n588), .Z(n582) );
  NAND U1606 ( .A(n627), .B(n523), .Z(n588) );
  XNOR U1607 ( .A(n586), .B(n628), .Z(n587) );
  ANDN U1608 ( .A(n554), .B(n629), .Z(n628) );
  MUX U1609 ( .IN0(o[25]), .IN1(n455), .SEL(n475), .F(\_MxM/n324 ) );
  XOR U1610 ( .A(n637), .B(\_MxM/Y0[26] ), .Z(n455) );
  XNOR U1611 ( .A(n638), .B(n639), .Z(n637) );
  AND U1612 ( .A(n487), .B(n641), .Z(n640) );
  XNOR U1613 ( .A(n635), .B(n639), .Z(n641) );
  XNOR U1614 ( .A(n603), .B(n602), .Z(n639) );
  IV U1615 ( .A(n601), .Z(n602) );
  XOR U1616 ( .A(n633), .B(n645), .Z(n603) );
  XNOR U1617 ( .A(n617), .B(n616), .Z(n645) );
  XOR U1618 ( .A(n646), .B(n611), .Z(n616) );
  XOR U1619 ( .A(n612), .B(n613), .Z(n611) );
  NANDN U1620 ( .B(n647), .A(n522), .Z(n613) );
  IV U1621 ( .A(n614), .Z(n612) );
  XOR U1622 ( .A(n607), .B(n615), .Z(n646) );
  XNOR U1623 ( .A(n626), .B(n625), .Z(n617) );
  XOR U1624 ( .A(n657), .B(n622), .Z(n625) );
  XNOR U1625 ( .A(n621), .B(n658), .Z(n622) );
  ANDN U1626 ( .A(n620), .B(n585), .Z(n658) );
  XOR U1627 ( .A(n659), .B(n660), .Z(n621) );
  AND U1628 ( .A(n661), .B(n662), .Z(n660) );
  XNOR U1629 ( .A(n663), .B(n659), .Z(n662) );
  AND U1630 ( .A(n583), .B(n579), .Z(n623) );
  XNOR U1631 ( .A(n631), .B(n632), .Z(n626) );
  NAND U1632 ( .A(n667), .B(n523), .Z(n632) );
  XNOR U1633 ( .A(n630), .B(n668), .Z(n631) );
  ANDN U1634 ( .A(n554), .B(n669), .Z(n668) );
  MUX U1635 ( .IN0(o[24]), .IN1(n452), .SEL(n475), .F(\_MxM/n323 ) );
  XOR U1636 ( .A(n677), .B(\_MxM/Y0[25] ), .Z(n452) );
  XNOR U1637 ( .A(n678), .B(n679), .Z(n677) );
  AND U1638 ( .A(n487), .B(n681), .Z(n680) );
  XNOR U1639 ( .A(n675), .B(n679), .Z(n681) );
  XNOR U1640 ( .A(n644), .B(n643), .Z(n679) );
  IV U1641 ( .A(n642), .Z(n643) );
  XOR U1642 ( .A(n673), .B(n685), .Z(n644) );
  XNOR U1643 ( .A(n653), .B(n652), .Z(n685) );
  XOR U1644 ( .A(n686), .B(n656), .Z(n652) );
  XNOR U1645 ( .A(n649), .B(n650), .Z(n656) );
  NANDN U1646 ( .B(n647), .A(n552), .Z(n650) );
  XNOR U1647 ( .A(n648), .B(n687), .Z(n649) );
  ANDN U1648 ( .A(n688), .B(n555), .Z(n687) );
  XNOR U1649 ( .A(n655), .B(n651), .Z(n686) );
  XNOR U1650 ( .A(n695), .B(n696), .Z(n655) );
  IV U1651 ( .A(n654), .Z(n696) );
  XNOR U1652 ( .A(n666), .B(n665), .Z(n653) );
  XOR U1653 ( .A(n703), .B(n661), .Z(n665) );
  XNOR U1654 ( .A(n659), .B(n704), .Z(n661) );
  ANDN U1655 ( .A(n620), .B(n629), .Z(n704) );
  AND U1656 ( .A(n627), .B(n579), .Z(n663) );
  XNOR U1657 ( .A(n671), .B(n672), .Z(n666) );
  NAND U1658 ( .A(n711), .B(n523), .Z(n672) );
  XNOR U1659 ( .A(n670), .B(n712), .Z(n671) );
  ANDN U1660 ( .A(n554), .B(n713), .Z(n712) );
  MUX U1661 ( .IN0(o[23]), .IN1(n449), .SEL(n475), .F(\_MxM/n322 ) );
  XOR U1662 ( .A(n721), .B(\_MxM/Y0[24] ), .Z(n449) );
  XNOR U1663 ( .A(n722), .B(n723), .Z(n721) );
  AND U1664 ( .A(n487), .B(n725), .Z(n724) );
  XNOR U1665 ( .A(n719), .B(n723), .Z(n725) );
  XNOR U1666 ( .A(n684), .B(n683), .Z(n723) );
  IV U1667 ( .A(n682), .Z(n683) );
  XOR U1668 ( .A(n717), .B(n728), .Z(n684) );
  XNOR U1669 ( .A(n694), .B(n693), .Z(n728) );
  XOR U1670 ( .A(n729), .B(n699), .Z(n693) );
  XNOR U1671 ( .A(n690), .B(n691), .Z(n699) );
  NANDN U1672 ( .B(n647), .A(n583), .Z(n691) );
  XNOR U1673 ( .A(n689), .B(n730), .Z(n690) );
  ANDN U1674 ( .A(n688), .B(n585), .Z(n730) );
  XNOR U1675 ( .A(n698), .B(n692), .Z(n729) );
  XNOR U1676 ( .A(n737), .B(n700), .Z(n698) );
  IV U1677 ( .A(n702), .Z(n700) );
  AND U1678 ( .A(n741), .B(n522), .Z(n701) );
  XNOR U1679 ( .A(n710), .B(n709), .Z(n694) );
  XOR U1680 ( .A(n745), .B(n706), .Z(n709) );
  XNOR U1681 ( .A(n705), .B(n746), .Z(n706) );
  ANDN U1682 ( .A(n620), .B(n669), .Z(n746) );
  AND U1683 ( .A(n667), .B(n579), .Z(n707) );
  XNOR U1684 ( .A(n715), .B(n716), .Z(n710) );
  NAND U1685 ( .A(n753), .B(n523), .Z(n716) );
  XNOR U1686 ( .A(n714), .B(n754), .Z(n715) );
  ANDN U1687 ( .A(n554), .B(n755), .Z(n754) );
  MUX U1688 ( .IN0(o[22]), .IN1(n446), .SEL(n475), .F(\_MxM/n321 ) );
  XOR U1689 ( .A(n765), .B(\_MxM/Y0[23] ), .Z(n446) );
  XNOR U1690 ( .A(n766), .B(n727), .Z(n765) );
  AND U1691 ( .A(n487), .B(n768), .Z(n767) );
  XNOR U1692 ( .A(n763), .B(n727), .Z(n768) );
  XOR U1693 ( .A(n726), .B(n769), .Z(n727) );
  XNOR U1694 ( .A(n761), .B(n760), .Z(n769) );
  XOR U1695 ( .A(n770), .B(n771), .Z(n760) );
  XOR U1696 ( .A(n772), .B(n773), .Z(n771) );
  XOR U1697 ( .A(n776), .B(n777), .Z(n772) );
  ANDN U1698 ( .A(n775), .B(n778), .Z(n777) );
  XNOR U1699 ( .A(n781), .B(n759), .Z(n770) );
  XOR U1700 ( .A(n780), .B(n778), .Z(n781) );
  XNOR U1701 ( .A(n736), .B(n735), .Z(n761) );
  XOR U1702 ( .A(n785), .B(n744), .Z(n735) );
  XNOR U1703 ( .A(n732), .B(n733), .Z(n744) );
  NANDN U1704 ( .B(n647), .A(n627), .Z(n733) );
  XNOR U1705 ( .A(n731), .B(n786), .Z(n732) );
  ANDN U1706 ( .A(n688), .B(n629), .Z(n786) );
  XNOR U1707 ( .A(n743), .B(n734), .Z(n785) );
  XOR U1708 ( .A(n793), .B(n739), .Z(n743) );
  XNOR U1709 ( .A(n738), .B(n794), .Z(n739) );
  ANDN U1710 ( .A(n795), .B(n555), .Z(n794) );
  XOR U1711 ( .A(n796), .B(n797), .Z(n738) );
  AND U1712 ( .A(n798), .B(n799), .Z(n797) );
  XNOR U1713 ( .A(n800), .B(n796), .Z(n799) );
  AND U1714 ( .A(n552), .B(n741), .Z(n740) );
  XNOR U1715 ( .A(n752), .B(n751), .Z(n736) );
  XOR U1716 ( .A(n804), .B(n748), .Z(n751) );
  XNOR U1717 ( .A(n747), .B(n805), .Z(n748) );
  ANDN U1718 ( .A(n620), .B(n713), .Z(n805) );
  AND U1719 ( .A(n711), .B(n579), .Z(n749) );
  XNOR U1720 ( .A(n757), .B(n758), .Z(n752) );
  NAND U1721 ( .A(n812), .B(n523), .Z(n758) );
  XNOR U1722 ( .A(n756), .B(n813), .Z(n757) );
  ANDN U1723 ( .A(n554), .B(n814), .Z(n813) );
  MUX U1724 ( .IN0(o[21]), .IN1(n443), .SEL(n475), .F(\_MxM/n320 ) );
  XOR U1725 ( .A(n824), .B(\_MxM/Y0[22] ), .Z(n443) );
  XNOR U1726 ( .A(n825), .B(n826), .Z(n824) );
  AND U1727 ( .A(n487), .B(n828), .Z(n827) );
  XNOR U1728 ( .A(n822), .B(n826), .Z(n828) );
  XNOR U1729 ( .A(n820), .B(n819), .Z(n826) );
  IV U1730 ( .A(n818), .Z(n819) );
  XNOR U1731 ( .A(n784), .B(n783), .Z(n820) );
  XOR U1732 ( .A(n832), .B(n775), .Z(n783) );
  XNOR U1733 ( .A(n778), .B(n833), .Z(n775) );
  NANDN U1734 ( .B(n834), .A(n522), .Z(n779) );
  XOR U1735 ( .A(n774), .B(n782), .Z(n832) );
  XNOR U1736 ( .A(n792), .B(n791), .Z(n784) );
  XOR U1737 ( .A(n846), .B(n803), .Z(n791) );
  XNOR U1738 ( .A(n788), .B(n789), .Z(n803) );
  NANDN U1739 ( .B(n647), .A(n667), .Z(n789) );
  XNOR U1740 ( .A(n787), .B(n847), .Z(n788) );
  ANDN U1741 ( .A(n688), .B(n669), .Z(n847) );
  XOR U1742 ( .A(n848), .B(n849), .Z(n787) );
  AND U1743 ( .A(n850), .B(n851), .Z(n849) );
  XOR U1744 ( .A(n852), .B(n848), .Z(n851) );
  XNOR U1745 ( .A(n802), .B(n790), .Z(n846) );
  XOR U1746 ( .A(n856), .B(n798), .Z(n802) );
  XNOR U1747 ( .A(n796), .B(n857), .Z(n798) );
  ANDN U1748 ( .A(n795), .B(n585), .Z(n857) );
  XOR U1749 ( .A(n858), .B(n859), .Z(n796) );
  AND U1750 ( .A(n860), .B(n861), .Z(n859) );
  XNOR U1751 ( .A(n862), .B(n858), .Z(n861) );
  AND U1752 ( .A(n583), .B(n741), .Z(n800) );
  XNOR U1753 ( .A(n811), .B(n810), .Z(n792) );
  XOR U1754 ( .A(n866), .B(n807), .Z(n810) );
  XNOR U1755 ( .A(n806), .B(n867), .Z(n807) );
  ANDN U1756 ( .A(n620), .B(n755), .Z(n867) );
  XOR U1757 ( .A(n868), .B(n869), .Z(n806) );
  AND U1758 ( .A(n870), .B(n871), .Z(n869) );
  XNOR U1759 ( .A(n872), .B(n868), .Z(n871) );
  AND U1760 ( .A(n753), .B(n579), .Z(n808) );
  XNOR U1761 ( .A(n816), .B(n817), .Z(n811) );
  NAND U1762 ( .A(n876), .B(n523), .Z(n817) );
  XNOR U1763 ( .A(n815), .B(n877), .Z(n816) );
  ANDN U1764 ( .A(n554), .B(n878), .Z(n877) );
  XOR U1765 ( .A(n879), .B(n880), .Z(n815) );
  AND U1766 ( .A(n881), .B(n882), .Z(n880) );
  XOR U1767 ( .A(n883), .B(n879), .Z(n882) );
  MUX U1768 ( .IN0(o[20]), .IN1(n440), .SEL(n475), .F(\_MxM/n319 ) );
  XOR U1769 ( .A(n887), .B(\_MxM/Y0[21] ), .Z(n440) );
  XNOR U1770 ( .A(n888), .B(n889), .Z(n887) );
  AND U1771 ( .A(n487), .B(n891), .Z(n890) );
  XNOR U1772 ( .A(n885), .B(n889), .Z(n891) );
  XNOR U1773 ( .A(n831), .B(n830), .Z(n889) );
  IV U1774 ( .A(n829), .Z(n830) );
  XNOR U1775 ( .A(n843), .B(n842), .Z(n831) );
  XOR U1776 ( .A(n895), .B(n845), .Z(n842) );
  XNOR U1777 ( .A(n840), .B(n839), .Z(n845) );
  XNOR U1778 ( .A(n896), .B(n897), .Z(n839) );
  IV U1779 ( .A(n838), .Z(n897) );
  XNOR U1780 ( .A(n836), .B(n837), .Z(n840) );
  NANDN U1781 ( .B(n834), .A(n552), .Z(n837) );
  XNOR U1782 ( .A(n835), .B(n903), .Z(n836) );
  ANDN U1783 ( .A(n904), .B(n555), .Z(n903) );
  XNOR U1784 ( .A(n855), .B(n854), .Z(n843) );
  XOR U1785 ( .A(n914), .B(n865), .Z(n854) );
  XNOR U1786 ( .A(n850), .B(n852), .Z(n865) );
  NANDN U1787 ( .B(n647), .A(n711), .Z(n852) );
  XNOR U1788 ( .A(n848), .B(n915), .Z(n850) );
  ANDN U1789 ( .A(n688), .B(n713), .Z(n915) );
  XOR U1790 ( .A(n916), .B(n917), .Z(n848) );
  AND U1791 ( .A(n918), .B(n919), .Z(n917) );
  XOR U1792 ( .A(n920), .B(n916), .Z(n919) );
  XNOR U1793 ( .A(n864), .B(n853), .Z(n914) );
  XOR U1794 ( .A(n924), .B(n860), .Z(n864) );
  XNOR U1795 ( .A(n858), .B(n925), .Z(n860) );
  ANDN U1796 ( .A(n795), .B(n629), .Z(n925) );
  XOR U1797 ( .A(n926), .B(n927), .Z(n858) );
  AND U1798 ( .A(n928), .B(n929), .Z(n927) );
  XNOR U1799 ( .A(n930), .B(n926), .Z(n929) );
  AND U1800 ( .A(n627), .B(n741), .Z(n862) );
  XNOR U1801 ( .A(n875), .B(n874), .Z(n855) );
  XOR U1802 ( .A(n934), .B(n870), .Z(n874) );
  XNOR U1803 ( .A(n868), .B(n935), .Z(n870) );
  ANDN U1804 ( .A(n620), .B(n814), .Z(n935) );
  XOR U1805 ( .A(n936), .B(n937), .Z(n868) );
  AND U1806 ( .A(n938), .B(n939), .Z(n937) );
  XNOR U1807 ( .A(n940), .B(n936), .Z(n939) );
  AND U1808 ( .A(n812), .B(n579), .Z(n872) );
  XNOR U1809 ( .A(n881), .B(n883), .Z(n875) );
  NAND U1810 ( .A(n944), .B(n523), .Z(n883) );
  XNOR U1811 ( .A(n879), .B(n945), .Z(n881) );
  ANDN U1812 ( .A(n554), .B(n946), .Z(n945) );
  XOR U1813 ( .A(n947), .B(n948), .Z(n879) );
  AND U1814 ( .A(n949), .B(n950), .Z(n948) );
  XOR U1815 ( .A(n951), .B(n947), .Z(n950) );
  MUX U1816 ( .IN0(o[19]), .IN1(n437), .SEL(n475), .F(\_MxM/n318 ) );
  XOR U1817 ( .A(n955), .B(\_MxM/Y0[20] ), .Z(n437) );
  XNOR U1818 ( .A(n956), .B(n957), .Z(n955) );
  AND U1819 ( .A(n487), .B(n959), .Z(n958) );
  XNOR U1820 ( .A(n953), .B(n957), .Z(n959) );
  XNOR U1821 ( .A(n894), .B(n893), .Z(n957) );
  IV U1822 ( .A(n892), .Z(n893) );
  XNOR U1823 ( .A(n910), .B(n909), .Z(n894) );
  XOR U1824 ( .A(n963), .B(n913), .Z(n909) );
  XNOR U1825 ( .A(n900), .B(n899), .Z(n913) );
  XOR U1826 ( .A(n968), .B(n901), .Z(n964) );
  AND U1827 ( .A(n969), .B(n522), .Z(n901) );
  IV U1828 ( .A(n898), .Z(n968) );
  XNOR U1829 ( .A(n906), .B(n907), .Z(n900) );
  NANDN U1830 ( .B(n834), .A(n583), .Z(n907) );
  XNOR U1831 ( .A(n905), .B(n973), .Z(n906) );
  ANDN U1832 ( .A(n904), .B(n585), .Z(n973) );
  XNOR U1833 ( .A(n912), .B(n908), .Z(n963) );
  IV U1834 ( .A(n911), .Z(n912) );
  XNOR U1835 ( .A(n923), .B(n922), .Z(n910) );
  XOR U1836 ( .A(n983), .B(n933), .Z(n922) );
  XNOR U1837 ( .A(n918), .B(n920), .Z(n933) );
  NANDN U1838 ( .B(n647), .A(n753), .Z(n920) );
  XNOR U1839 ( .A(n916), .B(n984), .Z(n918) );
  ANDN U1840 ( .A(n688), .B(n755), .Z(n984) );
  XOR U1841 ( .A(n985), .B(n986), .Z(n916) );
  AND U1842 ( .A(n987), .B(n988), .Z(n986) );
  XOR U1843 ( .A(n989), .B(n985), .Z(n988) );
  XNOR U1844 ( .A(n932), .B(n921), .Z(n983) );
  XOR U1845 ( .A(n993), .B(n928), .Z(n932) );
  XNOR U1846 ( .A(n926), .B(n994), .Z(n928) );
  ANDN U1847 ( .A(n795), .B(n669), .Z(n994) );
  XOR U1848 ( .A(n995), .B(n996), .Z(n926) );
  AND U1849 ( .A(n997), .B(n998), .Z(n996) );
  XNOR U1850 ( .A(n999), .B(n995), .Z(n998) );
  AND U1851 ( .A(n667), .B(n741), .Z(n930) );
  XNOR U1852 ( .A(n943), .B(n942), .Z(n923) );
  XOR U1853 ( .A(n1003), .B(n938), .Z(n942) );
  XNOR U1854 ( .A(n936), .B(n1004), .Z(n938) );
  ANDN U1855 ( .A(n620), .B(n878), .Z(n1004) );
  AND U1856 ( .A(n876), .B(n579), .Z(n940) );
  XNOR U1857 ( .A(n949), .B(n951), .Z(n943) );
  NAND U1858 ( .A(n1011), .B(n523), .Z(n951) );
  XNOR U1859 ( .A(n947), .B(n1012), .Z(n949) );
  ANDN U1860 ( .A(n554), .B(n1013), .Z(n1012) );
  XOR U1861 ( .A(n1014), .B(n1015), .Z(n947) );
  AND U1862 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR U1863 ( .A(n1018), .B(n1014), .Z(n1017) );
  MUX U1864 ( .IN0(o[18]), .IN1(n434), .SEL(n475), .F(\_MxM/n317 ) );
  XOR U1865 ( .A(n1022), .B(\_MxM/Y0[19] ), .Z(n434) );
  XNOR U1866 ( .A(n1023), .B(n1024), .Z(n1022) );
  AND U1867 ( .A(n487), .B(n1026), .Z(n1025) );
  XOR U1868 ( .A(n1020), .B(n1024), .Z(n1026) );
  XOR U1869 ( .A(n1019), .B(n1024), .Z(n1020) );
  XNOR U1870 ( .A(n962), .B(n961), .Z(n1024) );
  IV U1871 ( .A(n960), .Z(n961) );
  XNOR U1872 ( .A(n979), .B(n978), .Z(n962) );
  XOR U1873 ( .A(n1029), .B(n982), .Z(n978) );
  XNOR U1874 ( .A(n972), .B(n971), .Z(n982) );
  XOR U1875 ( .A(n1030), .B(n966), .Z(n971) );
  XNOR U1876 ( .A(n965), .B(n1031), .Z(n966) );
  ANDN U1877 ( .A(n1032), .B(n555), .Z(n1031) );
  XOR U1878 ( .A(n1033), .B(n1034), .Z(n965) );
  AND U1879 ( .A(n1035), .B(n1036), .Z(n1034) );
  XNOR U1880 ( .A(n1037), .B(n1033), .Z(n1036) );
  AND U1881 ( .A(n552), .B(n969), .Z(n967) );
  XNOR U1882 ( .A(n975), .B(n976), .Z(n972) );
  NANDN U1883 ( .B(n834), .A(n627), .Z(n976) );
  XNOR U1884 ( .A(n974), .B(n1041), .Z(n975) );
  ANDN U1885 ( .A(n904), .B(n629), .Z(n1041) );
  XNOR U1886 ( .A(n981), .B(n977), .Z(n1029) );
  XNOR U1887 ( .A(n1048), .B(n1049), .Z(n981) );
  IV U1888 ( .A(n980), .Z(n1049) );
  XNOR U1889 ( .A(n992), .B(n991), .Z(n979) );
  XOR U1890 ( .A(n1055), .B(n1002), .Z(n991) );
  XNOR U1891 ( .A(n987), .B(n989), .Z(n1002) );
  NANDN U1892 ( .B(n647), .A(n812), .Z(n989) );
  XNOR U1893 ( .A(n985), .B(n1056), .Z(n987) );
  ANDN U1894 ( .A(n688), .B(n814), .Z(n1056) );
  XOR U1895 ( .A(n1057), .B(n1058), .Z(n985) );
  AND U1896 ( .A(n1059), .B(n1060), .Z(n1058) );
  XOR U1897 ( .A(n1061), .B(n1057), .Z(n1060) );
  XNOR U1898 ( .A(n1001), .B(n990), .Z(n1055) );
  XOR U1899 ( .A(n1065), .B(n997), .Z(n1001) );
  XNOR U1900 ( .A(n995), .B(n1066), .Z(n997) );
  ANDN U1901 ( .A(n795), .B(n713), .Z(n1066) );
  XOR U1902 ( .A(n1067), .B(n1068), .Z(n995) );
  AND U1903 ( .A(n1069), .B(n1070), .Z(n1068) );
  XNOR U1904 ( .A(n1071), .B(n1067), .Z(n1070) );
  AND U1905 ( .A(n711), .B(n741), .Z(n999) );
  XNOR U1906 ( .A(n1010), .B(n1009), .Z(n992) );
  XOR U1907 ( .A(n1075), .B(n1006), .Z(n1009) );
  XNOR U1908 ( .A(n1005), .B(n1076), .Z(n1006) );
  ANDN U1909 ( .A(n620), .B(n946), .Z(n1076) );
  XOR U1910 ( .A(n1077), .B(n1078), .Z(n1005) );
  AND U1911 ( .A(n1079), .B(n1080), .Z(n1078) );
  XNOR U1912 ( .A(n1081), .B(n1077), .Z(n1080) );
  AND U1913 ( .A(n944), .B(n579), .Z(n1007) );
  XNOR U1914 ( .A(n1016), .B(n1018), .Z(n1010) );
  NAND U1915 ( .A(n1085), .B(n523), .Z(n1018) );
  XNOR U1916 ( .A(n1014), .B(n1086), .Z(n1016) );
  ANDN U1917 ( .A(n554), .B(n1087), .Z(n1086) );
  NANDN U1918 ( .B(n1088), .A(n1089), .Z(n1014) );
  NAND U1919 ( .A(n1090), .B(n1091), .Z(n1089) );
  MUX U1920 ( .IN0(o[17]), .IN1(n431), .SEL(n475), .F(\_MxM/n316 ) );
  XOR U1921 ( .A(n1096), .B(\_MxM/Y0[18] ), .Z(n431) );
  XOR U1922 ( .A(n1097), .B(n1098), .Z(n1096) );
  AND U1923 ( .A(n487), .B(n1100), .Z(n1099) );
  XOR U1924 ( .A(n1094), .B(n1098), .Z(n1100) );
  XOR U1925 ( .A(n1093), .B(n1098), .Z(n1094) );
  XOR U1926 ( .A(n1028), .B(n1027), .Z(n1098) );
  XNOR U1927 ( .A(n1103), .B(n1052), .Z(n1046) );
  XNOR U1928 ( .A(n1040), .B(n1039), .Z(n1052) );
  XOR U1929 ( .A(n1104), .B(n1035), .Z(n1039) );
  XNOR U1930 ( .A(n1033), .B(n1105), .Z(n1035) );
  ANDN U1931 ( .A(n1032), .B(n585), .Z(n1105) );
  XOR U1932 ( .A(n1106), .B(n1107), .Z(n1033) );
  AND U1933 ( .A(n1108), .B(n1109), .Z(n1107) );
  XNOR U1934 ( .A(n1110), .B(n1106), .Z(n1109) );
  AND U1935 ( .A(n583), .B(n969), .Z(n1037) );
  XNOR U1936 ( .A(n1043), .B(n1044), .Z(n1040) );
  NANDN U1937 ( .B(n834), .A(n667), .Z(n1044) );
  XNOR U1938 ( .A(n1042), .B(n1114), .Z(n1043) );
  ANDN U1939 ( .A(n904), .B(n669), .Z(n1114) );
  XOR U1940 ( .A(n1115), .B(n1116), .Z(n1042) );
  AND U1941 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U1942 ( .A(n1119), .B(n1115), .Z(n1118) );
  XNOR U1943 ( .A(n1051), .B(n1045), .Z(n1103) );
  XOR U1944 ( .A(n1123), .B(n1053), .Z(n1051) );
  NAND U1945 ( .A(n1127), .B(n1128), .Z(n1054) );
  NANDN U1946 ( .B(n1129), .A(n522), .Z(n1128) );
  NANDN U1947 ( .B(n1130), .A(n1131), .Z(n1127) );
  XNOR U1948 ( .A(n1064), .B(n1063), .Z(n1047) );
  XOR U1949 ( .A(n1135), .B(n1074), .Z(n1063) );
  XNOR U1950 ( .A(n1059), .B(n1061), .Z(n1074) );
  NANDN U1951 ( .B(n647), .A(n876), .Z(n1061) );
  XNOR U1952 ( .A(n1057), .B(n1136), .Z(n1059) );
  ANDN U1953 ( .A(n688), .B(n878), .Z(n1136) );
  XOR U1954 ( .A(n1137), .B(n1138), .Z(n1057) );
  AND U1955 ( .A(n1139), .B(n1140), .Z(n1138) );
  XOR U1956 ( .A(n1141), .B(n1137), .Z(n1140) );
  XNOR U1957 ( .A(n1073), .B(n1062), .Z(n1135) );
  XOR U1958 ( .A(n1145), .B(n1069), .Z(n1073) );
  XNOR U1959 ( .A(n1067), .B(n1146), .Z(n1069) );
  ANDN U1960 ( .A(n795), .B(n755), .Z(n1146) );
  XOR U1961 ( .A(n1147), .B(n1148), .Z(n1067) );
  AND U1962 ( .A(n1149), .B(n1150), .Z(n1148) );
  XNOR U1963 ( .A(n1151), .B(n1147), .Z(n1150) );
  AND U1964 ( .A(n753), .B(n741), .Z(n1071) );
  XOR U1965 ( .A(n1084), .B(n1083), .Z(n1064) );
  XOR U1966 ( .A(n1155), .B(n1079), .Z(n1083) );
  XNOR U1967 ( .A(n1077), .B(n1156), .Z(n1079) );
  ANDN U1968 ( .A(n620), .B(n1013), .Z(n1156) );
  AND U1969 ( .A(n1011), .B(n579), .Z(n1081) );
  XOR U1970 ( .A(n1091), .B(n1090), .Z(n1084) );
  NAND U1971 ( .A(n1163), .B(n523), .Z(n1090) );
  XNOR U1972 ( .A(n1088), .B(n1164), .Z(n1091) );
  ANDN U1973 ( .A(n554), .B(n1165), .Z(n1164) );
  NANDN U1974 ( .B(n1166), .A(n1167), .Z(n1088) );
  NAND U1975 ( .A(n1168), .B(n1169), .Z(n1167) );
  IV U1976 ( .A(n1092), .Z(n1093) );
  MUX U1977 ( .IN0(o[16]), .IN1(n428), .SEL(n475), .F(\_MxM/n315 ) );
  XOR U1978 ( .A(n1174), .B(\_MxM/Y0[17] ), .Z(n428) );
  XOR U1979 ( .A(n1175), .B(n1176), .Z(n1174) );
  AND U1980 ( .A(n487), .B(n1178), .Z(n1177) );
  XOR U1981 ( .A(n1172), .B(n1176), .Z(n1178) );
  XOR U1982 ( .A(n1171), .B(n1176), .Z(n1172) );
  XOR U1983 ( .A(n1102), .B(n1101), .Z(n1176) );
  XNOR U1984 ( .A(n1181), .B(n1134), .Z(n1121) );
  XNOR U1985 ( .A(n1113), .B(n1112), .Z(n1134) );
  XOR U1986 ( .A(n1182), .B(n1108), .Z(n1112) );
  XNOR U1987 ( .A(n1106), .B(n1183), .Z(n1108) );
  ANDN U1988 ( .A(n1032), .B(n629), .Z(n1183) );
  XOR U1989 ( .A(n1184), .B(n1185), .Z(n1106) );
  AND U1990 ( .A(n1186), .B(n1187), .Z(n1185) );
  XNOR U1991 ( .A(n1188), .B(n1184), .Z(n1187) );
  AND U1992 ( .A(n627), .B(n969), .Z(n1110) );
  XNOR U1993 ( .A(n1117), .B(n1119), .Z(n1113) );
  NANDN U1994 ( .B(n834), .A(n711), .Z(n1119) );
  XNOR U1995 ( .A(n1115), .B(n1192), .Z(n1117) );
  ANDN U1996 ( .A(n904), .B(n713), .Z(n1192) );
  XOR U1997 ( .A(n1193), .B(n1194), .Z(n1115) );
  AND U1998 ( .A(n1195), .B(n1196), .Z(n1194) );
  XOR U1999 ( .A(n1197), .B(n1193), .Z(n1196) );
  XOR U2000 ( .A(n1133), .B(n1120), .Z(n1181) );
  XNOR U2001 ( .A(n1201), .B(n1125), .Z(n1133) );
  XNOR U2002 ( .A(n1202), .B(n1131), .Z(n1125) );
  AND U2003 ( .A(n552), .B(n1203), .Z(n1131) );
  NAND U2004 ( .A(n1204), .B(n1130), .Z(n1202) );
  XOR U2005 ( .A(n1205), .B(n1206), .Z(n1130) );
  AND U2006 ( .A(n1207), .B(n1208), .Z(n1206) );
  XOR U2007 ( .A(n1209), .B(n1205), .Z(n1208) );
  NANDN U2008 ( .B(n555), .A(n1210), .Z(n1204) );
  XNOR U2009 ( .A(n1124), .B(n1132), .Z(n1201) );
  IV U2010 ( .A(n1126), .Z(n1124) );
  XNOR U2011 ( .A(n1144), .B(n1143), .Z(n1122) );
  XOR U2012 ( .A(n1216), .B(n1154), .Z(n1143) );
  XNOR U2013 ( .A(n1139), .B(n1141), .Z(n1154) );
  NANDN U2014 ( .B(n647), .A(n944), .Z(n1141) );
  XNOR U2015 ( .A(n1137), .B(n1217), .Z(n1139) );
  ANDN U2016 ( .A(n688), .B(n946), .Z(n1217) );
  XNOR U2017 ( .A(n1153), .B(n1142), .Z(n1216) );
  XOR U2018 ( .A(n1224), .B(n1149), .Z(n1153) );
  XNOR U2019 ( .A(n1147), .B(n1225), .Z(n1149) );
  ANDN U2020 ( .A(n795), .B(n814), .Z(n1225) );
  XOR U2021 ( .A(n1226), .B(n1227), .Z(n1147) );
  AND U2022 ( .A(n1228), .B(n1229), .Z(n1227) );
  XNOR U2023 ( .A(n1230), .B(n1226), .Z(n1229) );
  AND U2024 ( .A(n812), .B(n741), .Z(n1151) );
  XOR U2025 ( .A(n1162), .B(n1161), .Z(n1144) );
  XOR U2026 ( .A(n1234), .B(n1158), .Z(n1161) );
  XNOR U2027 ( .A(n1157), .B(n1235), .Z(n1158) );
  ANDN U2028 ( .A(n620), .B(n1087), .Z(n1235) );
  XOR U2029 ( .A(n1236), .B(n1237), .Z(n1157) );
  AND U2030 ( .A(n1238), .B(n1239), .Z(n1237) );
  XNOR U2031 ( .A(n1240), .B(n1236), .Z(n1239) );
  AND U2032 ( .A(n1085), .B(n579), .Z(n1159) );
  XOR U2033 ( .A(n1169), .B(n1168), .Z(n1162) );
  NAND U2034 ( .A(n1244), .B(n523), .Z(n1168) );
  XNOR U2035 ( .A(n1166), .B(n1245), .Z(n1169) );
  ANDN U2036 ( .A(n554), .B(n1246), .Z(n1245) );
  NAND U2037 ( .A(n1247), .B(n1248), .Z(n1166) );
  NAND U2038 ( .A(n1249), .B(n1250), .Z(n1247) );
  IV U2039 ( .A(n1170), .Z(n1171) );
  MUX U2040 ( .IN0(o[15]), .IN1(n425), .SEL(n475), .F(\_MxM/n314 ) );
  XOR U2041 ( .A(n1255), .B(\_MxM/Y0[16] ), .Z(n425) );
  XOR U2042 ( .A(n1256), .B(n1257), .Z(n1255) );
  AND U2043 ( .A(n487), .B(n1259), .Z(n1258) );
  XOR U2044 ( .A(n1253), .B(n1257), .Z(n1259) );
  XOR U2045 ( .A(n1252), .B(n1257), .Z(n1253) );
  XOR U2046 ( .A(n1180), .B(n1179), .Z(n1257) );
  XNOR U2047 ( .A(n1263), .B(n1213), .Z(n1199) );
  XNOR U2048 ( .A(n1191), .B(n1190), .Z(n1213) );
  XOR U2049 ( .A(n1264), .B(n1186), .Z(n1190) );
  XNOR U2050 ( .A(n1184), .B(n1265), .Z(n1186) );
  ANDN U2051 ( .A(n1032), .B(n669), .Z(n1265) );
  XOR U2052 ( .A(n1266), .B(n1267), .Z(n1184) );
  AND U2053 ( .A(n1268), .B(n1269), .Z(n1267) );
  XNOR U2054 ( .A(n1270), .B(n1266), .Z(n1269) );
  AND U2055 ( .A(n667), .B(n969), .Z(n1188) );
  XNOR U2056 ( .A(n1195), .B(n1197), .Z(n1191) );
  NANDN U2057 ( .B(n834), .A(n753), .Z(n1197) );
  XNOR U2058 ( .A(n1193), .B(n1274), .Z(n1195) );
  ANDN U2059 ( .A(n904), .B(n755), .Z(n1274) );
  XNOR U2060 ( .A(n1212), .B(n1198), .Z(n1263) );
  XOR U2061 ( .A(n1281), .B(n1215), .Z(n1212) );
  XNOR U2062 ( .A(n1207), .B(n1209), .Z(n1215) );
  NAND U2063 ( .A(n583), .B(n1203), .Z(n1209) );
  XNOR U2064 ( .A(n1205), .B(n1282), .Z(n1207) );
  ANDN U2065 ( .A(n1210), .B(n585), .Z(n1282) );
  XOR U2066 ( .A(n1283), .B(n1284), .Z(n1205) );
  AND U2067 ( .A(n1285), .B(n1286), .Z(n1284) );
  XOR U2068 ( .A(n1287), .B(n1283), .Z(n1286) );
  XNOR U2069 ( .A(n1214), .B(n1211), .Z(n1281) );
  AND U2070 ( .A(n1292), .B(n1293), .Z(n1291) );
  NANDN U2071 ( .B(n1294), .A(n522), .Z(n1293) );
  NANDN U2072 ( .B(n1295), .A(n1296), .Z(n1292) );
  XNOR U2073 ( .A(n1223), .B(n1222), .Z(n1200) );
  XOR U2074 ( .A(n1300), .B(n1233), .Z(n1222) );
  XNOR U2075 ( .A(n1219), .B(n1220), .Z(n1233) );
  NANDN U2076 ( .B(n647), .A(n1011), .Z(n1220) );
  XNOR U2077 ( .A(n1218), .B(n1301), .Z(n1219) );
  ANDN U2078 ( .A(n688), .B(n1013), .Z(n1301) );
  XNOR U2079 ( .A(n1232), .B(n1221), .Z(n1300) );
  XOR U2080 ( .A(n1308), .B(n1228), .Z(n1232) );
  XNOR U2081 ( .A(n1226), .B(n1309), .Z(n1228) );
  ANDN U2082 ( .A(n795), .B(n878), .Z(n1309) );
  XOR U2083 ( .A(n1310), .B(n1311), .Z(n1226) );
  AND U2084 ( .A(n1312), .B(n1313), .Z(n1311) );
  XNOR U2085 ( .A(n1314), .B(n1310), .Z(n1313) );
  AND U2086 ( .A(n876), .B(n741), .Z(n1230) );
  XOR U2087 ( .A(n1243), .B(n1242), .Z(n1223) );
  XOR U2088 ( .A(n1318), .B(n1238), .Z(n1242) );
  XNOR U2089 ( .A(n1236), .B(n1319), .Z(n1238) );
  ANDN U2090 ( .A(n620), .B(n1165), .Z(n1319) );
  XOR U2091 ( .A(n1320), .B(n1321), .Z(n1236) );
  AND U2092 ( .A(n1322), .B(n1323), .Z(n1321) );
  XNOR U2093 ( .A(n1324), .B(n1320), .Z(n1323) );
  AND U2094 ( .A(n1163), .B(n579), .Z(n1240) );
  XOR U2095 ( .A(n1250), .B(n1249), .Z(n1243) );
  NAND U2096 ( .A(n1328), .B(n523), .Z(n1249) );
  XOR U2097 ( .A(n1248), .B(n1329), .Z(n1250) );
  ANDN U2098 ( .A(n554), .B(n1330), .Z(n1329) );
  ANDN U2099 ( .A(n1331), .B(n1332), .Z(n1248) );
  NAND U2100 ( .A(n1333), .B(n1334), .Z(n1331) );
  IV U2101 ( .A(n1251), .Z(n1252) );
  MUX U2102 ( .IN0(o[14]), .IN1(n422), .SEL(n475), .F(\_MxM/n313 ) );
  XOR U2103 ( .A(n1339), .B(\_MxM/Y0[15] ), .Z(n422) );
  XOR U2104 ( .A(n1340), .B(n1341), .Z(n1339) );
  AND U2105 ( .A(n487), .B(n1343), .Z(n1342) );
  XOR U2106 ( .A(n1337), .B(n1341), .Z(n1343) );
  XOR U2107 ( .A(n1336), .B(n1341), .Z(n1337) );
  XNOR U2108 ( .A(n1262), .B(n1261), .Z(n1341) );
  XOR U2109 ( .A(n1344), .B(n1345), .Z(n1261) );
  XOR U2110 ( .A(n1346), .B(n1347), .Z(n1345) );
  XOR U2111 ( .A(n1348), .B(n1346), .Z(n1347) );
  XNOR U2112 ( .A(n1354), .B(n1290), .Z(n1279) );
  XNOR U2113 ( .A(n1273), .B(n1272), .Z(n1290) );
  XOR U2114 ( .A(n1355), .B(n1268), .Z(n1272) );
  XNOR U2115 ( .A(n1266), .B(n1356), .Z(n1268) );
  ANDN U2116 ( .A(n1032), .B(n713), .Z(n1356) );
  AND U2117 ( .A(n711), .B(n969), .Z(n1270) );
  XNOR U2118 ( .A(n1276), .B(n1277), .Z(n1273) );
  NANDN U2119 ( .B(n834), .A(n812), .Z(n1277) );
  XNOR U2120 ( .A(n1275), .B(n1363), .Z(n1276) );
  ANDN U2121 ( .A(n904), .B(n814), .Z(n1363) );
  XOR U2122 ( .A(n1364), .B(n1365), .Z(n1275) );
  AND U2123 ( .A(n1366), .B(n1367), .Z(n1365) );
  XOR U2124 ( .A(n1368), .B(n1364), .Z(n1367) );
  XNOR U2125 ( .A(n1289), .B(n1278), .Z(n1354) );
  XOR U2126 ( .A(n1372), .B(n1299), .Z(n1289) );
  XNOR U2127 ( .A(n1285), .B(n1287), .Z(n1299) );
  NAND U2128 ( .A(n627), .B(n1203), .Z(n1287) );
  XNOR U2129 ( .A(n1283), .B(n1373), .Z(n1285) );
  ANDN U2130 ( .A(n1210), .B(n629), .Z(n1373) );
  XOR U2131 ( .A(n1374), .B(n1375), .Z(n1283) );
  AND U2132 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR U2133 ( .A(n1378), .B(n1374), .Z(n1377) );
  XNOR U2134 ( .A(n1298), .B(n1288), .Z(n1372) );
  XOR U2135 ( .A(n1386), .B(n1296), .Z(n1382) );
  AND U2136 ( .A(n552), .B(n1387), .Z(n1296) );
  NAND U2137 ( .A(n1388), .B(n1295), .Z(n1386) );
  XOR U2138 ( .A(n1389), .B(n1390), .Z(n1295) );
  AND U2139 ( .A(n1391), .B(n1392), .Z(n1390) );
  XNOR U2140 ( .A(n1393), .B(n1389), .Z(n1392) );
  NANDN U2141 ( .B(n555), .A(n1394), .Z(n1388) );
  XNOR U2142 ( .A(n1307), .B(n1306), .Z(n1280) );
  XOR U2143 ( .A(n1395), .B(n1317), .Z(n1306) );
  XNOR U2144 ( .A(n1303), .B(n1304), .Z(n1317) );
  NANDN U2145 ( .B(n647), .A(n1085), .Z(n1304) );
  XNOR U2146 ( .A(n1302), .B(n1396), .Z(n1303) );
  ANDN U2147 ( .A(n688), .B(n1087), .Z(n1396) );
  XNOR U2148 ( .A(n1316), .B(n1305), .Z(n1395) );
  XOR U2149 ( .A(n1403), .B(n1312), .Z(n1316) );
  XNOR U2150 ( .A(n1310), .B(n1404), .Z(n1312) );
  ANDN U2151 ( .A(n795), .B(n946), .Z(n1404) );
  AND U2152 ( .A(n944), .B(n741), .Z(n1314) );
  XOR U2153 ( .A(n1327), .B(n1326), .Z(n1307) );
  XOR U2154 ( .A(n1411), .B(n1322), .Z(n1326) );
  XNOR U2155 ( .A(n1320), .B(n1412), .Z(n1322) );
  ANDN U2156 ( .A(n620), .B(n1246), .Z(n1412) );
  AND U2157 ( .A(n1244), .B(n579), .Z(n1324) );
  XOR U2158 ( .A(n1334), .B(n1333), .Z(n1327) );
  NAND U2159 ( .A(n1419), .B(n523), .Z(n1333) );
  XNOR U2160 ( .A(n1332), .B(n1420), .Z(n1334) );
  ANDN U2161 ( .A(n554), .B(n1421), .Z(n1420) );
  NAND U2162 ( .A(n1422), .B(n1423), .Z(n1332) );
  NAND U2163 ( .A(n1424), .B(n1425), .Z(n1422) );
  IV U2164 ( .A(n1335), .Z(n1336) );
  MUX U2165 ( .IN0(o[13]), .IN1(n419), .SEL(n475), .F(\_MxM/n312 ) );
  XOR U2166 ( .A(n1430), .B(\_MxM/Y0[14] ), .Z(n419) );
  XOR U2167 ( .A(n1431), .B(n1432), .Z(n1430) );
  AND U2168 ( .A(n487), .B(n1434), .Z(n1433) );
  XOR U2169 ( .A(n1428), .B(n1432), .Z(n1434) );
  XOR U2170 ( .A(n1427), .B(n1432), .Z(n1428) );
  XOR U2171 ( .A(n1435), .B(n1349), .Z(n1352) );
  NAND U2172 ( .A(n1346), .B(n1439), .Z(n1350) );
  AND U2173 ( .A(n1440), .B(n1441), .Z(n1439) );
  NANDN U2174 ( .B(n1442), .A(n522), .Z(n1441) );
  NANDN U2175 ( .B(n1443), .A(n1444), .Z(n1440) );
  AND U2176 ( .A(n1445), .B(n1446), .Z(n1346) );
  NANDN U2177 ( .B(n1447), .A(n1448), .Z(n1446) );
  OR U2178 ( .A(n1449), .B(n1450), .Z(n1445) );
  XNOR U2179 ( .A(n1371), .B(n1370), .Z(n1353) );
  XOR U2180 ( .A(n1454), .B(n1381), .Z(n1370) );
  XNOR U2181 ( .A(n1362), .B(n1361), .Z(n1381) );
  XOR U2182 ( .A(n1455), .B(n1358), .Z(n1361) );
  XNOR U2183 ( .A(n1357), .B(n1456), .Z(n1358) );
  ANDN U2184 ( .A(n1032), .B(n755), .Z(n1456) );
  XOR U2185 ( .A(n1457), .B(n1458), .Z(n1357) );
  AND U2186 ( .A(n1459), .B(n1460), .Z(n1458) );
  XNOR U2187 ( .A(n1461), .B(n1457), .Z(n1460) );
  AND U2188 ( .A(n753), .B(n969), .Z(n1359) );
  XNOR U2189 ( .A(n1366), .B(n1368), .Z(n1362) );
  NANDN U2190 ( .B(n834), .A(n876), .Z(n1368) );
  XNOR U2191 ( .A(n1364), .B(n1465), .Z(n1366) );
  ANDN U2192 ( .A(n904), .B(n878), .Z(n1465) );
  XNOR U2193 ( .A(n1380), .B(n1369), .Z(n1454) );
  XOR U2194 ( .A(n1472), .B(n1385), .Z(n1380) );
  XNOR U2195 ( .A(n1376), .B(n1378), .Z(n1385) );
  NAND U2196 ( .A(n667), .B(n1203), .Z(n1378) );
  XNOR U2197 ( .A(n1374), .B(n1473), .Z(n1376) );
  ANDN U2198 ( .A(n1210), .B(n669), .Z(n1473) );
  XOR U2199 ( .A(n1474), .B(n1475), .Z(n1374) );
  AND U2200 ( .A(n1476), .B(n1477), .Z(n1475) );
  XOR U2201 ( .A(n1478), .B(n1474), .Z(n1477) );
  XNOR U2202 ( .A(n1384), .B(n1379), .Z(n1472) );
  XOR U2203 ( .A(n1482), .B(n1391), .Z(n1384) );
  XNOR U2204 ( .A(n1389), .B(n1483), .Z(n1391) );
  ANDN U2205 ( .A(n1394), .B(n585), .Z(n1483) );
  XOR U2206 ( .A(n1484), .B(n1485), .Z(n1389) );
  AND U2207 ( .A(n1486), .B(n1487), .Z(n1485) );
  XNOR U2208 ( .A(n1488), .B(n1484), .Z(n1487) );
  AND U2209 ( .A(n583), .B(n1387), .Z(n1393) );
  XNOR U2210 ( .A(n1402), .B(n1401), .Z(n1371) );
  XOR U2211 ( .A(n1492), .B(n1410), .Z(n1401) );
  XNOR U2212 ( .A(n1398), .B(n1399), .Z(n1410) );
  NANDN U2213 ( .B(n647), .A(n1163), .Z(n1399) );
  XNOR U2214 ( .A(n1397), .B(n1493), .Z(n1398) );
  ANDN U2215 ( .A(n688), .B(n1165), .Z(n1493) );
  XNOR U2216 ( .A(n1409), .B(n1400), .Z(n1492) );
  XOR U2217 ( .A(n1500), .B(n1406), .Z(n1409) );
  XNOR U2218 ( .A(n1405), .B(n1501), .Z(n1406) );
  ANDN U2219 ( .A(n795), .B(n1013), .Z(n1501) );
  AND U2220 ( .A(n1011), .B(n741), .Z(n1407) );
  XOR U2221 ( .A(n1418), .B(n1417), .Z(n1402) );
  XOR U2222 ( .A(n1508), .B(n1414), .Z(n1417) );
  XNOR U2223 ( .A(n1413), .B(n1509), .Z(n1414) );
  ANDN U2224 ( .A(n620), .B(n1330), .Z(n1509) );
  AND U2225 ( .A(n1328), .B(n579), .Z(n1415) );
  XOR U2226 ( .A(n1425), .B(n1424), .Z(n1418) );
  NAND U2227 ( .A(n1516), .B(n523), .Z(n1424) );
  XOR U2228 ( .A(n1423), .B(n1517), .Z(n1425) );
  ANDN U2229 ( .A(n554), .B(n1518), .Z(n1517) );
  ANDN U2230 ( .A(n1519), .B(n1520), .Z(n1423) );
  NAND U2231 ( .A(n1521), .B(n1522), .Z(n1519) );
  IV U2232 ( .A(n1426), .Z(n1427) );
  MUX U2233 ( .IN0(o[12]), .IN1(n416), .SEL(n475), .F(\_MxM/n311 ) );
  XOR U2234 ( .A(n1527), .B(\_MxM/Y0[13] ), .Z(n416) );
  XNOR U2235 ( .A(n1528), .B(n1529), .Z(n1527) );
  AND U2236 ( .A(n487), .B(n1531), .Z(n1530) );
  XNOR U2237 ( .A(n1525), .B(n1529), .Z(n1531) );
  XNOR U2238 ( .A(n1524), .B(n1529), .Z(n1525) );
  XNOR U2239 ( .A(n1453), .B(n1452), .Z(n1529) );
  XOR U2240 ( .A(n1532), .B(n1437), .Z(n1452) );
  NANDN U2241 ( .B(n1533), .A(n1534), .Z(n1443) );
  XOR U2242 ( .A(n1537), .B(n1450), .Z(n1447) );
  NAND U2243 ( .A(n1538), .B(n552), .Z(n1450) );
  NAND U2244 ( .A(n1539), .B(n1449), .Z(n1537) );
  NANDN U2245 ( .B(n555), .A(n1543), .Z(n1539) );
  XNOR U2246 ( .A(n1436), .B(n1451), .Z(n1532) );
  IV U2247 ( .A(n1438), .Z(n1436) );
  XNOR U2248 ( .A(n1471), .B(n1470), .Z(n1453) );
  XOR U2249 ( .A(n1550), .B(n1481), .Z(n1470) );
  XNOR U2250 ( .A(n1464), .B(n1463), .Z(n1481) );
  XOR U2251 ( .A(n1551), .B(n1459), .Z(n1463) );
  XNOR U2252 ( .A(n1457), .B(n1552), .Z(n1459) );
  ANDN U2253 ( .A(n1032), .B(n814), .Z(n1552) );
  XOR U2254 ( .A(n1553), .B(n1554), .Z(n1457) );
  AND U2255 ( .A(n1555), .B(n1556), .Z(n1554) );
  XNOR U2256 ( .A(n1557), .B(n1553), .Z(n1556) );
  AND U2257 ( .A(n812), .B(n969), .Z(n1461) );
  XNOR U2258 ( .A(n1467), .B(n1468), .Z(n1464) );
  NANDN U2259 ( .B(n834), .A(n944), .Z(n1468) );
  XNOR U2260 ( .A(n1466), .B(n1561), .Z(n1467) );
  ANDN U2261 ( .A(n904), .B(n946), .Z(n1561) );
  XNOR U2262 ( .A(n1480), .B(n1469), .Z(n1550) );
  XOR U2263 ( .A(n1568), .B(n1491), .Z(n1480) );
  XNOR U2264 ( .A(n1476), .B(n1478), .Z(n1491) );
  NAND U2265 ( .A(n711), .B(n1203), .Z(n1478) );
  XNOR U2266 ( .A(n1474), .B(n1569), .Z(n1476) );
  ANDN U2267 ( .A(n1210), .B(n713), .Z(n1569) );
  XOR U2268 ( .A(n1570), .B(n1571), .Z(n1474) );
  AND U2269 ( .A(n1572), .B(n1573), .Z(n1571) );
  XOR U2270 ( .A(n1574), .B(n1570), .Z(n1573) );
  XNOR U2271 ( .A(n1490), .B(n1479), .Z(n1568) );
  XOR U2272 ( .A(n1578), .B(n1486), .Z(n1490) );
  XNOR U2273 ( .A(n1484), .B(n1579), .Z(n1486) );
  ANDN U2274 ( .A(n1394), .B(n629), .Z(n1579) );
  XOR U2275 ( .A(n1580), .B(n1581), .Z(n1484) );
  AND U2276 ( .A(n1582), .B(n1583), .Z(n1581) );
  XNOR U2277 ( .A(n1584), .B(n1580), .Z(n1583) );
  AND U2278 ( .A(n627), .B(n1387), .Z(n1488) );
  XNOR U2279 ( .A(n1499), .B(n1498), .Z(n1471) );
  XOR U2280 ( .A(n1588), .B(n1507), .Z(n1498) );
  XNOR U2281 ( .A(n1495), .B(n1496), .Z(n1507) );
  NANDN U2282 ( .B(n647), .A(n1244), .Z(n1496) );
  XNOR U2283 ( .A(n1494), .B(n1589), .Z(n1495) );
  ANDN U2284 ( .A(n688), .B(n1246), .Z(n1589) );
  XNOR U2285 ( .A(n1506), .B(n1497), .Z(n1588) );
  XOR U2286 ( .A(n1596), .B(n1503), .Z(n1506) );
  XNOR U2287 ( .A(n1502), .B(n1597), .Z(n1503) );
  ANDN U2288 ( .A(n795), .B(n1087), .Z(n1597) );
  AND U2289 ( .A(n1085), .B(n741), .Z(n1504) );
  XOR U2290 ( .A(n1515), .B(n1514), .Z(n1499) );
  XOR U2291 ( .A(n1604), .B(n1511), .Z(n1514) );
  XNOR U2292 ( .A(n1510), .B(n1605), .Z(n1511) );
  ANDN U2293 ( .A(n620), .B(n1421), .Z(n1605) );
  AND U2294 ( .A(n1419), .B(n579), .Z(n1512) );
  XOR U2295 ( .A(n1522), .B(n1521), .Z(n1515) );
  NAND U2296 ( .A(n1612), .B(n523), .Z(n1521) );
  XNOR U2297 ( .A(n1520), .B(n1613), .Z(n1522) );
  ANDN U2298 ( .A(n554), .B(n1614), .Z(n1613) );
  NAND U2299 ( .A(n1615), .B(n1616), .Z(n1520) );
  NAND U2300 ( .A(n1617), .B(n1618), .Z(n1615) );
  IV U2301 ( .A(n1523), .Z(n1524) );
  MUX U2302 ( .IN0(o[11]), .IN1(n413), .SEL(n475), .F(\_MxM/n310 ) );
  XOR U2303 ( .A(n1623), .B(\_MxM/Y0[12] ), .Z(n413) );
  XOR U2304 ( .A(n1624), .B(n1625), .Z(n1623) );
  AND U2305 ( .A(n487), .B(n1627), .Z(n1626) );
  XOR U2306 ( .A(n1621), .B(n1625), .Z(n1627) );
  XOR U2307 ( .A(n1620), .B(n1625), .Z(n1621) );
  XNOR U2308 ( .A(n1628), .B(n1549), .Z(n1545) );
  XOR U2309 ( .A(n1534), .B(n1533), .Z(n1549) );
  NANDN U2310 ( .B(n1629), .A(n1630), .Z(n1533) );
  AND U2311 ( .A(n1632), .B(n1633), .Z(n1631) );
  NANDN U2312 ( .B(n1634), .A(n522), .Z(n1633) );
  NANDN U2313 ( .B(n1635), .A(n1636), .Z(n1632) );
  XNOR U2314 ( .A(n1541), .B(n1542), .Z(n1536) );
  NAND U2315 ( .A(n1538), .B(n583), .Z(n1542) );
  XNOR U2316 ( .A(n1540), .B(n1640), .Z(n1541) );
  ANDN U2317 ( .A(n1543), .B(n585), .Z(n1640) );
  XNOR U2318 ( .A(n1548), .B(n1544), .Z(n1628) );
  IV U2319 ( .A(n1547), .Z(n1548) );
  XNOR U2320 ( .A(n1567), .B(n1566), .Z(n1546) );
  XOR U2321 ( .A(n1650), .B(n1577), .Z(n1566) );
  XNOR U2322 ( .A(n1560), .B(n1559), .Z(n1577) );
  XOR U2323 ( .A(n1651), .B(n1555), .Z(n1559) );
  XNOR U2324 ( .A(n1553), .B(n1652), .Z(n1555) );
  ANDN U2325 ( .A(n1032), .B(n878), .Z(n1652) );
  AND U2326 ( .A(n876), .B(n969), .Z(n1557) );
  XNOR U2327 ( .A(n1563), .B(n1564), .Z(n1560) );
  NANDN U2328 ( .B(n834), .A(n1011), .Z(n1564) );
  XNOR U2329 ( .A(n1562), .B(n1659), .Z(n1563) );
  ANDN U2330 ( .A(n904), .B(n1013), .Z(n1659) );
  XNOR U2331 ( .A(n1576), .B(n1565), .Z(n1650) );
  XOR U2332 ( .A(n1666), .B(n1587), .Z(n1576) );
  XNOR U2333 ( .A(n1572), .B(n1574), .Z(n1587) );
  NAND U2334 ( .A(n753), .B(n1203), .Z(n1574) );
  XNOR U2335 ( .A(n1570), .B(n1667), .Z(n1572) );
  ANDN U2336 ( .A(n1210), .B(n755), .Z(n1667) );
  XNOR U2337 ( .A(n1586), .B(n1575), .Z(n1666) );
  XOR U2338 ( .A(n1674), .B(n1582), .Z(n1586) );
  XNOR U2339 ( .A(n1580), .B(n1675), .Z(n1582) );
  ANDN U2340 ( .A(n1394), .B(n669), .Z(n1675) );
  XOR U2341 ( .A(n1676), .B(n1677), .Z(n1580) );
  AND U2342 ( .A(n1678), .B(n1679), .Z(n1677) );
  XNOR U2343 ( .A(n1680), .B(n1676), .Z(n1679) );
  AND U2344 ( .A(n667), .B(n1387), .Z(n1584) );
  XNOR U2345 ( .A(n1595), .B(n1594), .Z(n1567) );
  XOR U2346 ( .A(n1684), .B(n1603), .Z(n1594) );
  XNOR U2347 ( .A(n1591), .B(n1592), .Z(n1603) );
  NANDN U2348 ( .B(n647), .A(n1328), .Z(n1592) );
  XNOR U2349 ( .A(n1590), .B(n1685), .Z(n1591) );
  ANDN U2350 ( .A(n688), .B(n1330), .Z(n1685) );
  XNOR U2351 ( .A(n1602), .B(n1593), .Z(n1684) );
  XOR U2352 ( .A(n1692), .B(n1599), .Z(n1602) );
  XNOR U2353 ( .A(n1598), .B(n1693), .Z(n1599) );
  ANDN U2354 ( .A(n795), .B(n1165), .Z(n1693) );
  AND U2355 ( .A(n1163), .B(n741), .Z(n1600) );
  XOR U2356 ( .A(n1611), .B(n1610), .Z(n1595) );
  XOR U2357 ( .A(n1700), .B(n1607), .Z(n1610) );
  XNOR U2358 ( .A(n1606), .B(n1701), .Z(n1607) );
  ANDN U2359 ( .A(n620), .B(n1518), .Z(n1701) );
  AND U2360 ( .A(n1516), .B(n579), .Z(n1608) );
  XOR U2361 ( .A(n1618), .B(n1617), .Z(n1611) );
  NAND U2362 ( .A(n1708), .B(n523), .Z(n1617) );
  XOR U2363 ( .A(n1616), .B(n1709), .Z(n1618) );
  ANDN U2364 ( .A(n554), .B(n1710), .Z(n1709) );
  ANDN U2365 ( .A(n1711), .B(n1712), .Z(n1616) );
  NAND U2366 ( .A(n1713), .B(n1714), .Z(n1711) );
  IV U2367 ( .A(n1619), .Z(n1620) );
  MUX U2368 ( .IN0(o[10]), .IN1(n410), .SEL(n475), .F(\_MxM/n309 ) );
  XOR U2369 ( .A(n1719), .B(\_MxM/Y0[11] ), .Z(n410) );
  XNOR U2370 ( .A(n1720), .B(n1721), .Z(n1719) );
  AND U2371 ( .A(n487), .B(n1723), .Z(n1722) );
  XNOR U2372 ( .A(n1717), .B(n1721), .Z(n1723) );
  XNOR U2373 ( .A(n1716), .B(n1721), .Z(n1717) );
  XNOR U2374 ( .A(n1646), .B(n1645), .Z(n1721) );
  XOR U2375 ( .A(n1724), .B(n1649), .Z(n1645) );
  XOR U2376 ( .A(n1639), .B(n1638), .Z(n1629) );
  XOR U2377 ( .A(n1732), .B(n1636), .Z(n1728) );
  AND U2378 ( .A(n1733), .B(n552), .Z(n1636) );
  NAND U2379 ( .A(n1734), .B(n1635), .Z(n1732) );
  XOR U2380 ( .A(n1735), .B(n1736), .Z(n1635) );
  AND U2381 ( .A(n1737), .B(n1738), .Z(n1736) );
  XNOR U2382 ( .A(n1739), .B(n1735), .Z(n1738) );
  NANDN U2383 ( .B(n555), .A(n1740), .Z(n1734) );
  XNOR U2384 ( .A(n1642), .B(n1643), .Z(n1639) );
  NAND U2385 ( .A(n1538), .B(n627), .Z(n1643) );
  XNOR U2386 ( .A(n1641), .B(n1741), .Z(n1642) );
  ANDN U2387 ( .A(n1543), .B(n629), .Z(n1741) );
  XNOR U2388 ( .A(n1648), .B(n1644), .Z(n1724) );
  IV U2389 ( .A(n1647), .Z(n1648) );
  XNOR U2390 ( .A(n1665), .B(n1664), .Z(n1646) );
  XOR U2391 ( .A(n1751), .B(n1673), .Z(n1664) );
  XNOR U2392 ( .A(n1658), .B(n1657), .Z(n1673) );
  XOR U2393 ( .A(n1752), .B(n1654), .Z(n1657) );
  XNOR U2394 ( .A(n1653), .B(n1753), .Z(n1654) );
  ANDN U2395 ( .A(n1032), .B(n946), .Z(n1753) );
  AND U2396 ( .A(n944), .B(n969), .Z(n1655) );
  XNOR U2397 ( .A(n1661), .B(n1662), .Z(n1658) );
  NANDN U2398 ( .B(n834), .A(n1085), .Z(n1662) );
  XNOR U2399 ( .A(n1660), .B(n1760), .Z(n1661) );
  ANDN U2400 ( .A(n904), .B(n1087), .Z(n1760) );
  XNOR U2401 ( .A(n1672), .B(n1663), .Z(n1751) );
  XOR U2402 ( .A(n1767), .B(n1683), .Z(n1672) );
  XNOR U2403 ( .A(n1669), .B(n1670), .Z(n1683) );
  NAND U2404 ( .A(n812), .B(n1203), .Z(n1670) );
  XNOR U2405 ( .A(n1668), .B(n1768), .Z(n1669) );
  ANDN U2406 ( .A(n1210), .B(n814), .Z(n1768) );
  XNOR U2407 ( .A(n1682), .B(n1671), .Z(n1767) );
  XOR U2408 ( .A(n1775), .B(n1678), .Z(n1682) );
  XNOR U2409 ( .A(n1676), .B(n1776), .Z(n1678) );
  ANDN U2410 ( .A(n1394), .B(n713), .Z(n1776) );
  XOR U2411 ( .A(n1777), .B(n1778), .Z(n1676) );
  AND U2412 ( .A(n1779), .B(n1780), .Z(n1778) );
  XNOR U2413 ( .A(n1781), .B(n1777), .Z(n1780) );
  AND U2414 ( .A(n711), .B(n1387), .Z(n1680) );
  XNOR U2415 ( .A(n1691), .B(n1690), .Z(n1665) );
  XOR U2416 ( .A(n1785), .B(n1699), .Z(n1690) );
  XNOR U2417 ( .A(n1687), .B(n1688), .Z(n1699) );
  NANDN U2418 ( .B(n647), .A(n1419), .Z(n1688) );
  XNOR U2419 ( .A(n1686), .B(n1786), .Z(n1687) );
  ANDN U2420 ( .A(n688), .B(n1421), .Z(n1786) );
  XNOR U2421 ( .A(n1698), .B(n1689), .Z(n1785) );
  XOR U2422 ( .A(n1793), .B(n1695), .Z(n1698) );
  XNOR U2423 ( .A(n1694), .B(n1794), .Z(n1695) );
  ANDN U2424 ( .A(n795), .B(n1246), .Z(n1794) );
  AND U2425 ( .A(n1244), .B(n741), .Z(n1696) );
  XOR U2426 ( .A(n1707), .B(n1706), .Z(n1691) );
  XOR U2427 ( .A(n1801), .B(n1703), .Z(n1706) );
  XNOR U2428 ( .A(n1702), .B(n1802), .Z(n1703) );
  ANDN U2429 ( .A(n620), .B(n1614), .Z(n1802) );
  AND U2430 ( .A(n1612), .B(n579), .Z(n1704) );
  XOR U2431 ( .A(n1714), .B(n1713), .Z(n1707) );
  NAND U2432 ( .A(n1809), .B(n523), .Z(n1713) );
  XNOR U2433 ( .A(n1712), .B(n1810), .Z(n1714) );
  ANDN U2434 ( .A(n554), .B(n1811), .Z(n1810) );
  NAND U2435 ( .A(n1812), .B(n1813), .Z(n1712) );
  NAND U2436 ( .A(n1814), .B(n1815), .Z(n1812) );
  IV U2437 ( .A(n1715), .Z(n1716) );
  MUX U2438 ( .IN0(o[9]), .IN1(n407), .SEL(n475), .F(\_MxM/n308 ) );
  XOR U2439 ( .A(n1820), .B(\_MxM/Y0[10] ), .Z(n407) );
  XOR U2440 ( .A(n1821), .B(n1822), .Z(n1820) );
  AND U2441 ( .A(n487), .B(n1824), .Z(n1823) );
  XOR U2442 ( .A(n1818), .B(n1822), .Z(n1824) );
  XOR U2443 ( .A(n1817), .B(n1822), .Z(n1818) );
  XNOR U2444 ( .A(n1825), .B(n1750), .Z(n1746) );
  XNOR U2445 ( .A(n1727), .B(n1726), .Z(n1750) );
  XOR U2446 ( .A(n1725), .B(n1826), .Z(n1726) );
  AND U2447 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U2448 ( .B(n1829), .A(n1830), .Z(n1828) );
  AND U2449 ( .A(n1831), .B(n1832), .Z(n1827) );
  NANDN U2450 ( .B(n1833), .A(n522), .Z(n1832) );
  OR U2451 ( .A(n1834), .B(n1835), .Z(n1831) );
  XNOR U2452 ( .A(n1731), .B(n1730), .Z(n1727) );
  XOR U2453 ( .A(n1839), .B(n1737), .Z(n1730) );
  XNOR U2454 ( .A(n1735), .B(n1840), .Z(n1737) );
  ANDN U2455 ( .A(n1740), .B(n585), .Z(n1840) );
  XOR U2456 ( .A(n1841), .B(n1842), .Z(n1735) );
  AND U2457 ( .A(n1843), .B(n1844), .Z(n1842) );
  XNOR U2458 ( .A(n1845), .B(n1841), .Z(n1844) );
  AND U2459 ( .A(n1733), .B(n583), .Z(n1739) );
  XNOR U2460 ( .A(n1743), .B(n1744), .Z(n1731) );
  NAND U2461 ( .A(n1538), .B(n667), .Z(n1744) );
  XNOR U2462 ( .A(n1742), .B(n1849), .Z(n1743) );
  ANDN U2463 ( .A(n1543), .B(n669), .Z(n1849) );
  XNOR U2464 ( .A(n1749), .B(n1745), .Z(n1825) );
  IV U2465 ( .A(n1748), .Z(n1749) );
  XNOR U2466 ( .A(n1766), .B(n1765), .Z(n1747) );
  XOR U2467 ( .A(n1859), .B(n1774), .Z(n1765) );
  XNOR U2468 ( .A(n1759), .B(n1758), .Z(n1774) );
  XOR U2469 ( .A(n1860), .B(n1755), .Z(n1758) );
  XNOR U2470 ( .A(n1754), .B(n1861), .Z(n1755) );
  ANDN U2471 ( .A(n1032), .B(n1013), .Z(n1861) );
  AND U2472 ( .A(n1011), .B(n969), .Z(n1756) );
  XNOR U2473 ( .A(n1762), .B(n1763), .Z(n1759) );
  NANDN U2474 ( .B(n834), .A(n1163), .Z(n1763) );
  XNOR U2475 ( .A(n1761), .B(n1868), .Z(n1762) );
  ANDN U2476 ( .A(n904), .B(n1165), .Z(n1868) );
  XNOR U2477 ( .A(n1773), .B(n1764), .Z(n1859) );
  XOR U2478 ( .A(n1875), .B(n1784), .Z(n1773) );
  XNOR U2479 ( .A(n1770), .B(n1771), .Z(n1784) );
  NAND U2480 ( .A(n876), .B(n1203), .Z(n1771) );
  XNOR U2481 ( .A(n1769), .B(n1876), .Z(n1770) );
  ANDN U2482 ( .A(n1210), .B(n878), .Z(n1876) );
  XNOR U2483 ( .A(n1783), .B(n1772), .Z(n1875) );
  XOR U2484 ( .A(n1883), .B(n1779), .Z(n1783) );
  XNOR U2485 ( .A(n1777), .B(n1884), .Z(n1779) );
  ANDN U2486 ( .A(n1394), .B(n755), .Z(n1884) );
  AND U2487 ( .A(n753), .B(n1387), .Z(n1781) );
  XNOR U2488 ( .A(n1792), .B(n1791), .Z(n1766) );
  XOR U2489 ( .A(n1891), .B(n1800), .Z(n1791) );
  XNOR U2490 ( .A(n1788), .B(n1789), .Z(n1800) );
  NANDN U2491 ( .B(n647), .A(n1516), .Z(n1789) );
  XNOR U2492 ( .A(n1787), .B(n1892), .Z(n1788) );
  ANDN U2493 ( .A(n688), .B(n1518), .Z(n1892) );
  XNOR U2494 ( .A(n1799), .B(n1790), .Z(n1891) );
  XOR U2495 ( .A(n1899), .B(n1796), .Z(n1799) );
  XNOR U2496 ( .A(n1795), .B(n1900), .Z(n1796) );
  ANDN U2497 ( .A(n795), .B(n1330), .Z(n1900) );
  AND U2498 ( .A(n1328), .B(n741), .Z(n1797) );
  XOR U2499 ( .A(n1808), .B(n1807), .Z(n1792) );
  XOR U2500 ( .A(n1907), .B(n1804), .Z(n1807) );
  XNOR U2501 ( .A(n1803), .B(n1908), .Z(n1804) );
  ANDN U2502 ( .A(n620), .B(n1710), .Z(n1908) );
  AND U2503 ( .A(n1708), .B(n579), .Z(n1805) );
  XOR U2504 ( .A(n1815), .B(n1814), .Z(n1808) );
  NAND U2505 ( .A(n1915), .B(n523), .Z(n1814) );
  XOR U2506 ( .A(n1813), .B(n1916), .Z(n1815) );
  ANDN U2507 ( .A(n554), .B(n1917), .Z(n1916) );
  ANDN U2508 ( .A(n1918), .B(n1919), .Z(n1813) );
  NAND U2509 ( .A(n1920), .B(n1921), .Z(n1918) );
  IV U2510 ( .A(n1816), .Z(n1817) );
  MUX U2511 ( .IN0(o[8]), .IN1(n404), .SEL(n475), .F(\_MxM/n307 ) );
  XOR U2512 ( .A(n1926), .B(\_MxM/Y0[9] ), .Z(n404) );
  XOR U2513 ( .A(n1927), .B(n1928), .Z(n1926) );
  AND U2514 ( .A(n487), .B(n1930), .Z(n1929) );
  XOR U2515 ( .A(n1924), .B(n1928), .Z(n1930) );
  XOR U2516 ( .A(n1923), .B(n1928), .Z(n1924) );
  XNOR U2517 ( .A(n1931), .B(n1858), .Z(n1854) );
  XNOR U2518 ( .A(n1838), .B(n1837), .Z(n1858) );
  XOR U2519 ( .A(n1932), .B(n1834), .Z(n1837) );
  XNOR U2520 ( .A(n1933), .B(n1830), .Z(n1834) );
  AND U2521 ( .A(n1934), .B(n552), .Z(n1830) );
  NAND U2522 ( .A(n1935), .B(n1829), .Z(n1933) );
  NANDN U2523 ( .B(n555), .A(n1939), .Z(n1935) );
  XNOR U2524 ( .A(n1835), .B(n1836), .Z(n1932) );
  XNOR U2525 ( .A(n1943), .B(n1946), .Z(n1945) );
  XNOR U2526 ( .A(n1848), .B(n1847), .Z(n1838) );
  XOR U2527 ( .A(n1947), .B(n1843), .Z(n1847) );
  XNOR U2528 ( .A(n1841), .B(n1948), .Z(n1843) );
  ANDN U2529 ( .A(n1740), .B(n629), .Z(n1948) );
  XOR U2530 ( .A(n1949), .B(n1950), .Z(n1841) );
  AND U2531 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR U2532 ( .A(n1953), .B(n1949), .Z(n1952) );
  AND U2533 ( .A(n1733), .B(n627), .Z(n1845) );
  XNOR U2534 ( .A(n1851), .B(n1852), .Z(n1848) );
  NAND U2535 ( .A(n1538), .B(n711), .Z(n1852) );
  XNOR U2536 ( .A(n1850), .B(n1957), .Z(n1851) );
  ANDN U2537 ( .A(n1543), .B(n713), .Z(n1957) );
  XNOR U2538 ( .A(n1857), .B(n1853), .Z(n1931) );
  IV U2539 ( .A(n1856), .Z(n1857) );
  XNOR U2540 ( .A(n1874), .B(n1873), .Z(n1855) );
  XOR U2541 ( .A(n1966), .B(n1882), .Z(n1873) );
  XNOR U2542 ( .A(n1867), .B(n1866), .Z(n1882) );
  XOR U2543 ( .A(n1967), .B(n1863), .Z(n1866) );
  XNOR U2544 ( .A(n1862), .B(n1968), .Z(n1863) );
  ANDN U2545 ( .A(n1032), .B(n1087), .Z(n1968) );
  AND U2546 ( .A(n1085), .B(n969), .Z(n1864) );
  XNOR U2547 ( .A(n1870), .B(n1871), .Z(n1867) );
  NANDN U2548 ( .B(n834), .A(n1244), .Z(n1871) );
  XNOR U2549 ( .A(n1869), .B(n1975), .Z(n1870) );
  ANDN U2550 ( .A(n904), .B(n1246), .Z(n1975) );
  XNOR U2551 ( .A(n1881), .B(n1872), .Z(n1966) );
  XOR U2552 ( .A(n1982), .B(n1890), .Z(n1881) );
  XNOR U2553 ( .A(n1878), .B(n1879), .Z(n1890) );
  NAND U2554 ( .A(n944), .B(n1203), .Z(n1879) );
  XNOR U2555 ( .A(n1877), .B(n1983), .Z(n1878) );
  ANDN U2556 ( .A(n1210), .B(n946), .Z(n1983) );
  XNOR U2557 ( .A(n1889), .B(n1880), .Z(n1982) );
  XOR U2558 ( .A(n1990), .B(n1886), .Z(n1889) );
  XNOR U2559 ( .A(n1885), .B(n1991), .Z(n1886) );
  ANDN U2560 ( .A(n1394), .B(n814), .Z(n1991) );
  AND U2561 ( .A(n812), .B(n1387), .Z(n1887) );
  XNOR U2562 ( .A(n1898), .B(n1897), .Z(n1874) );
  XOR U2563 ( .A(n1998), .B(n1906), .Z(n1897) );
  XNOR U2564 ( .A(n1894), .B(n1895), .Z(n1906) );
  NANDN U2565 ( .B(n647), .A(n1612), .Z(n1895) );
  XNOR U2566 ( .A(n1893), .B(n1999), .Z(n1894) );
  ANDN U2567 ( .A(n688), .B(n1614), .Z(n1999) );
  XNOR U2568 ( .A(n1905), .B(n1896), .Z(n1998) );
  XOR U2569 ( .A(n2006), .B(n1902), .Z(n1905) );
  XNOR U2570 ( .A(n1901), .B(n2007), .Z(n1902) );
  ANDN U2571 ( .A(n795), .B(n1421), .Z(n2007) );
  AND U2572 ( .A(n1419), .B(n741), .Z(n1903) );
  XOR U2573 ( .A(n1914), .B(n1913), .Z(n1898) );
  XOR U2574 ( .A(n2014), .B(n1910), .Z(n1913) );
  XNOR U2575 ( .A(n1909), .B(n2015), .Z(n1910) );
  ANDN U2576 ( .A(n620), .B(n1811), .Z(n2015) );
  AND U2577 ( .A(n1809), .B(n579), .Z(n1911) );
  XOR U2578 ( .A(n1921), .B(n1920), .Z(n1914) );
  NAND U2579 ( .A(n2022), .B(n523), .Z(n1920) );
  XNOR U2580 ( .A(n1919), .B(n2023), .Z(n1921) );
  ANDN U2581 ( .A(n554), .B(n2024), .Z(n2023) );
  NAND U2582 ( .A(n2025), .B(n2026), .Z(n1919) );
  NAND U2583 ( .A(n2027), .B(n2028), .Z(n2025) );
  IV U2584 ( .A(n1922), .Z(n1923) );
  MUX U2585 ( .IN0(o[7]), .IN1(n401), .SEL(n475), .F(\_MxM/n306 ) );
  XOR U2586 ( .A(n2033), .B(\_MxM/Y0[8] ), .Z(n401) );
  XOR U2587 ( .A(n2034), .B(n2035), .Z(n2033) );
  AND U2588 ( .A(n487), .B(n2037), .Z(n2036) );
  XOR U2589 ( .A(n2031), .B(n2035), .Z(n2037) );
  XOR U2590 ( .A(n2030), .B(n2035), .Z(n2031) );
  XNOR U2591 ( .A(n2038), .B(n1965), .Z(n1962) );
  XNOR U2592 ( .A(n1942), .B(n1941), .Z(n1965) );
  XOR U2593 ( .A(n2039), .B(n1946), .Z(n1941) );
  XNOR U2594 ( .A(n1937), .B(n1938), .Z(n1946) );
  NAND U2595 ( .A(n1934), .B(n583), .Z(n1938) );
  XNOR U2596 ( .A(n1936), .B(n2040), .Z(n1937) );
  ANDN U2597 ( .A(n1939), .B(n585), .Z(n2040) );
  XNOR U2598 ( .A(n1944), .B(n1940), .Z(n2039) );
  XOR U2599 ( .A(n1943), .B(n2047), .Z(n1944) );
  AND U2600 ( .A(n2048), .B(n2049), .Z(n2047) );
  NANDN U2601 ( .B(n2050), .A(n522), .Z(n2049) );
  NANDN U2602 ( .B(n2051), .A(n2052), .Z(n2048) );
  XNOR U2603 ( .A(n1956), .B(n1955), .Z(n1942) );
  XOR U2604 ( .A(n2056), .B(n1951), .Z(n1955) );
  XNOR U2605 ( .A(n1949), .B(n2057), .Z(n1951) );
  ANDN U2606 ( .A(n1740), .B(n669), .Z(n2057) );
  AND U2607 ( .A(n1733), .B(n667), .Z(n1953) );
  XNOR U2608 ( .A(n1959), .B(n1960), .Z(n1956) );
  NAND U2609 ( .A(n1538), .B(n753), .Z(n1960) );
  XNOR U2610 ( .A(n1958), .B(n2064), .Z(n1959) );
  ANDN U2611 ( .A(n1543), .B(n755), .Z(n2064) );
  XNOR U2612 ( .A(n1981), .B(n1980), .Z(n1963) );
  XOR U2613 ( .A(n2074), .B(n1989), .Z(n1980) );
  XNOR U2614 ( .A(n1974), .B(n1973), .Z(n1989) );
  XOR U2615 ( .A(n2075), .B(n1970), .Z(n1973) );
  XNOR U2616 ( .A(n1969), .B(n2076), .Z(n1970) );
  ANDN U2617 ( .A(n1032), .B(n1165), .Z(n2076) );
  AND U2618 ( .A(n1163), .B(n969), .Z(n1971) );
  XNOR U2619 ( .A(n1977), .B(n1978), .Z(n1974) );
  NANDN U2620 ( .B(n834), .A(n1328), .Z(n1978) );
  XNOR U2621 ( .A(n1976), .B(n2083), .Z(n1977) );
  ANDN U2622 ( .A(n904), .B(n1330), .Z(n2083) );
  XNOR U2623 ( .A(n1988), .B(n1979), .Z(n2074) );
  XOR U2624 ( .A(n2090), .B(n1997), .Z(n1988) );
  XNOR U2625 ( .A(n1985), .B(n1986), .Z(n1997) );
  NAND U2626 ( .A(n1011), .B(n1203), .Z(n1986) );
  XNOR U2627 ( .A(n1984), .B(n2091), .Z(n1985) );
  ANDN U2628 ( .A(n1210), .B(n1013), .Z(n2091) );
  XNOR U2629 ( .A(n1996), .B(n1987), .Z(n2090) );
  XOR U2630 ( .A(n2098), .B(n1993), .Z(n1996) );
  XNOR U2631 ( .A(n1992), .B(n2099), .Z(n1993) );
  ANDN U2632 ( .A(n1394), .B(n878), .Z(n2099) );
  AND U2633 ( .A(n876), .B(n1387), .Z(n1994) );
  XNOR U2634 ( .A(n2005), .B(n2004), .Z(n1981) );
  XOR U2635 ( .A(n2106), .B(n2013), .Z(n2004) );
  XNOR U2636 ( .A(n2001), .B(n2002), .Z(n2013) );
  NANDN U2637 ( .B(n647), .A(n1708), .Z(n2002) );
  XNOR U2638 ( .A(n2000), .B(n2107), .Z(n2001) );
  ANDN U2639 ( .A(n688), .B(n1710), .Z(n2107) );
  XNOR U2640 ( .A(n2012), .B(n2003), .Z(n2106) );
  XOR U2641 ( .A(n2114), .B(n2009), .Z(n2012) );
  XNOR U2642 ( .A(n2008), .B(n2115), .Z(n2009) );
  ANDN U2643 ( .A(n795), .B(n1518), .Z(n2115) );
  AND U2644 ( .A(n1516), .B(n741), .Z(n2010) );
  XOR U2645 ( .A(n2021), .B(n2020), .Z(n2005) );
  XOR U2646 ( .A(n2122), .B(n2017), .Z(n2020) );
  XNOR U2647 ( .A(n2016), .B(n2123), .Z(n2017) );
  ANDN U2648 ( .A(n620), .B(n1917), .Z(n2123) );
  AND U2649 ( .A(n1915), .B(n579), .Z(n2018) );
  XOR U2650 ( .A(n2028), .B(n2027), .Z(n2021) );
  NAND U2651 ( .A(n2130), .B(n523), .Z(n2027) );
  XOR U2652 ( .A(n2026), .B(n2131), .Z(n2028) );
  ANDN U2653 ( .A(n554), .B(n2132), .Z(n2131) );
  ANDN U2654 ( .A(n2133), .B(n2134), .Z(n2026) );
  NAND U2655 ( .A(n2135), .B(n2136), .Z(n2133) );
  IV U2656 ( .A(n2029), .Z(n2030) );
  MUX U2657 ( .IN0(o[6]), .IN1(n398), .SEL(n475), .F(\_MxM/n305 ) );
  XOR U2658 ( .A(n2141), .B(\_MxM/Y0[7] ), .Z(n398) );
  XOR U2659 ( .A(n2142), .B(n2143), .Z(n2141) );
  AND U2660 ( .A(n487), .B(n2145), .Z(n2144) );
  XOR U2661 ( .A(n2139), .B(n2143), .Z(n2145) );
  XOR U2662 ( .A(n2138), .B(n2143), .Z(n2139) );
  XNOR U2663 ( .A(n2146), .B(n2073), .Z(n2069) );
  XNOR U2664 ( .A(n2046), .B(n2045), .Z(n2073) );
  XOR U2665 ( .A(n2147), .B(n2055), .Z(n2045) );
  XNOR U2666 ( .A(n2042), .B(n2043), .Z(n2055) );
  NAND U2667 ( .A(n1934), .B(n627), .Z(n2043) );
  XNOR U2668 ( .A(n2041), .B(n2148), .Z(n2042) );
  ANDN U2669 ( .A(n1939), .B(n629), .Z(n2148) );
  XOR U2670 ( .A(n2149), .B(n2150), .Z(n2041) );
  AND U2671 ( .A(n2151), .B(n2152), .Z(n2150) );
  XOR U2672 ( .A(n2153), .B(n2149), .Z(n2152) );
  XNOR U2673 ( .A(n2054), .B(n2044), .Z(n2147) );
  XOR U2674 ( .A(n2161), .B(n2052), .Z(n2157) );
  AND U2675 ( .A(n2162), .B(n552), .Z(n2052) );
  NAND U2676 ( .A(n2163), .B(n2051), .Z(n2161) );
  XOR U2677 ( .A(n2164), .B(n2165), .Z(n2051) );
  AND U2678 ( .A(n2166), .B(n2167), .Z(n2165) );
  XNOR U2679 ( .A(n2168), .B(n2164), .Z(n2167) );
  NANDN U2680 ( .B(n555), .A(n2169), .Z(n2163) );
  XNOR U2681 ( .A(n2063), .B(n2062), .Z(n2046) );
  XOR U2682 ( .A(n2170), .B(n2059), .Z(n2062) );
  XNOR U2683 ( .A(n2058), .B(n2171), .Z(n2059) );
  ANDN U2684 ( .A(n1740), .B(n713), .Z(n2171) );
  AND U2685 ( .A(n1733), .B(n711), .Z(n2060) );
  XNOR U2686 ( .A(n2066), .B(n2067), .Z(n2063) );
  NAND U2687 ( .A(n1538), .B(n812), .Z(n2067) );
  XNOR U2688 ( .A(n2065), .B(n2178), .Z(n2066) );
  ANDN U2689 ( .A(n1543), .B(n814), .Z(n2178) );
  XNOR U2690 ( .A(n2072), .B(n2068), .Z(n2146) );
  XOR U2691 ( .A(n2189), .B(n2190), .Z(n2185) );
  NANDN U2692 ( .B(n2191), .A(n2192), .Z(n2189) );
  XNOR U2693 ( .A(n2089), .B(n2088), .Z(n2070) );
  XOR U2694 ( .A(n2193), .B(n2097), .Z(n2088) );
  XNOR U2695 ( .A(n2082), .B(n2081), .Z(n2097) );
  XOR U2696 ( .A(n2194), .B(n2078), .Z(n2081) );
  XNOR U2697 ( .A(n2077), .B(n2195), .Z(n2078) );
  ANDN U2698 ( .A(n1032), .B(n1246), .Z(n2195) );
  AND U2699 ( .A(n1244), .B(n969), .Z(n2079) );
  XNOR U2700 ( .A(n2085), .B(n2086), .Z(n2082) );
  NANDN U2701 ( .B(n834), .A(n1419), .Z(n2086) );
  XNOR U2702 ( .A(n2084), .B(n2202), .Z(n2085) );
  ANDN U2703 ( .A(n904), .B(n1421), .Z(n2202) );
  XNOR U2704 ( .A(n2096), .B(n2087), .Z(n2193) );
  XOR U2705 ( .A(n2209), .B(n2105), .Z(n2096) );
  XNOR U2706 ( .A(n2093), .B(n2094), .Z(n2105) );
  NAND U2707 ( .A(n1085), .B(n1203), .Z(n2094) );
  XNOR U2708 ( .A(n2092), .B(n2210), .Z(n2093) );
  ANDN U2709 ( .A(n1210), .B(n1087), .Z(n2210) );
  XNOR U2710 ( .A(n2104), .B(n2095), .Z(n2209) );
  XOR U2711 ( .A(n2217), .B(n2101), .Z(n2104) );
  XNOR U2712 ( .A(n2100), .B(n2218), .Z(n2101) );
  ANDN U2713 ( .A(n1394), .B(n946), .Z(n2218) );
  AND U2714 ( .A(n944), .B(n1387), .Z(n2102) );
  XNOR U2715 ( .A(n2113), .B(n2112), .Z(n2089) );
  XOR U2716 ( .A(n2225), .B(n2121), .Z(n2112) );
  XNOR U2717 ( .A(n2109), .B(n2110), .Z(n2121) );
  NANDN U2718 ( .B(n647), .A(n1809), .Z(n2110) );
  XNOR U2719 ( .A(n2108), .B(n2226), .Z(n2109) );
  ANDN U2720 ( .A(n688), .B(n1811), .Z(n2226) );
  XNOR U2721 ( .A(n2120), .B(n2111), .Z(n2225) );
  XOR U2722 ( .A(n2233), .B(n2117), .Z(n2120) );
  XNOR U2723 ( .A(n2116), .B(n2234), .Z(n2117) );
  ANDN U2724 ( .A(n795), .B(n1614), .Z(n2234) );
  AND U2725 ( .A(n1612), .B(n741), .Z(n2118) );
  XOR U2726 ( .A(n2129), .B(n2128), .Z(n2113) );
  XOR U2727 ( .A(n2241), .B(n2125), .Z(n2128) );
  XNOR U2728 ( .A(n2124), .B(n2242), .Z(n2125) );
  ANDN U2729 ( .A(n620), .B(n2024), .Z(n2242) );
  AND U2730 ( .A(n2022), .B(n579), .Z(n2126) );
  XOR U2731 ( .A(n2136), .B(n2135), .Z(n2129) );
  NAND U2732 ( .A(n2249), .B(n523), .Z(n2135) );
  XNOR U2733 ( .A(n2134), .B(n2250), .Z(n2136) );
  ANDN U2734 ( .A(n554), .B(n2251), .Z(n2250) );
  NAND U2735 ( .A(n2252), .B(n2253), .Z(n2134) );
  NAND U2736 ( .A(n2254), .B(n2255), .Z(n2252) );
  IV U2737 ( .A(n2137), .Z(n2138) );
  MUX U2738 ( .IN0(o[5]), .IN1(n395), .SEL(n475), .F(\_MxM/n304 ) );
  XOR U2739 ( .A(n2260), .B(\_MxM/Y0[6] ), .Z(n395) );
  XOR U2740 ( .A(n2261), .B(n2262), .Z(n2260) );
  AND U2741 ( .A(n487), .B(n2264), .Z(n2263) );
  XOR U2742 ( .A(n2258), .B(n2262), .Z(n2264) );
  XOR U2743 ( .A(n2257), .B(n2262), .Z(n2258) );
  XNOR U2744 ( .A(n2265), .B(n2188), .Z(n2183) );
  XNOR U2745 ( .A(n2156), .B(n2155), .Z(n2188) );
  XOR U2746 ( .A(n2266), .B(n2160), .Z(n2155) );
  XNOR U2747 ( .A(n2151), .B(n2153), .Z(n2160) );
  NAND U2748 ( .A(n1934), .B(n667), .Z(n2153) );
  XNOR U2749 ( .A(n2149), .B(n2267), .Z(n2151) );
  ANDN U2750 ( .A(n1939), .B(n669), .Z(n2267) );
  XNOR U2751 ( .A(n2159), .B(n2154), .Z(n2266) );
  XOR U2752 ( .A(n2274), .B(n2166), .Z(n2159) );
  XNOR U2753 ( .A(n2164), .B(n2275), .Z(n2166) );
  ANDN U2754 ( .A(n2169), .B(n585), .Z(n2275) );
  XOR U2755 ( .A(n2276), .B(n2277), .Z(n2164) );
  AND U2756 ( .A(n2278), .B(n2279), .Z(n2277) );
  XNOR U2757 ( .A(n2280), .B(n2276), .Z(n2279) );
  AND U2758 ( .A(n2162), .B(n583), .Z(n2168) );
  XNOR U2759 ( .A(n2177), .B(n2176), .Z(n2156) );
  XOR U2760 ( .A(n2284), .B(n2173), .Z(n2176) );
  XNOR U2761 ( .A(n2172), .B(n2285), .Z(n2173) );
  ANDN U2762 ( .A(n1740), .B(n755), .Z(n2285) );
  AND U2763 ( .A(n1733), .B(n753), .Z(n2174) );
  XNOR U2764 ( .A(n2180), .B(n2181), .Z(n2177) );
  NAND U2765 ( .A(n1538), .B(n876), .Z(n2181) );
  XNOR U2766 ( .A(n2179), .B(n2292), .Z(n2180) );
  ANDN U2767 ( .A(n1543), .B(n878), .Z(n2292) );
  XNOR U2768 ( .A(n2187), .B(n2182), .Z(n2265) );
  XOR U2769 ( .A(n2186), .B(n2299), .Z(n2187) );
  AND U2770 ( .A(n2190), .B(n2300), .Z(n2299) );
  AND U2771 ( .A(n2301), .B(n2302), .Z(n2300) );
  NANDN U2772 ( .B(n2303), .A(n522), .Z(n2302) );
  NAND U2773 ( .A(n2304), .B(n2305), .Z(n2301) );
  ANDN U2774 ( .A(n2192), .B(n2191), .Z(n2190) );
  ANDN U2775 ( .A(n2306), .B(n2307), .Z(n2191) );
  OR U2776 ( .A(n2308), .B(n2309), .Z(n2192) );
  XNOR U2777 ( .A(n2208), .B(n2207), .Z(n2184) );
  XOR U2778 ( .A(n2313), .B(n2216), .Z(n2207) );
  XNOR U2779 ( .A(n2201), .B(n2200), .Z(n2216) );
  XOR U2780 ( .A(n2314), .B(n2197), .Z(n2200) );
  XNOR U2781 ( .A(n2196), .B(n2315), .Z(n2197) );
  ANDN U2782 ( .A(n1032), .B(n1330), .Z(n2315) );
  AND U2783 ( .A(n1328), .B(n969), .Z(n2198) );
  XNOR U2784 ( .A(n2204), .B(n2205), .Z(n2201) );
  NANDN U2785 ( .B(n834), .A(n1516), .Z(n2205) );
  XNOR U2786 ( .A(n2203), .B(n2322), .Z(n2204) );
  ANDN U2787 ( .A(n904), .B(n1518), .Z(n2322) );
  XNOR U2788 ( .A(n2215), .B(n2206), .Z(n2313) );
  XOR U2789 ( .A(n2329), .B(n2224), .Z(n2215) );
  XNOR U2790 ( .A(n2212), .B(n2213), .Z(n2224) );
  NAND U2791 ( .A(n1163), .B(n1203), .Z(n2213) );
  XNOR U2792 ( .A(n2211), .B(n2330), .Z(n2212) );
  ANDN U2793 ( .A(n1210), .B(n1165), .Z(n2330) );
  XNOR U2794 ( .A(n2223), .B(n2214), .Z(n2329) );
  XOR U2795 ( .A(n2337), .B(n2220), .Z(n2223) );
  XNOR U2796 ( .A(n2219), .B(n2338), .Z(n2220) );
  ANDN U2797 ( .A(n1394), .B(n1013), .Z(n2338) );
  AND U2798 ( .A(n1011), .B(n1387), .Z(n2221) );
  XNOR U2799 ( .A(n2232), .B(n2231), .Z(n2208) );
  XOR U2800 ( .A(n2345), .B(n2240), .Z(n2231) );
  XNOR U2801 ( .A(n2228), .B(n2229), .Z(n2240) );
  NANDN U2802 ( .B(n647), .A(n1915), .Z(n2229) );
  XNOR U2803 ( .A(n2227), .B(n2346), .Z(n2228) );
  ANDN U2804 ( .A(n688), .B(n1917), .Z(n2346) );
  XNOR U2805 ( .A(n2239), .B(n2230), .Z(n2345) );
  XOR U2806 ( .A(n2353), .B(n2236), .Z(n2239) );
  XNOR U2807 ( .A(n2235), .B(n2354), .Z(n2236) );
  ANDN U2808 ( .A(n795), .B(n1710), .Z(n2354) );
  AND U2809 ( .A(n1708), .B(n741), .Z(n2237) );
  XOR U2810 ( .A(n2248), .B(n2247), .Z(n2232) );
  XOR U2811 ( .A(n2361), .B(n2244), .Z(n2247) );
  XNOR U2812 ( .A(n2243), .B(n2362), .Z(n2244) );
  ANDN U2813 ( .A(n620), .B(n2132), .Z(n2362) );
  AND U2814 ( .A(n2130), .B(n579), .Z(n2245) );
  XOR U2815 ( .A(n2255), .B(n2254), .Z(n2248) );
  NAND U2816 ( .A(n2369), .B(n523), .Z(n2254) );
  XOR U2817 ( .A(n2253), .B(n2370), .Z(n2255) );
  ANDN U2818 ( .A(n554), .B(n2371), .Z(n2370) );
  ANDN U2819 ( .A(n2372), .B(n2373), .Z(n2253) );
  NAND U2820 ( .A(n2374), .B(n2375), .Z(n2372) );
  IV U2821 ( .A(n2256), .Z(n2257) );
  MUX U2822 ( .IN0(o[4]), .IN1(n392), .SEL(n475), .F(\_MxM/n303 ) );
  XOR U2823 ( .A(n2380), .B(\_MxM/Y0[5] ), .Z(n392) );
  XOR U2824 ( .A(n2381), .B(n2382), .Z(n2380) );
  AND U2825 ( .A(n487), .B(n2384), .Z(n2383) );
  XOR U2826 ( .A(n2378), .B(n2382), .Z(n2384) );
  XOR U2827 ( .A(n2377), .B(n2382), .Z(n2378) );
  XNOR U2828 ( .A(n2385), .B(n2312), .Z(n2297) );
  XNOR U2829 ( .A(n2273), .B(n2272), .Z(n2312) );
  XOR U2830 ( .A(n2386), .B(n2283), .Z(n2272) );
  XNOR U2831 ( .A(n2269), .B(n2270), .Z(n2283) );
  NAND U2832 ( .A(n1934), .B(n711), .Z(n2270) );
  XNOR U2833 ( .A(n2268), .B(n2387), .Z(n2269) );
  ANDN U2834 ( .A(n1939), .B(n713), .Z(n2387) );
  XNOR U2835 ( .A(n2282), .B(n2271), .Z(n2386) );
  XOR U2836 ( .A(n2394), .B(n2278), .Z(n2282) );
  XNOR U2837 ( .A(n2276), .B(n2395), .Z(n2278) );
  ANDN U2838 ( .A(n2169), .B(n629), .Z(n2395) );
  XOR U2839 ( .A(n2396), .B(n2397), .Z(n2276) );
  AND U2840 ( .A(n2398), .B(n2399), .Z(n2397) );
  XNOR U2841 ( .A(n2400), .B(n2396), .Z(n2399) );
  AND U2842 ( .A(n2162), .B(n627), .Z(n2280) );
  XNOR U2843 ( .A(n2291), .B(n2290), .Z(n2273) );
  XOR U2844 ( .A(n2404), .B(n2287), .Z(n2290) );
  XNOR U2845 ( .A(n2286), .B(n2405), .Z(n2287) );
  ANDN U2846 ( .A(n1740), .B(n814), .Z(n2405) );
  AND U2847 ( .A(n1733), .B(n812), .Z(n2288) );
  XNOR U2848 ( .A(n2294), .B(n2295), .Z(n2291) );
  NAND U2849 ( .A(n1538), .B(n944), .Z(n2295) );
  XNOR U2850 ( .A(n2293), .B(n2412), .Z(n2294) );
  ANDN U2851 ( .A(n1543), .B(n946), .Z(n2412) );
  XOR U2852 ( .A(n2311), .B(n2296), .Z(n2385) );
  XOR U2853 ( .A(n2419), .B(n2304), .Z(n2311) );
  XOR U2854 ( .A(n2423), .B(n2309), .Z(n2307) );
  NAND U2855 ( .A(n2424), .B(n552), .Z(n2309) );
  NAND U2856 ( .A(n2425), .B(n2308), .Z(n2423) );
  NANDN U2857 ( .B(n555), .A(n2429), .Z(n2425) );
  ANDN U2858 ( .A(n2430), .B(n2431), .Z(n2305) );
  XNOR U2859 ( .A(n2328), .B(n2327), .Z(n2298) );
  XOR U2860 ( .A(n2435), .B(n2336), .Z(n2327) );
  XNOR U2861 ( .A(n2321), .B(n2320), .Z(n2336) );
  XOR U2862 ( .A(n2436), .B(n2317), .Z(n2320) );
  XNOR U2863 ( .A(n2316), .B(n2437), .Z(n2317) );
  ANDN U2864 ( .A(n1032), .B(n1421), .Z(n2437) );
  AND U2865 ( .A(n1419), .B(n969), .Z(n2318) );
  XNOR U2866 ( .A(n2324), .B(n2325), .Z(n2321) );
  NANDN U2867 ( .B(n834), .A(n1612), .Z(n2325) );
  XNOR U2868 ( .A(n2323), .B(n2444), .Z(n2324) );
  ANDN U2869 ( .A(n904), .B(n1614), .Z(n2444) );
  XNOR U2870 ( .A(n2335), .B(n2326), .Z(n2435) );
  XOR U2871 ( .A(n2451), .B(n2344), .Z(n2335) );
  XNOR U2872 ( .A(n2332), .B(n2333), .Z(n2344) );
  NAND U2873 ( .A(n1244), .B(n1203), .Z(n2333) );
  XNOR U2874 ( .A(n2331), .B(n2452), .Z(n2332) );
  ANDN U2875 ( .A(n1210), .B(n1246), .Z(n2452) );
  XNOR U2876 ( .A(n2343), .B(n2334), .Z(n2451) );
  XOR U2877 ( .A(n2459), .B(n2340), .Z(n2343) );
  XNOR U2878 ( .A(n2339), .B(n2460), .Z(n2340) );
  ANDN U2879 ( .A(n1394), .B(n1087), .Z(n2460) );
  AND U2880 ( .A(n1085), .B(n1387), .Z(n2341) );
  XNOR U2881 ( .A(n2352), .B(n2351), .Z(n2328) );
  XOR U2882 ( .A(n2467), .B(n2360), .Z(n2351) );
  XNOR U2883 ( .A(n2348), .B(n2349), .Z(n2360) );
  NANDN U2884 ( .B(n647), .A(n2022), .Z(n2349) );
  XNOR U2885 ( .A(n2347), .B(n2468), .Z(n2348) );
  ANDN U2886 ( .A(n688), .B(n2024), .Z(n2468) );
  XNOR U2887 ( .A(n2359), .B(n2350), .Z(n2467) );
  XOR U2888 ( .A(n2475), .B(n2356), .Z(n2359) );
  XNOR U2889 ( .A(n2355), .B(n2476), .Z(n2356) );
  ANDN U2890 ( .A(n795), .B(n1811), .Z(n2476) );
  AND U2891 ( .A(n1809), .B(n741), .Z(n2357) );
  XOR U2892 ( .A(n2368), .B(n2367), .Z(n2352) );
  XOR U2893 ( .A(n2483), .B(n2364), .Z(n2367) );
  XNOR U2894 ( .A(n2363), .B(n2484), .Z(n2364) );
  ANDN U2895 ( .A(n620), .B(n2251), .Z(n2484) );
  AND U2896 ( .A(n2249), .B(n579), .Z(n2365) );
  XOR U2897 ( .A(n2375), .B(n2374), .Z(n2368) );
  NAND U2898 ( .A(n2491), .B(n523), .Z(n2374) );
  XNOR U2899 ( .A(n2373), .B(n2492), .Z(n2375) );
  ANDN U2900 ( .A(n554), .B(n2493), .Z(n2492) );
  NAND U2901 ( .A(n2494), .B(n2495), .Z(n2373) );
  NAND U2902 ( .A(n2496), .B(n2497), .Z(n2494) );
  IV U2903 ( .A(n2376), .Z(n2377) );
  MUX U2904 ( .IN0(o[3]), .IN1(n389), .SEL(n475), .F(\_MxM/n302 ) );
  XNOR U2905 ( .A(n2501), .B(\_MxM/Y0[4] ), .Z(n389) );
  XNOR U2906 ( .A(n2503), .B(n2504), .Z(n2501) );
  XOR U2907 ( .A(n2502), .B(n2505), .Z(n2503) );
  AND U2908 ( .A(n487), .B(n2506), .Z(n2505) );
  XNOR U2909 ( .A(n2499), .B(n2504), .Z(n2506) );
  XOR U2910 ( .A(n2504), .B(n2498), .Z(n2499) );
  NOR U2911 ( .A(n2507), .B(n2508), .Z(n2498) );
  XNOR U2912 ( .A(n2509), .B(n2434), .Z(n2417) );
  XNOR U2913 ( .A(n2393), .B(n2392), .Z(n2434) );
  XOR U2914 ( .A(n2510), .B(n2403), .Z(n2392) );
  XNOR U2915 ( .A(n2389), .B(n2390), .Z(n2403) );
  NAND U2916 ( .A(n1934), .B(n753), .Z(n2390) );
  XNOR U2917 ( .A(n2388), .B(n2511), .Z(n2389) );
  ANDN U2918 ( .A(n1939), .B(n755), .Z(n2511) );
  XNOR U2919 ( .A(n2402), .B(n2391), .Z(n2510) );
  XOR U2920 ( .A(n2518), .B(n2398), .Z(n2402) );
  XNOR U2921 ( .A(n2396), .B(n2519), .Z(n2398) );
  ANDN U2922 ( .A(n2169), .B(n669), .Z(n2519) );
  AND U2923 ( .A(n2162), .B(n667), .Z(n2400) );
  XNOR U2924 ( .A(n2411), .B(n2410), .Z(n2393) );
  XOR U2925 ( .A(n2526), .B(n2407), .Z(n2410) );
  XNOR U2926 ( .A(n2406), .B(n2527), .Z(n2407) );
  ANDN U2927 ( .A(n1740), .B(n878), .Z(n2527) );
  AND U2928 ( .A(n1733), .B(n876), .Z(n2408) );
  XNOR U2929 ( .A(n2414), .B(n2415), .Z(n2411) );
  NAND U2930 ( .A(n1538), .B(n1011), .Z(n2415) );
  XNOR U2931 ( .A(n2413), .B(n2534), .Z(n2414) );
  ANDN U2932 ( .A(n1543), .B(n1013), .Z(n2534) );
  XNOR U2933 ( .A(n2433), .B(n2416), .Z(n2509) );
  XOR U2934 ( .A(n2541), .B(n2431), .Z(n2433) );
  XOR U2935 ( .A(n2422), .B(n2421), .Z(n2431) );
  XNOR U2936 ( .A(n2420), .B(n2542), .Z(n2421) );
  AND U2937 ( .A(n2543), .B(n2544), .Z(n2542) );
  NANDN U2938 ( .B(n2545), .A(n522), .Z(n2544) );
  NANDN U2939 ( .B(n2546), .A(n2547), .Z(n2543) );
  XNOR U2940 ( .A(n2427), .B(n2428), .Z(n2422) );
  NAND U2941 ( .A(n2424), .B(n583), .Z(n2428) );
  XNOR U2942 ( .A(n2426), .B(n2551), .Z(n2427) );
  ANDN U2943 ( .A(n2429), .B(n585), .Z(n2551) );
  NOR U2944 ( .A(n2555), .B(n2556), .Z(n2430) );
  XNOR U2945 ( .A(n2450), .B(n2449), .Z(n2418) );
  XOR U2946 ( .A(n2560), .B(n2458), .Z(n2449) );
  XNOR U2947 ( .A(n2443), .B(n2442), .Z(n2458) );
  XOR U2948 ( .A(n2561), .B(n2439), .Z(n2442) );
  XNOR U2949 ( .A(n2438), .B(n2562), .Z(n2439) );
  ANDN U2950 ( .A(n1032), .B(n1518), .Z(n2562) );
  AND U2951 ( .A(n1516), .B(n969), .Z(n2440) );
  XNOR U2952 ( .A(n2446), .B(n2447), .Z(n2443) );
  NANDN U2953 ( .B(n834), .A(n1708), .Z(n2447) );
  XNOR U2954 ( .A(n2445), .B(n2569), .Z(n2446) );
  ANDN U2955 ( .A(n904), .B(n1710), .Z(n2569) );
  XNOR U2956 ( .A(n2457), .B(n2448), .Z(n2560) );
  XOR U2957 ( .A(n2576), .B(n2466), .Z(n2457) );
  XNOR U2958 ( .A(n2454), .B(n2455), .Z(n2466) );
  NAND U2959 ( .A(n1328), .B(n1203), .Z(n2455) );
  XNOR U2960 ( .A(n2453), .B(n2577), .Z(n2454) );
  ANDN U2961 ( .A(n1210), .B(n1330), .Z(n2577) );
  XNOR U2962 ( .A(n2465), .B(n2456), .Z(n2576) );
  XOR U2963 ( .A(n2584), .B(n2462), .Z(n2465) );
  XNOR U2964 ( .A(n2461), .B(n2585), .Z(n2462) );
  ANDN U2965 ( .A(n1394), .B(n1165), .Z(n2585) );
  AND U2966 ( .A(n1163), .B(n1387), .Z(n2463) );
  XNOR U2967 ( .A(n2474), .B(n2473), .Z(n2450) );
  XOR U2968 ( .A(n2592), .B(n2482), .Z(n2473) );
  XNOR U2969 ( .A(n2470), .B(n2471), .Z(n2482) );
  NANDN U2970 ( .B(n647), .A(n2130), .Z(n2471) );
  XNOR U2971 ( .A(n2469), .B(n2593), .Z(n2470) );
  ANDN U2972 ( .A(n688), .B(n2132), .Z(n2593) );
  XNOR U2973 ( .A(n2481), .B(n2472), .Z(n2592) );
  XOR U2974 ( .A(n2600), .B(n2478), .Z(n2481) );
  XNOR U2975 ( .A(n2477), .B(n2601), .Z(n2478) );
  ANDN U2976 ( .A(n795), .B(n1917), .Z(n2601) );
  AND U2977 ( .A(n1915), .B(n741), .Z(n2479) );
  XOR U2978 ( .A(n2490), .B(n2489), .Z(n2474) );
  XOR U2979 ( .A(n2608), .B(n2486), .Z(n2489) );
  XNOR U2980 ( .A(n2485), .B(n2609), .Z(n2486) );
  ANDN U2981 ( .A(n620), .B(n2371), .Z(n2609) );
  AND U2982 ( .A(n2369), .B(n579), .Z(n2487) );
  XOR U2983 ( .A(n2497), .B(n2496), .Z(n2490) );
  NAND U2984 ( .A(n2616), .B(n523), .Z(n2496) );
  XOR U2985 ( .A(n2495), .B(n2617), .Z(n2497) );
  ANDN U2986 ( .A(n554), .B(n2618), .Z(n2617) );
  ANDN U2987 ( .A(n2619), .B(n2620), .Z(n2495) );
  NAND U2988 ( .A(n2621), .B(n2622), .Z(n2619) );
  IV U2989 ( .A(n2500), .Z(n2502) );
  MUX U2990 ( .IN0(o[2]), .IN1(n386), .SEL(n475), .F(\_MxM/n301 ) );
  IV U2991 ( .A(n2626), .Z(n475) );
  XNOR U2992 ( .A(n2624), .B(\_MxM/Y0[3] ), .Z(n386) );
  XNOR U2993 ( .A(n2627), .B(n2628), .Z(n2624) );
  XOR U2994 ( .A(n2625), .B(n2629), .Z(n2627) );
  AND U2995 ( .A(n487), .B(n2630), .Z(n2629) );
  XNOR U2996 ( .A(n2508), .B(n2628), .Z(n2630) );
  NANDN U2997 ( .B(n2631), .A(n2632), .Z(n2507) );
  XNOR U2998 ( .A(n2633), .B(n2559), .Z(n2539) );
  XNOR U2999 ( .A(n2517), .B(n2516), .Z(n2559) );
  XOR U3000 ( .A(n2634), .B(n2525), .Z(n2516) );
  XNOR U3001 ( .A(n2513), .B(n2514), .Z(n2525) );
  NAND U3002 ( .A(n1934), .B(n812), .Z(n2514) );
  XNOR U3003 ( .A(n2512), .B(n2635), .Z(n2513) );
  ANDN U3004 ( .A(n1939), .B(n814), .Z(n2635) );
  XNOR U3005 ( .A(n2524), .B(n2515), .Z(n2634) );
  XOR U3006 ( .A(n2642), .B(n2521), .Z(n2524) );
  XNOR U3007 ( .A(n2520), .B(n2643), .Z(n2521) );
  ANDN U3008 ( .A(n2169), .B(n713), .Z(n2643) );
  AND U3009 ( .A(n2162), .B(n711), .Z(n2522) );
  XNOR U3010 ( .A(n2533), .B(n2532), .Z(n2517) );
  XOR U3011 ( .A(n2650), .B(n2529), .Z(n2532) );
  XNOR U3012 ( .A(n2528), .B(n2651), .Z(n2529) );
  ANDN U3013 ( .A(n1740), .B(n946), .Z(n2651) );
  AND U3014 ( .A(n1733), .B(n944), .Z(n2530) );
  XNOR U3015 ( .A(n2536), .B(n2537), .Z(n2533) );
  NAND U3016 ( .A(n1538), .B(n1085), .Z(n2537) );
  XNOR U3017 ( .A(n2535), .B(n2658), .Z(n2536) );
  ANDN U3018 ( .A(n1543), .B(n1087), .Z(n2658) );
  XNOR U3019 ( .A(n2558), .B(n2538), .Z(n2633) );
  XOR U3020 ( .A(n2665), .B(n2556), .Z(n2558) );
  XOR U3021 ( .A(n2550), .B(n2549), .Z(n2556) );
  XOR U3022 ( .A(n2670), .B(n2547), .Z(n2666) );
  AND U3023 ( .A(n2671), .B(n552), .Z(n2547) );
  NAND U3024 ( .A(n2672), .B(n2546), .Z(n2670) );
  XOR U3025 ( .A(n2673), .B(n2674), .Z(n2546) );
  AND U3026 ( .A(n2675), .B(n2676), .Z(n2674) );
  XNOR U3027 ( .A(n2677), .B(n2673), .Z(n2676) );
  NANDN U3028 ( .B(n555), .A(n2678), .Z(n2672) );
  XNOR U3029 ( .A(n2553), .B(n2554), .Z(n2550) );
  NAND U3030 ( .A(n2424), .B(n627), .Z(n2554) );
  XNOR U3031 ( .A(n2552), .B(n2679), .Z(n2553) );
  ANDN U3032 ( .A(n2429), .B(n629), .Z(n2679) );
  XOR U3033 ( .A(n2680), .B(n2681), .Z(n2552) );
  AND U3034 ( .A(n2682), .B(n2683), .Z(n2681) );
  XOR U3035 ( .A(n2684), .B(n2680), .Z(n2683) );
  XNOR U3036 ( .A(n2555), .B(n2557), .Z(n2665) );
  XNOR U3037 ( .A(n2688), .B(n2691), .Z(n2690) );
  XNOR U3038 ( .A(n2575), .B(n2574), .Z(n2540) );
  XOR U3039 ( .A(n2692), .B(n2583), .Z(n2574) );
  XNOR U3040 ( .A(n2568), .B(n2567), .Z(n2583) );
  XOR U3041 ( .A(n2693), .B(n2564), .Z(n2567) );
  XNOR U3042 ( .A(n2563), .B(n2694), .Z(n2564) );
  ANDN U3043 ( .A(n1032), .B(n1614), .Z(n2694) );
  AND U3044 ( .A(n1612), .B(n969), .Z(n2565) );
  XNOR U3045 ( .A(n2571), .B(n2572), .Z(n2568) );
  NANDN U3046 ( .B(n834), .A(n1809), .Z(n2572) );
  XNOR U3047 ( .A(n2570), .B(n2701), .Z(n2571) );
  ANDN U3048 ( .A(n904), .B(n1811), .Z(n2701) );
  XNOR U3049 ( .A(n2582), .B(n2573), .Z(n2692) );
  XOR U3050 ( .A(n2708), .B(n2591), .Z(n2582) );
  XNOR U3051 ( .A(n2579), .B(n2580), .Z(n2591) );
  NAND U3052 ( .A(n1419), .B(n1203), .Z(n2580) );
  XNOR U3053 ( .A(n2578), .B(n2709), .Z(n2579) );
  ANDN U3054 ( .A(n1210), .B(n1421), .Z(n2709) );
  XNOR U3055 ( .A(n2590), .B(n2581), .Z(n2708) );
  XOR U3056 ( .A(n2716), .B(n2587), .Z(n2590) );
  XNOR U3057 ( .A(n2586), .B(n2717), .Z(n2587) );
  ANDN U3058 ( .A(n1394), .B(n1246), .Z(n2717) );
  AND U3059 ( .A(n1244), .B(n1387), .Z(n2588) );
  XNOR U3060 ( .A(n2599), .B(n2598), .Z(n2575) );
  XOR U3061 ( .A(n2724), .B(n2607), .Z(n2598) );
  XNOR U3062 ( .A(n2595), .B(n2596), .Z(n2607) );
  NANDN U3063 ( .B(n647), .A(n2249), .Z(n2596) );
  XNOR U3064 ( .A(n2594), .B(n2725), .Z(n2595) );
  ANDN U3065 ( .A(n688), .B(n2251), .Z(n2725) );
  XNOR U3066 ( .A(n2606), .B(n2597), .Z(n2724) );
  XOR U3067 ( .A(n2732), .B(n2603), .Z(n2606) );
  XNOR U3068 ( .A(n2602), .B(n2733), .Z(n2603) );
  ANDN U3069 ( .A(n795), .B(n2024), .Z(n2733) );
  AND U3070 ( .A(n2022), .B(n741), .Z(n2604) );
  XOR U3071 ( .A(n2615), .B(n2614), .Z(n2599) );
  XOR U3072 ( .A(n2740), .B(n2611), .Z(n2614) );
  XNOR U3073 ( .A(n2610), .B(n2741), .Z(n2611) );
  ANDN U3074 ( .A(n620), .B(n2493), .Z(n2741) );
  AND U3075 ( .A(n2491), .B(n579), .Z(n2612) );
  XOR U3076 ( .A(n2622), .B(n2621), .Z(n2615) );
  NAND U3077 ( .A(n2748), .B(n523), .Z(n2621) );
  XNOR U3078 ( .A(n2620), .B(n2749), .Z(n2622) );
  ANDN U3079 ( .A(n554), .B(n2750), .Z(n2749) );
  NAND U3080 ( .A(n2751), .B(n2752), .Z(n2620) );
  NAND U3081 ( .A(n2753), .B(n2754), .Z(n2751) );
  IV U3082 ( .A(n2623), .Z(n2625) );
  MUX U3083 ( .IN0(n383), .IN1(o[1]), .SEL(n2626), .F(\_MxM/n300 ) );
  XNOR U3084 ( .A(n2756), .B(\_MxM/Y0[2] ), .Z(n383) );
  XNOR U3085 ( .A(n2757), .B(n2758), .Z(n2756) );
  XNOR U3086 ( .A(n2755), .B(n2759), .Z(n2757) );
  AND U3087 ( .A(n487), .B(n2760), .Z(n2759) );
  XNOR U3088 ( .A(n2631), .B(n2758), .Z(n2760) );
  XOR U3089 ( .A(n2758), .B(n2632), .Z(n2631) );
  ANDN U3090 ( .A(n2761), .B(n2762), .Z(n2632) );
  XNOR U3091 ( .A(n2763), .B(n2687), .Z(n2663) );
  XNOR U3092 ( .A(n2641), .B(n2640), .Z(n2687) );
  XOR U3093 ( .A(n2764), .B(n2649), .Z(n2640) );
  XNOR U3094 ( .A(n2637), .B(n2638), .Z(n2649) );
  NAND U3095 ( .A(n1934), .B(n876), .Z(n2638) );
  XNOR U3096 ( .A(n2636), .B(n2765), .Z(n2637) );
  ANDN U3097 ( .A(n1939), .B(n878), .Z(n2765) );
  XNOR U3098 ( .A(n2648), .B(n2639), .Z(n2764) );
  XOR U3099 ( .A(n2772), .B(n2645), .Z(n2648) );
  XNOR U3100 ( .A(n2644), .B(n2773), .Z(n2645) );
  ANDN U3101 ( .A(n2169), .B(n755), .Z(n2773) );
  AND U3102 ( .A(n2162), .B(n753), .Z(n2646) );
  XNOR U3103 ( .A(n2657), .B(n2656), .Z(n2641) );
  XOR U3104 ( .A(n2780), .B(n2653), .Z(n2656) );
  XNOR U3105 ( .A(n2652), .B(n2781), .Z(n2653) );
  ANDN U3106 ( .A(n1740), .B(n1013), .Z(n2781) );
  AND U3107 ( .A(n1733), .B(n1011), .Z(n2654) );
  XNOR U3108 ( .A(n2660), .B(n2661), .Z(n2657) );
  NAND U3109 ( .A(n1538), .B(n1163), .Z(n2661) );
  XNOR U3110 ( .A(n2659), .B(n2788), .Z(n2660) );
  ANDN U3111 ( .A(n1543), .B(n1165), .Z(n2788) );
  XOR U3112 ( .A(n2686), .B(n2662), .Z(n2763) );
  XNOR U3113 ( .A(n2795), .B(n2691), .Z(n2686) );
  XNOR U3114 ( .A(n2669), .B(n2668), .Z(n2691) );
  XOR U3115 ( .A(n2796), .B(n2675), .Z(n2668) );
  XNOR U3116 ( .A(n2673), .B(n2797), .Z(n2675) );
  ANDN U3117 ( .A(n2678), .B(n585), .Z(n2797) );
  AND U3118 ( .A(n2671), .B(n583), .Z(n2677) );
  XNOR U3119 ( .A(n2682), .B(n2684), .Z(n2669) );
  NAND U3120 ( .A(n2424), .B(n667), .Z(n2684) );
  XNOR U3121 ( .A(n2680), .B(n2804), .Z(n2682) );
  ANDN U3122 ( .A(n2429), .B(n669), .Z(n2804) );
  XNOR U3123 ( .A(n2689), .B(n2685), .Z(n2795) );
  XOR U3124 ( .A(n2688), .B(n2811), .Z(n2689) );
  AND U3125 ( .A(n2812), .B(n2813), .Z(n2811) );
  NANDN U3126 ( .B(n2814), .A(n2815), .Z(n2813) );
  AND U3127 ( .A(n2816), .B(n2817), .Z(n2812) );
  NANDN U3128 ( .B(n2818), .A(n522), .Z(n2817) );
  OR U3129 ( .A(n2819), .B(n2820), .Z(n2816) );
  XNOR U3130 ( .A(n2707), .B(n2706), .Z(n2664) );
  XOR U3131 ( .A(n2824), .B(n2715), .Z(n2706) );
  XNOR U3132 ( .A(n2700), .B(n2699), .Z(n2715) );
  XOR U3133 ( .A(n2825), .B(n2696), .Z(n2699) );
  XNOR U3134 ( .A(n2695), .B(n2826), .Z(n2696) );
  ANDN U3135 ( .A(n1032), .B(n1710), .Z(n2826) );
  AND U3136 ( .A(n1708), .B(n969), .Z(n2697) );
  XNOR U3137 ( .A(n2703), .B(n2704), .Z(n2700) );
  NANDN U3138 ( .B(n834), .A(n1915), .Z(n2704) );
  XNOR U3139 ( .A(n2702), .B(n2833), .Z(n2703) );
  ANDN U3140 ( .A(n904), .B(n1917), .Z(n2833) );
  XNOR U3141 ( .A(n2714), .B(n2705), .Z(n2824) );
  XOR U3142 ( .A(n2840), .B(n2723), .Z(n2714) );
  XNOR U3143 ( .A(n2711), .B(n2712), .Z(n2723) );
  NAND U3144 ( .A(n1516), .B(n1203), .Z(n2712) );
  XNOR U3145 ( .A(n2710), .B(n2841), .Z(n2711) );
  ANDN U3146 ( .A(n1210), .B(n1518), .Z(n2841) );
  XNOR U3147 ( .A(n2722), .B(n2713), .Z(n2840) );
  XOR U3148 ( .A(n2848), .B(n2719), .Z(n2722) );
  XNOR U3149 ( .A(n2718), .B(n2849), .Z(n2719) );
  ANDN U3150 ( .A(n1394), .B(n1330), .Z(n2849) );
  AND U3151 ( .A(n1328), .B(n1387), .Z(n2720) );
  XNOR U3152 ( .A(n2731), .B(n2730), .Z(n2707) );
  XOR U3153 ( .A(n2856), .B(n2739), .Z(n2730) );
  XNOR U3154 ( .A(n2727), .B(n2728), .Z(n2739) );
  NANDN U3155 ( .B(n647), .A(n2369), .Z(n2728) );
  XNOR U3156 ( .A(n2726), .B(n2857), .Z(n2727) );
  ANDN U3157 ( .A(n688), .B(n2371), .Z(n2857) );
  XNOR U3158 ( .A(n2738), .B(n2729), .Z(n2856) );
  XOR U3159 ( .A(n2864), .B(n2735), .Z(n2738) );
  XNOR U3160 ( .A(n2734), .B(n2865), .Z(n2735) );
  ANDN U3161 ( .A(n795), .B(n2132), .Z(n2865) );
  AND U3162 ( .A(n2130), .B(n741), .Z(n2736) );
  XOR U3163 ( .A(n2747), .B(n2746), .Z(n2731) );
  XOR U3164 ( .A(n2872), .B(n2743), .Z(n2746) );
  XNOR U3165 ( .A(n2742), .B(n2873), .Z(n2743) );
  ANDN U3166 ( .A(n620), .B(n2618), .Z(n2873) );
  AND U3167 ( .A(n2616), .B(n579), .Z(n2744) );
  XOR U3168 ( .A(n2754), .B(n2753), .Z(n2747) );
  NAND U3169 ( .A(n2880), .B(n523), .Z(n2753) );
  XOR U3170 ( .A(n2752), .B(n2881), .Z(n2754) );
  ANDN U3171 ( .A(n554), .B(n2882), .Z(n2881) );
  ANDN U3172 ( .A(n2883), .B(n2884), .Z(n2752) );
  NAND U3173 ( .A(n2885), .B(n2886), .Z(n2883) );
  MUX U3174 ( .IN0(n379), .IN1(o[0]), .SEL(n2626), .F(\_MxM/n299 ) );
  NANDN U3175 ( .B(rst), .A(n474), .Z(n2626) );
  AND U3176 ( .A(n2889), .B(n2890), .Z(n474) );
  AND U3177 ( .A(n2891), .B(n2892), .Z(n2890) );
  ANDN U3178 ( .A(n2893), .B(\_MxM/n[7] ), .Z(n2892) );
  NOR U3179 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n2893) );
  NOR U3180 ( .A(\_MxM/n[5] ), .B(\_MxM/n[6] ), .Z(n2891) );
  AND U3181 ( .A(n2894), .B(n2895), .Z(n2889) );
  NOR U3182 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n2895) );
  ANDN U3183 ( .A(n374), .B(\_MxM/n[0] ), .Z(n2894) );
  NOR U3184 ( .A(\_MxM/n[3] ), .B(\_MxM/n[4] ), .Z(n374) );
  XOR U3185 ( .A(n2888), .B(\_MxM/Y0[1] ), .Z(n379) );
  XOR U3186 ( .A(n2896), .B(n2897), .Z(n2888) );
  XOR U3187 ( .A(n2898), .B(n2887), .Z(n2896) );
  NAND U3188 ( .A(n2899), .B(n487), .Z(n2898) );
  XOR U3189 ( .A(e_input[31]), .B(g_input[31]), .Z(n487) );
  XOR U3190 ( .A(n2761), .B(n2897), .Z(n2899) );
  XOR U3191 ( .A(n2762), .B(n2897), .Z(n2761) );
  XNOR U3192 ( .A(n2900), .B(n2810), .Z(n2793) );
  XNOR U3193 ( .A(n2771), .B(n2770), .Z(n2810) );
  XOR U3194 ( .A(n2901), .B(n2779), .Z(n2770) );
  XNOR U3195 ( .A(n2767), .B(n2768), .Z(n2779) );
  NAND U3196 ( .A(n1934), .B(n944), .Z(n2768) );
  XNOR U3197 ( .A(n2766), .B(n2902), .Z(n2767) );
  ANDN U3198 ( .A(n1939), .B(n946), .Z(n2902) );
  XNOR U3199 ( .A(n2778), .B(n2769), .Z(n2901) );
  XOR U3200 ( .A(n2909), .B(n2775), .Z(n2778) );
  XNOR U3201 ( .A(n2774), .B(n2910), .Z(n2775) );
  ANDN U3202 ( .A(n2169), .B(n814), .Z(n2910) );
  AND U3203 ( .A(n2162), .B(n812), .Z(n2776) );
  XNOR U3204 ( .A(n2787), .B(n2786), .Z(n2771) );
  XOR U3205 ( .A(n2917), .B(n2783), .Z(n2786) );
  XNOR U3206 ( .A(n2782), .B(n2918), .Z(n2783) );
  ANDN U3207 ( .A(n1740), .B(n1087), .Z(n2918) );
  AND U3208 ( .A(n1733), .B(n1085), .Z(n2784) );
  XNOR U3209 ( .A(n2790), .B(n2791), .Z(n2787) );
  NAND U3210 ( .A(n1538), .B(n1244), .Z(n2791) );
  XNOR U3211 ( .A(n2789), .B(n2925), .Z(n2790) );
  ANDN U3212 ( .A(n1543), .B(n1246), .Z(n2925) );
  XOR U3213 ( .A(n2809), .B(n2792), .Z(n2900) );
  XNOR U3214 ( .A(n2932), .B(n2823), .Z(n2809) );
  XNOR U3215 ( .A(n2803), .B(n2802), .Z(n2823) );
  XOR U3216 ( .A(n2933), .B(n2799), .Z(n2802) );
  XNOR U3217 ( .A(n2798), .B(n2934), .Z(n2799) );
  ANDN U3218 ( .A(n2678), .B(n629), .Z(n2934) );
  AND U3219 ( .A(n2671), .B(n627), .Z(n2800) );
  XNOR U3220 ( .A(n2806), .B(n2807), .Z(n2803) );
  NAND U3221 ( .A(n2424), .B(n711), .Z(n2807) );
  XNOR U3222 ( .A(n2805), .B(n2941), .Z(n2806) );
  ANDN U3223 ( .A(n2429), .B(n713), .Z(n2941) );
  XOR U3224 ( .A(n2822), .B(n2808), .Z(n2932) );
  XNOR U3225 ( .A(n2948), .B(n2819), .Z(n2822) );
  XNOR U3226 ( .A(n2949), .B(n2815), .Z(n2819) );
  AND U3227 ( .A(n2950), .B(n552), .Z(n2815) );
  NAND U3228 ( .A(n2951), .B(n2814), .Z(n2949) );
  NANDN U3229 ( .B(n555), .A(n2955), .Z(n2951) );
  XNOR U3230 ( .A(n2820), .B(n2821), .Z(n2948) );
  XNOR U3231 ( .A(n2959), .B(n2962), .Z(n2961) );
  XNOR U3232 ( .A(n2839), .B(n2838), .Z(n2794) );
  XOR U3233 ( .A(n2963), .B(n2847), .Z(n2838) );
  XNOR U3234 ( .A(n2832), .B(n2831), .Z(n2847) );
  XOR U3235 ( .A(n2964), .B(n2828), .Z(n2831) );
  XNOR U3236 ( .A(n2827), .B(n2965), .Z(n2828) );
  ANDN U3237 ( .A(n1032), .B(n1811), .Z(n2965) );
  AND U3238 ( .A(n1809), .B(n969), .Z(n2829) );
  XNOR U3239 ( .A(n2835), .B(n2836), .Z(n2832) );
  NANDN U3240 ( .B(n834), .A(n2022), .Z(n2836) );
  XNOR U3241 ( .A(n2834), .B(n2972), .Z(n2835) );
  ANDN U3242 ( .A(n904), .B(n2024), .Z(n2972) );
  XNOR U3243 ( .A(n2846), .B(n2837), .Z(n2963) );
  XOR U3244 ( .A(n2979), .B(n2855), .Z(n2846) );
  XNOR U3245 ( .A(n2843), .B(n2844), .Z(n2855) );
  NAND U3246 ( .A(n1612), .B(n1203), .Z(n2844) );
  XNOR U3247 ( .A(n2842), .B(n2980), .Z(n2843) );
  ANDN U3248 ( .A(n1210), .B(n1614), .Z(n2980) );
  XNOR U3249 ( .A(n2854), .B(n2845), .Z(n2979) );
  XOR U3250 ( .A(n2987), .B(n2851), .Z(n2854) );
  XNOR U3251 ( .A(n2850), .B(n2988), .Z(n2851) );
  ANDN U3252 ( .A(n1394), .B(n1421), .Z(n2988) );
  AND U3253 ( .A(n1419), .B(n1387), .Z(n2852) );
  XNOR U3254 ( .A(n2863), .B(n2862), .Z(n2839) );
  XOR U3255 ( .A(n2995), .B(n2871), .Z(n2862) );
  XNOR U3256 ( .A(n2859), .B(n2860), .Z(n2871) );
  NANDN U3257 ( .B(n647), .A(n2491), .Z(n2860) );
  XNOR U3258 ( .A(n2858), .B(n2996), .Z(n2859) );
  ANDN U3259 ( .A(n688), .B(n2493), .Z(n2996) );
  XNOR U3260 ( .A(n2870), .B(n2861), .Z(n2995) );
  XOR U3261 ( .A(n3003), .B(n2867), .Z(n2870) );
  XNOR U3262 ( .A(n2866), .B(n3004), .Z(n2867) );
  ANDN U3263 ( .A(n795), .B(n2251), .Z(n3004) );
  AND U3264 ( .A(n2249), .B(n741), .Z(n2868) );
  XOR U3265 ( .A(n2879), .B(n2878), .Z(n2863) );
  XOR U3266 ( .A(n3011), .B(n2875), .Z(n2878) );
  XNOR U3267 ( .A(n2874), .B(n3012), .Z(n2875) );
  ANDN U3268 ( .A(n620), .B(n2750), .Z(n3012) );
  AND U3269 ( .A(n2748), .B(n579), .Z(n2876) );
  XOR U3270 ( .A(n2886), .B(n2885), .Z(n2879) );
  NAND U3271 ( .A(n3019), .B(n523), .Z(n2885) );
  XNOR U3272 ( .A(n2884), .B(n3020), .Z(n2886) );
  ANDN U3273 ( .A(n554), .B(n3021), .Z(n3020) );
  NAND U3274 ( .A(n3022), .B(n3023), .Z(n2884) );
  NAND U3275 ( .A(n3024), .B(n3025), .Z(n3022) );
  XNOR U3276 ( .A(n3026), .B(n2947), .Z(n2930) );
  XNOR U3277 ( .A(n2908), .B(n2907), .Z(n2947) );
  XOR U3278 ( .A(n3027), .B(n2916), .Z(n2907) );
  XNOR U3279 ( .A(n2904), .B(n2905), .Z(n2916) );
  NAND U3280 ( .A(n1934), .B(n1011), .Z(n2905) );
  XNOR U3281 ( .A(n2903), .B(n3028), .Z(n2904) );
  ANDN U3282 ( .A(n1939), .B(n1013), .Z(n3028) );
  XOR U3283 ( .A(n3029), .B(n3030), .Z(n2903) );
  AND U3284 ( .A(n3031), .B(n3032), .Z(n3030) );
  XOR U3285 ( .A(n3033), .B(n3029), .Z(n3032) );
  XNOR U3286 ( .A(n2915), .B(n2906), .Z(n3027) );
  XOR U3287 ( .A(n3037), .B(n2912), .Z(n2915) );
  XNOR U3288 ( .A(n2911), .B(n3038), .Z(n2912) );
  ANDN U3289 ( .A(n2169), .B(n878), .Z(n3038) );
  XOR U3290 ( .A(n3039), .B(n3040), .Z(n2911) );
  AND U3291 ( .A(n3041), .B(n3042), .Z(n3040) );
  XNOR U3292 ( .A(n3043), .B(n3039), .Z(n3042) );
  AND U3293 ( .A(n2162), .B(n876), .Z(n2913) );
  XNOR U3294 ( .A(n2924), .B(n2923), .Z(n2908) );
  XOR U3295 ( .A(n3047), .B(n2920), .Z(n2923) );
  XNOR U3296 ( .A(n2919), .B(n3048), .Z(n2920) );
  ANDN U3297 ( .A(n1740), .B(n1165), .Z(n3048) );
  AND U3298 ( .A(n1733), .B(n1163), .Z(n2921) );
  XNOR U3299 ( .A(n2927), .B(n2928), .Z(n2924) );
  NAND U3300 ( .A(n1538), .B(n1328), .Z(n2928) );
  XNOR U3301 ( .A(n2926), .B(n3055), .Z(n2927) );
  ANDN U3302 ( .A(n1543), .B(n1330), .Z(n3055) );
  XNOR U3303 ( .A(n2946), .B(n2929), .Z(n3026) );
  XNOR U3304 ( .A(n3059), .B(n3060), .Z(n2929) );
  XNOR U3305 ( .A(n3061), .B(n2958), .Z(n2946) );
  XNOR U3306 ( .A(n2940), .B(n2939), .Z(n2958) );
  XOR U3307 ( .A(n3062), .B(n2936), .Z(n2939) );
  XNOR U3308 ( .A(n2935), .B(n3063), .Z(n2936) );
  ANDN U3309 ( .A(n2678), .B(n669), .Z(n3063) );
  XOR U3310 ( .A(n3064), .B(n3065), .Z(n2935) );
  AND U3311 ( .A(n3066), .B(n3067), .Z(n3065) );
  XNOR U3312 ( .A(n3068), .B(n3064), .Z(n3067) );
  AND U3313 ( .A(n2671), .B(n667), .Z(n2937) );
  XNOR U3314 ( .A(n2943), .B(n2944), .Z(n2940) );
  NAND U3315 ( .A(n2424), .B(n753), .Z(n2944) );
  XNOR U3316 ( .A(n2942), .B(n3072), .Z(n2943) );
  ANDN U3317 ( .A(n2429), .B(n755), .Z(n3072) );
  XOR U3318 ( .A(n3073), .B(n3074), .Z(n2942) );
  AND U3319 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR U3320 ( .A(n3077), .B(n3073), .Z(n3076) );
  XNOR U3321 ( .A(n2957), .B(n2945), .Z(n3061) );
  XOR U3322 ( .A(n3078), .B(n3079), .Z(n2945) );
  AND U3323 ( .A(n3080), .B(n3081), .Z(n3079) );
  XOR U3324 ( .A(n3082), .B(n3083), .Z(n3081) );
  XNOR U3325 ( .A(n3084), .B(n3078), .Z(n3082) );
  XNOR U3326 ( .A(n3035), .B(n3085), .Z(n3080) );
  XNOR U3327 ( .A(n3078), .B(n3036), .Z(n3085) );
  XNOR U3328 ( .A(n3054), .B(n3053), .Z(n3036) );
  XOR U3329 ( .A(n3086), .B(n3050), .Z(n3053) );
  XNOR U3330 ( .A(n3049), .B(n3087), .Z(n3050) );
  ANDN U3331 ( .A(n1740), .B(n1246), .Z(n3087) );
  AND U3332 ( .A(n1733), .B(n1244), .Z(n3051) );
  XNOR U3333 ( .A(n3057), .B(n3058), .Z(n3054) );
  NAND U3334 ( .A(n1419), .B(n1538), .Z(n3058) );
  XNOR U3335 ( .A(n3056), .B(n3094), .Z(n3057) );
  ANDN U3336 ( .A(n1543), .B(n1421), .Z(n3094) );
  XOR U3337 ( .A(n3098), .B(n3046), .Z(n3035) );
  XNOR U3338 ( .A(n3031), .B(n3033), .Z(n3046) );
  NAND U3339 ( .A(n1934), .B(n1085), .Z(n3033) );
  XNOR U3340 ( .A(n3029), .B(n3099), .Z(n3031) );
  ANDN U3341 ( .A(n1939), .B(n1087), .Z(n3099) );
  XNOR U3342 ( .A(n3045), .B(n3034), .Z(n3098) );
  XOR U3343 ( .A(n3106), .B(n3041), .Z(n3045) );
  XNOR U3344 ( .A(n3039), .B(n3107), .Z(n3041) );
  ANDN U3345 ( .A(n2169), .B(n946), .Z(n3107) );
  XOR U3346 ( .A(n3108), .B(n3109), .Z(n3039) );
  AND U3347 ( .A(n3110), .B(n3111), .Z(n3109) );
  XNOR U3348 ( .A(n3112), .B(n3108), .Z(n3111) );
  AND U3349 ( .A(n2162), .B(n944), .Z(n3043) );
  XOR U3350 ( .A(n3116), .B(n3117), .Z(n3078) );
  AND U3351 ( .A(n3118), .B(n3119), .Z(n3117) );
  XOR U3352 ( .A(n3120), .B(n3121), .Z(n3119) );
  XOR U3353 ( .A(n3116), .B(n3122), .Z(n3121) );
  XNOR U3354 ( .A(n3104), .B(n3123), .Z(n3118) );
  XNOR U3355 ( .A(n3116), .B(n3105), .Z(n3123) );
  XNOR U3356 ( .A(n3093), .B(n3092), .Z(n3105) );
  XOR U3357 ( .A(n3124), .B(n3089), .Z(n3092) );
  XNOR U3358 ( .A(n3088), .B(n3125), .Z(n3089) );
  ANDN U3359 ( .A(n1740), .B(n1330), .Z(n3125) );
  XOR U3360 ( .A(n3126), .B(n3127), .Z(n3088) );
  AND U3361 ( .A(n3128), .B(n3129), .Z(n3127) );
  XNOR U3362 ( .A(n3130), .B(n3126), .Z(n3129) );
  AND U3363 ( .A(n1733), .B(n1328), .Z(n3090) );
  XNOR U3364 ( .A(n3096), .B(n3097), .Z(n3093) );
  NAND U3365 ( .A(n1516), .B(n1538), .Z(n3097) );
  XNOR U3366 ( .A(n3095), .B(n3134), .Z(n3096) );
  ANDN U3367 ( .A(n1543), .B(n1518), .Z(n3134) );
  XOR U3368 ( .A(n3135), .B(n3136), .Z(n3095) );
  AND U3369 ( .A(n3137), .B(n3138), .Z(n3136) );
  XOR U3370 ( .A(n3139), .B(n3135), .Z(n3138) );
  XOR U3371 ( .A(n3140), .B(n3115), .Z(n3104) );
  XNOR U3372 ( .A(n3101), .B(n3102), .Z(n3115) );
  NAND U3373 ( .A(n1934), .B(n1163), .Z(n3102) );
  XNOR U3374 ( .A(n3100), .B(n3141), .Z(n3101) );
  ANDN U3375 ( .A(n1939), .B(n1165), .Z(n3141) );
  XOR U3376 ( .A(n3142), .B(n3143), .Z(n3100) );
  AND U3377 ( .A(n3144), .B(n3145), .Z(n3143) );
  XOR U3378 ( .A(n3146), .B(n3142), .Z(n3145) );
  XNOR U3379 ( .A(n3114), .B(n3103), .Z(n3140) );
  XOR U3380 ( .A(n3150), .B(n3110), .Z(n3114) );
  XNOR U3381 ( .A(n3108), .B(n3151), .Z(n3110) );
  ANDN U3382 ( .A(n2169), .B(n1013), .Z(n3151) );
  XOR U3383 ( .A(n3152), .B(n3153), .Z(n3108) );
  AND U3384 ( .A(n3154), .B(n3155), .Z(n3153) );
  XNOR U3385 ( .A(n3156), .B(n3152), .Z(n3155) );
  XOR U3386 ( .A(n3157), .B(n3112), .Z(n3150) );
  AND U3387 ( .A(n2162), .B(n1011), .Z(n3112) );
  IV U3388 ( .A(n3113), .Z(n3157) );
  XOR U3389 ( .A(n3161), .B(n3162), .Z(n3116) );
  AND U3390 ( .A(n3163), .B(n3164), .Z(n3162) );
  XOR U3391 ( .A(n3165), .B(n3166), .Z(n3164) );
  XOR U3392 ( .A(n3161), .B(n3167), .Z(n3166) );
  XNOR U3393 ( .A(n3148), .B(n3168), .Z(n3163) );
  XNOR U3394 ( .A(n3161), .B(n3149), .Z(n3168) );
  XNOR U3395 ( .A(n3133), .B(n3132), .Z(n3149) );
  XOR U3396 ( .A(n3169), .B(n3128), .Z(n3132) );
  XNOR U3397 ( .A(n3126), .B(n3170), .Z(n3128) );
  ANDN U3398 ( .A(n1740), .B(n1421), .Z(n3170) );
  XOR U3399 ( .A(n3171), .B(n3172), .Z(n3126) );
  AND U3400 ( .A(n3173), .B(n3174), .Z(n3172) );
  XNOR U3401 ( .A(n3175), .B(n3171), .Z(n3174) );
  AND U3402 ( .A(n1419), .B(n1733), .Z(n3130) );
  XNOR U3403 ( .A(n3137), .B(n3139), .Z(n3133) );
  NAND U3404 ( .A(n1612), .B(n1538), .Z(n3139) );
  XNOR U3405 ( .A(n3135), .B(n3179), .Z(n3137) );
  ANDN U3406 ( .A(n1543), .B(n1614), .Z(n3179) );
  XOR U3407 ( .A(n3183), .B(n3160), .Z(n3148) );
  XNOR U3408 ( .A(n3144), .B(n3146), .Z(n3160) );
  NAND U3409 ( .A(n1934), .B(n1244), .Z(n3146) );
  XNOR U3410 ( .A(n3142), .B(n3184), .Z(n3144) );
  ANDN U3411 ( .A(n1939), .B(n1246), .Z(n3184) );
  XOR U3412 ( .A(n3185), .B(n3186), .Z(n3142) );
  AND U3413 ( .A(n3187), .B(n3188), .Z(n3186) );
  XOR U3414 ( .A(n3189), .B(n3185), .Z(n3188) );
  XNOR U3415 ( .A(n3159), .B(n3147), .Z(n3183) );
  XOR U3416 ( .A(n3193), .B(n3154), .Z(n3159) );
  XNOR U3417 ( .A(n3152), .B(n3194), .Z(n3154) );
  ANDN U3418 ( .A(n2169), .B(n1087), .Z(n3194) );
  XOR U3419 ( .A(n3195), .B(n3196), .Z(n3152) );
  AND U3420 ( .A(n3197), .B(n3198), .Z(n3196) );
  XNOR U3421 ( .A(n3199), .B(n3195), .Z(n3198) );
  AND U3422 ( .A(n2162), .B(n1085), .Z(n3156) );
  XOR U3423 ( .A(n3203), .B(n3204), .Z(n3161) );
  AND U3424 ( .A(n3205), .B(n3206), .Z(n3204) );
  XOR U3425 ( .A(n3207), .B(n3208), .Z(n3206) );
  XOR U3426 ( .A(n3203), .B(n3209), .Z(n3208) );
  XNOR U3427 ( .A(n3191), .B(n3210), .Z(n3205) );
  XNOR U3428 ( .A(n3203), .B(n3192), .Z(n3210) );
  XNOR U3429 ( .A(n3178), .B(n3177), .Z(n3192) );
  XOR U3430 ( .A(n3211), .B(n3173), .Z(n3177) );
  XNOR U3431 ( .A(n3171), .B(n3212), .Z(n3173) );
  ANDN U3432 ( .A(n1740), .B(n1518), .Z(n3212) );
  XOR U3433 ( .A(n3213), .B(n3214), .Z(n3171) );
  AND U3434 ( .A(n3215), .B(n3216), .Z(n3214) );
  XNOR U3435 ( .A(n3217), .B(n3213), .Z(n3216) );
  AND U3436 ( .A(n1516), .B(n1733), .Z(n3175) );
  XNOR U3437 ( .A(n3181), .B(n3182), .Z(n3178) );
  NAND U3438 ( .A(n1708), .B(n1538), .Z(n3182) );
  XNOR U3439 ( .A(n3180), .B(n3221), .Z(n3181) );
  ANDN U3440 ( .A(n1543), .B(n1710), .Z(n3221) );
  XOR U3441 ( .A(n3222), .B(n3223), .Z(n3180) );
  AND U3442 ( .A(n3224), .B(n3225), .Z(n3223) );
  XOR U3443 ( .A(n3226), .B(n3222), .Z(n3225) );
  XOR U3444 ( .A(n3227), .B(n3202), .Z(n3191) );
  XNOR U3445 ( .A(n3187), .B(n3189), .Z(n3202) );
  NAND U3446 ( .A(n1934), .B(n1328), .Z(n3189) );
  XNOR U3447 ( .A(n3185), .B(n3228), .Z(n3187) );
  ANDN U3448 ( .A(n1939), .B(n1330), .Z(n3228) );
  XNOR U3449 ( .A(n3201), .B(n3190), .Z(n3227) );
  XOR U3450 ( .A(n3235), .B(n3197), .Z(n3201) );
  XNOR U3451 ( .A(n3195), .B(n3236), .Z(n3197) );
  ANDN U3452 ( .A(n2169), .B(n1165), .Z(n3236) );
  XOR U3453 ( .A(n3237), .B(n3238), .Z(n3195) );
  AND U3454 ( .A(n3239), .B(n3240), .Z(n3238) );
  XNOR U3455 ( .A(n3241), .B(n3237), .Z(n3240) );
  XOR U3456 ( .A(n3242), .B(n3199), .Z(n3235) );
  AND U3457 ( .A(n2162), .B(n1163), .Z(n3199) );
  IV U3458 ( .A(n3200), .Z(n3242) );
  XOR U3459 ( .A(n3246), .B(n3247), .Z(n3203) );
  AND U3460 ( .A(n3248), .B(n3249), .Z(n3247) );
  XOR U3461 ( .A(n3250), .B(n3251), .Z(n3249) );
  XOR U3462 ( .A(n3246), .B(n3252), .Z(n3251) );
  XNOR U3463 ( .A(n3233), .B(n3253), .Z(n3248) );
  XNOR U3464 ( .A(n3246), .B(n3234), .Z(n3253) );
  XNOR U3465 ( .A(n3220), .B(n3219), .Z(n3234) );
  XOR U3466 ( .A(n3254), .B(n3215), .Z(n3219) );
  XNOR U3467 ( .A(n3213), .B(n3255), .Z(n3215) );
  ANDN U3468 ( .A(n1740), .B(n1614), .Z(n3255) );
  XOR U3469 ( .A(n3256), .B(n3257), .Z(n3213) );
  AND U3470 ( .A(n3258), .B(n3259), .Z(n3257) );
  XNOR U3471 ( .A(n3260), .B(n3256), .Z(n3259) );
  AND U3472 ( .A(n1612), .B(n1733), .Z(n3217) );
  XNOR U3473 ( .A(n3224), .B(n3226), .Z(n3220) );
  NAND U3474 ( .A(n1809), .B(n1538), .Z(n3226) );
  XNOR U3475 ( .A(n3222), .B(n3264), .Z(n3224) );
  ANDN U3476 ( .A(n1543), .B(n1811), .Z(n3264) );
  XOR U3477 ( .A(n3268), .B(n3245), .Z(n3233) );
  XNOR U3478 ( .A(n3230), .B(n3231), .Z(n3245) );
  NAND U3479 ( .A(n1419), .B(n1934), .Z(n3231) );
  XNOR U3480 ( .A(n3229), .B(n3269), .Z(n3230) );
  ANDN U3481 ( .A(n1939), .B(n1421), .Z(n3269) );
  XOR U3482 ( .A(n3270), .B(n3271), .Z(n3229) );
  AND U3483 ( .A(n3272), .B(n3273), .Z(n3271) );
  XOR U3484 ( .A(n3274), .B(n3270), .Z(n3273) );
  XNOR U3485 ( .A(n3244), .B(n3232), .Z(n3268) );
  XOR U3486 ( .A(n3278), .B(n3239), .Z(n3244) );
  XNOR U3487 ( .A(n3237), .B(n3279), .Z(n3239) );
  ANDN U3488 ( .A(n2169), .B(n1246), .Z(n3279) );
  XOR U3489 ( .A(n3280), .B(n3281), .Z(n3237) );
  AND U3490 ( .A(n3282), .B(n3283), .Z(n3281) );
  XNOR U3491 ( .A(n3284), .B(n3280), .Z(n3283) );
  AND U3492 ( .A(n2162), .B(n1244), .Z(n3241) );
  XOR U3493 ( .A(n3288), .B(n3289), .Z(n3246) );
  AND U3494 ( .A(n3290), .B(n3291), .Z(n3289) );
  XOR U3495 ( .A(n3292), .B(n3293), .Z(n3291) );
  XOR U3496 ( .A(n3288), .B(n3294), .Z(n3293) );
  XNOR U3497 ( .A(n3276), .B(n3295), .Z(n3290) );
  XNOR U3498 ( .A(n3288), .B(n3277), .Z(n3295) );
  XNOR U3499 ( .A(n3263), .B(n3262), .Z(n3277) );
  XOR U3500 ( .A(n3296), .B(n3258), .Z(n3262) );
  XNOR U3501 ( .A(n3256), .B(n3297), .Z(n3258) );
  ANDN U3502 ( .A(n1740), .B(n1710), .Z(n3297) );
  XOR U3503 ( .A(n3298), .B(n3299), .Z(n3256) );
  AND U3504 ( .A(n3300), .B(n3301), .Z(n3299) );
  XNOR U3505 ( .A(n3302), .B(n3298), .Z(n3301) );
  XOR U3506 ( .A(n3303), .B(n3260), .Z(n3296) );
  AND U3507 ( .A(n1708), .B(n1733), .Z(n3260) );
  IV U3508 ( .A(n3261), .Z(n3303) );
  XNOR U3509 ( .A(n3266), .B(n3267), .Z(n3263) );
  NAND U3510 ( .A(n1915), .B(n1538), .Z(n3267) );
  XNOR U3511 ( .A(n3265), .B(n3307), .Z(n3266) );
  ANDN U3512 ( .A(n1543), .B(n1917), .Z(n3307) );
  XOR U3513 ( .A(n3308), .B(n3309), .Z(n3265) );
  AND U3514 ( .A(n3310), .B(n3311), .Z(n3309) );
  XOR U3515 ( .A(n3312), .B(n3308), .Z(n3311) );
  XOR U3516 ( .A(n3313), .B(n3287), .Z(n3276) );
  XNOR U3517 ( .A(n3272), .B(n3274), .Z(n3287) );
  NAND U3518 ( .A(n1516), .B(n1934), .Z(n3274) );
  XNOR U3519 ( .A(n3270), .B(n3314), .Z(n3272) );
  ANDN U3520 ( .A(n1939), .B(n1518), .Z(n3314) );
  XOR U3521 ( .A(n3315), .B(n3316), .Z(n3270) );
  AND U3522 ( .A(n3317), .B(n3318), .Z(n3316) );
  XOR U3523 ( .A(n3319), .B(n3315), .Z(n3318) );
  XNOR U3524 ( .A(n3286), .B(n3275), .Z(n3313) );
  XOR U3525 ( .A(n3323), .B(n3282), .Z(n3286) );
  XNOR U3526 ( .A(n3280), .B(n3324), .Z(n3282) );
  ANDN U3527 ( .A(n2169), .B(n1330), .Z(n3324) );
  XOR U3528 ( .A(n3325), .B(n3326), .Z(n3280) );
  AND U3529 ( .A(n3327), .B(n3328), .Z(n3326) );
  XNOR U3530 ( .A(n3329), .B(n3325), .Z(n3328) );
  XOR U3531 ( .A(n3330), .B(n3284), .Z(n3323) );
  AND U3532 ( .A(n2162), .B(n1328), .Z(n3284) );
  IV U3533 ( .A(n3285), .Z(n3330) );
  XOR U3534 ( .A(n3334), .B(n3335), .Z(n3288) );
  AND U3535 ( .A(n3336), .B(n3337), .Z(n3335) );
  XOR U3536 ( .A(n3338), .B(n3339), .Z(n3337) );
  XOR U3537 ( .A(n3334), .B(n3340), .Z(n3339) );
  XNOR U3538 ( .A(n3321), .B(n3341), .Z(n3336) );
  XNOR U3539 ( .A(n3334), .B(n3322), .Z(n3341) );
  XNOR U3540 ( .A(n3306), .B(n3305), .Z(n3322) );
  XOR U3541 ( .A(n3342), .B(n3300), .Z(n3305) );
  XNOR U3542 ( .A(n3298), .B(n3343), .Z(n3300) );
  ANDN U3543 ( .A(n1740), .B(n1811), .Z(n3343) );
  XOR U3544 ( .A(n3344), .B(n3345), .Z(n3298) );
  AND U3545 ( .A(n3346), .B(n3347), .Z(n3345) );
  XNOR U3546 ( .A(n3348), .B(n3344), .Z(n3347) );
  XOR U3547 ( .A(n3349), .B(n3302), .Z(n3342) );
  AND U3548 ( .A(n1809), .B(n1733), .Z(n3302) );
  IV U3549 ( .A(n3304), .Z(n3349) );
  XNOR U3550 ( .A(n3310), .B(n3312), .Z(n3306) );
  NAND U3551 ( .A(n2022), .B(n1538), .Z(n3312) );
  XNOR U3552 ( .A(n3308), .B(n3353), .Z(n3310) );
  ANDN U3553 ( .A(n1543), .B(n2024), .Z(n3353) );
  XOR U3554 ( .A(n3354), .B(n3355), .Z(n3308) );
  AND U3555 ( .A(n3356), .B(n3357), .Z(n3355) );
  XOR U3556 ( .A(n3358), .B(n3354), .Z(n3357) );
  XOR U3557 ( .A(n3359), .B(n3333), .Z(n3321) );
  XNOR U3558 ( .A(n3317), .B(n3319), .Z(n3333) );
  NAND U3559 ( .A(n1612), .B(n1934), .Z(n3319) );
  XNOR U3560 ( .A(n3315), .B(n3360), .Z(n3317) );
  ANDN U3561 ( .A(n1939), .B(n1614), .Z(n3360) );
  XNOR U3562 ( .A(n3332), .B(n3320), .Z(n3359) );
  XOR U3563 ( .A(n3367), .B(n3327), .Z(n3332) );
  XNOR U3564 ( .A(n3325), .B(n3368), .Z(n3327) );
  ANDN U3565 ( .A(n2169), .B(n1421), .Z(n3368) );
  XOR U3566 ( .A(n3369), .B(n3370), .Z(n3325) );
  AND U3567 ( .A(n3371), .B(n3372), .Z(n3370) );
  XNOR U3568 ( .A(n3373), .B(n3369), .Z(n3372) );
  XOR U3569 ( .A(n3374), .B(n3329), .Z(n3367) );
  AND U3570 ( .A(n1419), .B(n2162), .Z(n3329) );
  IV U3571 ( .A(n3331), .Z(n3374) );
  XOR U3572 ( .A(n3378), .B(n3379), .Z(n3334) );
  AND U3573 ( .A(n3380), .B(n3381), .Z(n3379) );
  XOR U3574 ( .A(n3382), .B(n3383), .Z(n3381) );
  XOR U3575 ( .A(n3378), .B(n3384), .Z(n3383) );
  XNOR U3576 ( .A(n3365), .B(n3385), .Z(n3380) );
  XNOR U3577 ( .A(n3378), .B(n3366), .Z(n3385) );
  XNOR U3578 ( .A(n3352), .B(n3351), .Z(n3366) );
  XOR U3579 ( .A(n3386), .B(n3346), .Z(n3351) );
  XNOR U3580 ( .A(n3344), .B(n3387), .Z(n3346) );
  ANDN U3581 ( .A(n1740), .B(n1917), .Z(n3387) );
  XOR U3582 ( .A(n3388), .B(n3389), .Z(n3344) );
  AND U3583 ( .A(n3390), .B(n3391), .Z(n3389) );
  XNOR U3584 ( .A(n3392), .B(n3388), .Z(n3391) );
  XOR U3585 ( .A(n3393), .B(n3348), .Z(n3386) );
  AND U3586 ( .A(n1915), .B(n1733), .Z(n3348) );
  IV U3587 ( .A(n3350), .Z(n3393) );
  XNOR U3588 ( .A(n3356), .B(n3358), .Z(n3352) );
  NAND U3589 ( .A(n2130), .B(n1538), .Z(n3358) );
  XNOR U3590 ( .A(n3354), .B(n3397), .Z(n3356) );
  ANDN U3591 ( .A(n1543), .B(n2132), .Z(n3397) );
  XOR U3592 ( .A(n3398), .B(n3399), .Z(n3354) );
  AND U3593 ( .A(n3400), .B(n3401), .Z(n3399) );
  XOR U3594 ( .A(n3402), .B(n3398), .Z(n3401) );
  XOR U3595 ( .A(n3403), .B(n3377), .Z(n3365) );
  XNOR U3596 ( .A(n3362), .B(n3363), .Z(n3377) );
  NAND U3597 ( .A(n1708), .B(n1934), .Z(n3363) );
  XNOR U3598 ( .A(n3361), .B(n3404), .Z(n3362) );
  ANDN U3599 ( .A(n1939), .B(n1710), .Z(n3404) );
  XOR U3600 ( .A(n3405), .B(n3406), .Z(n3361) );
  AND U3601 ( .A(n3407), .B(n3408), .Z(n3406) );
  XOR U3602 ( .A(n3409), .B(n3405), .Z(n3408) );
  XNOR U3603 ( .A(n3376), .B(n3364), .Z(n3403) );
  XOR U3604 ( .A(n3413), .B(n3371), .Z(n3376) );
  XNOR U3605 ( .A(n3369), .B(n3414), .Z(n3371) );
  ANDN U3606 ( .A(n2169), .B(n1518), .Z(n3414) );
  XOR U3607 ( .A(n3415), .B(n3416), .Z(n3369) );
  AND U3608 ( .A(n3417), .B(n3418), .Z(n3416) );
  XNOR U3609 ( .A(n3419), .B(n3415), .Z(n3418) );
  XOR U3610 ( .A(n3420), .B(n3373), .Z(n3413) );
  AND U3611 ( .A(n1516), .B(n2162), .Z(n3373) );
  IV U3612 ( .A(n3375), .Z(n3420) );
  XOR U3613 ( .A(n3424), .B(n3425), .Z(n3378) );
  AND U3614 ( .A(n3426), .B(n3427), .Z(n3425) );
  XOR U3615 ( .A(n3428), .B(n3429), .Z(n3427) );
  XOR U3616 ( .A(n3424), .B(n3430), .Z(n3429) );
  XNOR U3617 ( .A(n3411), .B(n3431), .Z(n3426) );
  XNOR U3618 ( .A(n3424), .B(n3412), .Z(n3431) );
  XNOR U3619 ( .A(n3396), .B(n3395), .Z(n3412) );
  XOR U3620 ( .A(n3432), .B(n3390), .Z(n3395) );
  XNOR U3621 ( .A(n3388), .B(n3433), .Z(n3390) );
  ANDN U3622 ( .A(n1740), .B(n2024), .Z(n3433) );
  XOR U3623 ( .A(n3434), .B(n3435), .Z(n3388) );
  AND U3624 ( .A(n3436), .B(n3437), .Z(n3435) );
  XNOR U3625 ( .A(n3438), .B(n3434), .Z(n3437) );
  XOR U3626 ( .A(n3439), .B(n3392), .Z(n3432) );
  AND U3627 ( .A(n2022), .B(n1733), .Z(n3392) );
  IV U3628 ( .A(n3394), .Z(n3439) );
  XNOR U3629 ( .A(n3400), .B(n3402), .Z(n3396) );
  NAND U3630 ( .A(n2249), .B(n1538), .Z(n3402) );
  XNOR U3631 ( .A(n3398), .B(n3443), .Z(n3400) );
  ANDN U3632 ( .A(n1543), .B(n2251), .Z(n3443) );
  XOR U3633 ( .A(n3444), .B(n3445), .Z(n3398) );
  AND U3634 ( .A(n3446), .B(n3447), .Z(n3445) );
  XOR U3635 ( .A(n3448), .B(n3444), .Z(n3447) );
  XOR U3636 ( .A(n3449), .B(n3423), .Z(n3411) );
  XNOR U3637 ( .A(n3407), .B(n3409), .Z(n3423) );
  NAND U3638 ( .A(n1809), .B(n1934), .Z(n3409) );
  XNOR U3639 ( .A(n3405), .B(n3450), .Z(n3407) );
  ANDN U3640 ( .A(n1939), .B(n1811), .Z(n3450) );
  XOR U3641 ( .A(n3451), .B(n3452), .Z(n3405) );
  AND U3642 ( .A(n3453), .B(n3454), .Z(n3452) );
  XOR U3643 ( .A(n3455), .B(n3451), .Z(n3454) );
  XNOR U3644 ( .A(n3422), .B(n3410), .Z(n3449) );
  XOR U3645 ( .A(n3459), .B(n3417), .Z(n3422) );
  XNOR U3646 ( .A(n3415), .B(n3460), .Z(n3417) );
  ANDN U3647 ( .A(n2169), .B(n1614), .Z(n3460) );
  XOR U3648 ( .A(n3461), .B(n3462), .Z(n3415) );
  AND U3649 ( .A(n3463), .B(n3464), .Z(n3462) );
  XNOR U3650 ( .A(n3465), .B(n3461), .Z(n3464) );
  XOR U3651 ( .A(n3466), .B(n3419), .Z(n3459) );
  AND U3652 ( .A(n1612), .B(n2162), .Z(n3419) );
  IV U3653 ( .A(n3421), .Z(n3466) );
  XOR U3654 ( .A(n3470), .B(n3471), .Z(n3424) );
  AND U3655 ( .A(n3472), .B(n3473), .Z(n3471) );
  XOR U3656 ( .A(n3474), .B(n3475), .Z(n3473) );
  XOR U3657 ( .A(n3470), .B(n3476), .Z(n3475) );
  XNOR U3658 ( .A(n3457), .B(n3477), .Z(n3472) );
  XNOR U3659 ( .A(n3470), .B(n3458), .Z(n3477) );
  XNOR U3660 ( .A(n3442), .B(n3441), .Z(n3458) );
  XOR U3661 ( .A(n3478), .B(n3436), .Z(n3441) );
  XNOR U3662 ( .A(n3434), .B(n3479), .Z(n3436) );
  ANDN U3663 ( .A(n1740), .B(n2132), .Z(n3479) );
  XOR U3664 ( .A(n3480), .B(n3481), .Z(n3434) );
  AND U3665 ( .A(n3482), .B(n3483), .Z(n3481) );
  XNOR U3666 ( .A(n3484), .B(n3480), .Z(n3483) );
  XOR U3667 ( .A(n3485), .B(n3438), .Z(n3478) );
  AND U3668 ( .A(n2130), .B(n1733), .Z(n3438) );
  IV U3669 ( .A(n3440), .Z(n3485) );
  XNOR U3670 ( .A(n3446), .B(n3448), .Z(n3442) );
  NAND U3671 ( .A(n2369), .B(n1538), .Z(n3448) );
  XNOR U3672 ( .A(n3444), .B(n3489), .Z(n3446) );
  ANDN U3673 ( .A(n1543), .B(n2371), .Z(n3489) );
  XOR U3674 ( .A(n3490), .B(n3491), .Z(n3444) );
  AND U3675 ( .A(n3492), .B(n3493), .Z(n3491) );
  XOR U3676 ( .A(n3494), .B(n3490), .Z(n3493) );
  XOR U3677 ( .A(n3495), .B(n3469), .Z(n3457) );
  XNOR U3678 ( .A(n3453), .B(n3455), .Z(n3469) );
  NAND U3679 ( .A(n1915), .B(n1934), .Z(n3455) );
  XNOR U3680 ( .A(n3451), .B(n3496), .Z(n3453) );
  ANDN U3681 ( .A(n1939), .B(n1917), .Z(n3496) );
  XOR U3682 ( .A(n3497), .B(n3498), .Z(n3451) );
  AND U3683 ( .A(n3499), .B(n3500), .Z(n3498) );
  XOR U3684 ( .A(n3501), .B(n3497), .Z(n3500) );
  XNOR U3685 ( .A(n3468), .B(n3456), .Z(n3495) );
  XOR U3686 ( .A(n3505), .B(n3463), .Z(n3468) );
  XNOR U3687 ( .A(n3461), .B(n3506), .Z(n3463) );
  ANDN U3688 ( .A(n2169), .B(n1710), .Z(n3506) );
  XOR U3689 ( .A(n3507), .B(n3508), .Z(n3461) );
  AND U3690 ( .A(n3509), .B(n3510), .Z(n3508) );
  XNOR U3691 ( .A(n3511), .B(n3507), .Z(n3510) );
  XOR U3692 ( .A(n3512), .B(n3465), .Z(n3505) );
  AND U3693 ( .A(n1708), .B(n2162), .Z(n3465) );
  IV U3694 ( .A(n3467), .Z(n3512) );
  XOR U3695 ( .A(n3516), .B(n3517), .Z(n3470) );
  AND U3696 ( .A(n3518), .B(n3519), .Z(n3517) );
  XOR U3697 ( .A(n3520), .B(n3521), .Z(n3519) );
  XOR U3698 ( .A(n3516), .B(n3522), .Z(n3521) );
  XNOR U3699 ( .A(n3503), .B(n3523), .Z(n3518) );
  XNOR U3700 ( .A(n3516), .B(n3504), .Z(n3523) );
  XNOR U3701 ( .A(n3488), .B(n3487), .Z(n3504) );
  XOR U3702 ( .A(n3524), .B(n3482), .Z(n3487) );
  XNOR U3703 ( .A(n3480), .B(n3525), .Z(n3482) );
  ANDN U3704 ( .A(n1740), .B(n2251), .Z(n3525) );
  XOR U3705 ( .A(n3526), .B(n3527), .Z(n3480) );
  AND U3706 ( .A(n3528), .B(n3529), .Z(n3527) );
  XNOR U3707 ( .A(n3530), .B(n3526), .Z(n3529) );
  XOR U3708 ( .A(n3531), .B(n3484), .Z(n3524) );
  AND U3709 ( .A(n2249), .B(n1733), .Z(n3484) );
  IV U3710 ( .A(n3486), .Z(n3531) );
  XNOR U3711 ( .A(n3492), .B(n3494), .Z(n3488) );
  NAND U3712 ( .A(n2491), .B(n1538), .Z(n3494) );
  XNOR U3713 ( .A(n3490), .B(n3535), .Z(n3492) );
  ANDN U3714 ( .A(n1543), .B(n2493), .Z(n3535) );
  XOR U3715 ( .A(n3539), .B(n3515), .Z(n3503) );
  XNOR U3716 ( .A(n3499), .B(n3501), .Z(n3515) );
  NAND U3717 ( .A(n2022), .B(n1934), .Z(n3501) );
  XNOR U3718 ( .A(n3497), .B(n3540), .Z(n3499) );
  ANDN U3719 ( .A(n1939), .B(n2024), .Z(n3540) );
  XOR U3720 ( .A(n3541), .B(n3542), .Z(n3497) );
  AND U3721 ( .A(n3543), .B(n3544), .Z(n3542) );
  XOR U3722 ( .A(n3545), .B(n3541), .Z(n3544) );
  XNOR U3723 ( .A(n3514), .B(n3502), .Z(n3539) );
  XOR U3724 ( .A(n3549), .B(n3509), .Z(n3514) );
  XNOR U3725 ( .A(n3507), .B(n3550), .Z(n3509) );
  ANDN U3726 ( .A(n2169), .B(n1811), .Z(n3550) );
  XOR U3727 ( .A(n3551), .B(n3552), .Z(n3507) );
  AND U3728 ( .A(n3553), .B(n3554), .Z(n3552) );
  XNOR U3729 ( .A(n3555), .B(n3551), .Z(n3554) );
  XOR U3730 ( .A(n3556), .B(n3511), .Z(n3549) );
  AND U3731 ( .A(n1809), .B(n2162), .Z(n3511) );
  IV U3732 ( .A(n3513), .Z(n3556) );
  XOR U3733 ( .A(n3560), .B(n3561), .Z(n3516) );
  AND U3734 ( .A(n3562), .B(n3563), .Z(n3561) );
  XOR U3735 ( .A(n3564), .B(n3565), .Z(n3563) );
  XOR U3736 ( .A(n3560), .B(n3566), .Z(n3565) );
  XNOR U3737 ( .A(n3547), .B(n3567), .Z(n3562) );
  XNOR U3738 ( .A(n3560), .B(n3548), .Z(n3567) );
  XNOR U3739 ( .A(n3534), .B(n3533), .Z(n3548) );
  XOR U3740 ( .A(n3568), .B(n3528), .Z(n3533) );
  XNOR U3741 ( .A(n3526), .B(n3569), .Z(n3528) );
  ANDN U3742 ( .A(n1740), .B(n2371), .Z(n3569) );
  XOR U3743 ( .A(n3570), .B(n3571), .Z(n3526) );
  AND U3744 ( .A(n3572), .B(n3573), .Z(n3571) );
  XNOR U3745 ( .A(n3574), .B(n3570), .Z(n3573) );
  XOR U3746 ( .A(n3575), .B(n3530), .Z(n3568) );
  AND U3747 ( .A(n2369), .B(n1733), .Z(n3530) );
  IV U3748 ( .A(n3532), .Z(n3575) );
  XNOR U3749 ( .A(n3537), .B(n3538), .Z(n3534) );
  NAND U3750 ( .A(n2616), .B(n1538), .Z(n3538) );
  XNOR U3751 ( .A(n3536), .B(n3579), .Z(n3537) );
  ANDN U3752 ( .A(n1543), .B(n2618), .Z(n3579) );
  XOR U3753 ( .A(n3580), .B(n3581), .Z(n3536) );
  AND U3754 ( .A(n3582), .B(n3583), .Z(n3581) );
  XOR U3755 ( .A(n3584), .B(n3580), .Z(n3583) );
  XOR U3756 ( .A(n3585), .B(n3559), .Z(n3547) );
  XNOR U3757 ( .A(n3543), .B(n3545), .Z(n3559) );
  NAND U3758 ( .A(n2130), .B(n1934), .Z(n3545) );
  XNOR U3759 ( .A(n3541), .B(n3586), .Z(n3543) );
  ANDN U3760 ( .A(n1939), .B(n2132), .Z(n3586) );
  XOR U3761 ( .A(n3587), .B(n3588), .Z(n3541) );
  AND U3762 ( .A(n3589), .B(n3590), .Z(n3588) );
  XOR U3763 ( .A(n3591), .B(n3587), .Z(n3590) );
  XNOR U3764 ( .A(n3558), .B(n3546), .Z(n3585) );
  XOR U3765 ( .A(n3595), .B(n3553), .Z(n3558) );
  XNOR U3766 ( .A(n3551), .B(n3596), .Z(n3553) );
  ANDN U3767 ( .A(n2169), .B(n1917), .Z(n3596) );
  XOR U3768 ( .A(n3597), .B(n3598), .Z(n3551) );
  AND U3769 ( .A(n3599), .B(n3600), .Z(n3598) );
  XNOR U3770 ( .A(n3601), .B(n3597), .Z(n3600) );
  XOR U3771 ( .A(n3602), .B(n3555), .Z(n3595) );
  AND U3772 ( .A(n1915), .B(n2162), .Z(n3555) );
  IV U3773 ( .A(n3557), .Z(n3602) );
  XOR U3774 ( .A(n3606), .B(n3607), .Z(n3560) );
  AND U3775 ( .A(n3608), .B(n3609), .Z(n3607) );
  XOR U3776 ( .A(n3610), .B(n3611), .Z(n3609) );
  XOR U3777 ( .A(n3606), .B(n3612), .Z(n3611) );
  XNOR U3778 ( .A(n3593), .B(n3613), .Z(n3608) );
  XNOR U3779 ( .A(n3606), .B(n3594), .Z(n3613) );
  XNOR U3780 ( .A(n3578), .B(n3577), .Z(n3594) );
  XOR U3781 ( .A(n3614), .B(n3572), .Z(n3577) );
  XNOR U3782 ( .A(n3570), .B(n3615), .Z(n3572) );
  ANDN U3783 ( .A(n1740), .B(n2493), .Z(n3615) );
  XOR U3784 ( .A(n3616), .B(n3617), .Z(n3570) );
  AND U3785 ( .A(n3618), .B(n3619), .Z(n3617) );
  XNOR U3786 ( .A(n3620), .B(n3616), .Z(n3619) );
  XOR U3787 ( .A(n3621), .B(n3574), .Z(n3614) );
  AND U3788 ( .A(n2491), .B(n1733), .Z(n3574) );
  IV U3789 ( .A(n3576), .Z(n3621) );
  XNOR U3790 ( .A(n3582), .B(n3584), .Z(n3578) );
  NAND U3791 ( .A(n2748), .B(n1538), .Z(n3584) );
  XNOR U3792 ( .A(n3580), .B(n3625), .Z(n3582) );
  ANDN U3793 ( .A(n1543), .B(n2750), .Z(n3625) );
  XOR U3794 ( .A(n3626), .B(n3627), .Z(n3580) );
  AND U3795 ( .A(n3628), .B(n3629), .Z(n3627) );
  XOR U3796 ( .A(n3630), .B(n3626), .Z(n3629) );
  XOR U3797 ( .A(n3631), .B(n3605), .Z(n3593) );
  XNOR U3798 ( .A(n3589), .B(n3591), .Z(n3605) );
  NAND U3799 ( .A(n2249), .B(n1934), .Z(n3591) );
  XNOR U3800 ( .A(n3587), .B(n3632), .Z(n3589) );
  ANDN U3801 ( .A(n1939), .B(n2251), .Z(n3632) );
  XOR U3802 ( .A(n3633), .B(n3634), .Z(n3587) );
  AND U3803 ( .A(n3635), .B(n3636), .Z(n3634) );
  XOR U3804 ( .A(n3637), .B(n3633), .Z(n3636) );
  XNOR U3805 ( .A(n3604), .B(n3592), .Z(n3631) );
  XOR U3806 ( .A(n3641), .B(n3599), .Z(n3604) );
  XNOR U3807 ( .A(n3597), .B(n3642), .Z(n3599) );
  ANDN U3808 ( .A(n2169), .B(n2024), .Z(n3642) );
  XOR U3809 ( .A(n3643), .B(n3644), .Z(n3597) );
  AND U3810 ( .A(n3645), .B(n3646), .Z(n3644) );
  XNOR U3811 ( .A(n3647), .B(n3643), .Z(n3646) );
  XOR U3812 ( .A(n3648), .B(n3601), .Z(n3641) );
  AND U3813 ( .A(n2022), .B(n2162), .Z(n3601) );
  IV U3814 ( .A(n3603), .Z(n3648) );
  XOR U3815 ( .A(n3652), .B(n3653), .Z(n3606) );
  AND U3816 ( .A(n3654), .B(n3655), .Z(n3653) );
  XOR U3817 ( .A(n3656), .B(n3657), .Z(n3655) );
  XOR U3818 ( .A(n3652), .B(n3658), .Z(n3657) );
  XNOR U3819 ( .A(n3639), .B(n3659), .Z(n3654) );
  XNOR U3820 ( .A(n3652), .B(n3640), .Z(n3659) );
  XNOR U3821 ( .A(n3624), .B(n3623), .Z(n3640) );
  XOR U3822 ( .A(n3660), .B(n3618), .Z(n3623) );
  XNOR U3823 ( .A(n3616), .B(n3661), .Z(n3618) );
  ANDN U3824 ( .A(n1740), .B(n2618), .Z(n3661) );
  XOR U3825 ( .A(n3662), .B(n3663), .Z(n3616) );
  AND U3826 ( .A(n3664), .B(n3665), .Z(n3663) );
  XNOR U3827 ( .A(n3666), .B(n3662), .Z(n3665) );
  XOR U3828 ( .A(n3667), .B(n3620), .Z(n3660) );
  AND U3829 ( .A(n2616), .B(n1733), .Z(n3620) );
  IV U3830 ( .A(n3622), .Z(n3667) );
  XNOR U3831 ( .A(n3628), .B(n3630), .Z(n3624) );
  NAND U3832 ( .A(n2880), .B(n1538), .Z(n3630) );
  XNOR U3833 ( .A(n3626), .B(n3671), .Z(n3628) );
  ANDN U3834 ( .A(n1543), .B(n2882), .Z(n3671) );
  XOR U3835 ( .A(n3672), .B(n3673), .Z(n3626) );
  AND U3836 ( .A(n3674), .B(n3675), .Z(n3673) );
  XOR U3837 ( .A(n3676), .B(n3672), .Z(n3675) );
  XOR U3838 ( .A(n3677), .B(n3651), .Z(n3639) );
  XNOR U3839 ( .A(n3635), .B(n3637), .Z(n3651) );
  NAND U3840 ( .A(n2369), .B(n1934), .Z(n3637) );
  XNOR U3841 ( .A(n3633), .B(n3678), .Z(n3635) );
  ANDN U3842 ( .A(n1939), .B(n2371), .Z(n3678) );
  XOR U3843 ( .A(n3679), .B(n3680), .Z(n3633) );
  AND U3844 ( .A(n3681), .B(n3682), .Z(n3680) );
  XOR U3845 ( .A(n3683), .B(n3679), .Z(n3682) );
  XNOR U3846 ( .A(n3650), .B(n3638), .Z(n3677) );
  XOR U3847 ( .A(n3687), .B(n3645), .Z(n3650) );
  XNOR U3848 ( .A(n3643), .B(n3688), .Z(n3645) );
  ANDN U3849 ( .A(n2169), .B(n2132), .Z(n3688) );
  XOR U3850 ( .A(n3689), .B(n3690), .Z(n3643) );
  AND U3851 ( .A(n3691), .B(n3692), .Z(n3690) );
  XNOR U3852 ( .A(n3693), .B(n3689), .Z(n3692) );
  XOR U3853 ( .A(n3694), .B(n3647), .Z(n3687) );
  AND U3854 ( .A(n2130), .B(n2162), .Z(n3647) );
  IV U3855 ( .A(n3649), .Z(n3694) );
  XOR U3856 ( .A(n3698), .B(n3699), .Z(n3652) );
  AND U3857 ( .A(n3700), .B(n3701), .Z(n3699) );
  XOR U3858 ( .A(n3702), .B(n3703), .Z(n3701) );
  XOR U3859 ( .A(n3698), .B(n3704), .Z(n3703) );
  XNOR U3860 ( .A(n3685), .B(n3705), .Z(n3700) );
  XNOR U3861 ( .A(n3698), .B(n3686), .Z(n3705) );
  XNOR U3862 ( .A(n3670), .B(n3669), .Z(n3686) );
  XOR U3863 ( .A(n3706), .B(n3664), .Z(n3669) );
  XNOR U3864 ( .A(n3662), .B(n3707), .Z(n3664) );
  ANDN U3865 ( .A(n1740), .B(n2750), .Z(n3707) );
  XOR U3866 ( .A(n3711), .B(n3666), .Z(n3706) );
  AND U3867 ( .A(n2748), .B(n1733), .Z(n3666) );
  IV U3868 ( .A(n3668), .Z(n3711) );
  XNOR U3869 ( .A(n3674), .B(n3676), .Z(n3670) );
  NAND U3870 ( .A(n3019), .B(n1538), .Z(n3676) );
  XNOR U3871 ( .A(n3672), .B(n3715), .Z(n3674) );
  ANDN U3872 ( .A(n1543), .B(n3021), .Z(n3715) );
  XOR U3873 ( .A(n3719), .B(n3697), .Z(n3685) );
  XNOR U3874 ( .A(n3681), .B(n3683), .Z(n3697) );
  NAND U3875 ( .A(n2491), .B(n1934), .Z(n3683) );
  XNOR U3876 ( .A(n3679), .B(n3720), .Z(n3681) );
  ANDN U3877 ( .A(n1939), .B(n2493), .Z(n3720) );
  XOR U3878 ( .A(n3721), .B(n3722), .Z(n3679) );
  AND U3879 ( .A(n3723), .B(n3724), .Z(n3722) );
  XOR U3880 ( .A(n3725), .B(n3721), .Z(n3724) );
  XNOR U3881 ( .A(n3696), .B(n3684), .Z(n3719) );
  XOR U3882 ( .A(n3729), .B(n3691), .Z(n3696) );
  XNOR U3883 ( .A(n3689), .B(n3730), .Z(n3691) );
  ANDN U3884 ( .A(n2169), .B(n2251), .Z(n3730) );
  XOR U3885 ( .A(n3731), .B(n3732), .Z(n3689) );
  AND U3886 ( .A(n3733), .B(n3734), .Z(n3732) );
  XNOR U3887 ( .A(n3735), .B(n3731), .Z(n3734) );
  XOR U3888 ( .A(n3736), .B(n3693), .Z(n3729) );
  AND U3889 ( .A(n2249), .B(n2162), .Z(n3693) );
  IV U3890 ( .A(n3695), .Z(n3736) );
  XOR U3891 ( .A(n3741), .B(n3742), .Z(n3060) );
  XOR U3892 ( .A(n3743), .B(n3740), .Z(n3741) );
  XNOR U3893 ( .A(n3728), .B(n3727), .Z(n3059) );
  XOR U3894 ( .A(n3744), .B(n3739), .Z(n3727) );
  XNOR U3895 ( .A(n3723), .B(n3725), .Z(n3739) );
  NAND U3896 ( .A(n2616), .B(n1934), .Z(n3725) );
  XNOR U3897 ( .A(n3721), .B(n3745), .Z(n3723) );
  ANDN U3898 ( .A(n1939), .B(n2618), .Z(n3745) );
  XOR U3899 ( .A(n3738), .B(n3726), .Z(n3744) );
  XOR U3900 ( .A(n3749), .B(n3750), .Z(n3726) );
  XOR U3901 ( .A(n3751), .B(n3733), .Z(n3738) );
  XNOR U3902 ( .A(n3731), .B(n3752), .Z(n3733) );
  ANDN U3903 ( .A(n2169), .B(n2371), .Z(n3752) );
  AND U3904 ( .A(n2369), .B(n2162), .Z(n3735) );
  XNOR U3905 ( .A(n3756), .B(n3757), .Z(n3737) );
  AND U3906 ( .A(n3758), .B(n3759), .Z(n3757) );
  XNOR U3907 ( .A(n3754), .B(n3760), .Z(n3759) );
  XNOR U3908 ( .A(n3755), .B(n3756), .Z(n3760) );
  AND U3909 ( .A(n2491), .B(n2162), .Z(n3755) );
  XOR U3910 ( .A(n3753), .B(n3761), .Z(n3754) );
  ANDN U3911 ( .A(n2169), .B(n2493), .Z(n3761) );
  XNOR U3912 ( .A(n3747), .B(n3765), .Z(n3758) );
  XNOR U3913 ( .A(n3748), .B(n3756), .Z(n3765) );
  AND U3914 ( .A(n2748), .B(n1934), .Z(n3748) );
  XOR U3915 ( .A(n3746), .B(n3766), .Z(n3747) );
  ANDN U3916 ( .A(n1939), .B(n2750), .Z(n3766) );
  XOR U3917 ( .A(n3770), .B(n3771), .Z(n3756) );
  AND U3918 ( .A(n3772), .B(n3773), .Z(n3771) );
  XNOR U3919 ( .A(n3763), .B(n3774), .Z(n3773) );
  XNOR U3920 ( .A(n3764), .B(n3770), .Z(n3774) );
  AND U3921 ( .A(n2616), .B(n2162), .Z(n3764) );
  XOR U3922 ( .A(n3762), .B(n3775), .Z(n3763) );
  ANDN U3923 ( .A(n2169), .B(n2618), .Z(n3775) );
  XNOR U3924 ( .A(n3768), .B(n3779), .Z(n3772) );
  XNOR U3925 ( .A(n3769), .B(n3770), .Z(n3779) );
  AND U3926 ( .A(n2880), .B(n1934), .Z(n3769) );
  XOR U3927 ( .A(n3767), .B(n3780), .Z(n3768) );
  ANDN U3928 ( .A(n1939), .B(n2882), .Z(n3780) );
  XOR U3929 ( .A(n3784), .B(n3785), .Z(n3770) );
  AND U3930 ( .A(n3786), .B(n3787), .Z(n3785) );
  XNOR U3931 ( .A(n3777), .B(n3788), .Z(n3787) );
  XNOR U3932 ( .A(n3778), .B(n3784), .Z(n3788) );
  AND U3933 ( .A(n2748), .B(n2162), .Z(n3778) );
  XOR U3934 ( .A(n3776), .B(n3789), .Z(n3777) );
  ANDN U3935 ( .A(n2169), .B(n2750), .Z(n3789) );
  XNOR U3936 ( .A(n3782), .B(n3793), .Z(n3786) );
  XNOR U3937 ( .A(n3783), .B(n3784), .Z(n3793) );
  AND U3938 ( .A(n3019), .B(n1934), .Z(n3783) );
  XOR U3939 ( .A(n3781), .B(n3794), .Z(n3782) );
  ANDN U3940 ( .A(n1939), .B(n3021), .Z(n3794) );
  XNOR U3941 ( .A(n3799), .B(n3791), .Z(n3750) );
  XNOR U3942 ( .A(n3790), .B(n3800), .Z(n3791) );
  ANDN U3943 ( .A(n2169), .B(n2882), .Z(n3800) );
  XNOR U3944 ( .A(n3803), .B(n3801), .Z(n3802) );
  ANDN U3945 ( .A(n2169), .B(n3021), .Z(n3803) );
  XNOR U3946 ( .A(n3798), .B(n3792), .Z(n3799) );
  AND U3947 ( .A(n2880), .B(n2162), .Z(n3792) );
  XNOR U3948 ( .A(n3796), .B(n3797), .Z(n3749) );
  NAND U3949 ( .A(n3807), .B(n1934), .Z(n3797) );
  XNOR U3950 ( .A(n3795), .B(n3808), .Z(n3796) );
  ANDN U3951 ( .A(n1939), .B(n3809), .Z(n3808) );
  NAND U3952 ( .A(g_input[0]), .B(n3810), .Z(n3795) );
  NANDN U3953 ( .B(n1934), .A(n3811), .Z(n3810) );
  NANDN U3954 ( .B(n3812), .A(n1939), .Z(n3811) );
  IV U3955 ( .A(n1833), .Z(n1934) );
  XNOR U3956 ( .A(n3805), .B(n3806), .Z(n3798) );
  NAND U3957 ( .A(n3807), .B(n2162), .Z(n3806) );
  XNOR U3958 ( .A(n3804), .B(n3815), .Z(n3805) );
  ANDN U3959 ( .A(n2169), .B(n3809), .Z(n3815) );
  NAND U3960 ( .A(g_input[0]), .B(n3816), .Z(n3804) );
  NANDN U3961 ( .B(n2162), .A(n3817), .Z(n3816) );
  NANDN U3962 ( .B(n3812), .A(n2169), .Z(n3817) );
  IV U3963 ( .A(n2050), .Z(n2162) );
  XNOR U3964 ( .A(n3714), .B(n3713), .Z(n3728) );
  XOR U3965 ( .A(n3820), .B(n3709), .Z(n3713) );
  XNOR U3966 ( .A(n3708), .B(n3821), .Z(n3709) );
  ANDN U3967 ( .A(n1740), .B(n2882), .Z(n3821) );
  XNOR U3968 ( .A(n3824), .B(n3822), .Z(n3823) );
  ANDN U3969 ( .A(n1740), .B(n3021), .Z(n3824) );
  XNOR U3970 ( .A(n3712), .B(n3710), .Z(n3820) );
  AND U3971 ( .A(n2880), .B(n1733), .Z(n3710) );
  XNOR U3972 ( .A(n3826), .B(n3827), .Z(n3712) );
  NAND U3973 ( .A(n3807), .B(n1733), .Z(n3827) );
  XNOR U3974 ( .A(n3825), .B(n3828), .Z(n3826) );
  ANDN U3975 ( .A(n1740), .B(n3809), .Z(n3828) );
  NAND U3976 ( .A(g_input[0]), .B(n3829), .Z(n3825) );
  NANDN U3977 ( .B(n1733), .A(n3830), .Z(n3829) );
  NANDN U3978 ( .B(n3812), .A(n1740), .Z(n3830) );
  IV U3979 ( .A(n1634), .Z(n1733) );
  XNOR U3980 ( .A(n3717), .B(n3718), .Z(n3714) );
  NAND U3981 ( .A(n3807), .B(n1538), .Z(n3718) );
  XNOR U3982 ( .A(n3716), .B(n3833), .Z(n3717) );
  ANDN U3983 ( .A(n1543), .B(n3809), .Z(n3833) );
  NAND U3984 ( .A(g_input[0]), .B(n3834), .Z(n3716) );
  NANDN U3985 ( .B(n1538), .A(n3835), .Z(n3834) );
  NANDN U3986 ( .B(n3812), .A(n1543), .Z(n3835) );
  IV U3987 ( .A(n1442), .Z(n1538) );
  XNOR U3988 ( .A(n3838), .B(n3839), .Z(n3740) );
  XOR U3989 ( .A(n3840), .B(n2962), .Z(n2957) );
  XNOR U3990 ( .A(n2953), .B(n2954), .Z(n2962) );
  NAND U3991 ( .A(n2950), .B(n583), .Z(n2954) );
  XNOR U3992 ( .A(n2952), .B(n3841), .Z(n2953) );
  ANDN U3993 ( .A(n2955), .B(n585), .Z(n3841) );
  XOR U3994 ( .A(n3842), .B(n3843), .Z(n2952) );
  AND U3995 ( .A(n3844), .B(n3845), .Z(n3843) );
  XOR U3996 ( .A(n3846), .B(n3842), .Z(n3845) );
  XNOR U3997 ( .A(n2960), .B(n2956), .Z(n3840) );
  XNOR U3998 ( .A(n3071), .B(n3070), .Z(n3083) );
  XOR U3999 ( .A(n3848), .B(n3066), .Z(n3070) );
  XNOR U4000 ( .A(n3064), .B(n3849), .Z(n3066) );
  ANDN U4001 ( .A(n2678), .B(n713), .Z(n3849) );
  XOR U4002 ( .A(n3850), .B(n3851), .Z(n3064) );
  AND U4003 ( .A(n3852), .B(n3853), .Z(n3851) );
  XNOR U4004 ( .A(n3854), .B(n3850), .Z(n3853) );
  AND U4005 ( .A(n2671), .B(n711), .Z(n3068) );
  XNOR U4006 ( .A(n3075), .B(n3077), .Z(n3071) );
  NAND U4007 ( .A(n2424), .B(n812), .Z(n3077) );
  XNOR U4008 ( .A(n3073), .B(n3858), .Z(n3075) );
  ANDN U4009 ( .A(n2429), .B(n814), .Z(n3858) );
  XOR U4010 ( .A(n3859), .B(n3860), .Z(n3073) );
  AND U4011 ( .A(n3861), .B(n3862), .Z(n3860) );
  XOR U4012 ( .A(n3863), .B(n3859), .Z(n3862) );
  XOR U4013 ( .A(n3864), .B(n3865), .Z(n3084) );
  XNOR U4014 ( .A(n3866), .B(n3847), .Z(n3864) );
  XOR U4015 ( .A(n3868), .B(n3869), .Z(n3122) );
  XOR U4016 ( .A(n3870), .B(n3867), .Z(n3868) );
  XNOR U4017 ( .A(n3857), .B(n3856), .Z(n3120) );
  XOR U4018 ( .A(n3871), .B(n3852), .Z(n3856) );
  XNOR U4019 ( .A(n3850), .B(n3872), .Z(n3852) );
  ANDN U4020 ( .A(n2678), .B(n755), .Z(n3872) );
  XOR U4021 ( .A(n3873), .B(n3874), .Z(n3850) );
  AND U4022 ( .A(n3875), .B(n3876), .Z(n3874) );
  XNOR U4023 ( .A(n3877), .B(n3873), .Z(n3876) );
  XOR U4024 ( .A(n3878), .B(n3854), .Z(n3871) );
  AND U4025 ( .A(n2671), .B(n753), .Z(n3854) );
  IV U4026 ( .A(n3855), .Z(n3878) );
  XNOR U4027 ( .A(n3861), .B(n3863), .Z(n3857) );
  NAND U4028 ( .A(n2424), .B(n876), .Z(n3863) );
  XNOR U4029 ( .A(n3859), .B(n3882), .Z(n3861) );
  ANDN U4030 ( .A(n2429), .B(n878), .Z(n3882) );
  XOR U4031 ( .A(n3883), .B(n3884), .Z(n3859) );
  AND U4032 ( .A(n3885), .B(n3886), .Z(n3884) );
  XOR U4033 ( .A(n3887), .B(n3883), .Z(n3886) );
  XOR U4034 ( .A(n3889), .B(n3890), .Z(n3167) );
  XOR U4035 ( .A(n3891), .B(n3888), .Z(n3889) );
  XNOR U4036 ( .A(n3881), .B(n3880), .Z(n3165) );
  XOR U4037 ( .A(n3892), .B(n3875), .Z(n3880) );
  XNOR U4038 ( .A(n3873), .B(n3893), .Z(n3875) );
  ANDN U4039 ( .A(n2678), .B(n814), .Z(n3893) );
  XOR U4040 ( .A(n3894), .B(n3895), .Z(n3873) );
  AND U4041 ( .A(n3896), .B(n3897), .Z(n3895) );
  XNOR U4042 ( .A(n3898), .B(n3894), .Z(n3897) );
  XOR U4043 ( .A(n3899), .B(n3877), .Z(n3892) );
  AND U4044 ( .A(n2671), .B(n812), .Z(n3877) );
  IV U4045 ( .A(n3879), .Z(n3899) );
  XNOR U4046 ( .A(n3885), .B(n3887), .Z(n3881) );
  NAND U4047 ( .A(n2424), .B(n944), .Z(n3887) );
  XNOR U4048 ( .A(n3883), .B(n3903), .Z(n3885) );
  ANDN U4049 ( .A(n2429), .B(n946), .Z(n3903) );
  XOR U4050 ( .A(n3904), .B(n3905), .Z(n3883) );
  AND U4051 ( .A(n3906), .B(n3907), .Z(n3905) );
  XOR U4052 ( .A(n3908), .B(n3904), .Z(n3907) );
  XOR U4053 ( .A(n3910), .B(n3911), .Z(n3209) );
  XOR U4054 ( .A(n3912), .B(n3909), .Z(n3910) );
  XNOR U4055 ( .A(n3902), .B(n3901), .Z(n3207) );
  XOR U4056 ( .A(n3913), .B(n3896), .Z(n3901) );
  XNOR U4057 ( .A(n3894), .B(n3914), .Z(n3896) );
  ANDN U4058 ( .A(n2678), .B(n878), .Z(n3914) );
  XOR U4059 ( .A(n3915), .B(n3916), .Z(n3894) );
  AND U4060 ( .A(n3917), .B(n3918), .Z(n3916) );
  XNOR U4061 ( .A(n3919), .B(n3915), .Z(n3918) );
  AND U4062 ( .A(n2671), .B(n876), .Z(n3898) );
  XNOR U4063 ( .A(n3906), .B(n3908), .Z(n3902) );
  NAND U4064 ( .A(n2424), .B(n1011), .Z(n3908) );
  XNOR U4065 ( .A(n3904), .B(n3923), .Z(n3906) );
  ANDN U4066 ( .A(n2429), .B(n1013), .Z(n3923) );
  XOR U4067 ( .A(n3924), .B(n3925), .Z(n3904) );
  AND U4068 ( .A(n3926), .B(n3927), .Z(n3925) );
  XOR U4069 ( .A(n3928), .B(n3924), .Z(n3927) );
  XOR U4070 ( .A(n3930), .B(n3931), .Z(n3252) );
  XOR U4071 ( .A(n3932), .B(n3929), .Z(n3930) );
  XNOR U4072 ( .A(n3922), .B(n3921), .Z(n3250) );
  XOR U4073 ( .A(n3933), .B(n3917), .Z(n3921) );
  XNOR U4074 ( .A(n3915), .B(n3934), .Z(n3917) );
  ANDN U4075 ( .A(n2678), .B(n946), .Z(n3934) );
  XOR U4076 ( .A(n3935), .B(n3936), .Z(n3915) );
  AND U4077 ( .A(n3937), .B(n3938), .Z(n3936) );
  XNOR U4078 ( .A(n3939), .B(n3935), .Z(n3938) );
  XOR U4079 ( .A(n3940), .B(n3919), .Z(n3933) );
  AND U4080 ( .A(n2671), .B(n944), .Z(n3919) );
  IV U4081 ( .A(n3920), .Z(n3940) );
  XNOR U4082 ( .A(n3926), .B(n3928), .Z(n3922) );
  NAND U4083 ( .A(n2424), .B(n1085), .Z(n3928) );
  XNOR U4084 ( .A(n3924), .B(n3944), .Z(n3926) );
  ANDN U4085 ( .A(n2429), .B(n1087), .Z(n3944) );
  XOR U4086 ( .A(n3945), .B(n3946), .Z(n3924) );
  AND U4087 ( .A(n3947), .B(n3948), .Z(n3946) );
  XOR U4088 ( .A(n3949), .B(n3945), .Z(n3948) );
  XOR U4089 ( .A(n3951), .B(n3952), .Z(n3294) );
  XOR U4090 ( .A(n3953), .B(n3950), .Z(n3951) );
  XNOR U4091 ( .A(n3943), .B(n3942), .Z(n3292) );
  XOR U4092 ( .A(n3954), .B(n3937), .Z(n3942) );
  XNOR U4093 ( .A(n3935), .B(n3955), .Z(n3937) );
  ANDN U4094 ( .A(n2678), .B(n1013), .Z(n3955) );
  XOR U4095 ( .A(n3956), .B(n3957), .Z(n3935) );
  AND U4096 ( .A(n3958), .B(n3959), .Z(n3957) );
  XNOR U4097 ( .A(n3960), .B(n3956), .Z(n3959) );
  XOR U4098 ( .A(n3961), .B(n3939), .Z(n3954) );
  AND U4099 ( .A(n2671), .B(n1011), .Z(n3939) );
  IV U4100 ( .A(n3941), .Z(n3961) );
  XNOR U4101 ( .A(n3947), .B(n3949), .Z(n3943) );
  NAND U4102 ( .A(n2424), .B(n1163), .Z(n3949) );
  XNOR U4103 ( .A(n3945), .B(n3965), .Z(n3947) );
  ANDN U4104 ( .A(n2429), .B(n1165), .Z(n3965) );
  XOR U4105 ( .A(n3966), .B(n3967), .Z(n3945) );
  AND U4106 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR U4107 ( .A(n3970), .B(n3966), .Z(n3969) );
  XOR U4108 ( .A(n3972), .B(n3973), .Z(n3340) );
  XOR U4109 ( .A(n3974), .B(n3971), .Z(n3972) );
  XNOR U4110 ( .A(n3964), .B(n3963), .Z(n3338) );
  XOR U4111 ( .A(n3975), .B(n3958), .Z(n3963) );
  XNOR U4112 ( .A(n3956), .B(n3976), .Z(n3958) );
  ANDN U4113 ( .A(n2678), .B(n1087), .Z(n3976) );
  XOR U4114 ( .A(n3977), .B(n3978), .Z(n3956) );
  AND U4115 ( .A(n3979), .B(n3980), .Z(n3978) );
  XNOR U4116 ( .A(n3981), .B(n3977), .Z(n3980) );
  XOR U4117 ( .A(n3982), .B(n3960), .Z(n3975) );
  AND U4118 ( .A(n2671), .B(n1085), .Z(n3960) );
  IV U4119 ( .A(n3962), .Z(n3982) );
  XNOR U4120 ( .A(n3968), .B(n3970), .Z(n3964) );
  NAND U4121 ( .A(n2424), .B(n1244), .Z(n3970) );
  XNOR U4122 ( .A(n3966), .B(n3986), .Z(n3968) );
  ANDN U4123 ( .A(n2429), .B(n1246), .Z(n3986) );
  XOR U4124 ( .A(n3987), .B(n3988), .Z(n3966) );
  AND U4125 ( .A(n3989), .B(n3990), .Z(n3988) );
  XOR U4126 ( .A(n3991), .B(n3987), .Z(n3990) );
  XOR U4127 ( .A(n3993), .B(n3994), .Z(n3384) );
  XOR U4128 ( .A(n3995), .B(n3992), .Z(n3993) );
  XNOR U4129 ( .A(n3985), .B(n3984), .Z(n3382) );
  XOR U4130 ( .A(n3996), .B(n3979), .Z(n3984) );
  XNOR U4131 ( .A(n3977), .B(n3997), .Z(n3979) );
  ANDN U4132 ( .A(n2678), .B(n1165), .Z(n3997) );
  XOR U4133 ( .A(n3998), .B(n3999), .Z(n3977) );
  AND U4134 ( .A(n4000), .B(n4001), .Z(n3999) );
  XNOR U4135 ( .A(n4002), .B(n3998), .Z(n4001) );
  XOR U4136 ( .A(n4003), .B(n3981), .Z(n3996) );
  AND U4137 ( .A(n2671), .B(n1163), .Z(n3981) );
  IV U4138 ( .A(n3983), .Z(n4003) );
  XNOR U4139 ( .A(n3989), .B(n3991), .Z(n3985) );
  NAND U4140 ( .A(n2424), .B(n1328), .Z(n3991) );
  XNOR U4141 ( .A(n3987), .B(n4007), .Z(n3989) );
  ANDN U4142 ( .A(n2429), .B(n1330), .Z(n4007) );
  XOR U4143 ( .A(n4008), .B(n4009), .Z(n3987) );
  AND U4144 ( .A(n4010), .B(n4011), .Z(n4009) );
  XOR U4145 ( .A(n4012), .B(n4008), .Z(n4011) );
  XOR U4146 ( .A(n4014), .B(n4015), .Z(n3430) );
  XOR U4147 ( .A(n4016), .B(n4013), .Z(n4014) );
  XNOR U4148 ( .A(n4006), .B(n4005), .Z(n3428) );
  XOR U4149 ( .A(n4017), .B(n4000), .Z(n4005) );
  XNOR U4150 ( .A(n3998), .B(n4018), .Z(n4000) );
  ANDN U4151 ( .A(n2678), .B(n1246), .Z(n4018) );
  XOR U4152 ( .A(n4019), .B(n4020), .Z(n3998) );
  AND U4153 ( .A(n4021), .B(n4022), .Z(n4020) );
  XNOR U4154 ( .A(n4023), .B(n4019), .Z(n4022) );
  XOR U4155 ( .A(n4024), .B(n4002), .Z(n4017) );
  AND U4156 ( .A(n2671), .B(n1244), .Z(n4002) );
  IV U4157 ( .A(n4004), .Z(n4024) );
  XNOR U4158 ( .A(n4010), .B(n4012), .Z(n4006) );
  NAND U4159 ( .A(n2424), .B(n1419), .Z(n4012) );
  XNOR U4160 ( .A(n4008), .B(n4028), .Z(n4010) );
  ANDN U4161 ( .A(n2429), .B(n1421), .Z(n4028) );
  XOR U4162 ( .A(n4029), .B(n4030), .Z(n4008) );
  AND U4163 ( .A(n4031), .B(n4032), .Z(n4030) );
  XOR U4164 ( .A(n4033), .B(n4029), .Z(n4032) );
  XOR U4165 ( .A(n4035), .B(n4036), .Z(n3476) );
  XOR U4166 ( .A(n4037), .B(n4034), .Z(n4035) );
  XNOR U4167 ( .A(n4027), .B(n4026), .Z(n3474) );
  XOR U4168 ( .A(n4038), .B(n4021), .Z(n4026) );
  XNOR U4169 ( .A(n4019), .B(n4039), .Z(n4021) );
  ANDN U4170 ( .A(n2678), .B(n1330), .Z(n4039) );
  XOR U4171 ( .A(n4040), .B(n4041), .Z(n4019) );
  AND U4172 ( .A(n4042), .B(n4043), .Z(n4041) );
  XNOR U4173 ( .A(n4044), .B(n4040), .Z(n4043) );
  XOR U4174 ( .A(n4045), .B(n4023), .Z(n4038) );
  AND U4175 ( .A(n2671), .B(n1328), .Z(n4023) );
  IV U4176 ( .A(n4025), .Z(n4045) );
  XNOR U4177 ( .A(n4031), .B(n4033), .Z(n4027) );
  NAND U4178 ( .A(n2424), .B(n1516), .Z(n4033) );
  XNOR U4179 ( .A(n4029), .B(n4049), .Z(n4031) );
  ANDN U4180 ( .A(n2429), .B(n1518), .Z(n4049) );
  XOR U4181 ( .A(n4050), .B(n4051), .Z(n4029) );
  AND U4182 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U4183 ( .A(n4054), .B(n4050), .Z(n4053) );
  XOR U4184 ( .A(n4056), .B(n4057), .Z(n3522) );
  XOR U4185 ( .A(n4058), .B(n4055), .Z(n4056) );
  XNOR U4186 ( .A(n4048), .B(n4047), .Z(n3520) );
  XOR U4187 ( .A(n4059), .B(n4042), .Z(n4047) );
  XNOR U4188 ( .A(n4040), .B(n4060), .Z(n4042) );
  ANDN U4189 ( .A(n2678), .B(n1421), .Z(n4060) );
  XOR U4190 ( .A(n4061), .B(n4062), .Z(n4040) );
  AND U4191 ( .A(n4063), .B(n4064), .Z(n4062) );
  XNOR U4192 ( .A(n4065), .B(n4061), .Z(n4064) );
  XOR U4193 ( .A(n4066), .B(n4044), .Z(n4059) );
  AND U4194 ( .A(n2671), .B(n1419), .Z(n4044) );
  IV U4195 ( .A(n4046), .Z(n4066) );
  XNOR U4196 ( .A(n4052), .B(n4054), .Z(n4048) );
  NAND U4197 ( .A(n2424), .B(n1612), .Z(n4054) );
  XNOR U4198 ( .A(n4050), .B(n4070), .Z(n4052) );
  ANDN U4199 ( .A(n2429), .B(n1614), .Z(n4070) );
  XOR U4200 ( .A(n4071), .B(n4072), .Z(n4050) );
  AND U4201 ( .A(n4073), .B(n4074), .Z(n4072) );
  XOR U4202 ( .A(n4075), .B(n4071), .Z(n4074) );
  XOR U4203 ( .A(n4077), .B(n4078), .Z(n3566) );
  XOR U4204 ( .A(n4079), .B(n4076), .Z(n4077) );
  XNOR U4205 ( .A(n4069), .B(n4068), .Z(n3564) );
  XOR U4206 ( .A(n4080), .B(n4063), .Z(n4068) );
  XNOR U4207 ( .A(n4061), .B(n4081), .Z(n4063) );
  ANDN U4208 ( .A(n2678), .B(n1518), .Z(n4081) );
  XOR U4209 ( .A(n4082), .B(n4083), .Z(n4061) );
  AND U4210 ( .A(n4084), .B(n4085), .Z(n4083) );
  XNOR U4211 ( .A(n4086), .B(n4082), .Z(n4085) );
  XOR U4212 ( .A(n4087), .B(n4065), .Z(n4080) );
  AND U4213 ( .A(n2671), .B(n1516), .Z(n4065) );
  IV U4214 ( .A(n4067), .Z(n4087) );
  XNOR U4215 ( .A(n4073), .B(n4075), .Z(n4069) );
  NAND U4216 ( .A(n2424), .B(n1708), .Z(n4075) );
  XNOR U4217 ( .A(n4071), .B(n4091), .Z(n4073) );
  ANDN U4218 ( .A(n2429), .B(n1710), .Z(n4091) );
  XOR U4219 ( .A(n4092), .B(n4093), .Z(n4071) );
  AND U4220 ( .A(n4094), .B(n4095), .Z(n4093) );
  XOR U4221 ( .A(n4096), .B(n4092), .Z(n4095) );
  XOR U4222 ( .A(n4098), .B(n4099), .Z(n3612) );
  XOR U4223 ( .A(n4100), .B(n4097), .Z(n4098) );
  XNOR U4224 ( .A(n4090), .B(n4089), .Z(n3610) );
  XOR U4225 ( .A(n4101), .B(n4084), .Z(n4089) );
  XNOR U4226 ( .A(n4082), .B(n4102), .Z(n4084) );
  ANDN U4227 ( .A(n2678), .B(n1614), .Z(n4102) );
  XOR U4228 ( .A(n4103), .B(n4104), .Z(n4082) );
  AND U4229 ( .A(n4105), .B(n4106), .Z(n4104) );
  XNOR U4230 ( .A(n4107), .B(n4103), .Z(n4106) );
  XOR U4231 ( .A(n4108), .B(n4086), .Z(n4101) );
  AND U4232 ( .A(n2671), .B(n1612), .Z(n4086) );
  IV U4233 ( .A(n4088), .Z(n4108) );
  XNOR U4234 ( .A(n4094), .B(n4096), .Z(n4090) );
  NAND U4235 ( .A(n2424), .B(n1809), .Z(n4096) );
  XNOR U4236 ( .A(n4092), .B(n4112), .Z(n4094) );
  ANDN U4237 ( .A(n2429), .B(n1811), .Z(n4112) );
  XOR U4238 ( .A(n4113), .B(n4114), .Z(n4092) );
  AND U4239 ( .A(n4115), .B(n4116), .Z(n4114) );
  XOR U4240 ( .A(n4117), .B(n4113), .Z(n4116) );
  XOR U4241 ( .A(n4119), .B(n4120), .Z(n3658) );
  XOR U4242 ( .A(n4121), .B(n4118), .Z(n4119) );
  XNOR U4243 ( .A(n4111), .B(n4110), .Z(n3656) );
  XOR U4244 ( .A(n4122), .B(n4105), .Z(n4110) );
  XNOR U4245 ( .A(n4103), .B(n4123), .Z(n4105) );
  ANDN U4246 ( .A(n2678), .B(n1710), .Z(n4123) );
  XOR U4247 ( .A(n4124), .B(n4125), .Z(n4103) );
  AND U4248 ( .A(n4126), .B(n4127), .Z(n4125) );
  XNOR U4249 ( .A(n4128), .B(n4124), .Z(n4127) );
  XOR U4250 ( .A(n4129), .B(n4107), .Z(n4122) );
  AND U4251 ( .A(n2671), .B(n1708), .Z(n4107) );
  IV U4252 ( .A(n4109), .Z(n4129) );
  XNOR U4253 ( .A(n4115), .B(n4117), .Z(n4111) );
  NAND U4254 ( .A(n2424), .B(n1915), .Z(n4117) );
  XNOR U4255 ( .A(n4113), .B(n4133), .Z(n4115) );
  ANDN U4256 ( .A(n2429), .B(n1917), .Z(n4133) );
  XOR U4257 ( .A(n4134), .B(n4135), .Z(n4113) );
  AND U4258 ( .A(n4136), .B(n4137), .Z(n4135) );
  XOR U4259 ( .A(n4138), .B(n4134), .Z(n4137) );
  XOR U4260 ( .A(n4140), .B(n4141), .Z(n3704) );
  XOR U4261 ( .A(n4142), .B(n4139), .Z(n4140) );
  XNOR U4262 ( .A(n4132), .B(n4131), .Z(n3702) );
  XOR U4263 ( .A(n4143), .B(n4126), .Z(n4131) );
  XNOR U4264 ( .A(n4124), .B(n4144), .Z(n4126) );
  ANDN U4265 ( .A(n2678), .B(n1811), .Z(n4144) );
  XOR U4266 ( .A(n4145), .B(n4146), .Z(n4124) );
  AND U4267 ( .A(n4147), .B(n4148), .Z(n4146) );
  XNOR U4268 ( .A(n4149), .B(n4145), .Z(n4148) );
  XOR U4269 ( .A(n4150), .B(n4128), .Z(n4143) );
  AND U4270 ( .A(n2671), .B(n1809), .Z(n4128) );
  IV U4271 ( .A(n4130), .Z(n4150) );
  XNOR U4272 ( .A(n4136), .B(n4138), .Z(n4132) );
  NAND U4273 ( .A(n2424), .B(n2022), .Z(n4138) );
  XNOR U4274 ( .A(n4134), .B(n4154), .Z(n4136) );
  ANDN U4275 ( .A(n2429), .B(n2024), .Z(n4154) );
  XOR U4276 ( .A(n4155), .B(n4156), .Z(n4134) );
  AND U4277 ( .A(n4157), .B(n4158), .Z(n4156) );
  XOR U4278 ( .A(n4159), .B(n4155), .Z(n4158) );
  XOR U4279 ( .A(n4161), .B(n4162), .Z(n3743) );
  XOR U4280 ( .A(n4163), .B(n4160), .Z(n4161) );
  XNOR U4281 ( .A(n4153), .B(n4152), .Z(n3742) );
  XOR U4282 ( .A(n4164), .B(n4147), .Z(n4152) );
  XNOR U4283 ( .A(n4145), .B(n4165), .Z(n4147) );
  ANDN U4284 ( .A(n2678), .B(n1917), .Z(n4165) );
  AND U4285 ( .A(n2671), .B(n1915), .Z(n4149) );
  XNOR U4286 ( .A(n4157), .B(n4159), .Z(n4153) );
  NAND U4287 ( .A(n2424), .B(n2130), .Z(n4159) );
  XNOR U4288 ( .A(n4155), .B(n4172), .Z(n4157) );
  ANDN U4289 ( .A(n2429), .B(n2132), .Z(n4172) );
  XOR U4290 ( .A(n4176), .B(n4177), .Z(n4160) );
  AND U4291 ( .A(n4178), .B(n4179), .Z(n4177) );
  XOR U4292 ( .A(n4180), .B(n4181), .Z(n4179) );
  XNOR U4293 ( .A(n4176), .B(n4182), .Z(n4181) );
  XNOR U4294 ( .A(n4170), .B(n4183), .Z(n4178) );
  XNOR U4295 ( .A(n4176), .B(n4171), .Z(n4183) );
  XNOR U4296 ( .A(n4174), .B(n4175), .Z(n4171) );
  NAND U4297 ( .A(n2249), .B(n2424), .Z(n4175) );
  XNOR U4298 ( .A(n4173), .B(n4184), .Z(n4174) );
  ANDN U4299 ( .A(n2429), .B(n2251), .Z(n4184) );
  XOR U4300 ( .A(n4188), .B(n4167), .Z(n4170) );
  XNOR U4301 ( .A(n4166), .B(n4189), .Z(n4167) );
  ANDN U4302 ( .A(n2678), .B(n2024), .Z(n4189) );
  AND U4303 ( .A(n2671), .B(n2022), .Z(n4168) );
  XOR U4304 ( .A(n4196), .B(n4197), .Z(n4176) );
  AND U4305 ( .A(n4198), .B(n4199), .Z(n4197) );
  XOR U4306 ( .A(n4200), .B(n4201), .Z(n4199) );
  XNOR U4307 ( .A(n4196), .B(n4202), .Z(n4201) );
  XNOR U4308 ( .A(n4194), .B(n4203), .Z(n4198) );
  XNOR U4309 ( .A(n4196), .B(n4195), .Z(n4203) );
  XNOR U4310 ( .A(n4186), .B(n4187), .Z(n4195) );
  NAND U4311 ( .A(n2369), .B(n2424), .Z(n4187) );
  XNOR U4312 ( .A(n4185), .B(n4204), .Z(n4186) );
  ANDN U4313 ( .A(n2429), .B(n2371), .Z(n4204) );
  XOR U4314 ( .A(n4208), .B(n4191), .Z(n4194) );
  XNOR U4315 ( .A(n4190), .B(n4209), .Z(n4191) );
  ANDN U4316 ( .A(n2678), .B(n2132), .Z(n4209) );
  AND U4317 ( .A(n2671), .B(n2130), .Z(n4192) );
  XOR U4318 ( .A(n4216), .B(n4217), .Z(n4196) );
  AND U4319 ( .A(n4218), .B(n4219), .Z(n4217) );
  XOR U4320 ( .A(n4220), .B(n4221), .Z(n4219) );
  XNOR U4321 ( .A(n4216), .B(n4222), .Z(n4221) );
  XNOR U4322 ( .A(n4214), .B(n4223), .Z(n4218) );
  XNOR U4323 ( .A(n4216), .B(n4215), .Z(n4223) );
  XNOR U4324 ( .A(n4206), .B(n4207), .Z(n4215) );
  NAND U4325 ( .A(n2491), .B(n2424), .Z(n4207) );
  XNOR U4326 ( .A(n4205), .B(n4224), .Z(n4206) );
  ANDN U4327 ( .A(n2429), .B(n2493), .Z(n4224) );
  XOR U4328 ( .A(n4228), .B(n4211), .Z(n4214) );
  XNOR U4329 ( .A(n4210), .B(n4229), .Z(n4211) );
  ANDN U4330 ( .A(n2678), .B(n2251), .Z(n4229) );
  AND U4331 ( .A(n2249), .B(n2671), .Z(n4212) );
  XOR U4332 ( .A(n4236), .B(n4237), .Z(n4216) );
  AND U4333 ( .A(n4238), .B(n4239), .Z(n4237) );
  XOR U4334 ( .A(n4240), .B(n4241), .Z(n4239) );
  XNOR U4335 ( .A(n4236), .B(n4242), .Z(n4241) );
  XNOR U4336 ( .A(n4234), .B(n4243), .Z(n4238) );
  XNOR U4337 ( .A(n4236), .B(n4235), .Z(n4243) );
  XNOR U4338 ( .A(n4226), .B(n4227), .Z(n4235) );
  NAND U4339 ( .A(n2616), .B(n2424), .Z(n4227) );
  XNOR U4340 ( .A(n4225), .B(n4244), .Z(n4226) );
  ANDN U4341 ( .A(n2429), .B(n2618), .Z(n4244) );
  XOR U4342 ( .A(n4248), .B(n4231), .Z(n4234) );
  XNOR U4343 ( .A(n4230), .B(n4249), .Z(n4231) );
  ANDN U4344 ( .A(n2678), .B(n2371), .Z(n4249) );
  AND U4345 ( .A(n2369), .B(n2671), .Z(n4232) );
  XOR U4346 ( .A(n4256), .B(n4257), .Z(n4236) );
  AND U4347 ( .A(n4258), .B(n4259), .Z(n4257) );
  XOR U4348 ( .A(n4260), .B(n4261), .Z(n4259) );
  XNOR U4349 ( .A(n4256), .B(n4262), .Z(n4261) );
  XNOR U4350 ( .A(n4254), .B(n4263), .Z(n4258) );
  XNOR U4351 ( .A(n4256), .B(n4255), .Z(n4263) );
  XNOR U4352 ( .A(n4246), .B(n4247), .Z(n4255) );
  NAND U4353 ( .A(n2748), .B(n2424), .Z(n4247) );
  XNOR U4354 ( .A(n4245), .B(n4264), .Z(n4246) );
  ANDN U4355 ( .A(n2429), .B(n2750), .Z(n4264) );
  XOR U4356 ( .A(n4268), .B(n4251), .Z(n4254) );
  XNOR U4357 ( .A(n4250), .B(n4269), .Z(n4251) );
  ANDN U4358 ( .A(n2678), .B(n2493), .Z(n4269) );
  AND U4359 ( .A(n2491), .B(n2671), .Z(n4252) );
  XOR U4360 ( .A(n4276), .B(n4277), .Z(n4256) );
  AND U4361 ( .A(n4278), .B(n4279), .Z(n4277) );
  XOR U4362 ( .A(n4280), .B(n4281), .Z(n4279) );
  XNOR U4363 ( .A(n4276), .B(n4282), .Z(n4281) );
  XNOR U4364 ( .A(n4274), .B(n4283), .Z(n4278) );
  XNOR U4365 ( .A(n4276), .B(n4275), .Z(n4283) );
  XNOR U4366 ( .A(n4266), .B(n4267), .Z(n4275) );
  NAND U4367 ( .A(n2880), .B(n2424), .Z(n4267) );
  XNOR U4368 ( .A(n4265), .B(n4284), .Z(n4266) );
  ANDN U4369 ( .A(n2429), .B(n2882), .Z(n4284) );
  XOR U4370 ( .A(n4285), .B(n4286), .Z(n4265) );
  AND U4371 ( .A(n4287), .B(n4288), .Z(n4286) );
  XOR U4372 ( .A(n4289), .B(n4285), .Z(n4288) );
  XOR U4373 ( .A(n4290), .B(n4271), .Z(n4274) );
  XNOR U4374 ( .A(n4270), .B(n4291), .Z(n4271) );
  ANDN U4375 ( .A(n2678), .B(n2618), .Z(n4291) );
  XOR U4376 ( .A(n4292), .B(n4293), .Z(n4270) );
  AND U4377 ( .A(n4294), .B(n4295), .Z(n4293) );
  XNOR U4378 ( .A(n4296), .B(n4292), .Z(n4295) );
  AND U4379 ( .A(n2616), .B(n2671), .Z(n4272) );
  XOR U4380 ( .A(n4300), .B(n4301), .Z(n4276) );
  AND U4381 ( .A(n4302), .B(n4303), .Z(n4301) );
  XOR U4382 ( .A(n4304), .B(n4305), .Z(n4303) );
  XNOR U4383 ( .A(n4300), .B(n4306), .Z(n4305) );
  XNOR U4384 ( .A(n4298), .B(n4307), .Z(n4302) );
  XNOR U4385 ( .A(n4300), .B(n4299), .Z(n4307) );
  XNOR U4386 ( .A(n4287), .B(n4289), .Z(n4299) );
  NAND U4387 ( .A(n3019), .B(n2424), .Z(n4289) );
  XNOR U4388 ( .A(n4285), .B(n4308), .Z(n4287) );
  ANDN U4389 ( .A(n2429), .B(n3021), .Z(n4308) );
  XOR U4390 ( .A(n4312), .B(n4294), .Z(n4298) );
  XNOR U4391 ( .A(n4292), .B(n4313), .Z(n4294) );
  ANDN U4392 ( .A(n2678), .B(n2750), .Z(n4313) );
  XOR U4393 ( .A(n4314), .B(n4315), .Z(n4292) );
  AND U4394 ( .A(n4316), .B(n4317), .Z(n4315) );
  XNOR U4395 ( .A(n4318), .B(n4314), .Z(n4317) );
  AND U4396 ( .A(n2748), .B(n2671), .Z(n4296) );
  XOR U4397 ( .A(n4323), .B(n4324), .Z(n3839) );
  XNOR U4398 ( .A(n4321), .B(n4320), .Z(n3838) );
  XOR U4399 ( .A(n4326), .B(n4316), .Z(n4320) );
  XNOR U4400 ( .A(n4314), .B(n4327), .Z(n4316) );
  ANDN U4401 ( .A(n2678), .B(n2882), .Z(n4327) );
  XNOR U4402 ( .A(n4330), .B(n4328), .Z(n4329) );
  ANDN U4403 ( .A(n2678), .B(n3021), .Z(n4330) );
  XNOR U4404 ( .A(n4319), .B(n4318), .Z(n4326) );
  AND U4405 ( .A(n2880), .B(n2671), .Z(n4318) );
  XNOR U4406 ( .A(n4332), .B(n4333), .Z(n4319) );
  NAND U4407 ( .A(n3807), .B(n2671), .Z(n4333) );
  XNOR U4408 ( .A(n4331), .B(n4334), .Z(n4332) );
  ANDN U4409 ( .A(n2678), .B(n3809), .Z(n4334) );
  NAND U4410 ( .A(g_input[0]), .B(n4335), .Z(n4331) );
  NANDN U4411 ( .B(n2671), .A(n4336), .Z(n4335) );
  NANDN U4412 ( .B(n3812), .A(n2678), .Z(n4336) );
  IV U4413 ( .A(n2545), .Z(n2671) );
  XNOR U4414 ( .A(n4310), .B(n4311), .Z(n4321) );
  NAND U4415 ( .A(n3807), .B(n2424), .Z(n4311) );
  XNOR U4416 ( .A(n4309), .B(n4339), .Z(n4310) );
  ANDN U4417 ( .A(n2429), .B(n3809), .Z(n4339) );
  NAND U4418 ( .A(g_input[0]), .B(n4340), .Z(n4309) );
  NANDN U4419 ( .B(n2424), .A(n4341), .Z(n4340) );
  NANDN U4420 ( .B(n3812), .A(n2429), .Z(n4341) );
  IV U4421 ( .A(n2303), .Z(n2424) );
  XOR U4422 ( .A(n4344), .B(n4345), .Z(n4322) );
  XOR U4423 ( .A(n2959), .B(n4346), .Z(n2960) );
  AND U4424 ( .A(n4347), .B(n4348), .Z(n4346) );
  NANDN U4425 ( .B(n4349), .A(n522), .Z(n4348) );
  NANDN U4426 ( .B(n4350), .A(n4351), .Z(n4347) );
  XNOR U4427 ( .A(n3844), .B(n3846), .Z(n3865) );
  NAND U4428 ( .A(n2950), .B(n627), .Z(n3846) );
  XNOR U4429 ( .A(n3842), .B(n4353), .Z(n3844) );
  ANDN U4430 ( .A(n2955), .B(n629), .Z(n4353) );
  XOR U4431 ( .A(n4354), .B(n4355), .Z(n3842) );
  AND U4432 ( .A(n4356), .B(n4357), .Z(n4355) );
  XOR U4433 ( .A(n4358), .B(n4354), .Z(n4357) );
  XNOR U4434 ( .A(n4359), .B(n4360), .Z(n3866) );
  IV U4435 ( .A(n4352), .Z(n4360) );
  XOR U4436 ( .A(n4361), .B(n4351), .Z(n4359) );
  AND U4437 ( .A(n4362), .B(n552), .Z(n4351) );
  IV U4438 ( .A(n585), .Z(n552) );
  NAND U4439 ( .A(n4363), .B(n4350), .Z(n4361) );
  XOR U4440 ( .A(n4364), .B(n4365), .Z(n4350) );
  AND U4441 ( .A(n4366), .B(n4367), .Z(n4365) );
  XNOR U4442 ( .A(n4368), .B(n4364), .Z(n4367) );
  NANDN U4443 ( .B(n555), .A(e_input[0]), .Z(n4363) );
  IV U4444 ( .A(n522), .Z(n555) );
  AND U4445 ( .A(n4369), .B(n4370), .Z(n522) );
  ANDN U4446 ( .A(g_input[31]), .B(n4371), .Z(n4369) );
  XNOR U4447 ( .A(n4356), .B(n4358), .Z(n3869) );
  NAND U4448 ( .A(n2950), .B(n667), .Z(n4358) );
  XNOR U4449 ( .A(n4354), .B(n4373), .Z(n4356) );
  ANDN U4450 ( .A(n2955), .B(n669), .Z(n4373) );
  XOR U4451 ( .A(n4374), .B(n4375), .Z(n4354) );
  AND U4452 ( .A(n4376), .B(n4377), .Z(n4375) );
  XOR U4453 ( .A(n4378), .B(n4374), .Z(n4377) );
  XNOR U4454 ( .A(n4379), .B(n4366), .Z(n3870) );
  XNOR U4455 ( .A(n4364), .B(n4380), .Z(n4366) );
  ANDN U4456 ( .A(e_input[0]), .B(n585), .Z(n4380) );
  XNOR U4457 ( .A(n4371), .B(g_input[30]), .Z(n4370) );
  NANDN U4458 ( .B(n4381), .A(n4382), .Z(n4371) );
  XOR U4459 ( .A(n4383), .B(n4384), .Z(n4364) );
  AND U4460 ( .A(n4385), .B(n4386), .Z(n4384) );
  XNOR U4461 ( .A(n4387), .B(n4383), .Z(n4386) );
  XOR U4462 ( .A(n4388), .B(n4368), .Z(n4379) );
  AND U4463 ( .A(n4362), .B(n583), .Z(n4368) );
  IV U4464 ( .A(n629), .Z(n583) );
  IV U4465 ( .A(n4372), .Z(n4388) );
  XNOR U4466 ( .A(n4376), .B(n4378), .Z(n3890) );
  NAND U4467 ( .A(n2950), .B(n711), .Z(n4378) );
  XNOR U4468 ( .A(n4374), .B(n4390), .Z(n4376) );
  ANDN U4469 ( .A(n2955), .B(n713), .Z(n4390) );
  XOR U4470 ( .A(n4391), .B(n4392), .Z(n4374) );
  AND U4471 ( .A(n4393), .B(n4394), .Z(n4392) );
  XOR U4472 ( .A(n4395), .B(n4391), .Z(n4394) );
  XNOR U4473 ( .A(n4396), .B(n4385), .Z(n3891) );
  XNOR U4474 ( .A(n4383), .B(n4397), .Z(n4385) );
  ANDN U4475 ( .A(e_input[0]), .B(n629), .Z(n4397) );
  XNOR U4476 ( .A(n4382), .B(g_input[29]), .Z(n4381) );
  ANDN U4477 ( .A(n4398), .B(n4399), .Z(n4382) );
  XOR U4478 ( .A(n4400), .B(n4401), .Z(n4383) );
  AND U4479 ( .A(n4402), .B(n4403), .Z(n4401) );
  XNOR U4480 ( .A(n4404), .B(n4400), .Z(n4403) );
  XOR U4481 ( .A(n4405), .B(n4387), .Z(n4396) );
  AND U4482 ( .A(n4362), .B(n627), .Z(n4387) );
  IV U4483 ( .A(n669), .Z(n627) );
  IV U4484 ( .A(n4389), .Z(n4405) );
  XNOR U4485 ( .A(n4393), .B(n4395), .Z(n3911) );
  NAND U4486 ( .A(n2950), .B(n753), .Z(n4395) );
  XNOR U4487 ( .A(n4391), .B(n4407), .Z(n4393) );
  ANDN U4488 ( .A(n2955), .B(n755), .Z(n4407) );
  XOR U4489 ( .A(n4408), .B(n4409), .Z(n4391) );
  AND U4490 ( .A(n4410), .B(n4411), .Z(n4409) );
  XOR U4491 ( .A(n4412), .B(n4408), .Z(n4411) );
  XNOR U4492 ( .A(n4413), .B(n4402), .Z(n3912) );
  XNOR U4493 ( .A(n4400), .B(n4414), .Z(n4402) );
  ANDN U4494 ( .A(e_input[0]), .B(n669), .Z(n4414) );
  XNOR U4495 ( .A(n4398), .B(g_input[28]), .Z(n4399) );
  ANDN U4496 ( .A(n4415), .B(n4416), .Z(n4398) );
  XOR U4497 ( .A(n4417), .B(n4418), .Z(n4400) );
  AND U4498 ( .A(n4419), .B(n4420), .Z(n4418) );
  XNOR U4499 ( .A(n4421), .B(n4417), .Z(n4420) );
  AND U4500 ( .A(n4362), .B(n667), .Z(n4404) );
  IV U4501 ( .A(n713), .Z(n667) );
  XNOR U4502 ( .A(n4410), .B(n4412), .Z(n3931) );
  NAND U4503 ( .A(n2950), .B(n812), .Z(n4412) );
  XNOR U4504 ( .A(n4408), .B(n4423), .Z(n4410) );
  ANDN U4505 ( .A(n2955), .B(n814), .Z(n4423) );
  XOR U4506 ( .A(n4424), .B(n4425), .Z(n4408) );
  AND U4507 ( .A(n4426), .B(n4427), .Z(n4425) );
  XOR U4508 ( .A(n4428), .B(n4424), .Z(n4427) );
  XNOR U4509 ( .A(n4429), .B(n4419), .Z(n3932) );
  XNOR U4510 ( .A(n4417), .B(n4430), .Z(n4419) );
  ANDN U4511 ( .A(e_input[0]), .B(n713), .Z(n4430) );
  ANDN U4512 ( .A(n4431), .B(n4432), .Z(n4415) );
  XOR U4513 ( .A(n4433), .B(n4434), .Z(n4417) );
  AND U4514 ( .A(n4435), .B(n4436), .Z(n4434) );
  XNOR U4515 ( .A(n4437), .B(n4433), .Z(n4436) );
  AND U4516 ( .A(n4362), .B(n711), .Z(n4421) );
  IV U4517 ( .A(n755), .Z(n711) );
  XNOR U4518 ( .A(n4426), .B(n4428), .Z(n3952) );
  NAND U4519 ( .A(n2950), .B(n876), .Z(n4428) );
  XNOR U4520 ( .A(n4424), .B(n4439), .Z(n4426) );
  ANDN U4521 ( .A(n2955), .B(n878), .Z(n4439) );
  XOR U4522 ( .A(n4440), .B(n4441), .Z(n4424) );
  AND U4523 ( .A(n4442), .B(n4443), .Z(n4441) );
  XOR U4524 ( .A(n4444), .B(n4440), .Z(n4443) );
  XNOR U4525 ( .A(n4445), .B(n4435), .Z(n3953) );
  XNOR U4526 ( .A(n4433), .B(n4446), .Z(n4435) );
  ANDN U4527 ( .A(e_input[0]), .B(n755), .Z(n4446) );
  XNOR U4528 ( .A(n4431), .B(g_input[26]), .Z(n4432) );
  ANDN U4529 ( .A(n4447), .B(n4448), .Z(n4431) );
  XOR U4530 ( .A(n4449), .B(n4450), .Z(n4433) );
  AND U4531 ( .A(n4451), .B(n4452), .Z(n4450) );
  XNOR U4532 ( .A(n4453), .B(n4449), .Z(n4452) );
  XOR U4533 ( .A(n4454), .B(n4437), .Z(n4445) );
  AND U4534 ( .A(n4362), .B(n753), .Z(n4437) );
  IV U4535 ( .A(n814), .Z(n753) );
  IV U4536 ( .A(n4438), .Z(n4454) );
  XNOR U4537 ( .A(n4442), .B(n4444), .Z(n3973) );
  NAND U4538 ( .A(n2950), .B(n944), .Z(n4444) );
  XNOR U4539 ( .A(n4440), .B(n4456), .Z(n4442) );
  ANDN U4540 ( .A(n2955), .B(n946), .Z(n4456) );
  XOR U4541 ( .A(n4457), .B(n4458), .Z(n4440) );
  AND U4542 ( .A(n4459), .B(n4460), .Z(n4458) );
  XOR U4543 ( .A(n4461), .B(n4457), .Z(n4460) );
  XNOR U4544 ( .A(n4462), .B(n4451), .Z(n3974) );
  XNOR U4545 ( .A(n4449), .B(n4463), .Z(n4451) );
  ANDN U4546 ( .A(e_input[0]), .B(n814), .Z(n4463) );
  ANDN U4547 ( .A(n4464), .B(n4465), .Z(n4447) );
  XOR U4548 ( .A(n4466), .B(n4467), .Z(n4449) );
  AND U4549 ( .A(n4468), .B(n4469), .Z(n4467) );
  XNOR U4550 ( .A(n4470), .B(n4466), .Z(n4469) );
  XOR U4551 ( .A(n4471), .B(n4453), .Z(n4462) );
  AND U4552 ( .A(n4362), .B(n812), .Z(n4453) );
  IV U4553 ( .A(n878), .Z(n812) );
  IV U4554 ( .A(n4455), .Z(n4471) );
  XNOR U4555 ( .A(n4459), .B(n4461), .Z(n3994) );
  NAND U4556 ( .A(n2950), .B(n1011), .Z(n4461) );
  XNOR U4557 ( .A(n4457), .B(n4473), .Z(n4459) );
  ANDN U4558 ( .A(n2955), .B(n1013), .Z(n4473) );
  XOR U4559 ( .A(n4474), .B(n4475), .Z(n4457) );
  AND U4560 ( .A(n4476), .B(n4477), .Z(n4475) );
  XOR U4561 ( .A(n4478), .B(n4474), .Z(n4477) );
  XNOR U4562 ( .A(n4479), .B(n4468), .Z(n3995) );
  XNOR U4563 ( .A(n4466), .B(n4480), .Z(n4468) );
  ANDN U4564 ( .A(e_input[0]), .B(n878), .Z(n4480) );
  XNOR U4565 ( .A(n4464), .B(g_input[24]), .Z(n4465) );
  ANDN U4566 ( .A(n4481), .B(n4482), .Z(n4464) );
  XOR U4567 ( .A(n4483), .B(n4484), .Z(n4466) );
  AND U4568 ( .A(n4485), .B(n4486), .Z(n4484) );
  XNOR U4569 ( .A(n4487), .B(n4483), .Z(n4486) );
  XOR U4570 ( .A(n4488), .B(n4470), .Z(n4479) );
  AND U4571 ( .A(n4362), .B(n876), .Z(n4470) );
  IV U4572 ( .A(n946), .Z(n876) );
  IV U4573 ( .A(n4472), .Z(n4488) );
  XNOR U4574 ( .A(n4476), .B(n4478), .Z(n4015) );
  NAND U4575 ( .A(n2950), .B(n1085), .Z(n4478) );
  XNOR U4576 ( .A(n4474), .B(n4490), .Z(n4476) );
  ANDN U4577 ( .A(n2955), .B(n1087), .Z(n4490) );
  XOR U4578 ( .A(n4491), .B(n4492), .Z(n4474) );
  AND U4579 ( .A(n4493), .B(n4494), .Z(n4492) );
  XOR U4580 ( .A(n4495), .B(n4491), .Z(n4494) );
  XNOR U4581 ( .A(n4496), .B(n4485), .Z(n4016) );
  XNOR U4582 ( .A(n4483), .B(n4497), .Z(n4485) );
  ANDN U4583 ( .A(e_input[0]), .B(n946), .Z(n4497) );
  ANDN U4584 ( .A(n4498), .B(n4499), .Z(n4481) );
  XOR U4585 ( .A(n4500), .B(n4501), .Z(n4483) );
  AND U4586 ( .A(n4502), .B(n4503), .Z(n4501) );
  XNOR U4587 ( .A(n4504), .B(n4500), .Z(n4503) );
  XOR U4588 ( .A(n4505), .B(n4487), .Z(n4496) );
  AND U4589 ( .A(n4362), .B(n944), .Z(n4487) );
  IV U4590 ( .A(n1013), .Z(n944) );
  IV U4591 ( .A(n4489), .Z(n4505) );
  XNOR U4592 ( .A(n4493), .B(n4495), .Z(n4036) );
  NAND U4593 ( .A(n2950), .B(n1163), .Z(n4495) );
  XNOR U4594 ( .A(n4491), .B(n4507), .Z(n4493) );
  ANDN U4595 ( .A(n2955), .B(n1165), .Z(n4507) );
  XOR U4596 ( .A(n4508), .B(n4509), .Z(n4491) );
  AND U4597 ( .A(n4510), .B(n4511), .Z(n4509) );
  XOR U4598 ( .A(n4512), .B(n4508), .Z(n4511) );
  XNOR U4599 ( .A(n4513), .B(n4502), .Z(n4037) );
  XNOR U4600 ( .A(n4500), .B(n4514), .Z(n4502) );
  ANDN U4601 ( .A(e_input[0]), .B(n1013), .Z(n4514) );
  XNOR U4602 ( .A(n4498), .B(g_input[22]), .Z(n4499) );
  ANDN U4603 ( .A(n4515), .B(n4516), .Z(n4498) );
  XOR U4604 ( .A(n4517), .B(n4518), .Z(n4500) );
  AND U4605 ( .A(n4519), .B(n4520), .Z(n4518) );
  XNOR U4606 ( .A(n4521), .B(n4517), .Z(n4520) );
  XOR U4607 ( .A(n4522), .B(n4504), .Z(n4513) );
  AND U4608 ( .A(n4362), .B(n1011), .Z(n4504) );
  IV U4609 ( .A(n1087), .Z(n1011) );
  IV U4610 ( .A(n4506), .Z(n4522) );
  XNOR U4611 ( .A(n4510), .B(n4512), .Z(n4057) );
  NAND U4612 ( .A(n2950), .B(n1244), .Z(n4512) );
  XNOR U4613 ( .A(n4508), .B(n4524), .Z(n4510) );
  ANDN U4614 ( .A(n2955), .B(n1246), .Z(n4524) );
  XOR U4615 ( .A(n4525), .B(n4526), .Z(n4508) );
  AND U4616 ( .A(n4527), .B(n4528), .Z(n4526) );
  XOR U4617 ( .A(n4529), .B(n4525), .Z(n4528) );
  XNOR U4618 ( .A(n4530), .B(n4519), .Z(n4058) );
  XNOR U4619 ( .A(n4517), .B(n4531), .Z(n4519) );
  ANDN U4620 ( .A(e_input[0]), .B(n1087), .Z(n4531) );
  ANDN U4621 ( .A(n4532), .B(n4533), .Z(n4515) );
  XOR U4622 ( .A(n4534), .B(n4535), .Z(n4517) );
  AND U4623 ( .A(n4536), .B(n4537), .Z(n4535) );
  XNOR U4624 ( .A(n4538), .B(n4534), .Z(n4537) );
  XOR U4625 ( .A(n4539), .B(n4521), .Z(n4530) );
  AND U4626 ( .A(n4362), .B(n1085), .Z(n4521) );
  IV U4627 ( .A(n1165), .Z(n1085) );
  IV U4628 ( .A(n4523), .Z(n4539) );
  XNOR U4629 ( .A(n4527), .B(n4529), .Z(n4078) );
  NAND U4630 ( .A(n2950), .B(n1328), .Z(n4529) );
  XNOR U4631 ( .A(n4525), .B(n4541), .Z(n4527) );
  ANDN U4632 ( .A(n2955), .B(n1330), .Z(n4541) );
  XOR U4633 ( .A(n4542), .B(n4543), .Z(n4525) );
  AND U4634 ( .A(n4544), .B(n4545), .Z(n4543) );
  XOR U4635 ( .A(n4546), .B(n4542), .Z(n4545) );
  XNOR U4636 ( .A(n4547), .B(n4536), .Z(n4079) );
  XNOR U4637 ( .A(n4534), .B(n4548), .Z(n4536) );
  ANDN U4638 ( .A(e_input[0]), .B(n1165), .Z(n4548) );
  XNOR U4639 ( .A(n4532), .B(g_input[20]), .Z(n4533) );
  ANDN U4640 ( .A(n4549), .B(n4550), .Z(n4532) );
  XOR U4641 ( .A(n4551), .B(n4552), .Z(n4534) );
  AND U4642 ( .A(n4553), .B(n4554), .Z(n4552) );
  XNOR U4643 ( .A(n4555), .B(n4551), .Z(n4554) );
  XOR U4644 ( .A(n4556), .B(n4538), .Z(n4547) );
  AND U4645 ( .A(n4362), .B(n1163), .Z(n4538) );
  IV U4646 ( .A(n1246), .Z(n1163) );
  IV U4647 ( .A(n4540), .Z(n4556) );
  XNOR U4648 ( .A(n4544), .B(n4546), .Z(n4099) );
  NAND U4649 ( .A(n2950), .B(n1419), .Z(n4546) );
  XNOR U4650 ( .A(n4542), .B(n4558), .Z(n4544) );
  ANDN U4651 ( .A(n2955), .B(n1421), .Z(n4558) );
  XOR U4652 ( .A(n4559), .B(n4560), .Z(n4542) );
  AND U4653 ( .A(n4561), .B(n4562), .Z(n4560) );
  XOR U4654 ( .A(n4563), .B(n4559), .Z(n4562) );
  XNOR U4655 ( .A(n4564), .B(n4553), .Z(n4100) );
  XNOR U4656 ( .A(n4551), .B(n4565), .Z(n4553) );
  ANDN U4657 ( .A(e_input[0]), .B(n1246), .Z(n4565) );
  ANDN U4658 ( .A(n4566), .B(n4567), .Z(n4549) );
  XOR U4659 ( .A(n4568), .B(n4569), .Z(n4551) );
  AND U4660 ( .A(n4570), .B(n4571), .Z(n4569) );
  XNOR U4661 ( .A(n4572), .B(n4568), .Z(n4571) );
  XOR U4662 ( .A(n4573), .B(n4555), .Z(n4564) );
  AND U4663 ( .A(n4362), .B(n1244), .Z(n4555) );
  IV U4664 ( .A(n1330), .Z(n1244) );
  IV U4665 ( .A(n4557), .Z(n4573) );
  XNOR U4666 ( .A(n4561), .B(n4563), .Z(n4120) );
  NAND U4667 ( .A(n2950), .B(n1516), .Z(n4563) );
  XNOR U4668 ( .A(n4559), .B(n4575), .Z(n4561) );
  ANDN U4669 ( .A(n2955), .B(n1518), .Z(n4575) );
  XOR U4670 ( .A(n4576), .B(n4577), .Z(n4559) );
  AND U4671 ( .A(n4578), .B(n4579), .Z(n4577) );
  XOR U4672 ( .A(n4580), .B(n4576), .Z(n4579) );
  XNOR U4673 ( .A(n4581), .B(n4570), .Z(n4121) );
  XNOR U4674 ( .A(n4568), .B(n4582), .Z(n4570) );
  ANDN U4675 ( .A(e_input[0]), .B(n1330), .Z(n4582) );
  XNOR U4676 ( .A(n4566), .B(g_input[18]), .Z(n4567) );
  ANDN U4677 ( .A(n4583), .B(n4584), .Z(n4566) );
  XOR U4678 ( .A(n4585), .B(n4586), .Z(n4568) );
  AND U4679 ( .A(n4587), .B(n4588), .Z(n4586) );
  XNOR U4680 ( .A(n4589), .B(n4585), .Z(n4588) );
  XOR U4681 ( .A(n4590), .B(n4572), .Z(n4581) );
  AND U4682 ( .A(n4362), .B(n1328), .Z(n4572) );
  IV U4683 ( .A(n1421), .Z(n1328) );
  IV U4684 ( .A(n4574), .Z(n4590) );
  XNOR U4685 ( .A(n4578), .B(n4580), .Z(n4141) );
  NAND U4686 ( .A(n2950), .B(n1612), .Z(n4580) );
  XNOR U4687 ( .A(n4576), .B(n4592), .Z(n4578) );
  ANDN U4688 ( .A(n2955), .B(n1614), .Z(n4592) );
  XOR U4689 ( .A(n4593), .B(n4594), .Z(n4576) );
  AND U4690 ( .A(n4595), .B(n4596), .Z(n4594) );
  XOR U4691 ( .A(n4597), .B(n4593), .Z(n4596) );
  XNOR U4692 ( .A(n4598), .B(n4587), .Z(n4142) );
  XNOR U4693 ( .A(n4585), .B(n4599), .Z(n4587) );
  ANDN U4694 ( .A(e_input[0]), .B(n1421), .Z(n4599) );
  ANDN U4695 ( .A(n4600), .B(n4601), .Z(n4583) );
  XOR U4696 ( .A(n4602), .B(n4603), .Z(n4585) );
  AND U4697 ( .A(n4604), .B(n4605), .Z(n4603) );
  XNOR U4698 ( .A(n4606), .B(n4602), .Z(n4605) );
  XOR U4699 ( .A(n4607), .B(n4589), .Z(n4598) );
  AND U4700 ( .A(n4362), .B(n1419), .Z(n4589) );
  IV U4701 ( .A(n1518), .Z(n1419) );
  IV U4702 ( .A(n4591), .Z(n4607) );
  XNOR U4703 ( .A(n4595), .B(n4597), .Z(n4162) );
  NAND U4704 ( .A(n2950), .B(n1708), .Z(n4597) );
  XNOR U4705 ( .A(n4593), .B(n4609), .Z(n4595) );
  ANDN U4706 ( .A(n2955), .B(n1710), .Z(n4609) );
  XNOR U4707 ( .A(n4613), .B(n4604), .Z(n4163) );
  XNOR U4708 ( .A(n4602), .B(n4614), .Z(n4604) );
  ANDN U4709 ( .A(e_input[0]), .B(n1518), .Z(n4614) );
  AND U4710 ( .A(n4362), .B(n1516), .Z(n4606) );
  XNOR U4711 ( .A(n4611), .B(n4612), .Z(n4180) );
  NAND U4712 ( .A(n2950), .B(n1809), .Z(n4612) );
  XNOR U4713 ( .A(n4610), .B(n4619), .Z(n4611) );
  ANDN U4714 ( .A(n2955), .B(n1811), .Z(n4619) );
  XNOR U4715 ( .A(n4623), .B(n4616), .Z(n4182) );
  XNOR U4716 ( .A(n4615), .B(n4624), .Z(n4616) );
  ANDN U4717 ( .A(e_input[0]), .B(n1614), .Z(n4624) );
  AND U4718 ( .A(n4362), .B(n1612), .Z(n4617) );
  XNOR U4719 ( .A(n4621), .B(n4622), .Z(n4200) );
  NAND U4720 ( .A(n2950), .B(n1915), .Z(n4622) );
  XNOR U4721 ( .A(n4620), .B(n4629), .Z(n4621) );
  ANDN U4722 ( .A(n2955), .B(n1917), .Z(n4629) );
  XNOR U4723 ( .A(n4633), .B(n4626), .Z(n4202) );
  XNOR U4724 ( .A(n4625), .B(n4634), .Z(n4626) );
  ANDN U4725 ( .A(e_input[0]), .B(n1710), .Z(n4634) );
  AND U4726 ( .A(n4362), .B(n1708), .Z(n4627) );
  XNOR U4727 ( .A(n4631), .B(n4632), .Z(n4220) );
  NAND U4728 ( .A(n2950), .B(n2022), .Z(n4632) );
  XNOR U4729 ( .A(n4630), .B(n4639), .Z(n4631) );
  ANDN U4730 ( .A(n2955), .B(n2024), .Z(n4639) );
  XNOR U4731 ( .A(n4643), .B(n4636), .Z(n4222) );
  XNOR U4732 ( .A(n4635), .B(n4644), .Z(n4636) );
  ANDN U4733 ( .A(e_input[0]), .B(n1811), .Z(n4644) );
  XOR U4734 ( .A(n4645), .B(n4646), .Z(n4635) );
  AND U4735 ( .A(n4647), .B(n4648), .Z(n4646) );
  XNOR U4736 ( .A(n4649), .B(n4645), .Z(n4648) );
  AND U4737 ( .A(n4362), .B(n1809), .Z(n4637) );
  XNOR U4738 ( .A(n4641), .B(n4642), .Z(n4240) );
  NAND U4739 ( .A(n2950), .B(n2130), .Z(n4642) );
  XNOR U4740 ( .A(n4640), .B(n4651), .Z(n4641) );
  ANDN U4741 ( .A(n2955), .B(n2132), .Z(n4651) );
  XOR U4742 ( .A(n4652), .B(n4653), .Z(n4640) );
  AND U4743 ( .A(n4654), .B(n4655), .Z(n4653) );
  XOR U4744 ( .A(n4656), .B(n4652), .Z(n4655) );
  XNOR U4745 ( .A(n4657), .B(n4647), .Z(n4242) );
  XNOR U4746 ( .A(n4645), .B(n4658), .Z(n4647) );
  ANDN U4747 ( .A(e_input[0]), .B(n1917), .Z(n4658) );
  XOR U4748 ( .A(n4659), .B(n4660), .Z(n4645) );
  AND U4749 ( .A(n4661), .B(n4662), .Z(n4660) );
  XNOR U4750 ( .A(n4663), .B(n4659), .Z(n4662) );
  XOR U4751 ( .A(n4664), .B(n4649), .Z(n4657) );
  AND U4752 ( .A(n4362), .B(n1915), .Z(n4649) );
  IV U4753 ( .A(n4650), .Z(n4664) );
  XNOR U4754 ( .A(n4654), .B(n4656), .Z(n4260) );
  NAND U4755 ( .A(n2950), .B(n2249), .Z(n4656) );
  XNOR U4756 ( .A(n4652), .B(n4666), .Z(n4654) );
  ANDN U4757 ( .A(n2955), .B(n2251), .Z(n4666) );
  XOR U4758 ( .A(n4667), .B(n4668), .Z(n4652) );
  AND U4759 ( .A(n4669), .B(n4670), .Z(n4668) );
  XOR U4760 ( .A(n4671), .B(n4667), .Z(n4670) );
  XNOR U4761 ( .A(n4672), .B(n4661), .Z(n4262) );
  XNOR U4762 ( .A(n4659), .B(n4673), .Z(n4661) );
  ANDN U4763 ( .A(e_input[0]), .B(n2024), .Z(n4673) );
  XOR U4764 ( .A(n4674), .B(n4675), .Z(n4659) );
  AND U4765 ( .A(n4676), .B(n4677), .Z(n4675) );
  XNOR U4766 ( .A(n4678), .B(n4674), .Z(n4677) );
  XOR U4767 ( .A(n4679), .B(n4663), .Z(n4672) );
  AND U4768 ( .A(n4362), .B(n2022), .Z(n4663) );
  IV U4769 ( .A(n4665), .Z(n4679) );
  XNOR U4770 ( .A(n4669), .B(n4671), .Z(n4280) );
  NAND U4771 ( .A(n2950), .B(n2369), .Z(n4671) );
  XNOR U4772 ( .A(n4667), .B(n4681), .Z(n4669) );
  ANDN U4773 ( .A(n2955), .B(n2371), .Z(n4681) );
  XNOR U4774 ( .A(n4685), .B(n4676), .Z(n4282) );
  XNOR U4775 ( .A(n4674), .B(n4686), .Z(n4676) );
  ANDN U4776 ( .A(e_input[0]), .B(n2132), .Z(n4686) );
  XOR U4777 ( .A(n4687), .B(n4688), .Z(n4674) );
  AND U4778 ( .A(n4689), .B(n4690), .Z(n4688) );
  XNOR U4779 ( .A(n4691), .B(n4687), .Z(n4690) );
  AND U4780 ( .A(n4362), .B(n2130), .Z(n4678) );
  XNOR U4781 ( .A(n4683), .B(n4684), .Z(n4304) );
  NAND U4782 ( .A(n2950), .B(n2491), .Z(n4684) );
  XNOR U4783 ( .A(n4682), .B(n4693), .Z(n4683) );
  ANDN U4784 ( .A(n2955), .B(n2493), .Z(n4693) );
  XNOR U4785 ( .A(n4697), .B(n4689), .Z(n4306) );
  XNOR U4786 ( .A(n4687), .B(n4698), .Z(n4689) );
  ANDN U4787 ( .A(e_input[0]), .B(n2251), .Z(n4698) );
  XOR U4788 ( .A(n4699), .B(n4700), .Z(n4687) );
  AND U4789 ( .A(n4701), .B(n4702), .Z(n4700) );
  XNOR U4790 ( .A(n4703), .B(n4699), .Z(n4702) );
  AND U4791 ( .A(n4362), .B(n2249), .Z(n4691) );
  XNOR U4792 ( .A(n4695), .B(n4696), .Z(n4324) );
  NAND U4793 ( .A(n2950), .B(n2616), .Z(n4696) );
  XNOR U4794 ( .A(n4694), .B(n4705), .Z(n4695) );
  ANDN U4795 ( .A(n2955), .B(n2618), .Z(n4705) );
  XNOR U4796 ( .A(n4709), .B(n4701), .Z(n4325) );
  XNOR U4797 ( .A(n4699), .B(n4710), .Z(n4701) );
  ANDN U4798 ( .A(e_input[0]), .B(n2371), .Z(n4710) );
  AND U4799 ( .A(n4362), .B(n2369), .Z(n4703) );
  XNOR U4800 ( .A(n4714), .B(n4715), .Z(n4704) );
  AND U4801 ( .A(n4716), .B(n4717), .Z(n4715) );
  XNOR U4802 ( .A(n4712), .B(n4718), .Z(n4717) );
  XNOR U4803 ( .A(n4713), .B(n4714), .Z(n4718) );
  AND U4804 ( .A(n4362), .B(n2491), .Z(n4713) );
  XOR U4805 ( .A(n4711), .B(n4719), .Z(n4712) );
  ANDN U4806 ( .A(e_input[0]), .B(n2493), .Z(n4719) );
  XNOR U4807 ( .A(n4707), .B(n4723), .Z(n4716) );
  XNOR U4808 ( .A(n4708), .B(n4714), .Z(n4723) );
  AND U4809 ( .A(n2748), .B(n2950), .Z(n4708) );
  XOR U4810 ( .A(n4706), .B(n4724), .Z(n4707) );
  ANDN U4811 ( .A(n2955), .B(n2750), .Z(n4724) );
  XOR U4812 ( .A(n4728), .B(n4729), .Z(n4714) );
  AND U4813 ( .A(n4730), .B(n4731), .Z(n4729) );
  XNOR U4814 ( .A(n4721), .B(n4732), .Z(n4731) );
  XNOR U4815 ( .A(n4722), .B(n4728), .Z(n4732) );
  AND U4816 ( .A(n4362), .B(n2616), .Z(n4722) );
  XOR U4817 ( .A(n4720), .B(n4733), .Z(n4721) );
  ANDN U4818 ( .A(e_input[0]), .B(n2618), .Z(n4733) );
  XNOR U4819 ( .A(n4726), .B(n4737), .Z(n4730) );
  XNOR U4820 ( .A(n4727), .B(n4728), .Z(n4737) );
  AND U4821 ( .A(n2880), .B(n2950), .Z(n4727) );
  XOR U4822 ( .A(n4725), .B(n4738), .Z(n4726) );
  ANDN U4823 ( .A(n2955), .B(n2882), .Z(n4738) );
  XOR U4824 ( .A(n4739), .B(n4740), .Z(n4725) );
  ANDN U4825 ( .A(n4741), .B(n4742), .Z(n4740) );
  XNOR U4826 ( .A(n4743), .B(n4739), .Z(n4741) );
  XOR U4827 ( .A(n4744), .B(n4745), .Z(n4728) );
  AND U4828 ( .A(n4746), .B(n4747), .Z(n4745) );
  XNOR U4829 ( .A(n4735), .B(n4748), .Z(n4747) );
  XNOR U4830 ( .A(n4736), .B(n4744), .Z(n4748) );
  AND U4831 ( .A(n4362), .B(n2748), .Z(n4736) );
  XOR U4832 ( .A(n4734), .B(n4749), .Z(n4735) );
  ANDN U4833 ( .A(e_input[0]), .B(n2750), .Z(n4749) );
  XNOR U4834 ( .A(n4742), .B(n4753), .Z(n4746) );
  XNOR U4835 ( .A(n4743), .B(n4744), .Z(n4753) );
  AND U4836 ( .A(n3019), .B(n2950), .Z(n4743) );
  XOR U4837 ( .A(n4739), .B(n4754), .Z(n4742) );
  ANDN U4838 ( .A(n2955), .B(n3021), .Z(n4754) );
  XNOR U4839 ( .A(n4759), .B(n4751), .Z(n4345) );
  XNOR U4840 ( .A(n4750), .B(n4760), .Z(n4751) );
  ANDN U4841 ( .A(e_input[0]), .B(n2882), .Z(n4760) );
  XNOR U4842 ( .A(n4763), .B(n4761), .Z(n4762) );
  ANDN U4843 ( .A(e_input[0]), .B(n3021), .Z(n4763) );
  ANDN U4844 ( .A(n4362), .B(n3809), .Z(n4764) );
  XNOR U4845 ( .A(n4758), .B(n4752), .Z(n4759) );
  AND U4846 ( .A(n4362), .B(n2880), .Z(n4752) );
  XNOR U4847 ( .A(n4756), .B(n4757), .Z(n4344) );
  NAND U4848 ( .A(n3807), .B(n2950), .Z(n4757) );
  XNOR U4849 ( .A(n4755), .B(n4768), .Z(n4756) );
  ANDN U4850 ( .A(n2955), .B(n3809), .Z(n4768) );
  NAND U4851 ( .A(g_input[0]), .B(n4769), .Z(n4755) );
  NANDN U4852 ( .B(n2950), .A(n4770), .Z(n4769) );
  NANDN U4853 ( .B(n3812), .A(n2955), .Z(n4770) );
  IV U4854 ( .A(n2818), .Z(n2950) );
  XNOR U4855 ( .A(n4766), .B(n4767), .Z(n4758) );
  NAND U4856 ( .A(n3807), .B(n4362), .Z(n4767) );
  XNOR U4857 ( .A(n4765), .B(n4773), .Z(n4766) );
  ANDN U4858 ( .A(e_input[0]), .B(n3809), .Z(n4773) );
  NAND U4859 ( .A(g_input[0]), .B(n4774), .Z(n4765) );
  NANDN U4860 ( .B(n4362), .A(n4775), .Z(n4774) );
  NANDN U4861 ( .B(n3812), .A(e_input[0]), .Z(n4775) );
  IV U4862 ( .A(n4349), .Z(n4362) );
  XNOR U4863 ( .A(n2978), .B(n2977), .Z(n2931) );
  XOR U4864 ( .A(n4777), .B(n2986), .Z(n2977) );
  XNOR U4865 ( .A(n2971), .B(n2970), .Z(n2986) );
  XOR U4866 ( .A(n4778), .B(n2967), .Z(n2970) );
  XNOR U4867 ( .A(n2966), .B(n4779), .Z(n2967) );
  ANDN U4868 ( .A(n1032), .B(n1917), .Z(n4779) );
  AND U4869 ( .A(n1915), .B(n969), .Z(n2968) );
  XNOR U4870 ( .A(n2974), .B(n2975), .Z(n2971) );
  NANDN U4871 ( .B(n834), .A(n2130), .Z(n2975) );
  XNOR U4872 ( .A(n2973), .B(n4786), .Z(n2974) );
  ANDN U4873 ( .A(n904), .B(n2132), .Z(n4786) );
  XOR U4874 ( .A(n2985), .B(n2976), .Z(n4777) );
  XNOR U4875 ( .A(n4790), .B(n4791), .Z(n2976) );
  XOR U4876 ( .A(n4792), .B(n2994), .Z(n2985) );
  XNOR U4877 ( .A(n2982), .B(n2983), .Z(n2994) );
  NAND U4878 ( .A(n1708), .B(n1203), .Z(n2983) );
  XNOR U4879 ( .A(n2981), .B(n4793), .Z(n2982) );
  ANDN U4880 ( .A(n1210), .B(n1710), .Z(n4793) );
  XNOR U4881 ( .A(n2993), .B(n2984), .Z(n4792) );
  XOR U4882 ( .A(n4797), .B(n4798), .Z(n2984) );
  AND U4883 ( .A(n4799), .B(n4800), .Z(n4798) );
  XOR U4884 ( .A(n4801), .B(n4802), .Z(n4800) );
  XNOR U4885 ( .A(n4797), .B(n4803), .Z(n4802) );
  XNOR U4886 ( .A(n4784), .B(n4804), .Z(n4799) );
  XNOR U4887 ( .A(n4797), .B(n4785), .Z(n4804) );
  XNOR U4888 ( .A(n4788), .B(n4789), .Z(n4785) );
  NANDN U4889 ( .B(n834), .A(n2249), .Z(n4789) );
  XNOR U4890 ( .A(n4787), .B(n4805), .Z(n4788) );
  ANDN U4891 ( .A(n904), .B(n2251), .Z(n4805) );
  XOR U4892 ( .A(n4809), .B(n4781), .Z(n4784) );
  XNOR U4893 ( .A(n4780), .B(n4810), .Z(n4781) );
  ANDN U4894 ( .A(n1032), .B(n2024), .Z(n4810) );
  AND U4895 ( .A(n2022), .B(n969), .Z(n4782) );
  XOR U4896 ( .A(n4817), .B(n4818), .Z(n4797) );
  AND U4897 ( .A(n4819), .B(n4820), .Z(n4818) );
  XOR U4898 ( .A(n4821), .B(n4822), .Z(n4820) );
  XNOR U4899 ( .A(n4817), .B(n4823), .Z(n4822) );
  XNOR U4900 ( .A(n4815), .B(n4824), .Z(n4819) );
  XNOR U4901 ( .A(n4817), .B(n4816), .Z(n4824) );
  XNOR U4902 ( .A(n4807), .B(n4808), .Z(n4816) );
  NANDN U4903 ( .B(n834), .A(n2369), .Z(n4808) );
  XNOR U4904 ( .A(n4806), .B(n4825), .Z(n4807) );
  ANDN U4905 ( .A(n904), .B(n2371), .Z(n4825) );
  XOR U4906 ( .A(n4829), .B(n4812), .Z(n4815) );
  XNOR U4907 ( .A(n4811), .B(n4830), .Z(n4812) );
  ANDN U4908 ( .A(n1032), .B(n2132), .Z(n4830) );
  AND U4909 ( .A(n2130), .B(n969), .Z(n4813) );
  XOR U4910 ( .A(n4837), .B(n4838), .Z(n4817) );
  AND U4911 ( .A(n4839), .B(n4840), .Z(n4838) );
  XOR U4912 ( .A(n4841), .B(n4842), .Z(n4840) );
  XNOR U4913 ( .A(n4837), .B(n4843), .Z(n4842) );
  XNOR U4914 ( .A(n4835), .B(n4844), .Z(n4839) );
  XNOR U4915 ( .A(n4837), .B(n4836), .Z(n4844) );
  XNOR U4916 ( .A(n4827), .B(n4828), .Z(n4836) );
  NANDN U4917 ( .B(n834), .A(n2491), .Z(n4828) );
  XNOR U4918 ( .A(n4826), .B(n4845), .Z(n4827) );
  ANDN U4919 ( .A(n904), .B(n2493), .Z(n4845) );
  XOR U4920 ( .A(n4849), .B(n4832), .Z(n4835) );
  XNOR U4921 ( .A(n4831), .B(n4850), .Z(n4832) );
  ANDN U4922 ( .A(n1032), .B(n2251), .Z(n4850) );
  AND U4923 ( .A(n2249), .B(n969), .Z(n4833) );
  XOR U4924 ( .A(n4857), .B(n4858), .Z(n4837) );
  AND U4925 ( .A(n4859), .B(n4860), .Z(n4858) );
  XOR U4926 ( .A(n4861), .B(n4862), .Z(n4860) );
  XNOR U4927 ( .A(n4857), .B(n4863), .Z(n4862) );
  XNOR U4928 ( .A(n4855), .B(n4864), .Z(n4859) );
  XNOR U4929 ( .A(n4857), .B(n4856), .Z(n4864) );
  XNOR U4930 ( .A(n4847), .B(n4848), .Z(n4856) );
  NANDN U4931 ( .B(n834), .A(n2616), .Z(n4848) );
  XNOR U4932 ( .A(n4846), .B(n4865), .Z(n4847) );
  ANDN U4933 ( .A(n904), .B(n2618), .Z(n4865) );
  XOR U4934 ( .A(n4869), .B(n4852), .Z(n4855) );
  XNOR U4935 ( .A(n4851), .B(n4870), .Z(n4852) );
  ANDN U4936 ( .A(n1032), .B(n2371), .Z(n4870) );
  AND U4937 ( .A(n2369), .B(n969), .Z(n4853) );
  XOR U4938 ( .A(n4877), .B(n4878), .Z(n4857) );
  AND U4939 ( .A(n4879), .B(n4880), .Z(n4878) );
  XOR U4940 ( .A(n4881), .B(n4882), .Z(n4880) );
  XNOR U4941 ( .A(n4877), .B(n4883), .Z(n4882) );
  XNOR U4942 ( .A(n4875), .B(n4884), .Z(n4879) );
  XNOR U4943 ( .A(n4877), .B(n4876), .Z(n4884) );
  XNOR U4944 ( .A(n4867), .B(n4868), .Z(n4876) );
  NANDN U4945 ( .B(n834), .A(n2748), .Z(n4868) );
  XNOR U4946 ( .A(n4866), .B(n4885), .Z(n4867) );
  ANDN U4947 ( .A(n904), .B(n2750), .Z(n4885) );
  XOR U4948 ( .A(n4889), .B(n4872), .Z(n4875) );
  XNOR U4949 ( .A(n4871), .B(n4890), .Z(n4872) );
  ANDN U4950 ( .A(n1032), .B(n2493), .Z(n4890) );
  XOR U4951 ( .A(n4891), .B(n4892), .Z(n4871) );
  AND U4952 ( .A(n4893), .B(n4894), .Z(n4892) );
  XNOR U4953 ( .A(n4895), .B(n4891), .Z(n4894) );
  AND U4954 ( .A(n2491), .B(n969), .Z(n4873) );
  XOR U4955 ( .A(n4899), .B(n4900), .Z(n4877) );
  AND U4956 ( .A(n4901), .B(n4902), .Z(n4900) );
  XOR U4957 ( .A(n4903), .B(n4904), .Z(n4902) );
  XNOR U4958 ( .A(n4899), .B(n4905), .Z(n4904) );
  XNOR U4959 ( .A(n4897), .B(n4906), .Z(n4901) );
  XNOR U4960 ( .A(n4899), .B(n4898), .Z(n4906) );
  XNOR U4961 ( .A(n4887), .B(n4888), .Z(n4898) );
  NANDN U4962 ( .B(n834), .A(n2880), .Z(n4888) );
  XNOR U4963 ( .A(n4886), .B(n4907), .Z(n4887) );
  ANDN U4964 ( .A(n904), .B(n2882), .Z(n4907) );
  XOR U4965 ( .A(n4908), .B(n4909), .Z(n4886) );
  AND U4966 ( .A(n4910), .B(n4911), .Z(n4909) );
  XOR U4967 ( .A(n4912), .B(n4908), .Z(n4911) );
  XOR U4968 ( .A(n4913), .B(n4893), .Z(n4897) );
  XNOR U4969 ( .A(n4891), .B(n4914), .Z(n4893) );
  ANDN U4970 ( .A(n1032), .B(n2618), .Z(n4914) );
  XOR U4971 ( .A(n4915), .B(n4916), .Z(n4891) );
  AND U4972 ( .A(n4917), .B(n4918), .Z(n4916) );
  XNOR U4973 ( .A(n4919), .B(n4915), .Z(n4918) );
  AND U4974 ( .A(n2616), .B(n969), .Z(n4895) );
  XOR U4975 ( .A(n4923), .B(n4924), .Z(n4899) );
  AND U4976 ( .A(n4925), .B(n4926), .Z(n4924) );
  XOR U4977 ( .A(n4927), .B(n4928), .Z(n4926) );
  XNOR U4978 ( .A(n4923), .B(n4929), .Z(n4928) );
  XNOR U4979 ( .A(n4921), .B(n4930), .Z(n4925) );
  XNOR U4980 ( .A(n4923), .B(n4922), .Z(n4930) );
  XNOR U4981 ( .A(n4910), .B(n4912), .Z(n4922) );
  NANDN U4982 ( .B(n834), .A(n3019), .Z(n4912) );
  XNOR U4983 ( .A(n4908), .B(n4931), .Z(n4910) );
  ANDN U4984 ( .A(n904), .B(n3021), .Z(n4931) );
  XOR U4985 ( .A(n4935), .B(n4917), .Z(n4921) );
  XNOR U4986 ( .A(n4915), .B(n4936), .Z(n4917) );
  ANDN U4987 ( .A(n1032), .B(n2750), .Z(n4936) );
  AND U4988 ( .A(n2748), .B(n969), .Z(n4919) );
  XOR U4989 ( .A(n4944), .B(n4945), .Z(n4791) );
  XNOR U4990 ( .A(n4942), .B(n4941), .Z(n4790) );
  XOR U4991 ( .A(n4947), .B(n4938), .Z(n4941) );
  XNOR U4992 ( .A(n4937), .B(n4948), .Z(n4938) );
  ANDN U4993 ( .A(n1032), .B(n2882), .Z(n4948) );
  XNOR U4994 ( .A(n4951), .B(n4949), .Z(n4950) );
  ANDN U4995 ( .A(n1032), .B(n3021), .Z(n4951) );
  XNOR U4996 ( .A(n4940), .B(n4939), .Z(n4947) );
  AND U4997 ( .A(n2880), .B(n969), .Z(n4939) );
  XNOR U4998 ( .A(n4954), .B(n4955), .Z(n4940) );
  NAND U4999 ( .A(n3807), .B(n969), .Z(n4955) );
  XNOR U5000 ( .A(n4953), .B(n4956), .Z(n4954) );
  ANDN U5001 ( .A(n1032), .B(n3809), .Z(n4956) );
  NAND U5002 ( .A(g_input[0]), .B(n4957), .Z(n4953) );
  NANDN U5003 ( .B(n969), .A(n4958), .Z(n4957) );
  NANDN U5004 ( .B(n3812), .A(n1032), .Z(n4958) );
  IV U5005 ( .A(n4952), .Z(n969) );
  XNOR U5006 ( .A(n4933), .B(n4934), .Z(n4942) );
  NANDN U5007 ( .B(n834), .A(n3807), .Z(n4934) );
  XNOR U5008 ( .A(n4932), .B(n4961), .Z(n4933) );
  ANDN U5009 ( .A(n904), .B(n3809), .Z(n4961) );
  NAND U5010 ( .A(g_input[0]), .B(n4962), .Z(n4932) );
  NAND U5011 ( .A(n4963), .B(n834), .Z(n4962) );
  NANDN U5012 ( .B(n3812), .A(n904), .Z(n4963) );
  XOR U5013 ( .A(n4966), .B(n4967), .Z(n4943) );
  XOR U5014 ( .A(n4968), .B(n2990), .Z(n2993) );
  XNOR U5015 ( .A(n2989), .B(n4969), .Z(n2990) );
  ANDN U5016 ( .A(n1394), .B(n1518), .Z(n4969) );
  XNOR U5017 ( .A(n4600), .B(g_input[16]), .Z(n4601) );
  ANDN U5018 ( .A(n4970), .B(n4971), .Z(n4600) );
  AND U5019 ( .A(n1516), .B(n1387), .Z(n2991) );
  IV U5020 ( .A(n1614), .Z(n1516) );
  XNOR U5021 ( .A(n4795), .B(n4796), .Z(n4801) );
  NAND U5022 ( .A(n1809), .B(n1203), .Z(n4796) );
  XNOR U5023 ( .A(n4794), .B(n4976), .Z(n4795) );
  ANDN U5024 ( .A(n1210), .B(n1811), .Z(n4976) );
  XNOR U5025 ( .A(n4980), .B(n4973), .Z(n4803) );
  XNOR U5026 ( .A(n4972), .B(n4981), .Z(n4973) );
  ANDN U5027 ( .A(n1394), .B(n1614), .Z(n4981) );
  ANDN U5028 ( .A(n4982), .B(n4983), .Z(n4970) );
  AND U5029 ( .A(n1612), .B(n1387), .Z(n4974) );
  IV U5030 ( .A(n1710), .Z(n1612) );
  XNOR U5031 ( .A(n4978), .B(n4979), .Z(n4821) );
  NAND U5032 ( .A(n1915), .B(n1203), .Z(n4979) );
  XNOR U5033 ( .A(n4977), .B(n4988), .Z(n4978) );
  ANDN U5034 ( .A(n1210), .B(n1917), .Z(n4988) );
  XNOR U5035 ( .A(n4992), .B(n4985), .Z(n4823) );
  XNOR U5036 ( .A(n4984), .B(n4993), .Z(n4985) );
  ANDN U5037 ( .A(n1394), .B(n1710), .Z(n4993) );
  XNOR U5038 ( .A(n4982), .B(g_input[14]), .Z(n4983) );
  ANDN U5039 ( .A(n4994), .B(n4995), .Z(n4982) );
  AND U5040 ( .A(n1708), .B(n1387), .Z(n4986) );
  IV U5041 ( .A(n1811), .Z(n1708) );
  XNOR U5042 ( .A(n4990), .B(n4991), .Z(n4841) );
  NAND U5043 ( .A(n2022), .B(n1203), .Z(n4991) );
  XNOR U5044 ( .A(n4989), .B(n5000), .Z(n4990) );
  ANDN U5045 ( .A(n1210), .B(n2024), .Z(n5000) );
  XNOR U5046 ( .A(n5004), .B(n4997), .Z(n4843) );
  XNOR U5047 ( .A(n4996), .B(n5005), .Z(n4997) );
  ANDN U5048 ( .A(n1394), .B(n1811), .Z(n5005) );
  ANDN U5049 ( .A(n5006), .B(n5007), .Z(n4994) );
  AND U5050 ( .A(n1809), .B(n1387), .Z(n4998) );
  IV U5051 ( .A(n1917), .Z(n1809) );
  XNOR U5052 ( .A(n5002), .B(n5003), .Z(n4861) );
  NAND U5053 ( .A(n2130), .B(n1203), .Z(n5003) );
  XNOR U5054 ( .A(n5001), .B(n5012), .Z(n5002) );
  ANDN U5055 ( .A(n1210), .B(n2132), .Z(n5012) );
  XNOR U5056 ( .A(n5016), .B(n5009), .Z(n4863) );
  XNOR U5057 ( .A(n5008), .B(n5017), .Z(n5009) );
  ANDN U5058 ( .A(n1394), .B(n1917), .Z(n5017) );
  XNOR U5059 ( .A(n5006), .B(g_input[12]), .Z(n5007) );
  ANDN U5060 ( .A(n5018), .B(n5019), .Z(n5006) );
  AND U5061 ( .A(n1915), .B(n1387), .Z(n5010) );
  IV U5062 ( .A(n2024), .Z(n1915) );
  XNOR U5063 ( .A(n5014), .B(n5015), .Z(n4881) );
  NAND U5064 ( .A(n2249), .B(n1203), .Z(n5015) );
  XNOR U5065 ( .A(n5013), .B(n5024), .Z(n5014) );
  ANDN U5066 ( .A(n1210), .B(n2251), .Z(n5024) );
  XOR U5067 ( .A(n5025), .B(n5026), .Z(n5013) );
  AND U5068 ( .A(n5027), .B(n5028), .Z(n5026) );
  XOR U5069 ( .A(n5029), .B(n5025), .Z(n5028) );
  XNOR U5070 ( .A(n5030), .B(n5021), .Z(n4883) );
  XNOR U5071 ( .A(n5020), .B(n5031), .Z(n5021) );
  ANDN U5072 ( .A(n1394), .B(n2024), .Z(n5031) );
  ANDN U5073 ( .A(n5032), .B(n5033), .Z(n5018) );
  AND U5074 ( .A(n2022), .B(n1387), .Z(n5022) );
  IV U5075 ( .A(n2132), .Z(n2022) );
  XNOR U5076 ( .A(n5027), .B(n5029), .Z(n4903) );
  NAND U5077 ( .A(n2369), .B(n1203), .Z(n5029) );
  XNOR U5078 ( .A(n5025), .B(n5038), .Z(n5027) );
  ANDN U5079 ( .A(n1210), .B(n2371), .Z(n5038) );
  XOR U5080 ( .A(n5039), .B(n5040), .Z(n5025) );
  AND U5081 ( .A(n5041), .B(n5042), .Z(n5040) );
  XOR U5082 ( .A(n5043), .B(n5039), .Z(n5042) );
  XNOR U5083 ( .A(n5044), .B(n5035), .Z(n4905) );
  XNOR U5084 ( .A(n5034), .B(n5045), .Z(n5035) );
  ANDN U5085 ( .A(n1394), .B(n2132), .Z(n5045) );
  XNOR U5086 ( .A(n5032), .B(g_input[10]), .Z(n5033) );
  ANDN U5087 ( .A(n5046), .B(n5047), .Z(n5032) );
  XOR U5088 ( .A(n5048), .B(n5049), .Z(n5034) );
  AND U5089 ( .A(n5050), .B(n5051), .Z(n5049) );
  XNOR U5090 ( .A(n5052), .B(n5048), .Z(n5051) );
  XOR U5091 ( .A(n5053), .B(n5036), .Z(n5044) );
  AND U5092 ( .A(n2130), .B(n1387), .Z(n5036) );
  IV U5093 ( .A(n2251), .Z(n2130) );
  IV U5094 ( .A(n5037), .Z(n5053) );
  XNOR U5095 ( .A(n5041), .B(n5043), .Z(n4927) );
  NAND U5096 ( .A(n2491), .B(n1203), .Z(n5043) );
  XNOR U5097 ( .A(n5039), .B(n5055), .Z(n5041) );
  ANDN U5098 ( .A(n1210), .B(n2493), .Z(n5055) );
  XNOR U5099 ( .A(n5059), .B(n5050), .Z(n4929) );
  XNOR U5100 ( .A(n5048), .B(n5060), .Z(n5050) );
  ANDN U5101 ( .A(n1394), .B(n2251), .Z(n5060) );
  ANDN U5102 ( .A(n5061), .B(n5062), .Z(n5046) );
  XOR U5103 ( .A(n5063), .B(n5064), .Z(n5048) );
  AND U5104 ( .A(n5065), .B(n5066), .Z(n5064) );
  XNOR U5105 ( .A(n5067), .B(n5063), .Z(n5066) );
  AND U5106 ( .A(n2249), .B(n1387), .Z(n5052) );
  IV U5107 ( .A(n2371), .Z(n2249) );
  XNOR U5108 ( .A(n5057), .B(n5058), .Z(n4945) );
  NAND U5109 ( .A(n2616), .B(n1203), .Z(n5058) );
  XNOR U5110 ( .A(n5056), .B(n5069), .Z(n5057) );
  ANDN U5111 ( .A(n1210), .B(n2618), .Z(n5069) );
  XNOR U5112 ( .A(n5073), .B(n5065), .Z(n4946) );
  XNOR U5113 ( .A(n5063), .B(n5074), .Z(n5065) );
  ANDN U5114 ( .A(n1394), .B(n2371), .Z(n5074) );
  AND U5115 ( .A(n2369), .B(n1387), .Z(n5067) );
  XNOR U5116 ( .A(n5078), .B(n5079), .Z(n5068) );
  AND U5117 ( .A(n5080), .B(n5081), .Z(n5079) );
  XNOR U5118 ( .A(n5076), .B(n5082), .Z(n5081) );
  XNOR U5119 ( .A(n5077), .B(n5078), .Z(n5082) );
  AND U5120 ( .A(n2491), .B(n1387), .Z(n5077) );
  XOR U5121 ( .A(n5075), .B(n5083), .Z(n5076) );
  ANDN U5122 ( .A(n1394), .B(n2493), .Z(n5083) );
  XNOR U5123 ( .A(n5071), .B(n5087), .Z(n5080) );
  XNOR U5124 ( .A(n5072), .B(n5078), .Z(n5087) );
  AND U5125 ( .A(n2748), .B(n1203), .Z(n5072) );
  XOR U5126 ( .A(n5070), .B(n5088), .Z(n5071) );
  ANDN U5127 ( .A(n1210), .B(n2750), .Z(n5088) );
  XOR U5128 ( .A(n5092), .B(n5093), .Z(n5078) );
  AND U5129 ( .A(n5094), .B(n5095), .Z(n5093) );
  XNOR U5130 ( .A(n5085), .B(n5096), .Z(n5095) );
  XNOR U5131 ( .A(n5086), .B(n5092), .Z(n5096) );
  AND U5132 ( .A(n2616), .B(n1387), .Z(n5086) );
  XOR U5133 ( .A(n5084), .B(n5097), .Z(n5085) );
  ANDN U5134 ( .A(n1394), .B(n2618), .Z(n5097) );
  XNOR U5135 ( .A(n5090), .B(n5101), .Z(n5094) );
  XNOR U5136 ( .A(n5091), .B(n5092), .Z(n5101) );
  AND U5137 ( .A(n2880), .B(n1203), .Z(n5091) );
  XOR U5138 ( .A(n5089), .B(n5102), .Z(n5090) );
  ANDN U5139 ( .A(n1210), .B(n2882), .Z(n5102) );
  XOR U5140 ( .A(n5103), .B(n5104), .Z(n5089) );
  ANDN U5141 ( .A(n5105), .B(n5106), .Z(n5104) );
  XNOR U5142 ( .A(n5107), .B(n5103), .Z(n5105) );
  XOR U5143 ( .A(n5108), .B(n5109), .Z(n5092) );
  AND U5144 ( .A(n5110), .B(n5111), .Z(n5109) );
  XNOR U5145 ( .A(n5099), .B(n5112), .Z(n5111) );
  XNOR U5146 ( .A(n5100), .B(n5108), .Z(n5112) );
  AND U5147 ( .A(n2748), .B(n1387), .Z(n5100) );
  XOR U5148 ( .A(n5098), .B(n5113), .Z(n5099) );
  ANDN U5149 ( .A(n1394), .B(n2750), .Z(n5113) );
  XNOR U5150 ( .A(n5106), .B(n5117), .Z(n5110) );
  XNOR U5151 ( .A(n5107), .B(n5108), .Z(n5117) );
  AND U5152 ( .A(n3019), .B(n1203), .Z(n5107) );
  XOR U5153 ( .A(n5103), .B(n5118), .Z(n5106) );
  ANDN U5154 ( .A(n1210), .B(n3021), .Z(n5118) );
  XNOR U5155 ( .A(n5123), .B(n5115), .Z(n4967) );
  XNOR U5156 ( .A(n5114), .B(n5124), .Z(n5115) );
  ANDN U5157 ( .A(n1394), .B(n2882), .Z(n5124) );
  XNOR U5158 ( .A(n5127), .B(n5125), .Z(n5126) );
  ANDN U5159 ( .A(n1394), .B(n3021), .Z(n5127) );
  XNOR U5160 ( .A(n5122), .B(n5116), .Z(n5123) );
  AND U5161 ( .A(n2880), .B(n1387), .Z(n5116) );
  XNOR U5162 ( .A(n5120), .B(n5121), .Z(n4966) );
  NAND U5163 ( .A(n3807), .B(n1203), .Z(n5121) );
  XNOR U5164 ( .A(n5119), .B(n5131), .Z(n5120) );
  ANDN U5165 ( .A(n1210), .B(n3809), .Z(n5131) );
  NAND U5166 ( .A(g_input[0]), .B(n5132), .Z(n5119) );
  NANDN U5167 ( .B(n1203), .A(n5133), .Z(n5132) );
  NANDN U5168 ( .B(n3812), .A(n1210), .Z(n5133) );
  IV U5169 ( .A(n1129), .Z(n1203) );
  XNOR U5170 ( .A(n5129), .B(n5130), .Z(n5122) );
  NAND U5171 ( .A(n3807), .B(n1387), .Z(n5130) );
  XNOR U5172 ( .A(n5128), .B(n5136), .Z(n5129) );
  ANDN U5173 ( .A(n1394), .B(n3809), .Z(n5136) );
  NAND U5174 ( .A(g_input[0]), .B(n5137), .Z(n5128) );
  NANDN U5175 ( .B(n1387), .A(n5138), .Z(n5137) );
  NANDN U5176 ( .B(n3812), .A(n1394), .Z(n5138) );
  IV U5177 ( .A(n1294), .Z(n1387) );
  XNOR U5178 ( .A(n3002), .B(n3001), .Z(n2978) );
  XOR U5179 ( .A(n5141), .B(n3010), .Z(n3001) );
  XNOR U5180 ( .A(n2998), .B(n2999), .Z(n3010) );
  NANDN U5181 ( .B(n647), .A(n2616), .Z(n2999) );
  XNOR U5182 ( .A(n2997), .B(n5142), .Z(n2998) );
  ANDN U5183 ( .A(n688), .B(n2618), .Z(n5142) );
  XOR U5184 ( .A(n3009), .B(n3000), .Z(n5141) );
  XOR U5185 ( .A(n5146), .B(n5147), .Z(n3000) );
  XOR U5186 ( .A(n5148), .B(n3006), .Z(n3009) );
  XNOR U5187 ( .A(n3005), .B(n5149), .Z(n3006) );
  ANDN U5188 ( .A(n795), .B(n2371), .Z(n5149) );
  XNOR U5189 ( .A(n5061), .B(g_input[8]), .Z(n5062) );
  ANDN U5190 ( .A(n5150), .B(n5151), .Z(n5061) );
  AND U5191 ( .A(n2369), .B(n741), .Z(n3007) );
  IV U5192 ( .A(n2493), .Z(n2369) );
  XNOR U5193 ( .A(n5155), .B(n5156), .Z(n3008) );
  AND U5194 ( .A(n5157), .B(n5158), .Z(n5156) );
  XNOR U5195 ( .A(n5153), .B(n5159), .Z(n5158) );
  XNOR U5196 ( .A(n5154), .B(n5155), .Z(n5159) );
  AND U5197 ( .A(n2491), .B(n741), .Z(n5154) );
  IV U5198 ( .A(n2618), .Z(n2491) );
  XOR U5199 ( .A(n5152), .B(n5160), .Z(n5153) );
  ANDN U5200 ( .A(n795), .B(n2493), .Z(n5160) );
  ANDN U5201 ( .A(n5161), .B(n5162), .Z(n5150) );
  XNOR U5202 ( .A(n5144), .B(n5166), .Z(n5157) );
  XNOR U5203 ( .A(n5145), .B(n5155), .Z(n5166) );
  ANDN U5204 ( .A(n2748), .B(n647), .Z(n5145) );
  XOR U5205 ( .A(n5143), .B(n5167), .Z(n5144) );
  ANDN U5206 ( .A(n688), .B(n2750), .Z(n5167) );
  XOR U5207 ( .A(n5171), .B(n5172), .Z(n5155) );
  AND U5208 ( .A(n5173), .B(n5174), .Z(n5172) );
  XNOR U5209 ( .A(n5164), .B(n5175), .Z(n5174) );
  XNOR U5210 ( .A(n5165), .B(n5171), .Z(n5175) );
  AND U5211 ( .A(n2616), .B(n741), .Z(n5165) );
  IV U5212 ( .A(n2750), .Z(n2616) );
  XOR U5213 ( .A(n5163), .B(n5176), .Z(n5164) );
  ANDN U5214 ( .A(n795), .B(n2618), .Z(n5176) );
  XNOR U5215 ( .A(n5161), .B(g_input[6]), .Z(n5162) );
  ANDN U5216 ( .A(n5177), .B(n5178), .Z(n5161) );
  XNOR U5217 ( .A(n5169), .B(n5182), .Z(n5173) );
  XNOR U5218 ( .A(n5170), .B(n5171), .Z(n5182) );
  ANDN U5219 ( .A(n2880), .B(n647), .Z(n5170) );
  XOR U5220 ( .A(n5168), .B(n5183), .Z(n5169) );
  ANDN U5221 ( .A(n688), .B(n2882), .Z(n5183) );
  XOR U5222 ( .A(n5184), .B(n5185), .Z(n5168) );
  ANDN U5223 ( .A(n5186), .B(n5187), .Z(n5185) );
  XNOR U5224 ( .A(n5188), .B(n5184), .Z(n5186) );
  XOR U5225 ( .A(n5189), .B(n5190), .Z(n5171) );
  AND U5226 ( .A(n5191), .B(n5192), .Z(n5190) );
  XNOR U5227 ( .A(n5180), .B(n5193), .Z(n5192) );
  XNOR U5228 ( .A(n5181), .B(n5189), .Z(n5193) );
  AND U5229 ( .A(n2748), .B(n741), .Z(n5181) );
  XOR U5230 ( .A(n5179), .B(n5194), .Z(n5180) );
  ANDN U5231 ( .A(n795), .B(n2750), .Z(n5194) );
  ANDN U5232 ( .A(n5195), .B(n5196), .Z(n5177) );
  XNOR U5233 ( .A(n5187), .B(n5200), .Z(n5191) );
  XNOR U5234 ( .A(n5188), .B(n5189), .Z(n5200) );
  ANDN U5235 ( .A(n3019), .B(n647), .Z(n5188) );
  XOR U5236 ( .A(n5184), .B(n5201), .Z(n5187) );
  ANDN U5237 ( .A(n688), .B(n3021), .Z(n5201) );
  XNOR U5238 ( .A(n5206), .B(n5198), .Z(n5147) );
  XNOR U5239 ( .A(n5197), .B(n5207), .Z(n5198) );
  ANDN U5240 ( .A(n795), .B(n2882), .Z(n5207) );
  XNOR U5241 ( .A(n5210), .B(n5208), .Z(n5209) );
  ANDN U5242 ( .A(n795), .B(n3021), .Z(n5210) );
  XNOR U5243 ( .A(n5205), .B(n5199), .Z(n5206) );
  AND U5244 ( .A(n2880), .B(n741), .Z(n5199) );
  XNOR U5245 ( .A(n5203), .B(n5204), .Z(n5146) );
  NANDN U5246 ( .B(n647), .A(n3807), .Z(n5204) );
  XNOR U5247 ( .A(n5202), .B(n5215), .Z(n5203) );
  ANDN U5248 ( .A(n688), .B(n3809), .Z(n5215) );
  NAND U5249 ( .A(g_input[0]), .B(n5216), .Z(n5202) );
  NAND U5250 ( .A(n5217), .B(n647), .Z(n5216) );
  NANDN U5251 ( .B(n3812), .A(n688), .Z(n5217) );
  XNOR U5252 ( .A(n5213), .B(n5214), .Z(n5205) );
  NAND U5253 ( .A(n3807), .B(n741), .Z(n5214) );
  XNOR U5254 ( .A(n5212), .B(n5220), .Z(n5213) );
  ANDN U5255 ( .A(n795), .B(n3809), .Z(n5220) );
  NAND U5256 ( .A(g_input[0]), .B(n5221), .Z(n5212) );
  NANDN U5257 ( .B(n741), .A(n5222), .Z(n5221) );
  NANDN U5258 ( .B(n3812), .A(n795), .Z(n5222) );
  IV U5259 ( .A(n5211), .Z(n741) );
  XOR U5260 ( .A(n3018), .B(n3017), .Z(n3002) );
  XOR U5261 ( .A(n5225), .B(n3014), .Z(n3017) );
  XNOR U5262 ( .A(n3013), .B(n5226), .Z(n3014) );
  ANDN U5263 ( .A(n620), .B(n2882), .Z(n5226) );
  IV U5264 ( .A(n2748), .Z(n2882) );
  XNOR U5265 ( .A(n5195), .B(g_input[4]), .Z(n5196) );
  ANDN U5266 ( .A(n5227), .B(n5228), .Z(n5195) );
  XNOR U5267 ( .A(n5231), .B(n5229), .Z(n5230) );
  ANDN U5268 ( .A(n620), .B(n3021), .Z(n5231) );
  IV U5269 ( .A(n2880), .Z(n3021) );
  IV U5270 ( .A(n3809), .Z(n3019) );
  XNOR U5271 ( .A(n3016), .B(n3015), .Z(n5225) );
  AND U5272 ( .A(n2880), .B(n579), .Z(n3015) );
  ANDN U5273 ( .A(n5236), .B(n5237), .Z(n5227) );
  XNOR U5274 ( .A(n5234), .B(n5235), .Z(n3016) );
  NAND U5275 ( .A(n3807), .B(n579), .Z(n5235) );
  XNOR U5276 ( .A(n5233), .B(n5238), .Z(n5234) );
  ANDN U5277 ( .A(n620), .B(n3809), .Z(n5238) );
  NAND U5278 ( .A(g_input[0]), .B(n5239), .Z(n5233) );
  NANDN U5279 ( .B(n579), .A(n5240), .Z(n5239) );
  NANDN U5280 ( .B(n3812), .A(n620), .Z(n5240) );
  IV U5281 ( .A(n5232), .Z(n579) );
  XOR U5282 ( .A(n3025), .B(n3024), .Z(n3018) );
  NAND U5283 ( .A(n3807), .B(n523), .Z(n3024) );
  IV U5284 ( .A(n3812), .Z(n3807) );
  XOR U5285 ( .A(n3023), .B(n5243), .Z(n3025) );
  ANDN U5286 ( .A(n554), .B(n3809), .Z(n5243) );
  XNOR U5287 ( .A(n5236), .B(g_input[2]), .Z(n5237) );
  NOR U5288 ( .A(g_input[0]), .B(n5244), .Z(n5236) );
  NANDN U5289 ( .B(n523), .A(n5246), .Z(n5245) );
  NANDN U5290 ( .B(n3812), .A(n554), .Z(n5246) );
  XOR U5291 ( .A(g_input[0]), .B(g_input[1]), .Z(n5244) );
  AND U5292 ( .A(n5248), .B(n5247), .Z(n523) );
  ANDN U5293 ( .A(e_input[31]), .B(n5249), .Z(n5248) );
  NANDN U5294 ( .B(n5250), .A(n5242), .Z(n5249) );
  XNOR U5295 ( .A(n5250), .B(e_input[29]), .Z(n5242) );
  NAND U5296 ( .A(n5241), .B(n5251), .Z(n5250) );
  XOR U5297 ( .A(n5251), .B(e_input[28]), .Z(n5241) );
  ANDN U5298 ( .A(n5218), .B(n5252), .Z(n5251) );
  XNOR U5299 ( .A(n5252), .B(e_input[27]), .Z(n5218) );
  NAND U5300 ( .A(n5219), .B(n5253), .Z(n5252) );
  XOR U5301 ( .A(n5253), .B(e_input[26]), .Z(n5219) );
  ANDN U5302 ( .A(n5224), .B(n5254), .Z(n5253) );
  XNOR U5303 ( .A(n5254), .B(e_input[25]), .Z(n5224) );
  NAND U5304 ( .A(n5223), .B(n5255), .Z(n5254) );
  XOR U5305 ( .A(n5255), .B(e_input[24]), .Z(n5223) );
  ANDN U5306 ( .A(n4964), .B(n5256), .Z(n5255) );
  XNOR U5307 ( .A(n5256), .B(e_input[23]), .Z(n4964) );
  NAND U5308 ( .A(n4965), .B(n5257), .Z(n5256) );
  XOR U5309 ( .A(n5257), .B(e_input[22]), .Z(n4965) );
  ANDN U5310 ( .A(n4960), .B(n5258), .Z(n5257) );
  XNOR U5311 ( .A(n5258), .B(e_input[21]), .Z(n4960) );
  NAND U5312 ( .A(n4959), .B(n5259), .Z(n5258) );
  XOR U5313 ( .A(n5259), .B(e_input[20]), .Z(n4959) );
  ANDN U5314 ( .A(n5135), .B(n5260), .Z(n5259) );
  XNOR U5315 ( .A(n5260), .B(e_input[19]), .Z(n5135) );
  NAND U5316 ( .A(n5134), .B(n5261), .Z(n5260) );
  XOR U5317 ( .A(n5261), .B(e_input[18]), .Z(n5134) );
  ANDN U5318 ( .A(n5140), .B(n5262), .Z(n5261) );
  XNOR U5319 ( .A(n5262), .B(e_input[17]), .Z(n5140) );
  NAND U5320 ( .A(n5139), .B(n5263), .Z(n5262) );
  XOR U5321 ( .A(n5263), .B(e_input[16]), .Z(n5139) );
  ANDN U5322 ( .A(n3837), .B(n5264), .Z(n5263) );
  XNOR U5323 ( .A(n5264), .B(e_input[15]), .Z(n3837) );
  NAND U5324 ( .A(n3836), .B(n5265), .Z(n5264) );
  XOR U5325 ( .A(n5265), .B(e_input[14]), .Z(n3836) );
  ANDN U5326 ( .A(n3832), .B(n5266), .Z(n5265) );
  XNOR U5327 ( .A(n5266), .B(e_input[13]), .Z(n3832) );
  NAND U5328 ( .A(n3831), .B(n5267), .Z(n5266) );
  XOR U5329 ( .A(n5267), .B(e_input[12]), .Z(n3831) );
  ANDN U5330 ( .A(n3814), .B(n5268), .Z(n5267) );
  XNOR U5331 ( .A(n5268), .B(e_input[11]), .Z(n3814) );
  NAND U5332 ( .A(n3813), .B(n5269), .Z(n5268) );
  XOR U5333 ( .A(n5269), .B(e_input[10]), .Z(n3813) );
  ANDN U5334 ( .A(n3819), .B(n5270), .Z(n5269) );
  XNOR U5335 ( .A(n5270), .B(e_input[9]), .Z(n3819) );
  NAND U5336 ( .A(n3818), .B(n5271), .Z(n5270) );
  XOR U5337 ( .A(n5271), .B(e_input[8]), .Z(n3818) );
  ANDN U5338 ( .A(n4343), .B(n5272), .Z(n5271) );
  XNOR U5339 ( .A(n5272), .B(e_input[7]), .Z(n4343) );
  NAND U5340 ( .A(n4342), .B(n5273), .Z(n5272) );
  XOR U5341 ( .A(n5273), .B(e_input[6]), .Z(n4342) );
  ANDN U5342 ( .A(n4338), .B(n5274), .Z(n5273) );
  XNOR U5343 ( .A(n5274), .B(e_input[5]), .Z(n4338) );
  NAND U5344 ( .A(n4337), .B(n5275), .Z(n5274) );
  XOR U5345 ( .A(n5275), .B(e_input[4]), .Z(n4337) );
  ANDN U5346 ( .A(n4772), .B(n5276), .Z(n5275) );
  XNOR U5347 ( .A(n5276), .B(e_input[3]), .Z(n4772) );
  NAND U5348 ( .A(n4771), .B(n5277), .Z(n5276) );
  XOR U5349 ( .A(n5277), .B(e_input[2]), .Z(n4771) );
  NOR U5350 ( .A(n4776), .B(e_input[0]), .Z(n5277) );
  XOR U5351 ( .A(e_input[0]), .B(e_input[1]), .Z(n4776) );
endmodule

