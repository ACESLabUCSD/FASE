
module MxM_TG_W8_N100 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n51 , \_MxM/n48 , \_MxM/n45 , \_MxM/n42 , \_MxM/n39 ,
         \_MxM/n36 , \_MxM/n33 , \_MxM/n30 , \_MxM/N17 , \_MxM/N16 ,
         \_MxM/N15 , \_MxM/N14 , \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N9 ,
         \_MxM/N8 , \_MxM/N7 , \_MxM/N6 , \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/Y1[0] , \_MxM/Y1[1] , \_MxM/Y1[2] , \_MxM/Y1[3] , \_MxM/Y1[4] ,
         \_MxM/Y1[5] , \_MxM/Y1[6] , \_MxM/Y1[7] , \_MxM/Y0[7] , \_MxM/Y0[6] ,
         \_MxM/Y0[5] , \_MxM/Y0[4] , \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] ,
         \_MxM/Y0[0] , \_MxM/add_43/carry[6] , \_MxM/add_43/carry[5] ,
         \_MxM/add_43/carry[4] , \_MxM/add_43/carry[3] ,
         \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362;

  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n30 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n33 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n36 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n39 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n42 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n45 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n48 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n51 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N14 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N13 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N12 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N11 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  MUX U1 ( .IN0(n1), .IN1(n220), .SEL(n221), .F(n266) );
  IV U2 ( .A(n288), .Z(n1) );
  MUX U3 ( .IN0(n236), .IN1(n251), .SEL(n238), .F(n230) );
  XOR U4 ( .A(n170), .B(n208), .Z(n171) );
  MUX U5 ( .IN0(e_input[5]), .IN1(n345), .SEL(e_input[7]), .F(n87) );
  XNOR U6 ( .A(n113), .B(n114), .Z(n112) );
  NAND U7 ( .A(n145), .B(n181), .Z(n180) );
  MUX U8 ( .IN0(n2), .IN1(n98), .SEL(n99), .F(n72) );
  IV U9 ( .A(\_MxM/Y0[3] ), .Z(n2) );
  XOR U10 ( .A(n322), .B(g_input[3]), .Z(n323) );
  XNOR U11 ( .A(n191), .B(n222), .Z(n192) );
  MUX U12 ( .IN0(e_input[3]), .IN1(n296), .SEL(e_input[7]), .F(n148) );
  MUX U13 ( .IN0(e_input[6]), .IN1(n350), .SEL(e_input[7]), .F(n70) );
  XNOR U14 ( .A(n154), .B(n124), .Z(n116) );
  MUX U15 ( .IN0(n151), .IN1(n3), .SEL(n152), .F(n108) );
  IV U16 ( .A(n153), .Z(n3) );
  MUX U17 ( .IN0(n4), .IN1(n72), .SEL(n73), .F(n43) );
  IV U18 ( .A(\_MxM/Y0[4] ), .Z(n4) );
  XNOR U19 ( .A(n309), .B(n310), .Z(n288) );
  MUX U20 ( .IN0(n242), .IN1(n260), .SEL(n244), .F(n215) );
  XOR U21 ( .A(n95), .B(n127), .Z(n96) );
  MUX U22 ( .IN0(n193), .IN1(n191), .SEL(n192), .F(n5) );
  IV U23 ( .A(n5), .Z(n150) );
  XNOR U24 ( .A(n206), .B(n205), .Z(n190) );
  NAND U25 ( .A(n89), .B(n119), .Z(n118) );
  XNOR U26 ( .A(n166), .B(n165), .Z(n153) );
  XNOR U27 ( .A(n117), .B(n116), .Z(n110) );
  XNOR U28 ( .A(n43), .B(n44), .Z(n25) );
  NOR U29 ( .A(g_input[0]), .B(n347), .Z(n337) );
  XOR U30 ( .A(n286), .B(n287), .Z(n220) );
  XNOR U31 ( .A(n318), .B(n199), .Z(n205) );
  MUX U32 ( .IN0(n91), .IN1(n112), .SEL(n90), .F(n59) );
  MUX U33 ( .IN0(g_input[6]), .IN1(n226), .SEL(g_input[7]), .F(n71) );
  MUX U34 ( .IN0(n6), .IN1(n110), .SEL(n109), .F(n83) );
  IV U35 ( .A(n108), .Z(n6) );
  MUX U36 ( .IN0(n7), .IN1(n132), .SEL(n133), .F(n98) );
  IV U37 ( .A(\_MxM/Y0[2] ), .Z(n7) );
  MUX U38 ( .IN0(\_MxM/Y0[6] ), .IN1(n25), .SEL(n24), .F(n22) );
  MUX U39 ( .IN0(g_input[1]), .IN1(n347), .SEL(g_input[7]), .F(n289) );
  MUX U40 ( .IN0(g_input[2]), .IN1(n336), .SEL(g_input[7]), .F(n207) );
  MUX U41 ( .IN0(g_input[3]), .IN1(n323), .SEL(g_input[7]), .F(n8) );
  IV U42 ( .A(n8), .Z(n167) );
  XNOR U43 ( .A(n194), .B(n159), .Z(n165) );
  MUX U44 ( .IN0(n185), .IN1(n9), .SEL(n184), .F(n145) );
  IV U45 ( .A(n183), .Z(n9) );
  AND U46 ( .A(n65), .B(n34), .Z(n64) );
  MUX U47 ( .IN0(n10), .IN1(n173), .SEL(n174), .F(n132) );
  IV U48 ( .A(\_MxM/Y0[1] ), .Z(n10) );
  XNOR U49 ( .A(n82), .B(n83), .Z(n102) );
  MUX U50 ( .IN0(\_MxM/Y0[7] ), .IN1(n22), .SEL(n23), .F(n11) );
  IV U51 ( .A(n11), .Z(n19) );
  MUX U52 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n12), .F(\_MxM/n51 ) );
  MUX U53 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n12), .F(\_MxM/n48 ) );
  MUX U54 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n12), .F(\_MxM/n45 ) );
  MUX U55 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n12), .F(\_MxM/n42 ) );
  MUX U56 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n12), .F(\_MxM/n39 ) );
  MUX U57 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n12), .F(\_MxM/n36 ) );
  IV U58 ( .A(n13), .Z(n12) );
  MUX U59 ( .IN0(o[6]), .IN1(\_MxM/Y1[6] ), .SEL(n13), .F(\_MxM/n33 ) );
  MUX U60 ( .IN0(o[7]), .IN1(\_MxM/Y1[7] ), .SEL(n13), .F(\_MxM/n30 ) );
  AND U61 ( .A(n14), .B(n15), .Z(n13) );
  ANDN U62 ( .A(n16), .B(\_MxM/n[2] ), .Z(n15) );
  NOR U63 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n16) );
  ANDN U64 ( .A(n17), .B(n18), .Z(n14) );
  ANDN U65 ( .A(\_MxM/N11 ), .B(\_MxM/n[1] ), .Z(n17) );
  XNOR U66 ( .A(n19), .B(n20), .Z(\_MxM/Y1[7] ) );
  XNOR U67 ( .A(\_MxM/Y0[7] ), .B(n21), .Z(n20) );
  XNOR U68 ( .A(n23), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XOR U69 ( .A(n22), .B(n21), .Z(n23) );
  XNOR U70 ( .A(n24), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XOR U71 ( .A(n25), .B(n26), .Z(n24) );
  ANDN U72 ( .A(n21), .B(n27), .Z(n26) );
  NANDN U73 ( .B(n28), .A(n29), .Z(n21) );
  ANDN U74 ( .A(n30), .B(n27), .Z(n28) );
  NAND U75 ( .A(n31), .B(n32), .Z(n27) );
  OR U76 ( .A(n33), .B(n34), .Z(n32) );
  AND U77 ( .A(n35), .B(n36), .Z(n31) );
  OR U78 ( .A(n37), .B(n38), .Z(n36) );
  OR U79 ( .A(n39), .B(n40), .Z(n35) );
  NOR U80 ( .A(n41), .B(n42), .Z(n30) );
  ANDN U81 ( .A(n45), .B(n46), .Z(n44) );
  XOR U82 ( .A(\_MxM/Y0[5] ), .B(n47), .Z(n45) );
  XNOR U83 ( .A(n46), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U84 ( .A(n48), .B(n49), .Z(n46) );
  XNOR U85 ( .A(n47), .B(n50), .Z(n48) );
  AND U86 ( .A(n29), .B(n51), .Z(n50) );
  XOR U87 ( .A(n41), .B(n52), .Z(n51) );
  XOR U88 ( .A(n52), .B(n42), .Z(n41) );
  OR U89 ( .A(n53), .B(n54), .Z(n42) );
  IV U90 ( .A(n49), .Z(n52) );
  XNOR U91 ( .A(n40), .B(n39), .Z(n49) );
  OR U92 ( .A(n55), .B(n56), .Z(n39) );
  AND U93 ( .A(n57), .B(n58), .Z(n40) );
  XNOR U94 ( .A(n59), .B(n60), .Z(n58) );
  ANDN U95 ( .A(n61), .B(n62), .Z(n60) );
  XOR U96 ( .A(n59), .B(n63), .Z(n61) );
  XNOR U97 ( .A(n33), .B(n64), .Z(n57) );
  NAND U98 ( .A(n66), .B(n67), .Z(n34) );
  NANDN U99 ( .B(n68), .A(n69), .Z(n66) );
  NANDN U100 ( .B(n37), .A(n70), .Z(n65) );
  NANDN U101 ( .B(n38), .A(n71), .Z(n33) );
  IV U102 ( .A(n43), .Z(n47) );
  XNOR U103 ( .A(n73), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U104 ( .A(n75), .B(n76), .Z(n73) );
  XNOR U105 ( .A(n74), .B(n77), .Z(n75) );
  AND U106 ( .A(n29), .B(n78), .Z(n77) );
  XOR U107 ( .A(n53), .B(n79), .Z(n78) );
  XOR U108 ( .A(n79), .B(n54), .Z(n53) );
  OR U109 ( .A(n80), .B(n81), .Z(n54) );
  IV U110 ( .A(n76), .Z(n79) );
  XNOR U111 ( .A(n56), .B(n55), .Z(n76) );
  OR U112 ( .A(n82), .B(n83), .Z(n55) );
  XOR U113 ( .A(n63), .B(n62), .Z(n56) );
  XOR U114 ( .A(n59), .B(n84), .Z(n62) );
  AND U115 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U116 ( .B(n37), .A(n87), .Z(n86) );
  OR U117 ( .A(n88), .B(n89), .Z(n85) );
  XOR U118 ( .A(n68), .B(n69), .Z(n63) );
  NANDN U119 ( .B(n38), .A(n92), .Z(n69) );
  XNOR U120 ( .A(n67), .B(n93), .Z(n68) );
  AND U121 ( .A(n71), .B(n70), .Z(n93) );
  ANDN U122 ( .A(n94), .B(n95), .Z(n67) );
  NANDN U123 ( .B(n96), .A(n97), .Z(n94) );
  IV U124 ( .A(n72), .Z(n74) );
  XNOR U125 ( .A(n99), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U126 ( .A(n101), .B(n102), .Z(n99) );
  XNOR U127 ( .A(n100), .B(n103), .Z(n101) );
  AND U128 ( .A(n29), .B(n104), .Z(n103) );
  XOR U129 ( .A(n80), .B(n105), .Z(n104) );
  XOR U130 ( .A(n105), .B(n81), .Z(n80) );
  OR U131 ( .A(n106), .B(n107), .Z(n81) );
  IV U132 ( .A(n102), .Z(n105) );
  XOR U133 ( .A(n91), .B(n90), .Z(n82) );
  XNOR U134 ( .A(n111), .B(n112), .Z(n90) );
  ANDN U135 ( .A(n115), .B(n116), .Z(n114) );
  XOR U136 ( .A(n113), .B(n117), .Z(n115) );
  XNOR U137 ( .A(n118), .B(n88), .Z(n111) );
  NAND U138 ( .A(n87), .B(n71), .Z(n88) );
  NANDN U139 ( .B(n37), .A(n120), .Z(n119) );
  XNOR U140 ( .A(n121), .B(n122), .Z(n89) );
  ANDN U141 ( .A(n123), .B(n124), .Z(n122) );
  XNOR U142 ( .A(n125), .B(n121), .Z(n123) );
  XOR U143 ( .A(n96), .B(n97), .Z(n91) );
  OR U144 ( .A(n126), .B(n38), .Z(n97) );
  AND U145 ( .A(n92), .B(n70), .Z(n127) );
  NAND U146 ( .A(n128), .B(n129), .Z(n95) );
  NANDN U147 ( .B(n130), .A(n131), .Z(n128) );
  IV U148 ( .A(n98), .Z(n100) );
  XNOR U149 ( .A(n133), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U150 ( .A(n134), .B(n135), .Z(n133) );
  XOR U151 ( .A(n132), .B(n136), .Z(n134) );
  AND U152 ( .A(n29), .B(n137), .Z(n136) );
  XOR U153 ( .A(n106), .B(n138), .Z(n137) );
  XOR U154 ( .A(n138), .B(n107), .Z(n106) );
  NANDN U155 ( .B(n139), .A(n140), .Z(n107) );
  IV U156 ( .A(n135), .Z(n138) );
  XOR U157 ( .A(n110), .B(n109), .Z(n135) );
  XNOR U158 ( .A(n108), .B(n141), .Z(n109) );
  AND U159 ( .A(n142), .B(n143), .Z(n141) );
  OR U160 ( .A(n144), .B(n145), .Z(n143) );
  AND U161 ( .A(n146), .B(n147), .Z(n142) );
  NANDN U162 ( .B(n37), .A(n148), .Z(n147) );
  NAND U163 ( .A(n149), .B(n150), .Z(n146) );
  XNOR U164 ( .A(n121), .B(n155), .Z(n124) );
  AND U165 ( .A(n71), .B(n120), .Z(n155) );
  XOR U166 ( .A(n156), .B(n157), .Z(n121) );
  ANDN U167 ( .A(n158), .B(n159), .Z(n157) );
  XNOR U168 ( .A(n160), .B(n156), .Z(n158) );
  XOR U169 ( .A(n161), .B(n125), .Z(n154) );
  NAND U170 ( .A(n87), .B(n92), .Z(n125) );
  IV U171 ( .A(n113), .Z(n161) );
  XOR U172 ( .A(n162), .B(n163), .Z(n113) );
  ANDN U173 ( .A(n164), .B(n165), .Z(n163) );
  XOR U174 ( .A(n162), .B(n166), .Z(n164) );
  XNOR U175 ( .A(n130), .B(n131), .Z(n117) );
  OR U176 ( .A(n167), .B(n38), .Z(n131) );
  XNOR U177 ( .A(n129), .B(n168), .Z(n130) );
  ANDN U178 ( .A(n70), .B(n126), .Z(n168) );
  ANDN U179 ( .A(n169), .B(n170), .Z(n129) );
  NANDN U180 ( .B(n171), .A(n172), .Z(n169) );
  XNOR U181 ( .A(n174), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U182 ( .A(n175), .B(n176), .Z(n174) );
  XNOR U183 ( .A(n177), .B(n173), .Z(n175) );
  NAND U184 ( .A(\_MxM/Y0[0] ), .B(n139), .Z(n173) );
  NAND U185 ( .A(n178), .B(n29), .Z(n177) );
  XOR U186 ( .A(e_input[7]), .B(g_input[7]), .Z(n29) );
  XNOR U187 ( .A(n140), .B(n176), .Z(n178) );
  XNOR U188 ( .A(n139), .B(n176), .Z(n140) );
  XNOR U189 ( .A(n153), .B(n152), .Z(n176) );
  XNOR U190 ( .A(n179), .B(n149), .Z(n152) );
  XNOR U191 ( .A(n180), .B(n144), .Z(n149) );
  NAND U192 ( .A(n71), .B(n148), .Z(n144) );
  NANDN U193 ( .B(n37), .A(n182), .Z(n181) );
  XNOR U194 ( .A(n150), .B(n151), .Z(n179) );
  XOR U195 ( .A(n186), .B(n187), .Z(n151) );
  AND U196 ( .A(n188), .B(n189), .Z(n187) );
  XNOR U197 ( .A(n186), .B(n190), .Z(n189) );
  XNOR U198 ( .A(n156), .B(n195), .Z(n159) );
  AND U199 ( .A(n92), .B(n120), .Z(n195) );
  XOR U200 ( .A(n196), .B(n197), .Z(n156) );
  ANDN U201 ( .A(n198), .B(n199), .Z(n197) );
  XNOR U202 ( .A(n200), .B(n196), .Z(n198) );
  XOR U203 ( .A(n201), .B(n160), .Z(n194) );
  NANDN U204 ( .B(n126), .A(n87), .Z(n160) );
  IV U205 ( .A(n162), .Z(n201) );
  XOR U206 ( .A(n202), .B(n203), .Z(n162) );
  ANDN U207 ( .A(n204), .B(n205), .Z(n203) );
  XOR U208 ( .A(n202), .B(n206), .Z(n204) );
  XNOR U209 ( .A(n171), .B(n172), .Z(n166) );
  NANDN U210 ( .B(n38), .A(n207), .Z(n172) );
  ANDN U211 ( .A(n70), .B(n167), .Z(n208) );
  NAND U212 ( .A(n209), .B(n210), .Z(n170) );
  NANDN U213 ( .B(n211), .A(n212), .Z(n209) );
  XNOR U214 ( .A(n190), .B(n188), .Z(n139) );
  XNOR U215 ( .A(n213), .B(n193), .Z(n188) );
  XNOR U216 ( .A(n184), .B(n185), .Z(n193) );
  NAND U217 ( .A(n92), .B(n148), .Z(n185) );
  XNOR U218 ( .A(n183), .B(n214), .Z(n184) );
  AND U219 ( .A(n182), .B(n71), .Z(n214) );
  XOR U220 ( .A(n215), .B(n216), .Z(n183) );
  AND U221 ( .A(n217), .B(n218), .Z(n216) );
  XNOR U222 ( .A(n219), .B(n215), .Z(n218) );
  XNOR U223 ( .A(n192), .B(n186), .Z(n213) );
  XOR U224 ( .A(n220), .B(n221), .Z(n186) );
  AND U225 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U226 ( .B(n37), .A(n225), .Z(n224) );
  NANDN U227 ( .B(n226), .A(n227), .Z(n37) );
  AND U228 ( .A(n228), .B(g_input[7]), .Z(n227) );
  NANDN U229 ( .B(n229), .A(n230), .Z(n223) );
  XNOR U230 ( .A(n231), .B(n232), .Z(n191) );
  AND U231 ( .A(n233), .B(n234), .Z(n232) );
  XOR U232 ( .A(n230), .B(n235), .Z(n234) );
  XNOR U233 ( .A(n229), .B(n231), .Z(n235) );
  NAND U234 ( .A(n71), .B(n225), .Z(n229) );
  XNOR U235 ( .A(n239), .B(n236), .Z(n238) );
  XOR U236 ( .A(n217), .B(n240), .Z(n233) );
  XNOR U237 ( .A(n219), .B(n231), .Z(n240) );
  NANDN U238 ( .B(n126), .A(n148), .Z(n219) );
  XOR U239 ( .A(n215), .B(n241), .Z(n217) );
  AND U240 ( .A(n182), .B(n92), .Z(n241) );
  XNOR U241 ( .A(n245), .B(n242), .Z(n244) );
  XOR U242 ( .A(n246), .B(n247), .Z(n231) );
  AND U243 ( .A(n248), .B(n249), .Z(n247) );
  XOR U244 ( .A(n237), .B(n250), .Z(n249) );
  XNOR U245 ( .A(n239), .B(n246), .Z(n250) );
  NAND U246 ( .A(n92), .B(n225), .Z(n239) );
  XOR U247 ( .A(n236), .B(n251), .Z(n237) );
  AND U248 ( .A(n71), .B(e_input[0]), .Z(n251) );
  XNOR U249 ( .A(n228), .B(g_input[6]), .Z(n226) );
  NOR U250 ( .A(n252), .B(n253), .Z(n228) );
  XOR U251 ( .A(n254), .B(n255), .Z(n236) );
  AND U252 ( .A(n256), .B(n257), .Z(n255) );
  XNOR U253 ( .A(n258), .B(n254), .Z(n257) );
  XOR U254 ( .A(n243), .B(n259), .Z(n248) );
  XNOR U255 ( .A(n245), .B(n246), .Z(n259) );
  NANDN U256 ( .B(n167), .A(n148), .Z(n245) );
  XOR U257 ( .A(n242), .B(n260), .Z(n243) );
  ANDN U258 ( .A(n182), .B(n126), .Z(n260) );
  XOR U259 ( .A(n261), .B(n262), .Z(n242) );
  AND U260 ( .A(n263), .B(n264), .Z(n262) );
  XNOR U261 ( .A(n265), .B(n261), .Z(n264) );
  XOR U262 ( .A(n266), .B(n267), .Z(n246) );
  AND U263 ( .A(n268), .B(n269), .Z(n267) );
  XOR U264 ( .A(n256), .B(n270), .Z(n269) );
  XNOR U265 ( .A(n258), .B(n266), .Z(n270) );
  NANDN U266 ( .B(n126), .A(n225), .Z(n258) );
  XOR U267 ( .A(n254), .B(n271), .Z(n256) );
  AND U268 ( .A(n92), .B(e_input[0]), .Z(n271) );
  XNOR U269 ( .A(n272), .B(g_input[5]), .Z(n92) );
  NAND U270 ( .A(n273), .B(g_input[7]), .Z(n272) );
  XOR U271 ( .A(n253), .B(g_input[5]), .Z(n273) );
  XOR U272 ( .A(n252), .B(g_input[5]), .Z(n253) );
  NANDN U273 ( .B(n274), .A(n275), .Z(n252) );
  XOR U274 ( .A(n276), .B(n277), .Z(n254) );
  ANDN U275 ( .A(n278), .B(n279), .Z(n277) );
  XNOR U276 ( .A(n280), .B(n276), .Z(n278) );
  XOR U277 ( .A(n263), .B(n281), .Z(n268) );
  XNOR U278 ( .A(n265), .B(n266), .Z(n281) );
  NAND U279 ( .A(n148), .B(n207), .Z(n265) );
  XOR U280 ( .A(n261), .B(n282), .Z(n263) );
  ANDN U281 ( .A(n182), .B(n167), .Z(n282) );
  XOR U282 ( .A(n283), .B(n284), .Z(n261) );
  ANDN U283 ( .A(n285), .B(n286), .Z(n284) );
  XNOR U284 ( .A(n287), .B(n283), .Z(n285) );
  NAND U285 ( .A(n148), .B(n289), .Z(n287) );
  XNOR U286 ( .A(n283), .B(n290), .Z(n286) );
  AND U287 ( .A(n207), .B(n182), .Z(n290) );
  AND U288 ( .A(n291), .B(g_input[0]), .Z(n283) );
  NANDN U289 ( .B(n148), .A(n292), .Z(n291) );
  NAND U290 ( .A(n289), .B(n182), .Z(n292) );
  XNOR U291 ( .A(n293), .B(e_input[2]), .Z(n182) );
  NAND U292 ( .A(n294), .B(e_input[7]), .Z(n293) );
  XOR U293 ( .A(n295), .B(e_input[2]), .Z(n294) );
  XNOR U294 ( .A(n297), .B(n298), .Z(n221) );
  IV U295 ( .A(n279), .Z(n298) );
  XNOR U296 ( .A(n276), .B(n299), .Z(n279) );
  ANDN U297 ( .A(e_input[0]), .B(n126), .Z(n299) );
  XOR U298 ( .A(n300), .B(n301), .Z(n276) );
  AND U299 ( .A(n302), .B(n303), .Z(n301) );
  XOR U300 ( .A(n304), .B(n300), .Z(n303) );
  ANDN U301 ( .A(e_input[0]), .B(n167), .Z(n304) );
  XOR U302 ( .A(n305), .B(n300), .Z(n302) );
  AND U303 ( .A(n225), .B(n207), .Z(n305) );
  XOR U304 ( .A(n306), .B(n307), .Z(n300) );
  ANDN U305 ( .A(n308), .B(n309), .Z(n307) );
  XNOR U306 ( .A(n310), .B(n306), .Z(n308) );
  XOR U307 ( .A(n311), .B(n280), .Z(n297) );
  NANDN U308 ( .B(n167), .A(n225), .Z(n280) );
  IV U309 ( .A(n288), .Z(n311) );
  NAND U310 ( .A(n225), .B(n289), .Z(n310) );
  XNOR U311 ( .A(n306), .B(n312), .Z(n309) );
  AND U312 ( .A(n207), .B(e_input[0]), .Z(n312) );
  AND U313 ( .A(n313), .B(g_input[0]), .Z(n306) );
  NANDN U314 ( .B(n225), .A(n314), .Z(n313) );
  NAND U315 ( .A(n289), .B(e_input[0]), .Z(n314) );
  XNOR U316 ( .A(n315), .B(e_input[1]), .Z(n225) );
  NAND U317 ( .A(n316), .B(e_input[7]), .Z(n315) );
  XNOR U318 ( .A(e_input[1]), .B(n317), .Z(n316) );
  XNOR U319 ( .A(n196), .B(n319), .Z(n199) );
  ANDN U320 ( .A(n120), .B(n126), .Z(n319) );
  XOR U321 ( .A(n320), .B(g_input[4]), .Z(n126) );
  NAND U322 ( .A(n321), .B(g_input[7]), .Z(n320) );
  XOR U323 ( .A(n274), .B(g_input[4]), .Z(n321) );
  XNOR U324 ( .A(n275), .B(g_input[4]), .Z(n274) );
  NOR U325 ( .A(n322), .B(n323), .Z(n275) );
  XOR U326 ( .A(n324), .B(n325), .Z(n196) );
  AND U327 ( .A(n326), .B(n327), .Z(n325) );
  XOR U328 ( .A(n328), .B(n324), .Z(n327) );
  ANDN U329 ( .A(n120), .B(n167), .Z(n328) );
  XOR U330 ( .A(n329), .B(n324), .Z(n326) );
  AND U331 ( .A(n207), .B(n87), .Z(n329) );
  XOR U332 ( .A(n330), .B(n331), .Z(n324) );
  ANDN U333 ( .A(n332), .B(n333), .Z(n331) );
  XNOR U334 ( .A(n334), .B(n330), .Z(n332) );
  XOR U335 ( .A(n335), .B(n200), .Z(n318) );
  NANDN U336 ( .B(n167), .A(n87), .Z(n200) );
  NANDN U337 ( .B(n336), .A(n337), .Z(n322) );
  IV U338 ( .A(n202), .Z(n335) );
  XOR U339 ( .A(n338), .B(n334), .Z(n202) );
  NAND U340 ( .A(n87), .B(n289), .Z(n334) );
  IV U341 ( .A(n333), .Z(n338) );
  XNOR U342 ( .A(n330), .B(n339), .Z(n333) );
  AND U343 ( .A(n207), .B(n120), .Z(n339) );
  AND U344 ( .A(n340), .B(g_input[0]), .Z(n330) );
  NANDN U345 ( .B(n87), .A(n341), .Z(n340) );
  NAND U346 ( .A(n289), .B(n120), .Z(n341) );
  XNOR U347 ( .A(n342), .B(e_input[4]), .Z(n120) );
  NAND U348 ( .A(n343), .B(e_input[7]), .Z(n342) );
  XOR U349 ( .A(n344), .B(e_input[4]), .Z(n343) );
  XNOR U350 ( .A(n211), .B(n212), .Z(n206) );
  NANDN U351 ( .B(n38), .A(n289), .Z(n212) );
  XNOR U352 ( .A(n210), .B(n346), .Z(n211) );
  AND U353 ( .A(n207), .B(n70), .Z(n346) );
  XNOR U354 ( .A(n337), .B(g_input[2]), .Z(n336) );
  AND U355 ( .A(n348), .B(g_input[0]), .Z(n210) );
  NAND U356 ( .A(n349), .B(n38), .Z(n348) );
  NANDN U357 ( .B(n350), .A(n351), .Z(n38) );
  ANDN U358 ( .A(e_input[7]), .B(n352), .Z(n351) );
  NAND U359 ( .A(n289), .B(n70), .Z(n349) );
  XOR U360 ( .A(n352), .B(e_input[6]), .Z(n350) );
  OR U361 ( .A(n345), .B(n353), .Z(n352) );
  XOR U362 ( .A(n353), .B(e_input[5]), .Z(n345) );
  OR U363 ( .A(n344), .B(n354), .Z(n353) );
  XOR U364 ( .A(n354), .B(e_input[4]), .Z(n344) );
  OR U365 ( .A(n296), .B(n355), .Z(n354) );
  XOR U366 ( .A(n355), .B(e_input[3]), .Z(n296) );
  OR U367 ( .A(n295), .B(n356), .Z(n355) );
  XOR U368 ( .A(n356), .B(e_input[2]), .Z(n295) );
  NANDN U369 ( .B(e_input[0]), .A(n317), .Z(n356) );
  XNOR U370 ( .A(e_input[0]), .B(e_input[1]), .Z(n317) );
  XOR U371 ( .A(g_input[0]), .B(g_input[1]), .Z(n347) );
  AND U372 ( .A(n357), .B(n358), .Z(\_MxM/N17 ) );
  XOR U373 ( .A(\_MxM/n[6] ), .B(\_MxM/add_43/carry[6] ), .Z(n358) );
  AND U374 ( .A(\_MxM/N9 ), .B(n357), .Z(\_MxM/N16 ) );
  AND U375 ( .A(\_MxM/N8 ), .B(n357), .Z(\_MxM/N15 ) );
  AND U376 ( .A(\_MxM/N7 ), .B(n357), .Z(\_MxM/N14 ) );
  AND U377 ( .A(\_MxM/N6 ), .B(n357), .Z(\_MxM/N13 ) );
  AND U378 ( .A(\_MxM/N5 ), .B(n357), .Z(\_MxM/N12 ) );
  NAND U379 ( .A(n359), .B(n360), .Z(n357) );
  ANDN U380 ( .A(n361), .B(n18), .Z(n360) );
  OR U381 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n18) );
  NOR U382 ( .A(\_MxM/N11 ), .B(\_MxM/n[2] ), .Z(n361) );
  AND U383 ( .A(\_MxM/n[6] ), .B(n362), .Z(n359) );
  AND U384 ( .A(\_MxM/n[5] ), .B(\_MxM/n[1] ), .Z(n362) );
  IV U385 ( .A(\_MxM/n[0] ), .Z(\_MxM/N11 ) );
endmodule

