
module MxM_TG_W32_N10000 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MxM/n390 , \_MxM/n389 , \_MxM/n388 , \_MxM/n387 , \_MxM/n386 ,
         \_MxM/n385 , \_MxM/n384 , \_MxM/n383 , \_MxM/n382 , \_MxM/n381 ,
         \_MxM/n380 , \_MxM/n379 , \_MxM/n378 , \_MxM/n377 , \_MxM/n376 ,
         \_MxM/n375 , \_MxM/n374 , \_MxM/n373 , \_MxM/n372 , \_MxM/n371 ,
         \_MxM/n370 , \_MxM/n369 , \_MxM/n368 , \_MxM/n367 , \_MxM/n366 ,
         \_MxM/n365 , \_MxM/n364 , \_MxM/n363 , \_MxM/n362 , \_MxM/n361 ,
         \_MxM/n360 , \_MxM/n359 , \_MxM/n358 , \_MxM/n357 , \_MxM/n356 ,
         \_MxM/n355 , \_MxM/n354 , \_MxM/n353 , \_MxM/n352 , \_MxM/n351 ,
         \_MxM/n350 , \_MxM/n349 , \_MxM/n348 , \_MxM/n347 , \_MxM/n346 ,
         \_MxM/n345 , \_MxM/n344 , \_MxM/n343 , \_MxM/n342 , \_MxM/n341 ,
         \_MxM/n340 , \_MxM/n339 , \_MxM/n338 , \_MxM/n337 , \_MxM/n336 ,
         \_MxM/n335 , \_MxM/n334 , \_MxM/n333 , \_MxM/n332 , \_MxM/n331 ,
         \_MxM/n330 , \_MxM/n329 , \_MxM/n328 , \_MxM/n327 , \_MxM/n326 ,
         \_MxM/n325 , \_MxM/n324 , \_MxM/n323 , \_MxM/n322 , \_MxM/n321 ,
         \_MxM/n320 , \_MxM/n319 , \_MxM/n318 , \_MxM/n317 , \_MxM/n316 ,
         \_MxM/n315 , \_MxM/n314 , \_MxM/n313 , \_MxM/N19 , \_MxM/N18 ,
         \_MxM/N17 , \_MxM/N16 , \_MxM/N15 , \_MxM/N14 , \_MxM/N13 ,
         \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/n[0] ,
         \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] ,
         \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/n[10] ,
         \_MxM/n[11] , \_MxM/n[12] , \_MxM/n[13] , \_MxM/Y0[0] , \_MxM/Y0[1] ,
         \_MxM/Y0[2] , \_MxM/Y0[3] , \_MxM/Y0[4] , \_MxM/Y0[5] , \_MxM/Y0[6] ,
         \_MxM/Y0[7] , \_MxM/Y0[8] , \_MxM/Y0[9] , \_MxM/Y0[10] ,
         \_MxM/Y0[11] , \_MxM/Y0[12] , \_MxM/Y0[13] , \_MxM/Y0[14] ,
         \_MxM/Y0[15] , \_MxM/Y0[16] , \_MxM/Y0[17] , \_MxM/Y0[18] ,
         \_MxM/Y0[19] , \_MxM/Y0[20] , \_MxM/Y0[21] , \_MxM/Y0[22] ,
         \_MxM/Y0[23] , \_MxM/Y0[24] , \_MxM/Y0[25] , \_MxM/Y0[26] ,
         \_MxM/Y0[27] , \_MxM/Y0[28] , \_MxM/Y0[29] , \_MxM/Y0[30] ,
         \_MxM/Y0[31] , \_MxM/add_39/carry[13] , \_MxM/add_39/carry[12] ,
         \_MxM/add_39/carry[11] , \_MxM/add_39/carry[10] ,
         \_MxM/add_39/carry[9] , \_MxM/add_39/carry[8] ,
         \_MxM/add_39/carry[7] , \_MxM/add_39/carry[6] ,
         \_MxM/add_39/carry[5] , \_MxM/add_39/carry[4] ,
         \_MxM/add_39/carry[3] , \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n313 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n314 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n315 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n316 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n317 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n318 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n319 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n320 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n321 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n322 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n323 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n324 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n325 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n326 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n327 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n328 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y_reg[16]  ( .D(\_MxM/n329 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[16]) );
  DFF \_MxM/Y_reg[17]  ( .D(\_MxM/n330 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[17]) );
  DFF \_MxM/Y_reg[18]  ( .D(\_MxM/n331 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[18]) );
  DFF \_MxM/Y_reg[19]  ( .D(\_MxM/n332 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[19]) );
  DFF \_MxM/Y_reg[20]  ( .D(\_MxM/n333 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[20]) );
  DFF \_MxM/Y_reg[21]  ( .D(\_MxM/n334 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[21]) );
  DFF \_MxM/Y_reg[22]  ( .D(\_MxM/n335 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[22]) );
  DFF \_MxM/Y_reg[23]  ( .D(\_MxM/n336 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[23]) );
  DFF \_MxM/Y_reg[24]  ( .D(\_MxM/n337 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[24]) );
  DFF \_MxM/Y_reg[25]  ( .D(\_MxM/n338 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[25]) );
  DFF \_MxM/Y_reg[26]  ( .D(\_MxM/n339 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[26]) );
  DFF \_MxM/Y_reg[27]  ( .D(\_MxM/n340 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[27]) );
  DFF \_MxM/Y_reg[28]  ( .D(\_MxM/n341 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[28]) );
  DFF \_MxM/Y_reg[29]  ( .D(\_MxM/n342 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[29]) );
  DFF \_MxM/Y_reg[30]  ( .D(\_MxM/n343 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[30]) );
  DFF \_MxM/Y_reg[31]  ( .D(\_MxM/n344 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[31]) );
  DFF \_MxM/Y0_reg[31]  ( .D(\_MxM/n345 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[31] ) );
  DFF \_MxM/Y0_reg[30]  ( .D(\_MxM/n346 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[30] ) );
  DFF \_MxM/Y0_reg[29]  ( .D(\_MxM/n347 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[29] ) );
  DFF \_MxM/Y0_reg[28]  ( .D(\_MxM/n348 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[28] ) );
  DFF \_MxM/Y0_reg[27]  ( .D(\_MxM/n349 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[27] ) );
  DFF \_MxM/Y0_reg[26]  ( .D(\_MxM/n350 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[26] ) );
  DFF \_MxM/Y0_reg[25]  ( .D(\_MxM/n351 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[25] ) );
  DFF \_MxM/Y0_reg[24]  ( .D(\_MxM/n352 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[24] ) );
  DFF \_MxM/Y0_reg[23]  ( .D(\_MxM/n353 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[23] ) );
  DFF \_MxM/Y0_reg[22]  ( .D(\_MxM/n354 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[22] ) );
  DFF \_MxM/Y0_reg[21]  ( .D(\_MxM/n355 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[21] ) );
  DFF \_MxM/Y0_reg[20]  ( .D(\_MxM/n356 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[20] ) );
  DFF \_MxM/Y0_reg[19]  ( .D(\_MxM/n357 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[19] ) );
  DFF \_MxM/Y0_reg[18]  ( .D(\_MxM/n358 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[18] ) );
  DFF \_MxM/Y0_reg[17]  ( .D(\_MxM/n359 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[17] ) );
  DFF \_MxM/Y0_reg[16]  ( .D(\_MxM/n360 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[16] ) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/n361 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/n362 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/n363 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/n364 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/n365 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/n366 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/n367 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/n368 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n369 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n370 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n371 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n372 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n373 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n374 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n375 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n376 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[13]  ( .D(\_MxM/n377 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[13] ) );
  DFF \_MxM/n_reg[12]  ( .D(\_MxM/n378 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[12] ) );
  DFF \_MxM/n_reg[11]  ( .D(\_MxM/n379 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[11] ) );
  DFF \_MxM/n_reg[10]  ( .D(\_MxM/n380 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[10] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/n381 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/n382 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/n383 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n384 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n385 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n386 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n387 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n388 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n389 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n390 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N14 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N15 ) );
  HADDER \_MxM/add_39/U1_1_9  ( .IN0(\_MxM/n[9] ), .IN1(\_MxM/add_39/carry[9] ), .COUT(\_MxM/add_39/carry[10] ), .SUM(\_MxM/N16 ) );
  HADDER \_MxM/add_39/U1_1_10  ( .IN0(\_MxM/n[10] ), .IN1(
        \_MxM/add_39/carry[10] ), .COUT(\_MxM/add_39/carry[11] ), .SUM(
        \_MxM/N17 ) );
  HADDER \_MxM/add_39/U1_1_11  ( .IN0(\_MxM/n[11] ), .IN1(
        \_MxM/add_39/carry[11] ), .COUT(\_MxM/add_39/carry[12] ), .SUM(
        \_MxM/N18 ) );
  HADDER \_MxM/add_39/U1_1_12  ( .IN0(\_MxM/n[12] ), .IN1(
        \_MxM/add_39/carry[12] ), .COUT(\_MxM/add_39/carry[13] ), .SUM(
        \_MxM/N19 ) );
  MUX U1 ( .IN0(n3714), .IN1(n1), .SEL(n3715), .F(n3668) );
  IV U2 ( .A(n3716), .Z(n1) );
  MUX U3 ( .IN0(n3542), .IN1(n3544), .SEL(n3543), .F(n3496) );
  MUX U4 ( .IN0(n4315), .IN1(n4317), .SEL(n4316), .F(n4291) );
  MUX U5 ( .IN0(n3367), .IN1(n3369), .SEL(n3368), .F(n3321) );
  XNOR U6 ( .A(n4303), .B(n4302), .Z(n4318) );
  XNOR U7 ( .A(n4686), .B(n4684), .Z(n4691) );
  MUX U8 ( .IN0(n3271), .IN1(n3273), .SEL(n3272), .F(n3228) );
  MUX U9 ( .IN0(n5019), .IN1(n5021), .SEL(n5020), .F(n5007) );
  MUX U10 ( .IN0(n4877), .IN1(n2), .SEL(n4878), .F(n4857) );
  IV U11 ( .A(n4879), .Z(n2) );
  MUX U12 ( .IN0(n5026), .IN1(n3), .SEL(n5027), .F(n5014) );
  IV U13 ( .A(n5028), .Z(n3) );
  MUX U14 ( .IN0(n4236), .IN1(n4), .SEL(n4237), .F(n4216) );
  IV U15 ( .A(n4238), .Z(n4) );
  XNOR U16 ( .A(n3224), .B(n3223), .Z(n3260) );
  MUX U17 ( .IN0(n4641), .IN1(n5), .SEL(n4642), .F(n4631) );
  IV U18 ( .A(n4643), .Z(n5) );
  XNOR U19 ( .A(n3249), .B(n3247), .Z(n3284) );
  XNOR U20 ( .A(n4412), .B(n4410), .Z(n4419) );
  NANDN U21 ( .B(n1298), .A(n3025), .Z(n18) );
  MUX U22 ( .IN0(n3101), .IN1(n3103), .SEL(n3102), .F(n3062) );
  MUX U23 ( .IN0(n3094), .IN1(n6), .SEL(n3095), .F(n3055) );
  IV U24 ( .A(n3096), .Z(n6) );
  MUX U25 ( .IN0(n3106), .IN1(n3108), .SEL(n3107), .F(n3035) );
  MUX U26 ( .IN0(n1009), .IN1(n7), .SEL(n1010), .F(n940) );
  IV U27 ( .A(n1011), .Z(n7) );
  MUX U28 ( .IN0(n1306), .IN1(n1308), .SEL(n1307), .F(n1222) );
  MUX U29 ( .IN0(n1361), .IN1(n8), .SEL(n1362), .F(n1270) );
  IV U30 ( .A(n1363), .Z(n8) );
  MUX U31 ( .IN0(n1409), .IN1(n9), .SEL(n1410), .F(n1314) );
  IV U32 ( .A(n1411), .Z(n9) );
  MUX U33 ( .IN0(n1514), .IN1(n10), .SEL(n1515), .F(n1417) );
  IV U34 ( .A(n1516), .Z(n10) );
  MUX U35 ( .IN0(n1773), .IN1(n1775), .SEL(n1774), .F(n1672) );
  MUX U36 ( .IN0(n1889), .IN1(n11), .SEL(n1890), .F(n1781) );
  IV U37 ( .A(n1891), .Z(n11) );
  MUX U38 ( .IN0(n2062), .IN1(n12), .SEL(n2063), .F(n1953) );
  IV U39 ( .A(n2064), .Z(n12) );
  MUX U40 ( .IN0(g_input[29]), .IN1(n4387), .SEL(g_input[31]), .F(n13) );
  IV U41 ( .A(n13), .Z(n633) );
  MUX U42 ( .IN0(n14), .IN1(n4376), .SEL(g_input[31]), .F(n589) );
  IV U43 ( .A(g_input[30]), .Z(n14) );
  MUX U44 ( .IN0(n4938), .IN1(n4940), .SEL(n4939), .F(n4914) );
  MUX U45 ( .IN0(n4688), .IN1(n4690), .SEL(n4689), .F(n4673) );
  XNOR U46 ( .A(n5060), .B(n5058), .Z(n5065) );
  MUX U47 ( .IN0(n4271), .IN1(n4273), .SEL(n4272), .F(n4251) );
  MUX U48 ( .IN0(n4276), .IN1(n15), .SEL(n4277), .F(n4256) );
  IV U49 ( .A(n4278), .Z(n15) );
  XNOR U50 ( .A(n4926), .B(n4925), .Z(n4941) );
  MUX U51 ( .IN0(n5007), .IN1(n5009), .SEL(n5008), .F(n4995) );
  MUX U52 ( .IN0(n4857), .IN1(n16), .SEL(n4858), .F(n4837) );
  IV U53 ( .A(n4859), .Z(n16) );
  MUX U54 ( .IN0(n5014), .IN1(n17), .SEL(n5015), .F(n5002) );
  IV U55 ( .A(n5016), .Z(n17) );
  MUX U56 ( .IN0(n3186), .IN1(n3188), .SEL(n3187), .F(n3141) );
  XNOR U57 ( .A(n4644), .B(n4643), .Z(n4649) );
  MUX U58 ( .IN0(n4636), .IN1(n4638), .SEL(n4637), .F(n4626) );
  MUX U59 ( .IN0(n5131), .IN1(n18), .SEL(n5132), .F(n5120) );
  XNOR U60 ( .A(n3137), .B(n3136), .Z(n3175) );
  MUX U61 ( .IN0(n4621), .IN1(n19), .SEL(n4622), .F(n4608) );
  IV U62 ( .A(n4623), .Z(n19) );
  MUX U63 ( .IN0(n3055), .IN1(n20), .SEL(n3056), .F(n2925) );
  IV U64 ( .A(n3057), .Z(n20) );
  MUX U65 ( .IN0(n1161), .IN1(n21), .SEL(n1162), .F(n1081) );
  IV U66 ( .A(n1163), .Z(n21) );
  MUX U67 ( .IN0(n1222), .IN1(n1224), .SEL(n1223), .F(n1141) );
  MUX U68 ( .IN0(n1279), .IN1(n1281), .SEL(n1280), .F(n1197) );
  MUX U69 ( .IN0(n1594), .IN1(n1596), .SEL(n1595), .F(n1498) );
  MUX U70 ( .IN0(n1602), .IN1(n22), .SEL(n1603), .F(n1506) );
  IV U71 ( .A(n1604), .Z(n22) );
  MUX U72 ( .IN0(n1610), .IN1(n23), .SEL(n1611), .F(n1514) );
  IV U73 ( .A(n1612), .Z(n23) );
  MUX U74 ( .IN0(n1657), .IN1(n24), .SEL(n1658), .F(n1557) );
  IV U75 ( .A(n1659), .Z(n24) );
  MUX U76 ( .IN0(n1854), .IN1(n1856), .SEL(n1855), .F(n1746) );
  MUX U77 ( .IN0(n1996), .IN1(n25), .SEL(n1997), .F(n1889) );
  IV U78 ( .A(n1998), .Z(n25) );
  MUX U79 ( .IN0(n2176), .IN1(n26), .SEL(n2177), .F(n2062) );
  IV U80 ( .A(n2178), .Z(n26) );
  MUX U81 ( .IN0(n2802), .IN1(n27), .SEL(n2803), .F(n2677) );
  IV U82 ( .A(n2804), .Z(n27) );
  MUX U83 ( .IN0(n709), .IN1(n28), .SEL(n710), .F(n663) );
  IV U84 ( .A(n711), .Z(n28) );
  MUX U85 ( .IN0(n2958), .IN1(n2960), .SEL(n2959), .F(n2818) );
  MUX U86 ( .IN0(n29), .IN1(n744), .SEL(n743), .F(n706) );
  IV U87 ( .A(n742), .Z(n29) );
  MUX U88 ( .IN0(n3722), .IN1(n3724), .SEL(n3723), .F(n3678) );
  MUX U89 ( .IN0(n4700), .IN1(n4702), .SEL(n4701), .F(n4688) );
  XNOR U90 ( .A(n4698), .B(n4697), .Z(n4703) );
  MUX U91 ( .IN0(n4892), .IN1(n4894), .SEL(n4893), .F(n4872) );
  MUX U92 ( .IN0(n5040), .IN1(n30), .SEL(n5041), .F(n5026) );
  IV U93 ( .A(n5042), .Z(n30) );
  MUX U94 ( .IN0(n4251), .IN1(n4253), .SEL(n4252), .F(n4231) );
  MUX U95 ( .IN0(n4256), .IN1(n31), .SEL(n4257), .F(n4236) );
  IV U96 ( .A(n4258), .Z(n31) );
  MUX U97 ( .IN0(n3235), .IN1(n3237), .SEL(n3236), .F(n3191) );
  XNOR U98 ( .A(n4860), .B(n4859), .Z(n4875) );
  MUX U99 ( .IN0(n4995), .IN1(n4997), .SEL(n4996), .F(n4983) );
  XNOR U100 ( .A(n5005), .B(n5004), .Z(n5010) );
  NANDN U101 ( .B(n2054), .A(n3025), .Z(n44) );
  MUX U102 ( .IN0(n4631), .IN1(n32), .SEL(n4632), .F(n4621) );
  IV U103 ( .A(n4633), .Z(n32) );
  MUX U104 ( .IN0(n4626), .IN1(n4628), .SEL(n4627), .F(n4616) );
  XNOR U105 ( .A(n3097), .B(n3096), .Z(n3130) );
  MUX U106 ( .IN0(n1401), .IN1(n1403), .SEL(n1402), .F(n1306) );
  MUX U107 ( .IN0(n1698), .IN1(n33), .SEL(n1699), .F(n1602) );
  IV U108 ( .A(n1700), .Z(n33) );
  MUX U109 ( .IN0(n1706), .IN1(n34), .SEL(n1707), .F(n1610) );
  IV U110 ( .A(n1708), .Z(n34) );
  MUX U111 ( .IN0(n1664), .IN1(n1666), .SEL(n1665), .F(n1566) );
  MUX U112 ( .IN0(n1672), .IN1(n1674), .SEL(n1673), .F(n1574) );
  MUX U113 ( .IN0(n1758), .IN1(n35), .SEL(n1759), .F(n1657) );
  IV U114 ( .A(n1760), .Z(n35) );
  MUX U115 ( .IN0(n1791), .IN1(n1793), .SEL(n1792), .F(n1690) );
  MUX U116 ( .IN0(n1962), .IN1(n1964), .SEL(n1963), .F(n1854) );
  MUX U117 ( .IN0(n2104), .IN1(n36), .SEL(n2105), .F(n1996) );
  IV U118 ( .A(n2106), .Z(n36) );
  MUX U119 ( .IN0(n2272), .IN1(n2274), .SEL(n2273), .F(n2153) );
  MUX U120 ( .IN0(n2410), .IN1(n37), .SEL(n2411), .F(n2290) );
  IV U121 ( .A(n2412), .Z(n37) );
  MUX U122 ( .IN0(n2941), .IN1(n38), .SEL(n2942), .F(n2802) );
  IV U123 ( .A(n2943), .Z(n38) );
  MUX U124 ( .IN0(n735), .IN1(n737), .SEL(n736), .F(n693) );
  MUX U125 ( .IN0(n625), .IN1(n39), .SEL(n626), .F(n579) );
  IV U126 ( .A(n627), .Z(n39) );
  MUX U127 ( .IN0(n40), .IN1(n971), .SEL(n970), .F(n906) );
  IV U128 ( .A(n969), .Z(n40) );
  MUX U129 ( .IN0(n5062), .IN1(n5064), .SEL(n5063), .F(n5045) );
  MUX U130 ( .IN0(n4943), .IN1(n41), .SEL(n4944), .F(n4921) );
  IV U131 ( .A(n4945), .Z(n41) );
  MUX U132 ( .IN0(n4761), .IN1(n4763), .SEL(n4762), .F(n4745) );
  MUX U133 ( .IN0(n4872), .IN1(n4874), .SEL(n4873), .F(n4852) );
  MUX U134 ( .IN0(n4646), .IN1(n4648), .SEL(n4647), .F(n4636) );
  XNOR U135 ( .A(n4428), .B(n4427), .Z(n4435) );
  MUX U136 ( .IN0(n4211), .IN1(n4213), .SEL(n4212), .F(n4191) );
  XNOR U137 ( .A(n4239), .B(n4238), .Z(n4254) );
  MUX U138 ( .IN0(n4837), .IN1(n42), .SEL(n4838), .F(n4817) );
  IV U139 ( .A(n4839), .Z(n42) );
  MUX U140 ( .IN0(n5002), .IN1(n43), .SEL(n5003), .F(n4990) );
  IV U141 ( .A(n5004), .Z(n43) );
  MUX U142 ( .IN0(n3807), .IN1(n44), .SEL(n3808), .F(n3796) );
  MUX U143 ( .IN0(n4983), .IN1(n4985), .SEL(n4984), .F(n4800) );
  MUX U144 ( .IN0(n4172), .IN1(n45), .SEL(n4173), .F(n4151) );
  IV U145 ( .A(n4174), .Z(n45) );
  XNOR U146 ( .A(n4624), .B(n4623), .Z(n4629) );
  MUX U147 ( .IN0(n3062), .IN1(n3064), .SEL(n3063), .F(n2932) );
  MUX U148 ( .IN0(n1470), .IN1(n1472), .SEL(n1471), .F(n1368) );
  MUX U149 ( .IN0(n1506), .IN1(n46), .SEL(n1507), .F(n1409) );
  IV U150 ( .A(n1508), .Z(n46) );
  MUX U151 ( .IN0(n1498), .IN1(n1500), .SEL(n1499), .F(n1401) );
  MUX U152 ( .IN0(n1807), .IN1(n47), .SEL(n1808), .F(n1706) );
  IV U153 ( .A(n1809), .Z(n47) );
  MUX U154 ( .IN0(n1980), .IN1(n1982), .SEL(n1981), .F(n1873) );
  MUX U155 ( .IN0(n1973), .IN1(n48), .SEL(n1974), .F(n1866) );
  IV U156 ( .A(n1975), .Z(n48) );
  MUX U157 ( .IN0(n2012), .IN1(n49), .SEL(n2013), .F(n1905) );
  IV U158 ( .A(n2014), .Z(n49) );
  MUX U159 ( .IN0(n2069), .IN1(n2071), .SEL(n2070), .F(n1962) );
  MUX U160 ( .IN0(n2223), .IN1(n50), .SEL(n2224), .F(n2104) );
  IV U161 ( .A(n2225), .Z(n50) );
  MUX U162 ( .IN0(n2640), .IN1(n2642), .SEL(n2641), .F(n2516) );
  MUX U163 ( .IN0(n2648), .IN1(n51), .SEL(n2649), .F(n2524) );
  IV U164 ( .A(n2650), .Z(n51) );
  MUX U165 ( .IN0(g_input[28]), .IN1(n4405), .SEL(g_input[31]), .F(n52) );
  IV U166 ( .A(n52), .Z(n673) );
  MUX U167 ( .IN0(n693), .IN1(n695), .SEL(n694), .F(n652) );
  XNOR U168 ( .A(n974), .B(n971), .Z(n1034) );
  MUX U169 ( .IN0(n5125), .IN1(n5127), .SEL(n5126), .F(n5109) );
  MUX U170 ( .IN0(n53), .IN1(n4740), .SEL(n4741), .F(n4726) );
  IV U171 ( .A(n4742), .Z(n53) );
  XNOR U172 ( .A(n4259), .B(n4258), .Z(n4274) );
  MUX U173 ( .IN0(n5203), .IN1(n54), .SEL(n5204), .F(n5185) );
  IV U174 ( .A(n5205), .Z(n54) );
  MUX U175 ( .IN0(n4852), .IN1(n4854), .SEL(n4853), .F(n4832) );
  MUX U176 ( .IN0(n4191), .IN1(n4193), .SEL(n4192), .F(n4179) );
  NANDN U177 ( .B(n2549), .A(n3025), .Z(n67) );
  MUX U178 ( .IN0(n4196), .IN1(n55), .SEL(n4197), .F(n4172) );
  IV U179 ( .A(n4198), .Z(n55) );
  XNOR U180 ( .A(n3906), .B(n3904), .Z(n3919) );
  XNOR U181 ( .A(n4840), .B(n4839), .Z(n4855) );
  MUX U182 ( .IN0(n4990), .IN1(n56), .SEL(n4991), .F(n4978) );
  IV U183 ( .A(n4992), .Z(n56) );
  MUX U184 ( .IN0(n4616), .IN1(n4618), .SEL(n4617), .F(n4599) );
  MUX U185 ( .IN0(n4786), .IN1(n57), .SEL(n4787), .F(n2972) );
  IV U186 ( .A(n4788), .Z(n57) );
  MUX U187 ( .IN0(n1417), .IN1(n58), .SEL(n1418), .F(n1324) );
  IV U188 ( .A(n1419), .Z(n58) );
  MUX U189 ( .IN0(n1566), .IN1(n1568), .SEL(n1567), .F(n1470) );
  MUX U190 ( .IN0(n1690), .IN1(n1692), .SEL(n1691), .F(n1594) );
  MUX U191 ( .IN0(n1866), .IN1(n59), .SEL(n1867), .F(n1758) );
  IV U192 ( .A(n1868), .Z(n59) );
  MUX U193 ( .IN0(n2020), .IN1(n60), .SEL(n2021), .F(n1913) );
  IV U194 ( .A(n2022), .Z(n60) );
  MUX U195 ( .IN0(n2120), .IN1(n61), .SEL(n2121), .F(n2012) );
  IV U196 ( .A(n2122), .Z(n61) );
  MUX U197 ( .IN0(n2215), .IN1(n2217), .SEL(n2216), .F(n2096) );
  MUX U198 ( .IN0(n2207), .IN1(n2209), .SEL(n2208), .F(n2088) );
  MUX U199 ( .IN0(n2297), .IN1(n2299), .SEL(n2298), .F(n2183) );
  MUX U200 ( .IN0(n2590), .IN1(n62), .SEL(n2591), .F(n2465) );
  IV U201 ( .A(n2592), .Z(n62) );
  MUX U202 ( .IN0(n674), .IN1(n676), .SEL(n675), .F(n634) );
  MUX U203 ( .IN0(n1046), .IN1(n1048), .SEL(n1047), .F(n978) );
  MUX U204 ( .IN0(g_input[25]), .IN1(n4454), .SEL(g_input[31]), .F(n63) );
  IV U205 ( .A(n63), .Z(n818) );
  MUX U206 ( .IN0(n2045), .IN1(n2047), .SEL(n2046), .F(n1940) );
  XNOR U207 ( .A(n805), .B(n804), .Z(n860) );
  XNOR U208 ( .A(n290), .B(n1295), .Z(n1218) );
  AND U209 ( .A(n574), .B(n576), .Z(n545) );
  MUX U210 ( .IN0(n4756), .IN1(n64), .SEL(n4757), .F(n4740) );
  IV U211 ( .A(n4758), .Z(n64) );
  XNOR U212 ( .A(n4902), .B(n4901), .Z(n4919) );
  MUX U213 ( .IN0(n3801), .IN1(n3803), .SEL(n3802), .F(n3787) );
  MUX U214 ( .IN0(n4216), .IN1(n65), .SEL(n4217), .F(n4196) );
  IV U215 ( .A(n4218), .Z(n65) );
  XNOR U216 ( .A(n3182), .B(n3181), .Z(n3217) );
  MUX U217 ( .IN0(n66), .IN1(n5185), .SEL(n5186), .F(n5169) );
  IV U218 ( .A(n5187), .Z(n66) );
  MUX U219 ( .IN0(n4832), .IN1(n4834), .SEL(n4833), .F(n4812) );
  MUX U220 ( .IN0(n4334), .IN1(n67), .SEL(n4335), .F(n4320) );
  XNOR U221 ( .A(n4634), .B(n4633), .Z(n4639) );
  MUX U222 ( .IN0(n4817), .IN1(n68), .SEL(n4818), .F(n4786) );
  IV U223 ( .A(n4819), .Z(n68) );
  XNOR U224 ( .A(n3164), .B(n3162), .Z(n3199) );
  MUX U225 ( .IN0(n4978), .IN1(n69), .SEL(n4979), .F(n2995) );
  IV U226 ( .A(n4980), .Z(n69) );
  MUX U227 ( .IN0(n1913), .IN1(n70), .SEL(n1914), .F(n1807) );
  IV U228 ( .A(n1915), .Z(n70) );
  MUX U229 ( .IN0(n2351), .IN1(n2353), .SEL(n2352), .F(n2231) );
  MUX U230 ( .IN0(n2481), .IN1(n71), .SEL(n2482), .F(n2359) );
  IV U231 ( .A(n2483), .Z(n71) );
  MUX U232 ( .IN0(n2489), .IN1(n72), .SEL(n2490), .F(n2367) );
  IV U233 ( .A(n2491), .Z(n72) );
  MUX U234 ( .IN0(g_input[22]), .IN1(n4505), .SEL(g_input[31]), .F(n73) );
  IV U235 ( .A(n73), .Z(n1017) );
  MUX U236 ( .IN0(g_input[24]), .IN1(n4471), .SEL(g_input[31]), .F(n74) );
  IV U237 ( .A(n74), .Z(n882) );
  MUX U238 ( .IN0(g_input[17]), .IN1(n4590), .SEL(g_input[31]), .F(n75) );
  IV U239 ( .A(n75), .Z(n1425) );
  MUX U240 ( .IN0(g_input[19]), .IN1(n4556), .SEL(g_input[31]), .F(n76) );
  IV U241 ( .A(n76), .Z(n1250) );
  MUX U242 ( .IN0(g_input[26]), .IN1(n4438), .SEL(g_input[31]), .F(n77) );
  IV U243 ( .A(n77), .Z(n759) );
  MUX U244 ( .IN0(g_input[27]), .IN1(n4422), .SEL(g_input[31]), .F(n78) );
  IV U245 ( .A(n78), .Z(n717) );
  MUX U246 ( .IN0(n879), .IN1(n877), .SEL(n878), .F(n813) );
  MUX U247 ( .IN0(n2556), .IN1(n2558), .SEL(n2557), .F(n2430) );
  XNOR U248 ( .A(n1042), .B(n1041), .Z(n1108) );
  XOR U249 ( .A(n1386), .B(n1301), .Z(n1302) );
  ANDN U250 ( .A(n596), .B(n576), .Z(n565) );
  XNOR U251 ( .A(n5029), .B(n5028), .Z(n5036) );
  MUX U252 ( .IN0(n3796), .IN1(n79), .SEL(n3797), .F(n3782) );
  IV U253 ( .A(n3798), .Z(n79) );
  MUX U254 ( .IN0(n4771), .IN1(n4773), .SEL(n4772), .F(n4767) );
  MUX U255 ( .IN0(n80), .IN1(n5104), .SEL(n5105), .F(n5090) );
  IV U256 ( .A(n5106), .Z(n80) );
  MUX U257 ( .IN0(n81), .IN1(n4726), .SEL(n4727), .F(n4717) );
  IV U258 ( .A(n4728), .Z(n81) );
  XNOR U259 ( .A(n4219), .B(n4218), .Z(n4234) );
  NANDN U260 ( .B(n5217), .A(n3025), .Z(n97) );
  MUX U261 ( .IN0(n4812), .IN1(n4814), .SEL(n4813), .F(n4793) );
  XNOR U262 ( .A(n4993), .B(n4992), .Z(n4998) );
  XNOR U263 ( .A(n4820), .B(n4819), .Z(n4835) );
  XNOR U264 ( .A(n3058), .B(n3057), .Z(n3092) );
  MUX U265 ( .IN0(n1905), .IN1(n82), .SEL(n1906), .F(n1799) );
  IV U266 ( .A(n1907), .Z(n82) );
  MUX U267 ( .IN0(n2200), .IN1(n83), .SEL(n2201), .F(n2081) );
  IV U268 ( .A(n2202), .Z(n83) );
  MUX U269 ( .IN0(n2392), .IN1(n2394), .SEL(n2393), .F(n2272) );
  MUX U270 ( .IN0(n2614), .IN1(n84), .SEL(n2615), .F(n2489) );
  IV U271 ( .A(n2616), .Z(n84) );
  MUX U272 ( .IN0(g_input[12]), .IN1(n5013), .SEL(g_input[31]), .F(n85) );
  IV U273 ( .A(n85), .Z(n1921) );
  MUX U274 ( .IN0(n2809), .IN1(n2811), .SEL(n2810), .F(n2684) );
  MUX U275 ( .IN0(g_input[20]), .IN1(n4539), .SEL(g_input[31]), .F(n86) );
  IV U276 ( .A(n86), .Z(n1169) );
  MUX U277 ( .IN0(n2778), .IN1(n87), .SEL(n2779), .F(n2648) );
  IV U278 ( .A(n2780), .Z(n87) );
  MUX U279 ( .IN0(g_input[15]), .IN1(n4977), .SEL(g_input[31]), .F(n88) );
  IV U280 ( .A(n88), .Z(n1618) );
  MUX U281 ( .IN0(g_input[23]), .IN1(n4488), .SEL(g_input[31]), .F(n89) );
  IV U282 ( .A(n89), .Z(n950) );
  MUX U283 ( .IN0(g_input[21]), .IN1(n4522), .SEL(g_input[31]), .F(n90) );
  IV U284 ( .A(n90), .Z(n1091) );
  MUX U285 ( .IN0(n791), .IN1(n793), .SEL(n792), .F(n735) );
  MUX U286 ( .IN0(n947), .IN1(n945), .SEL(n946), .F(n877) );
  MUX U287 ( .IN0(n1006), .IN1(n1004), .SEL(n1005), .F(n935) );
  MUX U288 ( .IN0(n1195), .IN1(n1193), .SEL(n1194), .F(n1115) );
  MUX U289 ( .IN0(n91), .IN1(n1329), .SEL(n1330), .F(n1245) );
  IV U290 ( .A(n1331), .Z(n91) );
  MUX U291 ( .IN0(n1960), .IN1(n1958), .SEL(n1959), .F(n1850) );
  MUX U292 ( .IN0(n92), .IN1(n2250), .SEL(n2251), .F(n2131) );
  IV U293 ( .A(n2252), .Z(n92) );
  MUX U294 ( .IN0(n670), .IN1(n668), .SEL(n669), .F(n628) );
  MUX U295 ( .IN0(n978), .IN1(n980), .SEL(n979), .F(n909) );
  MUX U296 ( .IN0(n93), .IN1(n1146), .SEL(n1147), .F(n1066) );
  IV U297 ( .A(n1148), .Z(n93) );
  XOR U298 ( .A(n348), .B(n1635), .Z(n1539) );
  MUX U299 ( .IN0(n1940), .IN1(n1942), .SEL(n1941), .F(n1833) );
  ANDN U300 ( .A(n565), .B(n547), .Z(n536) );
  AND U301 ( .A(n605), .B(n607), .Z(n574) );
  MUX U302 ( .IN0(n1357), .IN1(n1355), .SEL(n1356), .F(n1264) );
  MUX U303 ( .IN0(n5120), .IN1(n94), .SEL(n5121), .F(n5104) );
  IV U304 ( .A(n5122), .Z(n94) );
  MUX U305 ( .IN0(n4231), .IN1(n4233), .SEL(n4232), .F(n4211) );
  MUX U306 ( .IN0(n5208), .IN1(n5210), .SEL(n5209), .F(n5190) );
  XNOR U307 ( .A(n5017), .B(n5016), .Z(n5022) );
  MUX U308 ( .IN0(n95), .IN1(n3782), .SEL(n3783), .F(n3768) );
  IV U309 ( .A(n3784), .Z(n95) );
  MUX U310 ( .IN0(n96), .IN1(n4717), .SEL(n4718), .F(n4705) );
  IV U311 ( .A(n4719), .Z(n96) );
  MUX U312 ( .IN0(n5214), .IN1(n97), .SEL(n5215), .F(n5203) );
  MUX U313 ( .IN0(n4793), .IN1(n4795), .SEL(n4794), .F(n2979) );
  MUX U314 ( .IN0(n2128), .IN1(n98), .SEL(n2129), .F(n2020) );
  IV U315 ( .A(n2130), .Z(n98) );
  MUX U316 ( .IN0(n2096), .IN1(n2098), .SEL(n2097), .F(n1988) );
  MUX U317 ( .IN0(n2290), .IN1(n99), .SEL(n2291), .F(n2176) );
  IV U318 ( .A(n2292), .Z(n99) );
  MUX U319 ( .IN0(n2465), .IN1(n100), .SEL(n2466), .F(n2343) );
  IV U320 ( .A(n2467), .Z(n100) );
  MUX U321 ( .IN0(n2417), .IN1(n2419), .SEL(n2418), .F(n2297) );
  MUX U322 ( .IN0(n2730), .IN1(n2732), .SEL(n2731), .F(n2598) );
  MUX U323 ( .IN0(n2738), .IN1(n101), .SEL(n2739), .F(n2606) );
  IV U324 ( .A(n2740), .Z(n101) );
  MUX U325 ( .IN0(g_input[16]), .IN1(n4607), .SEL(g_input[31]), .F(n102) );
  IV U326 ( .A(n102), .Z(n1522) );
  MUX U327 ( .IN0(g_input[18]), .IN1(n4573), .SEL(g_input[31]), .F(n103) );
  IV U328 ( .A(n103), .Z(n1334) );
  MUX U329 ( .IN0(g_input[14]), .IN1(n4989), .SEL(g_input[31]), .F(n104) );
  IV U330 ( .A(n104), .Z(n1714) );
  MUX U331 ( .IN0(n2770), .IN1(n2772), .SEL(n2771), .F(n2640) );
  MUX U332 ( .IN0(g_input[13]), .IN1(n5001), .SEL(g_input[31]), .F(n105) );
  IV U333 ( .A(n105), .Z(n1815) );
  MUX U334 ( .IN0(n2917), .IN1(n106), .SEL(n2918), .F(n2778) );
  IV U335 ( .A(n2919), .Z(n106) );
  XNOR U336 ( .A(n3075), .B(n3074), .Z(n3854) );
  MUX U337 ( .IN0(n810), .IN1(n107), .SEL(n811), .F(n751) );
  IV U338 ( .A(n812), .Z(n107) );
  MUX U339 ( .IN0(n1044), .IN1(n1042), .SEL(n1043), .F(n974) );
  MUX U340 ( .IN0(n108), .IN1(n1086), .SEL(n1087), .F(n1012) );
  IV U341 ( .A(n1088), .Z(n108) );
  MUX U342 ( .IN0(n1746), .IN1(n1748), .SEL(n1747), .F(n1645) );
  MUX U343 ( .IN0(n1366), .IN1(n1364), .SEL(n1365), .F(n1275) );
  MUX U344 ( .IN0(n1414), .IN1(n1412), .SEL(n1413), .F(n1319) );
  MUX U345 ( .IN0(n1910), .IN1(n1908), .SEL(n1909), .F(n1802) );
  MUX U346 ( .IN0(n1871), .IN1(n1869), .SEL(n1870), .F(n1761) );
  MUX U347 ( .IN0(n1894), .IN1(n1892), .SEL(n1893), .F(n1786) );
  MUX U348 ( .IN0(n2325), .IN1(n2323), .SEL(n2324), .F(n2203) );
  MUX U349 ( .IN0(n2486), .IN1(n2484), .SEL(n2485), .F(n2362) );
  MUX U350 ( .IN0(n109), .IN1(n2492), .SEL(n2493), .F(n2370) );
  IV U351 ( .A(n2494), .Z(n109) );
  MUX U352 ( .IN0(n703), .IN1(n701), .SEL(n702), .F(n658) );
  MUX U353 ( .IN0(n714), .IN1(n712), .SEL(n713), .F(n668) );
  XNOR U354 ( .A(n867), .B(n866), .Z(n928) );
  MUX U355 ( .IN0(n110), .IN1(n1309), .SEL(n1310), .F(n1225) );
  IV U356 ( .A(n1311), .Z(n110) );
  XNOR U357 ( .A(n1387), .B(n1397), .Z(n1486) );
  MUX U358 ( .IN0(n1840), .IN1(n111), .SEL(n1841), .F(n1729) );
  IV U359 ( .A(n1842), .Z(n111) );
  XOR U360 ( .A(n578), .B(n555), .Z(n552) );
  MUX U361 ( .IN0(n652), .IN1(n654), .SEL(n653), .F(n112) );
  IV U362 ( .A(n112), .Z(n618) );
  AND U363 ( .A(n686), .B(n688), .Z(n646) );
  NOR U364 ( .A(n1353), .B(n1354), .Z(n1352) );
  NANDN U365 ( .B(n524), .A(n536), .Z(n504) );
  MUX U366 ( .IN0(n539), .IN1(\_MxM/Y0[29] ), .SEL(n540), .F(n516) );
  MUX U367 ( .IN0(n4138), .IN1(n4136), .SEL(n4137), .F(n4115) );
  MUX U368 ( .IN0(n5074), .IN1(n4951), .SEL(n4952), .F(n5060) );
  MUX U369 ( .IN0(n5134), .IN1(n5136), .SEL(n5135), .F(n5131) );
  MUX U370 ( .IN0(n113), .IN1(n4731), .SEL(n4732), .F(n4712) );
  IV U371 ( .A(n4733), .Z(n113) );
  MUX U372 ( .IN0(n114), .IN1(n5090), .SEL(n5091), .F(n5081) );
  IV U373 ( .A(n5092), .Z(n114) );
  NANDN U374 ( .B(n4958), .A(n3025), .Z(n135) );
  MUX U375 ( .IN0(n4179), .IN1(n4181), .SEL(n4180), .F(n4161) );
  XNOR U376 ( .A(n4199), .B(n4198), .Z(n4214) );
  MUX U377 ( .IN0(n115), .IN1(n5158), .SEL(n5159), .F(n3011) );
  IV U378 ( .A(n5160), .Z(n115) );
  XNOR U379 ( .A(n4981), .B(n4980), .Z(n4986) );
  XNOR U380 ( .A(n4710), .B(n4709), .Z(n4715) );
  MUX U381 ( .IN0(n1873), .IN1(n1875), .SEL(n1874), .F(n1765) );
  MUX U382 ( .IN0(n1988), .IN1(n1990), .SEL(n1989), .F(n1881) );
  MUX U383 ( .IN0(n2231), .IN1(n2233), .SEL(n2232), .F(n2112) );
  MUX U384 ( .IN0(n2239), .IN1(n116), .SEL(n2240), .F(n2120) );
  IV U385 ( .A(n2241), .Z(n116) );
  MUX U386 ( .IN0(n2183), .IN1(n2185), .SEL(n2184), .F(n2069) );
  MUX U387 ( .IN0(n2320), .IN1(n117), .SEL(n2321), .F(n2200) );
  IV U388 ( .A(n2322), .Z(n117) );
  MUX U389 ( .IN0(n2516), .IN1(n2518), .SEL(n2517), .F(n2392) );
  MUX U390 ( .IN0(n2524), .IN1(n118), .SEL(n2525), .F(n2400) );
  IV U391 ( .A(n2526), .Z(n118) );
  MUX U392 ( .IN0(n2663), .IN1(n2665), .SEL(n2664), .F(n2539) );
  MUX U393 ( .IN0(n2714), .IN1(n2716), .SEL(n2715), .F(n2582) );
  MUX U394 ( .IN0(n2722), .IN1(n119), .SEL(n2723), .F(n2590) );
  IV U395 ( .A(n2724), .Z(n119) );
  MUX U396 ( .IN0(n2838), .IN1(n2840), .SEL(n2839), .F(n2706) );
  MUX U397 ( .IN0(n2831), .IN1(n120), .SEL(n2832), .F(n2699) );
  IV U398 ( .A(n2833), .Z(n120) );
  MUX U399 ( .IN0(n2878), .IN1(n121), .SEL(n2879), .F(n2746) );
  IV U400 ( .A(n2880), .Z(n121) );
  MUX U401 ( .IN0(n2786), .IN1(n122), .SEL(n2787), .F(n2656) );
  IV U402 ( .A(n2788), .Z(n122) );
  MUX U403 ( .IN0(n4791), .IN1(n4789), .SEL(n4790), .F(n2975) );
  MUX U404 ( .IN0(n3060), .IN1(n3058), .SEL(n3059), .F(n2928) );
  XNOR U405 ( .A(n3050), .B(n3049), .Z(n3112) );
  MUX U406 ( .IN0(n718), .IN1(n720), .SEL(n719), .F(n674) );
  MUX U407 ( .IN0(n1321), .IN1(n1319), .SEL(n1320), .F(n1235) );
  MUX U408 ( .IN0(n123), .IN1(n1709), .SEL(n1710), .F(n1613) );
  IV U409 ( .A(n1711), .Z(n123) );
  MUX U410 ( .IN0(n1687), .IN1(n1685), .SEL(n1686), .F(n1589) );
  MUX U411 ( .IN0(n1978), .IN1(n1976), .SEL(n1977), .F(n1869) );
  MUX U412 ( .IN0(n2017), .IN1(n2015), .SEL(n2016), .F(n1908) );
  MUX U413 ( .IN0(n2057), .IN1(n2059), .SEL(n2058), .F(n124) );
  IV U414 ( .A(n124), .Z(n1947) );
  MUX U415 ( .IN0(n2228), .IN1(n2226), .SEL(n2227), .F(n2107) );
  MUX U416 ( .IN0(n2415), .IN1(n2413), .SEL(n2414), .F(n2293) );
  MUX U417 ( .IN0(n125), .IN1(n2617), .SEL(n2618), .F(n2492) );
  IV U418 ( .A(n2619), .Z(n125) );
  MUX U419 ( .IN0(n2611), .IN1(n2609), .SEL(n2610), .F(n2484) );
  MUX U420 ( .IN0(n2572), .IN1(n2570), .SEL(n2571), .F(n2445) );
  MUX U421 ( .IN0(n2554), .IN1(n2552), .SEL(n2553), .F(n126) );
  IV U422 ( .A(n126), .Z(n2424) );
  MUX U423 ( .IN0(n2653), .IN1(n2651), .SEL(n2652), .F(n2527) );
  XNOR U424 ( .A(n2944), .B(n2943), .Z(n3068) );
  MUX U425 ( .IN0(n630), .IN1(n628), .SEL(n629), .F(n584) );
  MUX U426 ( .IN0(n815), .IN1(n813), .SEL(n814), .F(n754) );
  MUX U427 ( .IN0(n986), .IN1(n984), .SEL(n985), .F(n915) );
  MUX U428 ( .IN0(n127), .IN1(n994), .SEL(n995), .F(n925) );
  IV U429 ( .A(n996), .Z(n127) );
  XNOR U430 ( .A(n1115), .B(n1114), .Z(n1186) );
  MUX U431 ( .IN0(n128), .IN1(n1404), .SEL(n1405), .F(n1309) );
  IV U432 ( .A(n1406), .Z(n128) );
  XNOR U433 ( .A(n1732), .B(n1641), .Z(n1642) );
  MUX U434 ( .IN0(n1944), .IN1(n129), .SEL(n1945), .F(n1840) );
  IV U435 ( .A(n1946), .Z(n129) );
  MUX U436 ( .IN0(n2430), .IN1(n2432), .SEL(n2431), .F(n2312) );
  ANDN U437 ( .A(n611), .B(n615), .Z(n614) );
  MUX U438 ( .IN0(n130), .IN1(n845), .SEL(n846), .F(n786) );
  IV U439 ( .A(n847), .Z(n130) );
  ANDN U440 ( .A(n1551), .B(n1553), .Z(n1442) );
  MUX U441 ( .IN0(n178), .IN1(n2192), .SEL(n2191), .F(n2075) );
  NANDN U442 ( .B(n597), .A(n598), .Z(n566) );
  AND U443 ( .A(n646), .B(n648), .Z(n605) );
  NANDN U444 ( .B(n766), .A(n767), .Z(n722) );
  AND U445 ( .A(n964), .B(n966), .Z(n896) );
  MUX U446 ( .IN0(n1457), .IN1(n131), .SEL(n1456), .F(n1355) );
  IV U447 ( .A(n1455), .Z(n131) );
  AND U448 ( .A(n512), .B(n513), .Z(n507) );
  MUX U449 ( .IN0(n568), .IN1(\_MxM/Y0[28] ), .SEL(n569), .F(n539) );
  MUX U450 ( .IN0(n3745), .IN1(n3743), .SEL(n3744), .F(n3701) );
  MUX U451 ( .IN0(n3810), .IN1(n3812), .SEL(n3811), .F(n3807) );
  MUX U452 ( .IN0(n132), .IN1(n5095), .SEL(n5096), .F(n5076) );
  IV U453 ( .A(n5097), .Z(n132) );
  MUX U454 ( .IN0(n133), .IN1(n3768), .SEL(n3769), .F(n3759) );
  IV U455 ( .A(n3770), .Z(n133) );
  MUX U456 ( .IN0(n134), .IN1(n4712), .SEL(n4713), .F(n4700) );
  IV U457 ( .A(n4714), .Z(n134) );
  MUX U458 ( .IN0(n4955), .IN1(n135), .SEL(n4956), .F(n4943) );
  MUX U459 ( .IN0(n136), .IN1(n5081), .SEL(n5082), .F(n5069) );
  IV U460 ( .A(n5083), .Z(n136) );
  XNOR U461 ( .A(n4175), .B(n4174), .Z(n4194) );
  MUX U462 ( .IN0(n1765), .IN1(n1767), .SEL(n1766), .F(n1664) );
  MUX U463 ( .IN0(n1799), .IN1(n137), .SEL(n1800), .F(n1698) );
  IV U464 ( .A(n1801), .Z(n137) );
  MUX U465 ( .IN0(n2247), .IN1(n138), .SEL(n2248), .F(n2128) );
  IV U466 ( .A(n2249), .Z(n138) );
  MUX U467 ( .IN0(n2359), .IN1(n139), .SEL(n2360), .F(n2239) );
  IV U468 ( .A(n2361), .Z(n139) );
  MUX U469 ( .IN0(n2335), .IN1(n2337), .SEL(n2336), .F(n2215) );
  MUX U470 ( .IN0(n2449), .IN1(n2451), .SEL(n2450), .F(n2327) );
  MUX U471 ( .IN0(n2442), .IN1(n140), .SEL(n2443), .F(n2320) );
  IV U472 ( .A(n2444), .Z(n140) );
  MUX U473 ( .IN0(n2598), .IN1(n2600), .SEL(n2599), .F(n2473) );
  MUX U474 ( .IN0(n2532), .IN1(n141), .SEL(n2533), .F(n2410) );
  IV U475 ( .A(n2534), .Z(n141) );
  MUX U476 ( .IN0(n2846), .IN1(n2848), .SEL(n2847), .F(n2714) );
  MUX U477 ( .IN0(n2854), .IN1(n142), .SEL(n2855), .F(n2722) );
  IV U478 ( .A(n2856), .Z(n142) );
  MUX U479 ( .IN0(n3011), .IN1(n143), .SEL(n3012), .F(n2870) );
  IV U480 ( .A(n3013), .Z(n143) );
  MUX U481 ( .IN0(n2972), .IN1(n144), .SEL(n2973), .F(n2831) );
  IV U482 ( .A(n2974), .Z(n144) );
  MUX U483 ( .IN0(n2909), .IN1(n2911), .SEL(n2910), .F(n2770) );
  MUX U484 ( .IN0(n4981), .IN1(n4807), .SEL(n4809), .F(n2998) );
  MUX U485 ( .IN0(n760), .IN1(n762), .SEL(n761), .F(n718) );
  MUX U486 ( .IN0(n1564), .IN1(n1562), .SEL(n1563), .F(n1466) );
  MUX U487 ( .IN0(n1607), .IN1(n1605), .SEL(n1606), .F(n1509) );
  MUX U488 ( .IN0(n145), .IN1(n1613), .SEL(n1614), .F(n1517) );
  IV U489 ( .A(n1615), .Z(n145) );
  MUX U490 ( .IN0(n2001), .IN1(n1999), .SEL(n2000), .F(n1892) );
  MUX U491 ( .IN0(n146), .IN1(n2023), .SEL(n2024), .F(n1916) );
  IV U492 ( .A(n2025), .Z(n146) );
  MUX U493 ( .IN0(n2125), .IN1(n2123), .SEL(n2124), .F(n2015) );
  MUX U494 ( .IN0(n2086), .IN1(n2084), .SEL(n2085), .F(n1976) );
  MUX U495 ( .IN0(n2181), .IN1(n2179), .SEL(n2180), .F(n2065) );
  MUX U496 ( .IN0(n2595), .IN1(n2593), .SEL(n2594), .F(n2468) );
  MUX U497 ( .IN0(n2529), .IN1(n2527), .SEL(n2528), .F(n2405) );
  MUX U498 ( .IN0(n2743), .IN1(n2741), .SEL(n2742), .F(n2609) );
  MUX U499 ( .IN0(n147), .IN1(n2749), .SEL(n2750), .F(n2617) );
  IV U500 ( .A(n2751), .Z(n147) );
  MUX U501 ( .IN0(n2704), .IN1(n2702), .SEL(n2703), .F(n2570) );
  MUX U502 ( .IN0(n2791), .IN1(n2789), .SEL(n2790), .F(n2659) );
  XNOR U503 ( .A(n2920), .B(n2919), .Z(n3043) );
  MUX U504 ( .IN0(n748), .IN1(n746), .SEL(n747), .F(n701) );
  XNOR U505 ( .A(n813), .B(n812), .Z(n870) );
  MUX U506 ( .IN0(n1054), .IN1(n1056), .SEL(n1055), .F(n984) );
  XNOR U507 ( .A(n1004), .B(n1003), .Z(n1069) );
  XNOR U508 ( .A(n1164), .B(n1163), .Z(n1238) );
  XNOR U509 ( .A(n1193), .B(n1192), .Z(n1268) );
  MUX U510 ( .IN0(n1645), .IN1(n1647), .SEL(n1646), .F(n1544) );
  MUX U511 ( .IN0(n148), .IN1(n1383), .SEL(n1384), .F(n1292) );
  IV U512 ( .A(n1385), .Z(n148) );
  XNOR U513 ( .A(n1733), .B(n1743), .Z(n1843) );
  XOR U514 ( .A(n2161), .B(n2057), .Z(n2058) );
  MUX U515 ( .IN0(n149), .IN1(n2354), .SEL(n2355), .F(n2234) );
  IV U516 ( .A(n2356), .Z(n149) );
  MUX U517 ( .IN0(n2426), .IN1(n150), .SEL(n2425), .F(n2310) );
  IV U518 ( .A(n2424), .Z(n150) );
  MUX U519 ( .IN0(n621), .IN1(n151), .SEL(n620), .F(n593) );
  IV U520 ( .A(n619), .Z(n151) );
  XNOR U521 ( .A(n784), .B(n783), .Z(n837) );
  AND U522 ( .A(n1174), .B(n1176), .Z(n1096) );
  MUX U523 ( .IN0(n152), .IN1(n1282), .SEL(n1283), .F(n1202) );
  IV U524 ( .A(n1284), .Z(n152) );
  MUX U525 ( .IN0(n2436), .IN1(n2438), .SEL(n2437), .F(n2314) );
  NANDN U526 ( .B(n638), .A(n639), .Z(n597) );
  ANDN U527 ( .A(n677), .B(n648), .Z(n637) );
  NANDN U528 ( .B(n825), .A(n826), .Z(n766) );
  NAND U529 ( .A(n1442), .B(n1441), .Z(n1353) );
  MUX U530 ( .IN0(n153), .IN1(n1965), .SEL(n1966), .F(n1857) );
  IV U531 ( .A(n1967), .Z(n153) );
  ANDN U532 ( .A(n1105), .B(n1106), .Z(n1031) );
  MUX U533 ( .IN0(\_MxM/Y0[3] ), .IN1(n2627), .SEL(n2628), .F(n2504) );
  MUX U534 ( .IN0(n504), .IN1(n506), .SEL(n505), .F(n154) );
  IV U535 ( .A(n154), .Z(n503) );
  MUX U536 ( .IN0(n599), .IN1(\_MxM/Y0[27] ), .SEL(n600), .F(n568) );
  MUX U537 ( .IN0(n768), .IN1(\_MxM/Y0[23] ), .SEL(n769), .F(n724) );
  MUX U538 ( .IN0(n1025), .IN1(\_MxM/Y0[19] ), .SEL(n1026), .F(n958) );
  MUX U539 ( .IN0(n1342), .IN1(\_MxM/Y0[15] ), .SEL(n1343), .F(n1258) );
  MUX U540 ( .IN0(n1722), .IN1(\_MxM/Y0[11] ), .SEL(n1723), .F(n1626) );
  MUX U541 ( .IN0(n2144), .IN1(\_MxM/Y0[7] ), .SEL(n2145), .F(n2036) );
  MUX U542 ( .IN0(n4614), .IN1(n4168), .SEL(n4169), .F(n4597) );
  MUX U543 ( .IN0(n155), .IN1(n4145), .SEL(n3710), .F(n4124) );
  IV U544 ( .A(n3708), .Z(n155) );
  MUX U545 ( .IN0(n3584), .IN1(n3582), .SEL(n3583), .F(n3538) );
  MUX U546 ( .IN0(n4305), .IN1(n4303), .SEL(n4304), .F(n4279) );
  XNOR U547 ( .A(n4880), .B(n4879), .Z(n4895) );
  MUX U548 ( .IN0(n4337), .IN1(n4339), .SEL(n4338), .F(n4334) );
  MUX U549 ( .IN0(n156), .IN1(n3773), .SEL(n3774), .F(n3752) );
  IV U550 ( .A(n3775), .Z(n156) );
  NANDN U551 ( .B(n1638), .A(n3025), .Z(n188) );
  MUX U552 ( .IN0(n157), .IN1(n5149), .SEL(n5150), .F(n3003) );
  IV U553 ( .A(n5151), .Z(n157) );
  MUX U554 ( .IN0(n4800), .IN1(n4802), .SEL(n4801), .F(n2987) );
  MUX U555 ( .IN0(n3863), .IN1(n3861), .SEL(n3862), .F(n3075) );
  MUX U556 ( .IN0(n1881), .IN1(n1883), .SEL(n1882), .F(n1773) );
  MUX U557 ( .IN0(n2004), .IN1(n2006), .SEL(n2005), .F(n1897) );
  MUX U558 ( .IN0(n2088), .IN1(n2090), .SEL(n2089), .F(n1980) );
  MUX U559 ( .IN0(n2081), .IN1(n158), .SEL(n2082), .F(n1973) );
  IV U560 ( .A(n2083), .Z(n158) );
  MUX U561 ( .IN0(n2343), .IN1(n159), .SEL(n2344), .F(n2223) );
  IV U562 ( .A(n2345), .Z(n159) );
  MUX U563 ( .IN0(n2457), .IN1(n2459), .SEL(n2458), .F(n2335) );
  MUX U564 ( .IN0(n2473), .IN1(n2475), .SEL(n2474), .F(n2351) );
  MUX U565 ( .IN0(n2606), .IN1(n160), .SEL(n2607), .F(n2481) );
  IV U566 ( .A(n2608), .Z(n160) );
  MUX U567 ( .IN0(n2567), .IN1(n161), .SEL(n2568), .F(n2442) );
  IV U568 ( .A(n2569), .Z(n161) );
  MUX U569 ( .IN0(n2656), .IN1(n162), .SEL(n2657), .F(n2532) );
  IV U570 ( .A(n2658), .Z(n162) );
  MUX U571 ( .IN0(n2746), .IN1(n163), .SEL(n2747), .F(n2614) );
  IV U572 ( .A(n2748), .Z(n163) );
  MUX U573 ( .IN0(n2706), .IN1(n2708), .SEL(n2707), .F(n2574) );
  MUX U574 ( .IN0(g_input[8]), .IN1(n5068), .SEL(g_input[31]), .F(n164) );
  IV U575 ( .A(n164), .Z(n2375) );
  MUX U576 ( .IN0(n2995), .IN1(n165), .SEL(n2996), .F(n2854) );
  IV U577 ( .A(n2997), .Z(n165) );
  MUX U578 ( .IN0(n2948), .IN1(n2950), .SEL(n2949), .F(n2809) );
  MUX U579 ( .IN0(n869), .IN1(n867), .SEL(n868), .F(n805) );
  MUX U580 ( .IN0(n1763), .IN1(n1761), .SEL(n1762), .F(n1660) );
  MUX U581 ( .IN0(n1804), .IN1(n1802), .SEL(n1803), .F(n1701) );
  MUX U582 ( .IN0(n1735), .IN1(n1733), .SEL(n1734), .F(n1641) );
  MUX U583 ( .IN0(n166), .IN1(n1916), .SEL(n1917), .F(n1810) );
  IV U584 ( .A(n1918), .Z(n166) );
  MUX U585 ( .IN0(n2109), .IN1(n2107), .SEL(n2108), .F(n1999) );
  MUX U586 ( .IN0(n2205), .IN1(n2203), .SEL(n2204), .F(n2084) );
  MUX U587 ( .IN0(n2244), .IN1(n2242), .SEL(n2243), .F(n2123) );
  MUX U588 ( .IN0(n2164), .IN1(n2162), .SEL(n2163), .F(n2057) );
  MUX U589 ( .IN0(n2295), .IN1(n2293), .SEL(n2294), .F(n2179) );
  MUX U590 ( .IN0(n167), .IN1(n2370), .SEL(n2371), .F(n2250) );
  IV U591 ( .A(n2372), .Z(n167) );
  MUX U592 ( .IN0(n2673), .IN1(n2671), .SEL(n2672), .F(n2552) );
  MUX U593 ( .IN0(n2727), .IN1(n2725), .SEL(n2726), .F(n2593) );
  MUX U594 ( .IN0(n2836), .IN1(n2834), .SEL(n2835), .F(n2702) );
  MUX U595 ( .IN0(n2875), .IN1(n2873), .SEL(n2874), .F(n2741) );
  MUX U596 ( .IN0(n168), .IN1(n2881), .SEL(n2882), .F(n2749) );
  IV U597 ( .A(n2883), .Z(n168) );
  MUX U598 ( .IN0(n2783), .IN1(n2781), .SEL(n2782), .F(n2651) );
  MUX U599 ( .IN0(n2930), .IN1(n2928), .SEL(n2929), .F(n2789) );
  MUX U600 ( .IN0(n634), .IN1(n636), .SEL(n635), .F(n590) );
  MUX U601 ( .IN0(n756), .IN1(n754), .SEL(n755), .F(n712) );
  XNOR U602 ( .A(n945), .B(n944), .Z(n1007) );
  XNOR U603 ( .A(n1156), .B(n1155), .Z(n1228) );
  XNOR U604 ( .A(n1245), .B(n1244), .Z(n1322) );
  XNOR U605 ( .A(n1275), .B(n1274), .Z(n1359) );
  MUX U606 ( .IN0(n169), .IN1(n1501), .SEL(n1502), .F(n1404) );
  IV U607 ( .A(n1503), .Z(n169) );
  XNOR U608 ( .A(n1493), .B(n1492), .Z(n1582) );
  MUX U609 ( .IN0(n2048), .IN1(n170), .SEL(n2049), .F(n1944) );
  IV U610 ( .A(n2050), .Z(n170) );
  MUX U611 ( .IN0(n171), .IN1(n2115), .SEL(n2116), .F(n2007) );
  IV U612 ( .A(n2117), .Z(n171) );
  MUX U613 ( .IN0(n172), .IN1(n2338), .SEL(n2339), .F(n2218) );
  IV U614 ( .A(n2340), .Z(n172) );
  MUX U615 ( .IN0(n173), .IN1(n2601), .SEL(n2602), .F(n2476) );
  IV U616 ( .A(n2603), .Z(n173) );
  MUX U617 ( .IN0(n174), .IN1(n2519), .SEL(n2520), .F(n2395) );
  IV U618 ( .A(n2521), .Z(n174) );
  MUX U619 ( .IN0(n175), .IN1(n581), .SEL(n580), .F(n555) );
  IV U620 ( .A(n579), .Z(n175) );
  AND U621 ( .A(n617), .B(n618), .Z(n613) );
  MUX U622 ( .IN0(n904), .IN1(n902), .SEL(n903), .F(n842) );
  MUX U623 ( .IN0(n176), .IN1(n1049), .SEL(n1050), .F(n981) );
  IV U624 ( .A(n1051), .Z(n176) );
  AND U625 ( .A(n1255), .B(n1257), .Z(n1174) );
  MUX U626 ( .IN0(n1544), .IN1(n1546), .SEL(n1545), .F(n1453) );
  MUX U627 ( .IN0(n177), .IN1(n1768), .SEL(n1769), .F(n1667) );
  IV U628 ( .A(n1770), .Z(n177) );
  ANDN U629 ( .A(n1752), .B(n1754), .Z(n1651) );
  AND U630 ( .A(n2033), .B(n2035), .Z(n1926) );
  MUX U631 ( .IN0(n2316), .IN1(n2314), .SEL(n2315), .F(n178) );
  IV U632 ( .A(n178), .Z(n2190) );
  NANDN U633 ( .B(n678), .A(n679), .Z(n638) );
  MUX U634 ( .IN0(n765), .IN1(n179), .SEL(n764), .F(n721) );
  IV U635 ( .A(n763), .Z(n179) );
  AND U636 ( .A(n833), .B(n835), .Z(n822) );
  NANDN U637 ( .B(n888), .A(n889), .Z(n825) );
  MUX U638 ( .IN0(n180), .IN1(n1548), .SEL(n1549), .F(n1455) );
  IV U639 ( .A(n1550), .Z(n180) );
  MUX U640 ( .IN0(n181), .IN1(n2072), .SEL(n2073), .F(n1965) );
  IV U641 ( .A(n2074), .Z(n181) );
  MUX U642 ( .IN0(n2544), .IN1(n208), .SEL(n2543), .F(n182) );
  IV U643 ( .A(n182), .Z(n2420) );
  AND U644 ( .A(n545), .B(n547), .Z(n522) );
  ANDN U645 ( .A(n1183), .B(n1184), .Z(n1105) );
  NAND U646 ( .A(n493), .B(n495), .Z(n492) );
  MUX U647 ( .IN0(n640), .IN1(\_MxM/Y0[26] ), .SEL(n641), .F(n599) );
  MUX U648 ( .IN0(n827), .IN1(\_MxM/Y0[22] ), .SEL(n828), .F(n768) );
  MUX U649 ( .IN0(n1099), .IN1(\_MxM/Y0[18] ), .SEL(n1100), .F(n1025) );
  MUX U650 ( .IN0(n1433), .IN1(\_MxM/Y0[14] ), .SEL(n1434), .F(n1342) );
  MUX U651 ( .IN0(n1823), .IN1(\_MxM/Y0[10] ), .SEL(n1824), .F(n1722) );
  MUX U652 ( .IN0(n2263), .IN1(\_MxM/Y0[6] ), .SEL(n2264), .F(n2144) );
  MUX U653 ( .IN0(n4159), .IN1(n4157), .SEL(n4158), .F(n4136) );
  MUX U654 ( .IN0(n3734), .IN1(n3732), .SEL(n3733), .F(n183) );
  IV U655 ( .A(n183), .Z(n3690) );
  MUX U656 ( .IN0(n3657), .IN1(n3655), .SEL(n3656), .F(n3609) );
  MUX U657 ( .IN0(n4580), .IN1(n4126), .SEL(n4127), .F(n4563) );
  MUX U658 ( .IN0(n184), .IN1(n4061), .SEL(n3528), .F(n4040) );
  IV U659 ( .A(n3526), .Z(n184) );
  MUX U660 ( .IN0(n4710), .IN1(n4330), .SEL(n4331), .F(n4698) );
  MUX U661 ( .IN0(n4948), .IN1(n4946), .SEL(n4947), .F(n4926) );
  XNOR U662 ( .A(n4279), .B(n4278), .Z(n4296) );
  MUX U663 ( .IN0(n185), .IN1(n3977), .SEL(n3346), .F(n3956) );
  IV U664 ( .A(n3344), .Z(n185) );
  MUX U665 ( .IN0(n4656), .IN1(n4246), .SEL(n4248), .F(n4644) );
  MUX U666 ( .IN0(n5218), .IN1(n5220), .SEL(n5219), .F(n5214) );
  MUX U667 ( .IN0(n4862), .IN1(n4860), .SEL(n4861), .F(n4840) );
  MUX U668 ( .IN0(n186), .IN1(n5174), .SEL(n5175), .F(n5149) );
  IV U669 ( .A(n5176), .Z(n186) );
  MUX U670 ( .IN0(n187), .IN1(n5076), .SEL(n5077), .F(n5062) );
  IV U671 ( .A(n5078), .Z(n187) );
  MUX U672 ( .IN0(n3828), .IN1(n188), .SEL(n3829), .F(n3714) );
  MUX U673 ( .IN0(n189), .IN1(n3894), .SEL(n3173), .F(n3873) );
  IV U674 ( .A(n3171), .Z(n189) );
  MUX U675 ( .IN0(n1897), .IN1(n1899), .SEL(n1898), .F(n1791) );
  MUX U676 ( .IN0(n2870), .IN1(n190), .SEL(n2871), .F(n2738) );
  IV U677 ( .A(n2872), .Z(n190) );
  MUX U678 ( .IN0(g_input[7]), .IN1(n5157), .SEL(g_input[31]), .F(n191) );
  IV U679 ( .A(n191), .Z(n2497) );
  MUX U680 ( .IN0(g_input[11]), .IN1(n5025), .SEL(g_input[31]), .F(n192) );
  IV U681 ( .A(n192), .Z(n2028) );
  MUX U682 ( .IN0(n2932), .IN1(n2934), .SEL(n2933), .F(n2793) );
  MUX U683 ( .IN0(n2925), .IN1(n193), .SEL(n2926), .F(n2786) );
  IV U684 ( .A(n2927), .Z(n193) );
  MUX U685 ( .IN0(n3052), .IN1(n3050), .SEL(n3051), .F(n2920) );
  MUX U686 ( .IN0(n819), .IN1(n821), .SEL(n820), .F(n760) );
  MUX U687 ( .IN0(n1237), .IN1(n1235), .SEL(n1236), .F(n1156) );
  MUX U688 ( .IN0(n1389), .IN1(n1387), .SEL(n1388), .F(n1301) );
  MUX U689 ( .IN0(n1788), .IN1(n1786), .SEL(n1787), .F(n1685) );
  MUX U690 ( .IN0(n2348), .IN1(n2346), .SEL(n2347), .F(n2226) );
  MUX U691 ( .IN0(n2447), .IN1(n2445), .SEL(n2446), .F(n2323) );
  MUX U692 ( .IN0(n2661), .IN1(n2659), .SEL(n2660), .F(n2535) );
  MUX U693 ( .IN0(n2859), .IN1(n2857), .SEL(n2858), .F(n2725) );
  MUX U694 ( .IN0(n194), .IN1(n3022), .SEL(n3023), .F(n2881) );
  IV U695 ( .A(n3024), .Z(n194) );
  MUX U696 ( .IN0(n3016), .IN1(n3014), .SEL(n3015), .F(n2873) );
  MUX U697 ( .IN0(n2977), .IN1(n2975), .SEL(n2976), .F(n2834) );
  XNOR U698 ( .A(n877), .B(n876), .Z(n938) );
  XNOR U699 ( .A(n935), .B(n934), .Z(n997) );
  XNOR U700 ( .A(n1086), .B(n1085), .Z(n1159) );
  MUX U701 ( .IN0(n1215), .IN1(n195), .SEL(n1216), .F(n1136) );
  IV U702 ( .A(n1217), .Z(n195) );
  XNOR U703 ( .A(n1329), .B(n1328), .Z(n1415) );
  XNOR U704 ( .A(n1364), .B(n1363), .Z(n1459) );
  XNOR U705 ( .A(n1509), .B(n1508), .Z(n1600) );
  MUX U706 ( .IN0(n196), .IN1(n1693), .SEL(n1694), .F(n1597) );
  IV U707 ( .A(n1695), .Z(n196) );
  XNOR U708 ( .A(n1613), .B(n1612), .Z(n1704) );
  XNOR U709 ( .A(n1660), .B(n1659), .Z(n1756) );
  MUX U710 ( .IN0(n197), .IN1(n1884), .SEL(n1885), .F(n1776) );
  IV U711 ( .A(n1886), .Z(n197) );
  XNOR U712 ( .A(n1908), .B(n1907), .Z(n2010) );
  XNOR U713 ( .A(n1916), .B(n1915), .Z(n2018) );
  XNOR U714 ( .A(n2065), .B(n2064), .Z(n2174) );
  XNOR U715 ( .A(n2242), .B(n2241), .Z(n2357) );
  XNOR U716 ( .A(n2250), .B(n2249), .Z(n2365) );
  XNOR U717 ( .A(n2285), .B(n2284), .Z(n2398) );
  MUX U718 ( .IN0(n198), .IN1(n2585), .SEL(n2586), .F(n2460) );
  IV U719 ( .A(n2587), .Z(n198) );
  XNOR U720 ( .A(n2671), .B(n2681), .Z(n2800) );
  MUX U721 ( .IN0(n199), .IN1(n2773), .SEL(n2774), .F(n2643) );
  IV U722 ( .A(n2775), .Z(n199) );
  XNOR U723 ( .A(n584), .B(n581), .Z(n622) );
  MUX U724 ( .IN0(n660), .IN1(n658), .SEL(n659), .F(n611) );
  MUX U725 ( .IN0(n200), .IN1(n696), .SEL(n697), .F(n655) );
  IV U726 ( .A(n698), .Z(n200) );
  AND U727 ( .A(n915), .B(n917), .Z(n848) );
  MUX U728 ( .IN0(n201), .IN1(n1124), .SEL(n1125), .F(n1049) );
  IV U729 ( .A(n1126), .Z(n201) );
  MUX U730 ( .IN0(n1540), .IN1(n348), .SEL(n1539), .F(n1452) );
  AND U731 ( .A(n1623), .B(n1625), .Z(n1527) );
  ANDN U732 ( .A(n1860), .B(n1862), .Z(n1752) );
  MUX U733 ( .IN0(n202), .IN1(n1983), .SEL(n1984), .F(n1876) );
  IV U734 ( .A(n1985), .Z(n202) );
  AND U735 ( .A(n2260), .B(n2262), .Z(n2141) );
  MUX U736 ( .IN0(n203), .IN1(n2452), .SEL(n2453), .F(n2330) );
  IV U737 ( .A(n2454), .Z(n203) );
  MUX U738 ( .IN0(n204), .IN1(n2563), .SEL(n2562), .F(n2436) );
  IV U739 ( .A(n2561), .Z(n204) );
  NANDN U740 ( .B(n566), .A(n567), .Z(n537) );
  ANDN U741 ( .A(n721), .B(n688), .Z(n677) );
  NANDN U742 ( .B(n722), .A(n723), .Z(n678) );
  MUX U743 ( .IN0(n844), .IN1(n842), .SEL(n843), .F(n205) );
  IV U744 ( .A(n205), .Z(n782) );
  OR U745 ( .A(n1023), .B(n1024), .Z(n956) );
  MUX U746 ( .IN0(n206), .IN1(n1648), .SEL(n1649), .F(n1548) );
  IV U747 ( .A(n1650), .Z(n206) );
  MUX U748 ( .IN0(n207), .IN1(n2186), .SEL(n2187), .F(n2072) );
  IV U749 ( .A(n2188), .Z(n207) );
  MUX U750 ( .IN0(n2668), .IN1(n241), .SEL(n2667), .F(n208) );
  IV U751 ( .A(n208), .Z(n2542) );
  AND U752 ( .A(n822), .B(n824), .Z(n730) );
  MUX U753 ( .IN0(n209), .IN1(n1264), .SEL(n1265), .F(n1183) );
  IV U754 ( .A(n1266), .Z(n209) );
  ANDN U755 ( .A(n497), .B(n498), .Z(n489) );
  MUX U756 ( .IN0(n680), .IN1(\_MxM/Y0[25] ), .SEL(n681), .F(n640) );
  MUX U757 ( .IN0(n890), .IN1(\_MxM/Y0[21] ), .SEL(n891), .F(n827) );
  MUX U758 ( .IN0(n1177), .IN1(\_MxM/Y0[17] ), .SEL(n1178), .F(n1099) );
  MUX U759 ( .IN0(n1530), .IN1(\_MxM/Y0[13] ), .SEL(n1531), .F(n1433) );
  MUX U760 ( .IN0(n1929), .IN1(\_MxM/Y0[9] ), .SEL(n1930), .F(n1823) );
  MUX U761 ( .IN0(n2383), .IN1(\_MxM/Y0[5] ), .SEL(n2384), .F(n2263) );
  MUX U762 ( .IN0(n516), .IN1(\_MxM/Y0[30] ), .SEL(n517), .F(n482) );
  MUX U763 ( .IN0(n3065), .IN1(n3746), .SEL(n3066), .F(n210) );
  IV U764 ( .A(n210), .Z(n3704) );
  MUX U765 ( .IN0(n211), .IN1(n3690), .SEL(n3691), .F(n3644) );
  IV U766 ( .A(n3692), .Z(n211) );
  MUX U767 ( .IN0(n4096), .IN1(n4094), .SEL(n4095), .F(n4073) );
  MUX U768 ( .IN0(n3611), .IN1(n3609), .SEL(n3610), .F(n3563) );
  MUX U769 ( .IN0(n212), .IN1(n3508), .SEL(n3509), .F(n3462) );
  IV U770 ( .A(n3510), .Z(n212) );
  MUX U771 ( .IN0(n4512), .IN1(n4042), .SEL(n4043), .F(n4495) );
  MUX U772 ( .IN0(n3402), .IN1(n3400), .SEL(n3401), .F(n3356) );
  MUX U773 ( .IN0(n4012), .IN1(n4010), .SEL(n4011), .F(n3989) );
  MUX U774 ( .IN0(n3429), .IN1(n3427), .SEL(n3428), .F(n3381) );
  MUX U775 ( .IN0(n4796), .IN1(n4949), .SEL(n4797), .F(n213) );
  IV U776 ( .A(n213), .Z(n4929) );
  MUX U777 ( .IN0(n214), .IN1(n3326), .SEL(n3327), .F(n3281) );
  IV U778 ( .A(n3328), .Z(n214) );
  MUX U779 ( .IN0(n4444), .IN1(n3958), .SEL(n3959), .F(n4428) );
  MUX U780 ( .IN0(n5029), .IN1(n4887), .SEL(n4889), .F(n5017) );
  MUX U781 ( .IN0(n3226), .IN1(n3224), .SEL(n3225), .F(n3182) );
  MUX U782 ( .IN0(n4767), .IN1(n215), .SEL(n4768), .F(n4756) );
  IV U783 ( .A(n4770), .Z(n215) );
  MUX U784 ( .IN0(n3928), .IN1(n3926), .SEL(n3927), .F(n3906) );
  MUX U785 ( .IN0(n3251), .IN1(n3249), .SEL(n3250), .F(n3206) );
  MUX U786 ( .IN0(n4959), .IN1(n4961), .SEL(n4960), .F(n4955) );
  MUX U787 ( .IN0(n4221), .IN1(n4219), .SEL(n4220), .F(n4199) );
  NANDN U788 ( .B(n5238), .A(n3025), .Z(n250) );
  MUX U789 ( .IN0(n216), .IN1(n3153), .SEL(n3154), .F(n3109) );
  IV U790 ( .A(n3155), .Z(n216) );
  MUX U791 ( .IN0(n2327), .IN1(n2329), .SEL(n2328), .F(n2207) );
  MUX U792 ( .IN0(n2699), .IN1(n217), .SEL(n2700), .F(n2567) );
  IV U793 ( .A(n2701), .Z(n217) );
  MUX U794 ( .IN0(g_input[10]), .IN1(n5039), .SEL(g_input[31]), .F(n218) );
  IV U795 ( .A(n218), .Z(n2136) );
  MUX U796 ( .IN0(g_input[6]), .IN1(n5168), .SEL(g_input[31]), .F(n219) );
  IV U797 ( .A(n219), .Z(n2622) );
  MUX U798 ( .IN0(g_input[5]), .IN1(n5184), .SEL(g_input[31]), .F(n220) );
  IV U799 ( .A(n220), .Z(n2754) );
  MUX U800 ( .IN0(n4378), .IN1(n3875), .SEL(n3876), .F(n4358) );
  XNOR U801 ( .A(n4614), .B(n4612), .Z(n4619) );
  MUX U802 ( .IN0(n3077), .IN1(n3075), .SEL(n3076), .F(n2944) );
  MUX U803 ( .IN0(n751), .IN1(n221), .SEL(n752), .F(n709) );
  IV U804 ( .A(n753), .Z(n221) );
  MUX U805 ( .IN0(n290), .IN1(n1219), .SEL(n1218), .F(n1130) );
  MUX U806 ( .IN0(n1591), .IN1(n1589), .SEL(n1590), .F(n1493) );
  MUX U807 ( .IN0(n222), .IN1(n1810), .SEL(n1811), .F(n1709) );
  IV U808 ( .A(n1812), .Z(n222) );
  MUX U809 ( .IN0(n2470), .IN1(n2468), .SEL(n2469), .F(n2346) );
  MUX U810 ( .IN0(n2407), .IN1(n2405), .SEL(n2406), .F(n2285) );
  MUX U811 ( .IN0(n2537), .IN1(n2535), .SEL(n2536), .F(n2413) );
  MUX U812 ( .IN0(n3000), .IN1(n2998), .SEL(n2999), .F(n2857) );
  MUX U813 ( .IN0(n2922), .IN1(n2920), .SEL(n2921), .F(n2781) );
  XNOR U814 ( .A(n3014), .B(n3013), .Z(n5154) );
  XNOR U815 ( .A(n2975), .B(n2974), .Z(n4784) );
  XNOR U816 ( .A(n2928), .B(n2927), .Z(n3053) );
  MUX U817 ( .IN0(n976), .IN1(n974), .SEL(n975), .F(n902) );
  MUX U818 ( .IN0(n807), .IN1(n805), .SEL(n806), .F(n746) );
  XNOR U819 ( .A(n1012), .B(n1011), .Z(n1079) );
  MUX U820 ( .IN0(n1138), .IN1(n223), .SEL(n1137), .F(n1054) );
  IV U821 ( .A(n1136), .Z(n223) );
  XNOR U822 ( .A(n1076), .B(n1075), .Z(n1149) );
  XNOR U823 ( .A(n1412), .B(n1411), .Z(n1504) );
  XNOR U824 ( .A(n1420), .B(n1419), .Z(n1512) );
  XNOR U825 ( .A(n1466), .B(n1465), .Z(n1555) );
  MUX U826 ( .IN0(n224), .IN1(n1675), .SEL(n1676), .F(n1579) );
  IV U827 ( .A(n1677), .Z(n224) );
  XNOR U828 ( .A(n1701), .B(n1700), .Z(n1797) );
  MUX U829 ( .IN0(n225), .IN1(n1900), .SEL(n1901), .F(n1794) );
  IV U830 ( .A(n1902), .Z(n225) );
  XNOR U831 ( .A(n1869), .B(n1868), .Z(n1971) );
  XNOR U832 ( .A(n1958), .B(n1957), .Z(n2060) );
  XNOR U833 ( .A(n1999), .B(n1998), .Z(n2102) );
  MUX U834 ( .IN0(n226), .IN1(n2218), .SEL(n2219), .F(n2099) );
  IV U835 ( .A(n2220), .Z(n226) );
  MUX U836 ( .IN0(n227), .IN1(n2275), .SEL(n2276), .F(n2158) );
  IV U837 ( .A(n2277), .Z(n227) );
  XNOR U838 ( .A(n2323), .B(n2322), .Z(n2440) );
  XNOR U839 ( .A(n2362), .B(n2361), .Z(n2479) );
  XNOR U840 ( .A(n2370), .B(n2369), .Z(n2487) );
  XNOR U841 ( .A(n2670), .B(n2552), .Z(n2553) );
  MUX U842 ( .IN0(n228), .IN1(n2849), .SEL(n2850), .F(n2717) );
  IV U843 ( .A(n2851), .Z(n228) );
  MUX U844 ( .IN0(n2867), .IN1(n298), .SEL(n2866), .F(n229) );
  IV U845 ( .A(n229), .Z(n2733) );
  MUX U846 ( .IN0(n230), .IN1(n2825), .SEL(n2826), .F(n2692) );
  IV U847 ( .A(n2827), .Z(n230) );
  MUX U848 ( .IN0(n590), .IN1(n592), .SEL(n591), .F(n560) );
  XNOR U849 ( .A(n628), .B(n627), .Z(n661) );
  MUX U850 ( .IN0(n231), .IN1(n738), .SEL(n739), .F(n696) );
  IV U851 ( .A(n740), .Z(n231) );
  MUX U852 ( .IN0(n232), .IN1(n912), .SEL(n913), .F(n845) );
  IV U853 ( .A(n914), .Z(n232) );
  MUX U854 ( .IN0(n233), .IN1(n1202), .SEL(n1203), .F(n1124) );
  IV U855 ( .A(n1204), .Z(n233) );
  AND U856 ( .A(n1430), .B(n1432), .Z(n1339) );
  MUX U857 ( .IN0(n234), .IN1(n1569), .SEL(n1570), .F(n1473) );
  IV U858 ( .A(n1571), .Z(n234) );
  XNOR U859 ( .A(n1451), .B(n1452), .Z(n1448) );
  AND U860 ( .A(n1651), .B(n1653), .Z(n1551) );
  AND U861 ( .A(n1820), .B(n1822), .Z(n1719) );
  MUX U862 ( .IN0(n235), .IN1(n2091), .SEL(n2092), .F(n1983) );
  IV U863 ( .A(n2093), .Z(n235) );
  AND U864 ( .A(n2380), .B(n2382), .Z(n2260) );
  MUX U865 ( .IN0(n236), .IN1(n2577), .SEL(n2578), .F(n2452) );
  IV U866 ( .A(n2579), .Z(n236) );
  MUX U867 ( .IN0(n237), .IN1(n2689), .SEL(n2690), .F(n2561) );
  IV U868 ( .A(n2691), .Z(n237) );
  NAND U869 ( .A(n555), .B(n554), .Z(n549) );
  XNOR U870 ( .A(n593), .B(n618), .Z(n609) );
  ANDN U871 ( .A(n730), .B(n731), .Z(n686) );
  AND U872 ( .A(n778), .B(n779), .Z(n777) );
  ANDN U873 ( .A(n1031), .B(n1032), .Z(n964) );
  NAND U874 ( .A(n1096), .B(n1098), .Z(n1023) );
  MUX U875 ( .IN0(n238), .IN1(n1857), .SEL(n1858), .F(n1749) );
  IV U876 ( .A(n1859), .Z(n238) );
  MUX U877 ( .IN0(n239), .IN1(n2075), .SEL(n2076), .F(n1968) );
  IV U878 ( .A(n2077), .Z(n239) );
  MUX U879 ( .IN0(n240), .IN1(n2300), .SEL(n2301), .F(n2186) );
  IV U880 ( .A(n2302), .Z(n240) );
  MUX U881 ( .IN0(n2798), .IN1(n272), .SEL(n2797), .F(n241) );
  IV U882 ( .A(n241), .Z(n2666) );
  XNOR U883 ( .A(n566), .B(n571), .Z(n567) );
  XNOR U884 ( .A(n678), .B(n683), .Z(n679) );
  XNOR U885 ( .A(n825), .B(n830), .Z(n826) );
  XOR U886 ( .A(n1264), .B(n1353), .Z(n1348) );
  XNOR U887 ( .A(n2937), .B(n2936), .Z(n2766) );
  MUX U888 ( .IN0(n724), .IN1(\_MxM/Y0[24] ), .SEL(n725), .F(n680) );
  MUX U889 ( .IN0(n958), .IN1(\_MxM/Y0[20] ), .SEL(n959), .F(n890) );
  MUX U890 ( .IN0(n1258), .IN1(\_MxM/Y0[16] ), .SEL(n1259), .F(n1177) );
  MUX U891 ( .IN0(n1626), .IN1(\_MxM/Y0[12] ), .SEL(n1627), .F(n1530) );
  MUX U892 ( .IN0(n2036), .IN1(\_MxM/Y0[8] ), .SEL(n2037), .F(n1929) );
  MUX U893 ( .IN0(\_MxM/Y0[4] ), .IN1(n2504), .SEL(n2505), .F(n2383) );
  XNOR U894 ( .A(n516), .B(n520), .Z(n518) );
  MUX U895 ( .IN0(n3676), .IN1(n3674), .SEL(n3675), .F(n3628) );
  MUX U896 ( .IN0(n4597), .IN1(n4147), .SEL(n4148), .F(n4580) );
  MUX U897 ( .IN0(n242), .IN1(n4124), .SEL(n3664), .F(n4103) );
  IV U898 ( .A(n3662), .Z(n242) );
  MUX U899 ( .IN0(n4075), .IN1(n4073), .SEL(n4074), .F(n4052) );
  MUX U900 ( .IN0(n3565), .IN1(n3563), .SEL(n3564), .F(n3519) );
  MUX U901 ( .IN0(n243), .IN1(n3598), .SEL(n3599), .F(n3552) );
  IV U902 ( .A(n3600), .Z(n243) );
  MUX U903 ( .IN0(n3494), .IN1(n3492), .SEL(n3493), .F(n3446) );
  MUX U904 ( .IN0(n4529), .IN1(n4063), .SEL(n4064), .F(n4512) );
  MUX U905 ( .IN0(n4327), .IN1(n4325), .SEL(n4326), .F(n4303) );
  MUX U906 ( .IN0(n244), .IN1(n4040), .SEL(n3482), .F(n4019) );
  IV U907 ( .A(n3480), .Z(n244) );
  MUX U908 ( .IN0(n4698), .IN1(n4310), .SEL(n4312), .F(n4686) );
  MUX U909 ( .IN0(n3991), .IN1(n3989), .SEL(n3990), .F(n3968) );
  MUX U910 ( .IN0(n3383), .IN1(n3381), .SEL(n3382), .F(n3337) );
  MUX U911 ( .IN0(n245), .IN1(n3416), .SEL(n3417), .F(n3370) );
  IV U912 ( .A(n3418), .Z(n245) );
  MUX U913 ( .IN0(n3312), .IN1(n3310), .SEL(n3311), .F(n3267) );
  MUX U914 ( .IN0(n4461), .IN1(n3979), .SEL(n3980), .F(n4444) );
  MUX U915 ( .IN0(n4764), .IN1(n4350), .SEL(n4351), .F(n246) );
  IV U916 ( .A(n246), .Z(n4750) );
  MUX U917 ( .IN0(n4882), .IN1(n4880), .SEL(n4881), .F(n4860) );
  MUX U918 ( .IN0(n4241), .IN1(n4239), .SEL(n4240), .F(n4219) );
  MUX U919 ( .IN0(n247), .IN1(n3956), .SEL(n3300), .F(n3935) );
  IV U920 ( .A(n3298), .Z(n247) );
  MUX U921 ( .IN0(n5017), .IN1(n4867), .SEL(n4869), .F(n5005) );
  MUX U922 ( .IN0(n3831), .IN1(n3833), .SEL(n3832), .F(n3828) );
  MUX U923 ( .IN0(n4644), .IN1(n4226), .SEL(n4228), .F(n4634) );
  MUX U924 ( .IN0(n3908), .IN1(n3906), .SEL(n3907), .F(n3885) );
  MUX U925 ( .IN0(n3208), .IN1(n3206), .SEL(n3207), .F(n3164) );
  MUX U926 ( .IN0(n248), .IN1(n3238), .SEL(n3239), .F(n3196) );
  IV U927 ( .A(n3240), .Z(n248) );
  MUX U928 ( .IN0(n3139), .IN1(n3137), .SEL(n3138), .F(n3097) );
  MUX U929 ( .IN0(n249), .IN1(n3752), .SEL(n3753), .F(n3727) );
  IV U930 ( .A(n3754), .Z(n249) );
  XNOR U931 ( .A(n5233), .B(g_input[3]), .Z(n5234) );
  XNOR U932 ( .A(n4487), .B(g_input[23]), .Z(n4488) );
  MUX U933 ( .IN0(n4395), .IN1(n3896), .SEL(n3897), .F(n4378) );
  MUX U934 ( .IN0(n5235), .IN1(n250), .SEL(n5236), .F(n3019) );
  MUX U935 ( .IN0(n2112), .IN1(n2114), .SEL(n2113), .F(n2004) );
  MUX U936 ( .IN0(n2367), .IN1(n251), .SEL(n2368), .F(n2247) );
  IV U937 ( .A(n2369), .Z(n251) );
  MUX U938 ( .IN0(n2582), .IN1(n2584), .SEL(n2583), .F(n2457) );
  MUX U939 ( .IN0(n2539), .IN1(n2541), .SEL(n2540), .F(n2417) );
  MUX U940 ( .IN0(n2862), .IN1(n2864), .SEL(n2863), .F(n2730) );
  XNOR U941 ( .A(n5074), .B(n5073), .Z(n5079) );
  XNOR U942 ( .A(n4789), .B(n4788), .Z(n4815) );
  XNOR U943 ( .A(n4157), .B(n4155), .Z(n4170) );
  MUX U944 ( .IN0(n252), .IN1(n3873), .SEL(n3128), .F(n3853) );
  IV U945 ( .A(n3126), .Z(n252) );
  MUX U946 ( .IN0(n937), .IN1(n935), .SEL(n936), .F(n867) );
  MUX U947 ( .IN0(n1014), .IN1(n1012), .SEL(n1013), .F(n945) );
  MUX U948 ( .IN0(n253), .IN1(n5141), .SEL(e_input[31]), .F(n1133) );
  IV U949 ( .A(e_input[19]), .Z(n253) );
  MUX U950 ( .IN0(n254), .IN1(n1420), .SEL(n1421), .F(n1329) );
  IV U951 ( .A(n1422), .Z(n254) );
  MUX U952 ( .IN0(n255), .IN1(n3838), .SEL(e_input[31]), .F(n1638) );
  IV U953 ( .A(e_input[13]), .Z(n255) );
  MUX U954 ( .IN0(n1662), .IN1(n1660), .SEL(n1661), .F(n1562) );
  MUX U955 ( .IN0(n1852), .IN1(n1850), .SEL(n1851), .F(n1733) );
  MUX U956 ( .IN0(n256), .IN1(n2131), .SEL(n2132), .F(n2023) );
  IV U957 ( .A(n2133), .Z(n256) );
  MUX U958 ( .IN0(n2364), .IN1(n2362), .SEL(n2363), .F(n2242) );
  MUX U959 ( .IN0(n2946), .IN1(n2944), .SEL(n2945), .F(n2805) );
  XNOR U960 ( .A(n2998), .B(n2997), .Z(n4974) );
  MUX U961 ( .IN0(n257), .IN1(n3040), .SEL(n3041), .F(n2912) );
  IV U962 ( .A(n3042), .Z(n257) );
  XOR U963 ( .A(n968), .B(n906), .Z(n903) );
  MUX U964 ( .IN0(n258), .IN1(n1066), .SEL(n1067), .F(n994) );
  IV U965 ( .A(n1068), .Z(n258) );
  ANDN U966 ( .A(n1130), .B(n1129), .Z(n1057) );
  XNOR U967 ( .A(n1235), .B(n1234), .Z(n1312) );
  MUX U968 ( .IN0(n1292), .IN1(n259), .SEL(n1293), .F(n1215) );
  IV U969 ( .A(n1294), .Z(n259) );
  XNOR U970 ( .A(n1605), .B(n1604), .Z(n1696) );
  XNOR U971 ( .A(n1589), .B(n1588), .Z(n1678) );
  MUX U972 ( .IN0(n260), .IN1(n1776), .SEL(n1777), .F(n1675) );
  IV U973 ( .A(n1778), .Z(n260) );
  MUX U974 ( .IN0(n261), .IN1(n1794), .SEL(n1795), .F(n1693) );
  IV U975 ( .A(n1796), .Z(n261) );
  XNOR U976 ( .A(n1709), .B(n1708), .Z(n1805) );
  XNOR U977 ( .A(n1892), .B(n1891), .Z(n1994) );
  MUX U978 ( .IN0(n262), .IN1(n2234), .SEL(n2235), .F(n2115) );
  IV U979 ( .A(n2236), .Z(n262) );
  XNOR U980 ( .A(n2162), .B(n2172), .Z(n2278) );
  XNOR U981 ( .A(n2179), .B(n2178), .Z(n2288) );
  XNOR U982 ( .A(n2203), .B(n2202), .Z(n2318) );
  XNOR U983 ( .A(n2226), .B(n2225), .Z(n2341) );
  MUX U984 ( .IN0(n263), .IN1(n2460), .SEL(n2461), .F(n2338) );
  IV U985 ( .A(n2462), .Z(n263) );
  XNOR U986 ( .A(n2535), .B(n2534), .Z(n2654) );
  XNOR U987 ( .A(n2527), .B(n2526), .Z(n2646) );
  XNOR U988 ( .A(n2593), .B(n2592), .Z(n2720) );
  XNOR U989 ( .A(n2702), .B(n2701), .Z(n2829) );
  XNOR U990 ( .A(n2741), .B(n2740), .Z(n2868) );
  XNOR U991 ( .A(n2749), .B(n2748), .Z(n2876) );
  MUX U992 ( .IN0(n595), .IN1(n593), .SEL(n594), .F(n563) );
  NAND U993 ( .A(n706), .B(n705), .Z(n699) );
  XNOR U994 ( .A(n668), .B(n667), .Z(n707) );
  MUX U995 ( .IN0(n264), .IN1(n794), .SEL(n795), .F(n738) );
  IV U996 ( .A(n796), .Z(n264) );
  AND U997 ( .A(n1339), .B(n1341), .Z(n1255) );
  MUX U998 ( .IN0(n265), .IN1(n1373), .SEL(n1374), .F(n1282) );
  IV U999 ( .A(n1375), .Z(n265) );
  MUX U1000 ( .IN0(n266), .IN1(n1876), .SEL(n1877), .F(n1768) );
  IV U1001 ( .A(n1878), .Z(n266) );
  AND U1002 ( .A(n1926), .B(n1928), .Z(n1820) );
  MUX U1003 ( .IN0(n267), .IN1(n2330), .SEL(n2331), .F(n2210) );
  IV U1004 ( .A(n2332), .Z(n267) );
  XNOR U1005 ( .A(n2311), .B(n2310), .Z(n2308) );
  ANDN U1006 ( .A(n2502), .B(n2503), .Z(n2380) );
  MUX U1007 ( .IN0(n2692), .IN1(n2815), .SEL(n2694), .F(n2559) );
  MUX U1008 ( .IN0(n2843), .IN1(n361), .SEL(n2842), .F(n268) );
  IV U1009 ( .A(n268), .Z(n2709) );
  MUX U1010 ( .IN0(n269), .IN1(n2812), .SEL(n2813), .F(n2689) );
  IV U1011 ( .A(n2814), .Z(n269) );
  ANDN U1012 ( .A(n637), .B(n607), .Z(n596) );
  MUX U1013 ( .IN0(n839), .IN1(n841), .SEL(n840), .F(n270) );
  IV U1014 ( .A(n270), .Z(n784) );
  AND U1015 ( .A(n896), .B(n898), .Z(n833) );
  XOR U1016 ( .A(n848), .B(n845), .Z(n899) );
  NANDN U1017 ( .B(n956), .A(n957), .Z(n888) );
  XNOR U1018 ( .A(n1633), .B(n1634), .Z(n1653) );
  MUX U1019 ( .IN0(n271), .IN1(n2420), .SEL(n2421), .F(n2300) );
  IV U1020 ( .A(n2422), .Z(n271) );
  MUX U1021 ( .IN0(n2937), .IN1(n2935), .SEL(n2936), .F(n272) );
  IV U1022 ( .A(n272), .Z(n2796) );
  MUX U1023 ( .IN0(n533), .IN1(n531), .SEL(n532), .F(n273) );
  IV U1024 ( .A(n273), .Z(n510) );
  NANDN U1025 ( .B(n537), .A(n538), .Z(n494) );
  XOR U1026 ( .A(n1126), .B(n1125), .Z(n1106) );
  XOR U1027 ( .A(n1355), .B(n1354), .Z(n1439) );
  XOR U1028 ( .A(n1968), .B(n1965), .Z(n2042) );
  AND U1029 ( .A(n522), .B(n524), .Z(n497) );
  MUX U1030 ( .IN0(n2891), .IN1(\_MxM/Y0[1] ), .SEL(n2892), .F(n2759) );
  XNOR U1031 ( .A(n568), .B(n572), .Z(n570) );
  XNOR U1032 ( .A(n680), .B(n684), .Z(n682) );
  XNOR U1033 ( .A(n827), .B(n831), .Z(n829) );
  XNOR U1034 ( .A(n1025), .B(n1029), .Z(n1027) );
  XNOR U1035 ( .A(n1258), .B(n1262), .Z(n1260) );
  XNOR U1036 ( .A(n1530), .B(n1534), .Z(n1532) );
  XNOR U1037 ( .A(n1823), .B(n1827), .Z(n1825) );
  XNOR U1038 ( .A(n2144), .B(n2148), .Z(n2146) );
  MUX U1039 ( .IN0(n274), .IN1(n4166), .SEL(n3749), .F(n4145) );
  IV U1040 ( .A(n3748), .Z(n274) );
  MUX U1041 ( .IN0(n3630), .IN1(n3628), .SEL(n3629), .F(n3582) );
  MUX U1042 ( .IN0(n4117), .IN1(n4115), .SEL(n4116), .F(n4094) );
  MUX U1043 ( .IN0(n4563), .IN1(n4105), .SEL(n4106), .F(n4546) );
  MUX U1044 ( .IN0(n275), .IN1(n3552), .SEL(n3553), .F(n3508) );
  IV U1045 ( .A(n3554), .Z(n275) );
  MUX U1046 ( .IN0(n276), .IN1(n4082), .SEL(n3572), .F(n4061) );
  IV U1047 ( .A(n3570), .Z(n276) );
  MUX U1048 ( .IN0(n3448), .IN1(n3446), .SEL(n3447), .F(n3400) );
  MUX U1049 ( .IN0(n4033), .IN1(n4031), .SEL(n4032), .F(n4010) );
  MUX U1050 ( .IN0(n3475), .IN1(n3473), .SEL(n3474), .F(n3427) );
  MUX U1051 ( .IN0(n4495), .IN1(n4021), .SEL(n4022), .F(n4478) );
  MUX U1052 ( .IN0(n3844), .IN1(n4328), .SEL(n3845), .F(n277) );
  IV U1053 ( .A(n277), .Z(n4306) );
  MUX U1054 ( .IN0(n4686), .IN1(n4286), .SEL(n4288), .F(n4671) );
  MUX U1055 ( .IN0(n4281), .IN1(n4279), .SEL(n4280), .F(n4259) );
  MUX U1056 ( .IN0(n278), .IN1(n3370), .SEL(n3371), .F(n3326) );
  IV U1057 ( .A(n3372), .Z(n278) );
  MUX U1058 ( .IN0(n279), .IN1(n3998), .SEL(n3390), .F(n3977) );
  IV U1059 ( .A(n3388), .Z(n279) );
  MUX U1060 ( .IN0(n4904), .IN1(n4902), .SEL(n4903), .F(n4880) );
  MUX U1061 ( .IN0(n5043), .IN1(n4909), .SEL(n4911), .F(n5029) );
  MUX U1062 ( .IN0(n3269), .IN1(n3267), .SEL(n3268), .F(n3224) );
  MUX U1063 ( .IN0(n3949), .IN1(n3947), .SEL(n3948), .F(n3926) );
  MUX U1064 ( .IN0(n3293), .IN1(n3291), .SEL(n3292), .F(n3249) );
  MUX U1065 ( .IN0(n4428), .IN1(n3937), .SEL(n3938), .F(n4412) );
  MUX U1066 ( .IN0(g_input[1]), .IN1(n5250), .SEL(g_input[31]), .F(n280) );
  IV U1067 ( .A(n280), .Z(n3818) );
  MUX U1068 ( .IN0(n281), .IN1(n5169), .SEL(n5170), .F(n5158) );
  IV U1069 ( .A(n5171), .Z(n281) );
  MUX U1070 ( .IN0(n4634), .IN1(n4206), .SEL(n4208), .F(n4624) );
  MUX U1071 ( .IN0(n4201), .IN1(n4199), .SEL(n4200), .F(n4175) );
  MUX U1072 ( .IN0(n282), .IN1(n3196), .SEL(n3197), .F(n3153) );
  IV U1073 ( .A(n3198), .Z(n282) );
  MUX U1074 ( .IN0(n283), .IN1(n3915), .SEL(n3215), .F(n3894) );
  IV U1075 ( .A(n3213), .Z(n283) );
  XNOR U1076 ( .A(n5156), .B(g_input[7]), .Z(n5157) );
  XNOR U1077 ( .A(n5024), .B(g_input[11]), .Z(n5025) );
  XNOR U1078 ( .A(n4976), .B(g_input[15]), .Z(n4977) );
  XNOR U1079 ( .A(n4555), .B(g_input[19]), .Z(n4556) );
  MUX U1080 ( .IN0(g_input[2]), .IN1(n5243), .SEL(g_input[31]), .F(n284) );
  IV U1081 ( .A(n284), .Z(n3815) );
  MUX U1082 ( .IN0(n4822), .IN1(n4820), .SEL(n4821), .F(n4789) );
  MUX U1083 ( .IN0(n4993), .IN1(n4827), .SEL(n4829), .F(n4981) );
  MUX U1084 ( .IN0(n3099), .IN1(n3097), .SEL(n3098), .F(n3058) );
  MUX U1085 ( .IN0(n3121), .IN1(n3119), .SEL(n3120), .F(n3050) );
  XNOR U1086 ( .A(n4453), .B(g_input[25]), .Z(n4454) );
  MUX U1087 ( .IN0(n285), .IN1(n3825), .SEL(e_input[31]), .F(n2054) );
  IV U1088 ( .A(e_input[9]), .Z(n285) );
  MUX U1089 ( .IN0(n2574), .IN1(n2576), .SEL(n2575), .F(n2449) );
  MUX U1090 ( .IN0(n2793), .IN1(n2795), .SEL(n2794), .F(n2663) );
  MUX U1091 ( .IN0(g_input[4]), .IN1(n5202), .SEL(g_input[31]), .F(n2752) );
  MUX U1092 ( .IN0(n3019), .IN1(n286), .SEL(n3020), .F(n2878) );
  IV U1093 ( .A(n3021), .Z(n286) );
  MUX U1094 ( .IN0(g_input[9]), .IN1(n5053), .SEL(g_input[31]), .F(n287) );
  IV U1095 ( .A(n287), .Z(n2255) );
  MUX U1096 ( .IN0(n2987), .IN1(n2989), .SEL(n2988), .F(n2846) );
  MUX U1097 ( .IN0(e_input[1]), .IN1(n4782), .SEL(e_input[31]), .F(n288) );
  IV U1098 ( .A(n288), .Z(n4355) );
  XNOR U1099 ( .A(n3743), .B(n3741), .Z(n3757) );
  MUX U1100 ( .IN0(n1078), .IN1(n1076), .SEL(n1077), .F(n1004) );
  MUX U1101 ( .IN0(n289), .IN1(n1245), .SEL(n1246), .F(n1164) );
  IV U1102 ( .A(n1247), .Z(n289) );
  MUX U1103 ( .IN0(n1277), .IN1(n1275), .SEL(n1276), .F(n1193) );
  MUX U1104 ( .IN0(n1301), .IN1(n1303), .SEL(n1302), .F(n290) );
  MUX U1105 ( .IN0(n1703), .IN1(n1701), .SEL(n1702), .F(n1605) );
  MUX U1106 ( .IN0(n2287), .IN1(n2285), .SEL(n2286), .F(n2162) );
  MUX U1107 ( .IN0(n2807), .IN1(n2805), .SEL(n2806), .F(n2671) );
  MUX U1108 ( .IN0(n4358), .IN1(n3871), .SEL(n3872), .F(n291) );
  IV U1109 ( .A(n291), .Z(n2965) );
  XNOR U1110 ( .A(n4952), .B(n4949), .Z(n4950) );
  XNOR U1111 ( .A(n5255), .B(e_input[30]), .Z(n5253) );
  MUX U1112 ( .IN0(n292), .IN1(n857), .SEL(n858), .F(n794) );
  IV U1113 ( .A(n859), .Z(n292) );
  XNOR U1114 ( .A(n1319), .B(n1318), .Z(n1407) );
  MUX U1115 ( .IN0(n293), .IN1(n1483), .SEL(n1484), .F(n1383) );
  IV U1116 ( .A(n1485), .Z(n293) );
  MUX U1117 ( .IN0(n294), .IN1(n1597), .SEL(n1598), .F(n1501) );
  IV U1118 ( .A(n1599), .Z(n294) );
  XNOR U1119 ( .A(n1517), .B(n1516), .Z(n1608) );
  XNOR U1120 ( .A(n1562), .B(n1561), .Z(n1655) );
  XNOR U1121 ( .A(n1685), .B(n1684), .Z(n1779) );
  XNOR U1122 ( .A(n1850), .B(n1849), .Z(n1951) );
  XNOR U1123 ( .A(n2015), .B(n2014), .Z(n2118) );
  XNOR U1124 ( .A(n2023), .B(n2022), .Z(n2126) );
  XNOR U1125 ( .A(n1976), .B(n1975), .Z(n2079) );
  MUX U1126 ( .IN0(n295), .IN1(n2099), .SEL(n2100), .F(n1991) );
  IV U1127 ( .A(n2101), .Z(n295) );
  XNOR U1128 ( .A(n2346), .B(n2345), .Z(n2463) );
  MUX U1129 ( .IN0(n296), .IN1(n2476), .SEL(n2477), .F(n2354) );
  IV U1130 ( .A(n2478), .Z(n296) );
  XNOR U1131 ( .A(n2293), .B(n2292), .Z(n2408) );
  MUX U1132 ( .IN0(n297), .IN1(n2395), .SEL(n2396), .F(n2275) );
  IV U1133 ( .A(n2397), .Z(n297) );
  XNOR U1134 ( .A(n2609), .B(n2608), .Z(n2736) );
  XNOR U1135 ( .A(n2617), .B(n2616), .Z(n2744) );
  XNOR U1136 ( .A(n2570), .B(n2569), .Z(n2697) );
  XNOR U1137 ( .A(n2725), .B(n2724), .Z(n2852) );
  XNOR U1138 ( .A(n2659), .B(n2658), .Z(n2784) );
  XNOR U1139 ( .A(n2651), .B(n2650), .Z(n2776) );
  MUX U1140 ( .IN0(n3008), .IN1(n3006), .SEL(n3007), .F(n298) );
  IV U1141 ( .A(n298), .Z(n2865) );
  MUX U1142 ( .IN0(n299), .IN1(n2990), .SEL(n2991), .F(n2849) );
  IV U1143 ( .A(n2992), .Z(n299) );
  MUX U1144 ( .IN0(n300), .IN1(n2912), .SEL(n2913), .F(n2773) );
  IV U1145 ( .A(n2914), .Z(n300) );
  MUX U1146 ( .IN0(n2962), .IN1(n301), .SEL(n2963), .F(n2825) );
  IV U1147 ( .A(n2964), .Z(n301) );
  MUX U1148 ( .IN0(n586), .IN1(n584), .SEL(n585), .F(n551) );
  MUX U1149 ( .IN0(n302), .IN1(n655), .SEL(n656), .F(n619) );
  IV U1150 ( .A(n657), .Z(n302) );
  XNOR U1151 ( .A(n712), .B(n711), .Z(n749) );
  XNOR U1152 ( .A(n746), .B(n744), .Z(n797) );
  AND U1153 ( .A(n848), .B(n849), .Z(n778) );
  MUX U1154 ( .IN0(n303), .IN1(n981), .SEL(n982), .F(n912) );
  IV U1155 ( .A(n983), .Z(n303) );
  XOR U1156 ( .A(n1054), .B(n1058), .Z(n1127) );
  XNOR U1157 ( .A(n1540), .B(n1539), .Z(n1538) );
  MUX U1158 ( .IN0(n304), .IN1(n1667), .SEL(n1668), .F(n1569) );
  IV U1159 ( .A(n1669), .Z(n304) );
  AND U1160 ( .A(n1719), .B(n1721), .Z(n1623) );
  MUX U1161 ( .IN0(n305), .IN1(n1731), .SEL(n1730), .F(n1634) );
  IV U1162 ( .A(n1729), .Z(n305) );
  AND U1163 ( .A(n2141), .B(n2143), .Z(n2033) );
  MUX U1164 ( .IN0(n306), .IN1(n2210), .SEL(n2211), .F(n2091) );
  IV U1165 ( .A(n2212), .Z(n306) );
  MUX U1166 ( .IN0(n307), .IN1(n2709), .SEL(n2710), .F(n2577) );
  IV U1167 ( .A(n2711), .Z(n307) );
  MUX U1168 ( .IN0(n560), .IN1(n562), .SEL(n561), .F(n528) );
  AND U1169 ( .A(n783), .B(n784), .Z(n780) );
  MUX U1170 ( .IN0(n308), .IN1(n1749), .SEL(n1750), .F(n1648) );
  IV U1171 ( .A(n1751), .Z(n308) );
  XOR U1172 ( .A(n2189), .B(n2075), .Z(n2076) );
  XNOR U1173 ( .A(n2436), .B(n2434), .Z(n2545) );
  NANDN U1174 ( .B(n535), .A(n534), .Z(n506) );
  XNOR U1175 ( .A(n537), .B(n542), .Z(n538) );
  XNOR U1176 ( .A(n638), .B(n643), .Z(n639) );
  XNOR U1177 ( .A(n766), .B(n731), .Z(n767) );
  XNOR U1178 ( .A(n956), .B(n961), .Z(n957) );
  XOR U1179 ( .A(n1204), .B(n1203), .Z(n1184) );
  MUX U1180 ( .IN0(\_MxM/Y0[2] ), .IN1(n2759), .SEL(n2760), .F(n2627) );
  XOR U1181 ( .A(n1357), .B(n1356), .Z(n1436) );
  XOR U1182 ( .A(n1967), .B(n1966), .Z(n2039) );
  XOR U1183 ( .A(n2302), .B(n2301), .Z(n2386) );
  XNOR U1184 ( .A(n2632), .B(n2511), .Z(n2512) );
  XOR U1185 ( .A(n2798), .B(n2797), .Z(n2903) );
  XNOR U1186 ( .A(n599), .B(n603), .Z(n601) );
  XNOR U1187 ( .A(n724), .B(n728), .Z(n726) );
  XNOR U1188 ( .A(n890), .B(n894), .Z(n892) );
  XNOR U1189 ( .A(n1099), .B(n1103), .Z(n1101) );
  XNOR U1190 ( .A(n1342), .B(n1346), .Z(n1344) );
  XNOR U1191 ( .A(n1626), .B(n1630), .Z(n1628) );
  XNOR U1192 ( .A(n1929), .B(n1933), .Z(n1931) );
  XNOR U1193 ( .A(n2263), .B(n2267), .Z(n2265) );
  XOR U1194 ( .A(n482), .B(n483), .Z(n365) );
  MUX U1195 ( .IN0(n3720), .IN1(n3718), .SEL(n3719), .F(n3674) );
  MUX U1196 ( .IN0(n3703), .IN1(n3701), .SEL(n3702), .F(n3655) );
  MUX U1197 ( .IN0(n309), .IN1(n3644), .SEL(n3645), .F(n3598) );
  IV U1198 ( .A(n3646), .Z(n309) );
  MUX U1199 ( .IN0(n3540), .IN1(n3538), .SEL(n3539), .F(n3492) );
  MUX U1200 ( .IN0(n310), .IN1(n4103), .SEL(n3618), .F(n4082) );
  IV U1201 ( .A(n3616), .Z(n310) );
  MUX U1202 ( .IN0(n4546), .IN1(n4084), .SEL(n4085), .F(n4529) );
  MUX U1203 ( .IN0(n4054), .IN1(n4052), .SEL(n4053), .F(n4031) );
  MUX U1204 ( .IN0(n3521), .IN1(n3519), .SEL(n3520), .F(n3473) );
  MUX U1205 ( .IN0(n311), .IN1(n3462), .SEL(n3463), .F(n3416) );
  IV U1206 ( .A(n3464), .Z(n311) );
  MUX U1207 ( .IN0(n3358), .IN1(n3356), .SEL(n3357), .F(n3310) );
  MUX U1208 ( .IN0(n312), .IN1(n4019), .SEL(n3436), .F(n3998) );
  IV U1209 ( .A(n3434), .Z(n312) );
  MUX U1210 ( .IN0(n4478), .IN1(n4000), .SEL(n4001), .F(n4461) );
  MUX U1211 ( .IN0(n4928), .IN1(n4926), .SEL(n4927), .F(n4902) );
  MUX U1212 ( .IN0(n5060), .IN1(n4933), .SEL(n4935), .F(n5043) );
  MUX U1213 ( .IN0(n3970), .IN1(n3968), .SEL(n3969), .F(n3947) );
  MUX U1214 ( .IN0(n3339), .IN1(n3337), .SEL(n3338), .F(n3291) );
  MUX U1215 ( .IN0(n4671), .IN1(n4266), .SEL(n4268), .F(n4656) );
  MUX U1216 ( .IN0(n4261), .IN1(n4259), .SEL(n4260), .F(n4239) );
  MUX U1217 ( .IN0(n5128), .IN1(n4972), .SEL(n4973), .F(n313) );
  IV U1218 ( .A(n313), .Z(n5114) );
  MUX U1219 ( .IN0(n3804), .IN1(n3755), .SEL(n3756), .F(n314) );
  IV U1220 ( .A(n314), .Z(n3790) );
  MUX U1221 ( .IN0(n315), .IN1(n3787), .SEL(n3788), .F(n3773) );
  IV U1222 ( .A(n3789), .Z(n315) );
  MUX U1223 ( .IN0(n316), .IN1(n3281), .SEL(n3282), .F(n3238) );
  IV U1224 ( .A(n3283), .Z(n316) );
  MUX U1225 ( .IN0(n5211), .IN1(n5152), .SEL(n5153), .F(n317) );
  IV U1226 ( .A(n317), .Z(n5195) );
  MUX U1227 ( .IN0(n3184), .IN1(n3182), .SEL(n3183), .F(n3137) );
  MUX U1228 ( .IN0(n318), .IN1(n3935), .SEL(n3258), .F(n3915) );
  IV U1229 ( .A(n3256), .Z(n318) );
  MUX U1230 ( .IN0(n4412), .IN1(n3917), .SEL(n3918), .F(n4395) );
  MUX U1231 ( .IN0(n5239), .IN1(n5241), .SEL(n5240), .F(n5235) );
  MUX U1232 ( .IN0(n4842), .IN1(n4840), .SEL(n4841), .F(n4820) );
  MUX U1233 ( .IN0(n5005), .IN1(n4847), .SEL(n4849), .F(n4993) );
  MUX U1234 ( .IN0(n319), .IN1(n3759), .SEL(n3760), .F(n3737) );
  IV U1235 ( .A(n3761), .Z(n319) );
  MUX U1236 ( .IN0(n3887), .IN1(n3885), .SEL(n3886), .F(n3861) );
  MUX U1237 ( .IN0(n3166), .IN1(n3164), .SEL(n3165), .F(n3119) );
  XNOR U1238 ( .A(n5183), .B(g_input[5]), .Z(n5184) );
  XNOR U1239 ( .A(n5052), .B(g_input[9]), .Z(n5053) );
  MUX U1240 ( .IN0(n320), .IN1(n4966), .SEL(e_input[31]), .F(n4958) );
  IV U1241 ( .A(e_input[21]), .Z(n320) );
  XNOR U1242 ( .A(n5000), .B(g_input[13]), .Z(n5001) );
  XNOR U1243 ( .A(n4589), .B(g_input[17]), .Z(n4590) );
  XNOR U1244 ( .A(n4521), .B(g_input[21]), .Z(n4522) );
  AND U1245 ( .A(n5251), .B(g_input[0]), .Z(n3029) );
  MUX U1246 ( .IN0(n4177), .IN1(n4175), .SEL(n4176), .F(n4157) );
  MUX U1247 ( .IN0(n4624), .IN1(n4186), .SEL(n4188), .F(n4614) );
  MUX U1248 ( .IN0(n321), .IN1(n5230), .SEL(e_input[31]), .F(n5217) );
  IV U1249 ( .A(e_input[25]), .Z(n321) );
  MUX U1250 ( .IN0(n322), .IN1(n5248), .SEL(e_input[31]), .F(n5238) );
  IV U1251 ( .A(e_input[29]), .Z(n322) );
  XNOR U1252 ( .A(n4421), .B(g_input[27]), .Z(n4422) );
  MUX U1253 ( .IN0(g_input[3]), .IN1(n5234), .SEL(g_input[31]), .F(n2884) );
  MUX U1254 ( .IN0(n3003), .IN1(n3005), .SEL(n3004), .F(n2862) );
  MUX U1255 ( .IN0(n2979), .IN1(n2981), .SEL(n2980), .F(n2838) );
  MUX U1256 ( .IN0(e_input[20]), .IN1(n323), .SEL(e_input[31]), .F(n1036) );
  IV U1257 ( .A(n4965), .Z(n323) );
  MUX U1258 ( .IN0(e_input[16]), .IN1(n324), .SEL(e_input[31]), .F(n1398) );
  IV U1259 ( .A(n5145), .Z(n324) );
  MUX U1260 ( .IN0(e_input[8]), .IN1(n325), .SEL(e_input[31]), .F(n2173) );
  IV U1261 ( .A(n3824), .Z(n325) );
  MUX U1262 ( .IN0(e_input[12]), .IN1(n326), .SEL(e_input[31]), .F(n1744) );
  IV U1263 ( .A(n3837), .Z(n326) );
  MUX U1264 ( .IN0(e_input[4]), .IN1(n327), .SEL(e_input[31]), .F(n2682) );
  IV U1265 ( .A(n4343), .Z(n327) );
  XNOR U1266 ( .A(n4331), .B(n4328), .Z(n4329) );
  MUX U1267 ( .IN0(n328), .IN1(n3109), .SEL(n3110), .F(n3040) );
  IV U1268 ( .A(n3111), .Z(n328) );
  MUX U1269 ( .IN0(n329), .IN1(n5224), .SEL(e_input[31]), .F(n651) );
  IV U1270 ( .A(e_input[27]), .Z(n329) );
  MUX U1271 ( .IN0(e_input[26]), .IN1(n330), .SEL(e_input[31]), .F(n692) );
  IV U1272 ( .A(n5225), .Z(n330) );
  MUX U1273 ( .IN0(e_input[24]), .IN1(n331), .SEL(e_input[31]), .F(n799) );
  IV U1274 ( .A(n5229), .Z(n331) );
  MUX U1275 ( .IN0(e_input[28]), .IN1(n332), .SEL(e_input[31]), .F(n624) );
  IV U1276 ( .A(n5247), .Z(n332) );
  MUX U1277 ( .IN0(n1117), .IN1(n1115), .SEL(n1116), .F(n1042) );
  MUX U1278 ( .IN0(n333), .IN1(n1164), .SEL(n1165), .F(n1086) );
  IV U1279 ( .A(n1166), .Z(n333) );
  MUX U1280 ( .IN0(n1158), .IN1(n1156), .SEL(n1157), .F(n1076) );
  MUX U1281 ( .IN0(e_input[18]), .IN1(n334), .SEL(e_input[31]), .F(n1214) );
  IV U1282 ( .A(n5140), .Z(n334) );
  MUX U1283 ( .IN0(n335), .IN1(n5146), .SEL(e_input[31]), .F(n1298) );
  IV U1284 ( .A(e_input[17]), .Z(n335) );
  MUX U1285 ( .IN0(n1495), .IN1(n1493), .SEL(n1494), .F(n1387) );
  MUX U1286 ( .IN0(n1468), .IN1(n1466), .SEL(n1467), .F(n1364) );
  MUX U1287 ( .IN0(n1511), .IN1(n1509), .SEL(n1510), .F(n1412) );
  MUX U1288 ( .IN0(n336), .IN1(n1517), .SEL(n1518), .F(n1420) );
  IV U1289 ( .A(n1519), .Z(n336) );
  MUX U1290 ( .IN0(n337), .IN1(n3820), .SEL(e_input[31]), .F(n1837) );
  IV U1291 ( .A(e_input[11]), .Z(n337) );
  MUX U1292 ( .IN0(e_input[10]), .IN1(n338), .SEL(e_input[31]), .F(n1943) );
  IV U1293 ( .A(n3819), .Z(n338) );
  MUX U1294 ( .IN0(n2067), .IN1(n2065), .SEL(n2066), .F(n1958) );
  MUX U1295 ( .IN0(e_input[6]), .IN1(n339), .SEL(e_input[31]), .F(n2433) );
  IV U1296 ( .A(n4348), .Z(n339) );
  MUX U1297 ( .IN0(n340), .IN1(n4344), .SEL(e_input[31]), .F(n2549) );
  IV U1298 ( .A(e_input[5]), .Z(n340) );
  MUX U1299 ( .IN0(n341), .IN1(n4778), .SEL(e_input[31]), .F(n2822) );
  IV U1300 ( .A(e_input[3]), .Z(n341) );
  MUX U1301 ( .IN0(e_input[2]), .IN1(n342), .SEL(e_input[31]), .F(n2961) );
  IV U1302 ( .A(n4777), .Z(n342) );
  MUX U1303 ( .IN0(n3853), .IN1(n343), .SEL(n3090), .F(n2962) );
  IV U1304 ( .A(n3089), .Z(n343) );
  MUX U1305 ( .IN0(e_input[22]), .IN1(n344), .SEL(e_input[31]), .F(n908) );
  IV U1306 ( .A(n4971), .Z(n344) );
  MUX U1307 ( .IN0(n345), .IN1(n4970), .SEL(e_input[31]), .F(n838) );
  IV U1308 ( .A(e_input[23]), .Z(n345) );
  MUX U1309 ( .IN0(n346), .IN1(n925), .SEL(n926), .F(n857) );
  IV U1310 ( .A(n927), .Z(n346) );
  MUX U1311 ( .IN0(n347), .IN1(n1225), .SEL(n1226), .F(n1146) );
  IV U1312 ( .A(n1227), .Z(n347) );
  MUX U1313 ( .IN0(n1643), .IN1(n1641), .SEL(n1642), .F(n348) );
  MUX U1314 ( .IN0(e_input[14]), .IN1(n349), .SEL(e_input[31]), .F(n1547) );
  IV U1315 ( .A(n3842), .Z(n349) );
  MUX U1316 ( .IN0(n350), .IN1(n1579), .SEL(n1580), .F(n1483) );
  IV U1317 ( .A(n1581), .Z(n350) );
  XNOR U1318 ( .A(n1802), .B(n1801), .Z(n1903) );
  XNOR U1319 ( .A(n1810), .B(n1809), .Z(n1911) );
  XNOR U1320 ( .A(n1761), .B(n1760), .Z(n1864) );
  XNOR U1321 ( .A(n1786), .B(n1785), .Z(n1887) );
  MUX U1322 ( .IN0(n351), .IN1(n1991), .SEL(n1992), .F(n1884) );
  IV U1323 ( .A(n1993), .Z(n351) );
  MUX U1324 ( .IN0(n352), .IN1(n2007), .SEL(n2008), .F(n1900) );
  IV U1325 ( .A(n2009), .Z(n352) );
  MUX U1326 ( .IN0(n1947), .IN1(n2051), .SEL(n1949), .F(n1839) );
  XNOR U1327 ( .A(n2107), .B(n2106), .Z(n2221) );
  XNOR U1328 ( .A(n2084), .B(n2083), .Z(n2198) );
  XNOR U1329 ( .A(n2123), .B(n2122), .Z(n2237) );
  XNOR U1330 ( .A(n2131), .B(n2130), .Z(n2245) );
  MUX U1331 ( .IN0(n353), .IN1(n2158), .SEL(n2159), .F(n2048) );
  IV U1332 ( .A(n2160), .Z(n353) );
  MUX U1333 ( .IN0(n354), .IN1(n4349), .SEL(e_input[31]), .F(n2307) );
  IV U1334 ( .A(e_input[7]), .Z(n354) );
  XNOR U1335 ( .A(n2492), .B(n2491), .Z(n2612) );
  XNOR U1336 ( .A(n2484), .B(n2483), .Z(n2604) );
  XNOR U1337 ( .A(n2445), .B(n2444), .Z(n2565) );
  XNOR U1338 ( .A(n2468), .B(n2467), .Z(n2588) );
  XNOR U1339 ( .A(n2405), .B(n2404), .Z(n2522) );
  XNOR U1340 ( .A(n2413), .B(n2412), .Z(n2530) );
  MUX U1341 ( .IN0(n355), .IN1(n2643), .SEL(n2644), .F(n2519) );
  IV U1342 ( .A(n2645), .Z(n355) );
  MUX U1343 ( .IN0(n356), .IN1(n2733), .SEL(n2734), .F(n2601) );
  IV U1344 ( .A(n2735), .Z(n356) );
  MUX U1345 ( .IN0(n357), .IN1(n2717), .SEL(n2718), .F(n2585) );
  IV U1346 ( .A(n2719), .Z(n357) );
  XNOR U1347 ( .A(n2881), .B(n2880), .Z(n3017) );
  XNOR U1348 ( .A(n2873), .B(n2872), .Z(n3009) );
  XNOR U1349 ( .A(n2834), .B(n2833), .Z(n2970) );
  XNOR U1350 ( .A(n2857), .B(n2856), .Z(n2993) );
  XNOR U1351 ( .A(n2781), .B(n2780), .Z(n2915) );
  XNOR U1352 ( .A(n2789), .B(n2788), .Z(n2923) );
  MUX U1353 ( .IN0(n2965), .IN1(n4352), .SEL(n2967), .F(n2824) );
  XNOR U1354 ( .A(n2805), .B(n2804), .Z(n2939) );
  MUX U1355 ( .IN0(e_input[30]), .IN1(n358), .SEL(e_input[31]), .F(n558) );
  IV U1356 ( .A(n5253), .Z(n358) );
  XNOR U1357 ( .A(n701), .B(n705), .Z(n741) );
  NAND U1358 ( .A(n906), .B(n905), .Z(n900) );
  MUX U1359 ( .IN0(n909), .IN1(n911), .SEL(n910), .F(n839) );
  XNOR U1360 ( .A(n754), .B(n753), .Z(n808) );
  NAND U1361 ( .A(n1057), .B(n1058), .Z(n1052) );
  MUX U1362 ( .IN0(n359), .IN1(n1473), .SEL(n1474), .F(n1373) );
  IV U1363 ( .A(n1475), .Z(n359) );
  MUX U1364 ( .IN0(n360), .IN1(n3843), .SEL(e_input[31]), .F(n1446) );
  IV U1365 ( .A(e_input[15]), .Z(n360) );
  AND U1366 ( .A(n1527), .B(n1529), .Z(n1430) );
  ANDN U1367 ( .A(n1968), .B(n1969), .Z(n1860) );
  MUX U1368 ( .IN0(n2984), .IN1(n2982), .SEL(n2983), .F(n361) );
  IV U1369 ( .A(n361), .Z(n2841) );
  MUX U1370 ( .IN0(n362), .IN1(n2951), .SEL(n2952), .F(n2812) );
  IV U1371 ( .A(n2953), .Z(n362) );
  MUX U1372 ( .IN0(n553), .IN1(n551), .SEL(n552), .F(n531) );
  ANDN U1373 ( .A(n563), .B(n564), .Z(n534) );
  MUX U1374 ( .IN0(n363), .IN1(n786), .SEL(n787), .F(n763) );
  IV U1375 ( .A(n788), .Z(n363) );
  XNOR U1376 ( .A(n1448), .B(n1447), .Z(n1441) );
  XNOR U1377 ( .A(n2314), .B(n2309), .Z(n2423) );
  MUX U1378 ( .IN0(n528), .IN1(n530), .SEL(n529), .F(n364) );
  IV U1379 ( .A(n364), .Z(n513) );
  XNOR U1380 ( .A(n597), .B(n602), .Z(n598) );
  XNOR U1381 ( .A(n722), .B(n727), .Z(n723) );
  XNOR U1382 ( .A(n888), .B(n893), .Z(n889) );
  XOR U1383 ( .A(n1051), .B(n1050), .Z(n1032) );
  XOR U1384 ( .A(n1284), .B(n1283), .Z(n1266) );
  XOR U1385 ( .A(n1550), .B(n1549), .Z(n1629) );
  XOR U1386 ( .A(n1751), .B(n1750), .Z(n1826) );
  XOR U1387 ( .A(n1859), .B(n1858), .Z(n1932) );
  XOR U1388 ( .A(n2074), .B(n2073), .Z(n2147) );
  XOR U1389 ( .A(n2188), .B(n2187), .Z(n2266) );
  XOR U1390 ( .A(n2422), .B(n2421), .Z(n2508) );
  XOR U1391 ( .A(n2544), .B(n2543), .Z(n2632) );
  XOR U1392 ( .A(n2668), .B(n2667), .Z(n2762) );
  AND U1393 ( .A(\_MxM/Y0[0] ), .B(n2766), .Z(n2891) );
  XNOR U1394 ( .A(n539), .B(n543), .Z(n541) );
  XNOR U1395 ( .A(n640), .B(n644), .Z(n642) );
  XNOR U1396 ( .A(n768), .B(n771), .Z(n770) );
  XNOR U1397 ( .A(n958), .B(n962), .Z(n960) );
  XNOR U1398 ( .A(n1177), .B(n1181), .Z(n1179) );
  XNOR U1399 ( .A(n1433), .B(n1437), .Z(n1435) );
  XNOR U1400 ( .A(n1722), .B(n1726), .Z(n1724) );
  XNOR U1401 ( .A(n2036), .B(n2040), .Z(n2038) );
  XNOR U1402 ( .A(n2383), .B(n2387), .Z(n2385) );
  MUX U1403 ( .IN0(n365), .IN1(n474), .SEL(n480), .F(n477) );
  ANDN U1404 ( .A(n366), .B(\_MxM/n[0] ), .Z(\_MxM/n390 ) );
  AND U1405 ( .A(\_MxM/N8 ), .B(n366), .Z(\_MxM/n389 ) );
  AND U1406 ( .A(\_MxM/N9 ), .B(n366), .Z(\_MxM/n388 ) );
  AND U1407 ( .A(\_MxM/N10 ), .B(n366), .Z(\_MxM/n387 ) );
  AND U1408 ( .A(\_MxM/N11 ), .B(n366), .Z(\_MxM/n386 ) );
  AND U1409 ( .A(\_MxM/N12 ), .B(n366), .Z(\_MxM/n385 ) );
  AND U1410 ( .A(\_MxM/N13 ), .B(n366), .Z(\_MxM/n384 ) );
  AND U1411 ( .A(\_MxM/N14 ), .B(n366), .Z(\_MxM/n383 ) );
  AND U1412 ( .A(\_MxM/N15 ), .B(n366), .Z(\_MxM/n382 ) );
  AND U1413 ( .A(\_MxM/N16 ), .B(n366), .Z(\_MxM/n381 ) );
  AND U1414 ( .A(\_MxM/N17 ), .B(n366), .Z(\_MxM/n380 ) );
  AND U1415 ( .A(\_MxM/N18 ), .B(n366), .Z(\_MxM/n379 ) );
  AND U1416 ( .A(\_MxM/N19 ), .B(n366), .Z(\_MxM/n378 ) );
  AND U1417 ( .A(n366), .B(n367), .Z(\_MxM/n377 ) );
  XOR U1418 ( .A(\_MxM/n[13] ), .B(\_MxM/add_39/carry[13] ), .Z(n367) );
  ANDN U1419 ( .A(n368), .B(rst), .Z(n366) );
  NAND U1420 ( .A(n369), .B(n370), .Z(n368) );
  AND U1421 ( .A(n371), .B(n372), .Z(n370) );
  AND U1422 ( .A(n373), .B(n374), .Z(n372) );
  AND U1423 ( .A(n375), .B(n376), .Z(n374) );
  AND U1424 ( .A(\_MxM/n[13] ), .B(n377), .Z(n371) );
  AND U1425 ( .A(\_MxM/n[10] ), .B(\_MxM/n[0] ), .Z(n377) );
  AND U1426 ( .A(n378), .B(n379), .Z(n369) );
  AND U1427 ( .A(\_MxM/n[3] ), .B(n380), .Z(n379) );
  AND U1428 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n380) );
  AND U1429 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n378) );
  NAND U1430 ( .A(n381), .B(n382), .Z(\_MxM/n376 ) );
  NAND U1431 ( .A(n383), .B(n384), .Z(n382) );
  NAND U1432 ( .A(\_MxM/Y0[0] ), .B(rst), .Z(n381) );
  NAND U1433 ( .A(n385), .B(n386), .Z(\_MxM/n375 ) );
  NAND U1434 ( .A(n387), .B(n384), .Z(n386) );
  NAND U1435 ( .A(\_MxM/Y0[1] ), .B(rst), .Z(n385) );
  NAND U1436 ( .A(n388), .B(n389), .Z(\_MxM/n374 ) );
  NAND U1437 ( .A(n390), .B(n384), .Z(n389) );
  NAND U1438 ( .A(\_MxM/Y0[2] ), .B(rst), .Z(n388) );
  NAND U1439 ( .A(n391), .B(n392), .Z(\_MxM/n373 ) );
  NAND U1440 ( .A(n393), .B(n384), .Z(n392) );
  NAND U1441 ( .A(\_MxM/Y0[3] ), .B(rst), .Z(n391) );
  NAND U1442 ( .A(n394), .B(n395), .Z(\_MxM/n372 ) );
  NAND U1443 ( .A(n396), .B(n384), .Z(n395) );
  NAND U1444 ( .A(\_MxM/Y0[4] ), .B(rst), .Z(n394) );
  NAND U1445 ( .A(n397), .B(n398), .Z(\_MxM/n371 ) );
  NAND U1446 ( .A(n399), .B(n384), .Z(n398) );
  NAND U1447 ( .A(rst), .B(\_MxM/Y0[5] ), .Z(n397) );
  NAND U1448 ( .A(n400), .B(n401), .Z(\_MxM/n370 ) );
  NAND U1449 ( .A(n402), .B(n384), .Z(n401) );
  NAND U1450 ( .A(rst), .B(\_MxM/Y0[6] ), .Z(n400) );
  NAND U1451 ( .A(n403), .B(n404), .Z(\_MxM/n369 ) );
  NAND U1452 ( .A(n405), .B(n384), .Z(n404) );
  NAND U1453 ( .A(rst), .B(\_MxM/Y0[7] ), .Z(n403) );
  NAND U1454 ( .A(n406), .B(n407), .Z(\_MxM/n368 ) );
  NAND U1455 ( .A(n408), .B(n384), .Z(n407) );
  NAND U1456 ( .A(rst), .B(\_MxM/Y0[8] ), .Z(n406) );
  NAND U1457 ( .A(n409), .B(n410), .Z(\_MxM/n367 ) );
  NAND U1458 ( .A(n411), .B(n384), .Z(n410) );
  NAND U1459 ( .A(rst), .B(\_MxM/Y0[9] ), .Z(n409) );
  NAND U1460 ( .A(n412), .B(n413), .Z(\_MxM/n366 ) );
  NAND U1461 ( .A(n414), .B(n384), .Z(n413) );
  NAND U1462 ( .A(rst), .B(\_MxM/Y0[10] ), .Z(n412) );
  NAND U1463 ( .A(n415), .B(n416), .Z(\_MxM/n365 ) );
  NAND U1464 ( .A(n417), .B(n384), .Z(n416) );
  NAND U1465 ( .A(rst), .B(\_MxM/Y0[11] ), .Z(n415) );
  NAND U1466 ( .A(n418), .B(n419), .Z(\_MxM/n364 ) );
  NAND U1467 ( .A(n420), .B(n384), .Z(n419) );
  NAND U1468 ( .A(rst), .B(\_MxM/Y0[12] ), .Z(n418) );
  NAND U1469 ( .A(n421), .B(n422), .Z(\_MxM/n363 ) );
  NAND U1470 ( .A(n423), .B(n384), .Z(n422) );
  NAND U1471 ( .A(rst), .B(\_MxM/Y0[13] ), .Z(n421) );
  NAND U1472 ( .A(n424), .B(n425), .Z(\_MxM/n362 ) );
  NAND U1473 ( .A(n426), .B(n384), .Z(n425) );
  NAND U1474 ( .A(rst), .B(\_MxM/Y0[14] ), .Z(n424) );
  NAND U1475 ( .A(n427), .B(n428), .Z(\_MxM/n361 ) );
  NAND U1476 ( .A(n429), .B(n384), .Z(n428) );
  NAND U1477 ( .A(rst), .B(\_MxM/Y0[15] ), .Z(n427) );
  NAND U1478 ( .A(n430), .B(n431), .Z(\_MxM/n360 ) );
  NAND U1479 ( .A(n432), .B(n384), .Z(n431) );
  NAND U1480 ( .A(rst), .B(\_MxM/Y0[16] ), .Z(n430) );
  NAND U1481 ( .A(n433), .B(n434), .Z(\_MxM/n359 ) );
  NAND U1482 ( .A(n435), .B(n384), .Z(n434) );
  NAND U1483 ( .A(rst), .B(\_MxM/Y0[17] ), .Z(n433) );
  NAND U1484 ( .A(n436), .B(n437), .Z(\_MxM/n358 ) );
  NAND U1485 ( .A(n438), .B(n384), .Z(n437) );
  NAND U1486 ( .A(rst), .B(\_MxM/Y0[18] ), .Z(n436) );
  NAND U1487 ( .A(n439), .B(n440), .Z(\_MxM/n357 ) );
  NAND U1488 ( .A(n441), .B(n384), .Z(n440) );
  NAND U1489 ( .A(rst), .B(\_MxM/Y0[19] ), .Z(n439) );
  NAND U1490 ( .A(n442), .B(n443), .Z(\_MxM/n356 ) );
  NAND U1491 ( .A(n444), .B(n384), .Z(n443) );
  NAND U1492 ( .A(rst), .B(\_MxM/Y0[20] ), .Z(n442) );
  NAND U1493 ( .A(n445), .B(n446), .Z(\_MxM/n355 ) );
  NAND U1494 ( .A(n447), .B(n384), .Z(n446) );
  NAND U1495 ( .A(rst), .B(\_MxM/Y0[21] ), .Z(n445) );
  NAND U1496 ( .A(n448), .B(n449), .Z(\_MxM/n354 ) );
  NAND U1497 ( .A(n450), .B(n384), .Z(n449) );
  NAND U1498 ( .A(rst), .B(\_MxM/Y0[22] ), .Z(n448) );
  NAND U1499 ( .A(n451), .B(n452), .Z(\_MxM/n353 ) );
  NAND U1500 ( .A(n453), .B(n384), .Z(n452) );
  NAND U1501 ( .A(rst), .B(\_MxM/Y0[23] ), .Z(n451) );
  NAND U1502 ( .A(n454), .B(n455), .Z(\_MxM/n352 ) );
  NAND U1503 ( .A(n456), .B(n384), .Z(n455) );
  NAND U1504 ( .A(rst), .B(\_MxM/Y0[24] ), .Z(n454) );
  NAND U1505 ( .A(n457), .B(n458), .Z(\_MxM/n351 ) );
  NAND U1506 ( .A(n459), .B(n384), .Z(n458) );
  NAND U1507 ( .A(rst), .B(\_MxM/Y0[25] ), .Z(n457) );
  NAND U1508 ( .A(n460), .B(n461), .Z(\_MxM/n350 ) );
  NAND U1509 ( .A(n462), .B(n384), .Z(n461) );
  NAND U1510 ( .A(rst), .B(\_MxM/Y0[26] ), .Z(n460) );
  NAND U1511 ( .A(n463), .B(n464), .Z(\_MxM/n349 ) );
  NAND U1512 ( .A(n465), .B(n384), .Z(n464) );
  NAND U1513 ( .A(rst), .B(\_MxM/Y0[27] ), .Z(n463) );
  NAND U1514 ( .A(n466), .B(n467), .Z(\_MxM/n348 ) );
  NAND U1515 ( .A(n468), .B(n384), .Z(n467) );
  NAND U1516 ( .A(rst), .B(\_MxM/Y0[28] ), .Z(n466) );
  NAND U1517 ( .A(n469), .B(n470), .Z(\_MxM/n347 ) );
  NAND U1518 ( .A(n471), .B(n384), .Z(n470) );
  NAND U1519 ( .A(rst), .B(\_MxM/Y0[29] ), .Z(n469) );
  NAND U1520 ( .A(n472), .B(n473), .Z(\_MxM/n346 ) );
  NAND U1521 ( .A(n474), .B(n384), .Z(n473) );
  NAND U1522 ( .A(rst), .B(\_MxM/Y0[30] ), .Z(n472) );
  NAND U1523 ( .A(n475), .B(n476), .Z(\_MxM/n345 ) );
  NAND U1524 ( .A(n477), .B(n384), .Z(n476) );
  NOR U1525 ( .A(rst), .B(n478), .Z(n384) );
  NAND U1526 ( .A(\_MxM/Y0[31] ), .B(rst), .Z(n475) );
  MUX U1527 ( .IN0(o[31]), .IN1(n477), .SEL(n479), .F(\_MxM/n344 ) );
  XNOR U1528 ( .A(\_MxM/Y0[31] ), .B(n481), .Z(n480) );
  AND U1529 ( .A(n484), .B(n485), .Z(n483) );
  XNOR U1530 ( .A(\_MxM/Y0[31] ), .B(n486), .Z(n485) );
  MUX U1531 ( .IN0(o[30]), .IN1(n474), .SEL(n479), .F(\_MxM/n343 ) );
  XOR U1532 ( .A(n484), .B(\_MxM/Y0[31] ), .Z(n474) );
  XOR U1533 ( .A(n486), .B(n481), .Z(n484) );
  XOR U1534 ( .A(n487), .B(n488), .Z(n481) );
  XOR U1535 ( .A(n489), .B(n490), .Z(n488) );
  AND U1536 ( .A(n491), .B(n492), .Z(n490) );
  XOR U1537 ( .A(n499), .B(n497), .Z(n487) );
  XOR U1538 ( .A(n500), .B(n501), .Z(n499) );
  XOR U1539 ( .A(n502), .B(n503), .Z(n501) );
  XOR U1540 ( .A(n507), .B(n508), .Z(n502) );
  ANDN U1541 ( .A(n509), .B(n510), .Z(n508) );
  XOR U1542 ( .A(n514), .B(n515), .Z(n500) );
  XOR U1543 ( .A(n504), .B(n506), .Z(n515) );
  XOR U1544 ( .A(n513), .B(n510), .Z(n514) );
  IV U1545 ( .A(n482), .Z(n486) );
  MUX U1546 ( .IN0(o[29]), .IN1(n471), .SEL(n479), .F(\_MxM/n342 ) );
  XOR U1547 ( .A(n517), .B(\_MxM/Y0[30] ), .Z(n471) );
  XNOR U1548 ( .A(n518), .B(n519), .Z(n517) );
  AND U1549 ( .A(n491), .B(n521), .Z(n520) );
  XNOR U1550 ( .A(n495), .B(n519), .Z(n521) );
  XOR U1551 ( .A(n493), .B(n519), .Z(n495) );
  XNOR U1552 ( .A(n498), .B(n496), .Z(n519) );
  IV U1553 ( .A(n497), .Z(n496) );
  XNOR U1554 ( .A(n504), .B(n505), .Z(n498) );
  XNOR U1555 ( .A(n506), .B(n509), .Z(n505) );
  XNOR U1556 ( .A(n510), .B(n525), .Z(n509) );
  XOR U1557 ( .A(n511), .B(n512), .Z(n525) );
  NAND U1558 ( .A(n526), .B(n527), .Z(n512) );
  IV U1559 ( .A(n513), .Z(n511) );
  IV U1560 ( .A(n494), .Z(n493) );
  MUX U1561 ( .IN0(o[28]), .IN1(n468), .SEL(n479), .F(\_MxM/n341 ) );
  XOR U1562 ( .A(n540), .B(\_MxM/Y0[29] ), .Z(n468) );
  XNOR U1563 ( .A(n541), .B(n542), .Z(n540) );
  AND U1564 ( .A(n491), .B(n544), .Z(n543) );
  XNOR U1565 ( .A(n538), .B(n542), .Z(n544) );
  XNOR U1566 ( .A(n524), .B(n523), .Z(n542) );
  IV U1567 ( .A(n522), .Z(n523) );
  XOR U1568 ( .A(n536), .B(n535), .Z(n524) );
  XOR U1569 ( .A(n534), .B(n548), .Z(n535) );
  XNOR U1570 ( .A(n533), .B(n532), .Z(n548) );
  XNOR U1571 ( .A(n549), .B(n550), .Z(n532) );
  IV U1572 ( .A(n531), .Z(n550) );
  XNOR U1573 ( .A(n529), .B(n530), .Z(n533) );
  NAND U1574 ( .A(n556), .B(n527), .Z(n530) );
  XNOR U1575 ( .A(n528), .B(n557), .Z(n529) );
  ANDN U1576 ( .A(n558), .B(n559), .Z(n557) );
  MUX U1577 ( .IN0(o[27]), .IN1(n465), .SEL(n479), .F(\_MxM/n340 ) );
  XOR U1578 ( .A(n569), .B(\_MxM/Y0[28] ), .Z(n465) );
  XNOR U1579 ( .A(n570), .B(n571), .Z(n569) );
  AND U1580 ( .A(n491), .B(n573), .Z(n572) );
  XNOR U1581 ( .A(n567), .B(n571), .Z(n573) );
  XNOR U1582 ( .A(n547), .B(n546), .Z(n571) );
  IV U1583 ( .A(n545), .Z(n546) );
  XOR U1584 ( .A(n565), .B(n564), .Z(n547) );
  XOR U1585 ( .A(n563), .B(n577), .Z(n564) );
  XNOR U1586 ( .A(n553), .B(n552), .Z(n577) );
  XOR U1587 ( .A(n582), .B(n554), .Z(n578) );
  AND U1588 ( .A(n583), .B(n526), .Z(n554) );
  IV U1589 ( .A(n551), .Z(n582) );
  XNOR U1590 ( .A(n561), .B(n562), .Z(n553) );
  NAND U1591 ( .A(n587), .B(n527), .Z(n562) );
  XNOR U1592 ( .A(n560), .B(n588), .Z(n561) );
  ANDN U1593 ( .A(n558), .B(n589), .Z(n588) );
  MUX U1594 ( .IN0(o[26]), .IN1(n462), .SEL(n479), .F(\_MxM/n339 ) );
  XOR U1595 ( .A(n600), .B(\_MxM/Y0[27] ), .Z(n462) );
  XNOR U1596 ( .A(n601), .B(n602), .Z(n600) );
  AND U1597 ( .A(n491), .B(n604), .Z(n603) );
  XNOR U1598 ( .A(n598), .B(n602), .Z(n604) );
  XNOR U1599 ( .A(n576), .B(n575), .Z(n602) );
  IV U1600 ( .A(n574), .Z(n575) );
  XNOR U1601 ( .A(n596), .B(n608), .Z(n576) );
  XOR U1602 ( .A(n595), .B(n594), .Z(n608) );
  XOR U1603 ( .A(n609), .B(n610), .Z(n594) );
  XOR U1604 ( .A(n611), .B(n612), .Z(n610) );
  XOR U1605 ( .A(n613), .B(n614), .Z(n612) );
  XNOR U1606 ( .A(n586), .B(n585), .Z(n595) );
  XOR U1607 ( .A(n622), .B(n580), .Z(n585) );
  XNOR U1608 ( .A(n579), .B(n623), .Z(n580) );
  ANDN U1609 ( .A(n624), .B(n559), .Z(n623) );
  AND U1610 ( .A(n556), .B(n583), .Z(n581) );
  XNOR U1611 ( .A(n591), .B(n592), .Z(n586) );
  NAND U1612 ( .A(n631), .B(n527), .Z(n592) );
  XNOR U1613 ( .A(n590), .B(n632), .Z(n591) );
  ANDN U1614 ( .A(n558), .B(n633), .Z(n632) );
  MUX U1615 ( .IN0(o[25]), .IN1(n459), .SEL(n479), .F(\_MxM/n338 ) );
  XOR U1616 ( .A(n641), .B(\_MxM/Y0[26] ), .Z(n459) );
  XNOR U1617 ( .A(n642), .B(n643), .Z(n641) );
  AND U1618 ( .A(n491), .B(n645), .Z(n644) );
  XNOR U1619 ( .A(n639), .B(n643), .Z(n645) );
  XNOR U1620 ( .A(n607), .B(n606), .Z(n643) );
  IV U1621 ( .A(n605), .Z(n606) );
  XOR U1622 ( .A(n637), .B(n649), .Z(n607) );
  XNOR U1623 ( .A(n621), .B(n620), .Z(n649) );
  XOR U1624 ( .A(n650), .B(n615), .Z(n620) );
  XOR U1625 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U1626 ( .B(n651), .A(n526), .Z(n617) );
  IV U1627 ( .A(n618), .Z(n616) );
  XOR U1628 ( .A(n611), .B(n619), .Z(n650) );
  XNOR U1629 ( .A(n630), .B(n629), .Z(n621) );
  XOR U1630 ( .A(n661), .B(n626), .Z(n629) );
  XNOR U1631 ( .A(n625), .B(n662), .Z(n626) );
  ANDN U1632 ( .A(n624), .B(n589), .Z(n662) );
  XOR U1633 ( .A(n663), .B(n664), .Z(n625) );
  AND U1634 ( .A(n665), .B(n666), .Z(n664) );
  XNOR U1635 ( .A(n667), .B(n663), .Z(n666) );
  AND U1636 ( .A(n587), .B(n583), .Z(n627) );
  XNOR U1637 ( .A(n635), .B(n636), .Z(n630) );
  NAND U1638 ( .A(n671), .B(n527), .Z(n636) );
  XNOR U1639 ( .A(n634), .B(n672), .Z(n635) );
  ANDN U1640 ( .A(n558), .B(n673), .Z(n672) );
  MUX U1641 ( .IN0(o[24]), .IN1(n456), .SEL(n479), .F(\_MxM/n337 ) );
  XOR U1642 ( .A(n681), .B(\_MxM/Y0[25] ), .Z(n456) );
  XNOR U1643 ( .A(n682), .B(n683), .Z(n681) );
  AND U1644 ( .A(n491), .B(n685), .Z(n684) );
  XNOR U1645 ( .A(n679), .B(n683), .Z(n685) );
  XNOR U1646 ( .A(n648), .B(n647), .Z(n683) );
  IV U1647 ( .A(n646), .Z(n647) );
  XOR U1648 ( .A(n677), .B(n689), .Z(n648) );
  XNOR U1649 ( .A(n657), .B(n656), .Z(n689) );
  XOR U1650 ( .A(n690), .B(n660), .Z(n656) );
  XNOR U1651 ( .A(n653), .B(n654), .Z(n660) );
  NANDN U1652 ( .B(n651), .A(n556), .Z(n654) );
  XNOR U1653 ( .A(n652), .B(n691), .Z(n653) );
  ANDN U1654 ( .A(n692), .B(n559), .Z(n691) );
  XNOR U1655 ( .A(n659), .B(n655), .Z(n690) );
  XNOR U1656 ( .A(n699), .B(n700), .Z(n659) );
  IV U1657 ( .A(n658), .Z(n700) );
  XNOR U1658 ( .A(n670), .B(n669), .Z(n657) );
  XOR U1659 ( .A(n707), .B(n665), .Z(n669) );
  XNOR U1660 ( .A(n663), .B(n708), .Z(n665) );
  ANDN U1661 ( .A(n624), .B(n633), .Z(n708) );
  AND U1662 ( .A(n631), .B(n583), .Z(n667) );
  XNOR U1663 ( .A(n675), .B(n676), .Z(n670) );
  NAND U1664 ( .A(n715), .B(n527), .Z(n676) );
  XNOR U1665 ( .A(n674), .B(n716), .Z(n675) );
  ANDN U1666 ( .A(n558), .B(n717), .Z(n716) );
  MUX U1667 ( .IN0(o[23]), .IN1(n453), .SEL(n479), .F(\_MxM/n336 ) );
  XOR U1668 ( .A(n725), .B(\_MxM/Y0[24] ), .Z(n453) );
  XNOR U1669 ( .A(n726), .B(n727), .Z(n725) );
  AND U1670 ( .A(n491), .B(n729), .Z(n728) );
  XNOR U1671 ( .A(n723), .B(n727), .Z(n729) );
  XNOR U1672 ( .A(n688), .B(n687), .Z(n727) );
  IV U1673 ( .A(n686), .Z(n687) );
  XOR U1674 ( .A(n721), .B(n732), .Z(n688) );
  XNOR U1675 ( .A(n698), .B(n697), .Z(n732) );
  XOR U1676 ( .A(n733), .B(n703), .Z(n697) );
  XNOR U1677 ( .A(n694), .B(n695), .Z(n703) );
  NANDN U1678 ( .B(n651), .A(n587), .Z(n695) );
  XNOR U1679 ( .A(n693), .B(n734), .Z(n694) );
  ANDN U1680 ( .A(n692), .B(n589), .Z(n734) );
  XNOR U1681 ( .A(n702), .B(n696), .Z(n733) );
  XNOR U1682 ( .A(n741), .B(n704), .Z(n702) );
  IV U1683 ( .A(n706), .Z(n704) );
  AND U1684 ( .A(n745), .B(n526), .Z(n705) );
  XNOR U1685 ( .A(n714), .B(n713), .Z(n698) );
  XOR U1686 ( .A(n749), .B(n710), .Z(n713) );
  XNOR U1687 ( .A(n709), .B(n750), .Z(n710) );
  ANDN U1688 ( .A(n624), .B(n673), .Z(n750) );
  AND U1689 ( .A(n671), .B(n583), .Z(n711) );
  XNOR U1690 ( .A(n719), .B(n720), .Z(n714) );
  NAND U1691 ( .A(n757), .B(n527), .Z(n720) );
  XNOR U1692 ( .A(n718), .B(n758), .Z(n719) );
  ANDN U1693 ( .A(n558), .B(n759), .Z(n758) );
  MUX U1694 ( .IN0(o[22]), .IN1(n450), .SEL(n479), .F(\_MxM/n335 ) );
  XOR U1695 ( .A(n769), .B(\_MxM/Y0[23] ), .Z(n450) );
  XNOR U1696 ( .A(n770), .B(n731), .Z(n769) );
  AND U1697 ( .A(n491), .B(n772), .Z(n771) );
  XNOR U1698 ( .A(n767), .B(n731), .Z(n772) );
  XOR U1699 ( .A(n730), .B(n773), .Z(n731) );
  XNOR U1700 ( .A(n765), .B(n764), .Z(n773) );
  XOR U1701 ( .A(n774), .B(n775), .Z(n764) );
  XOR U1702 ( .A(n776), .B(n777), .Z(n775) );
  XOR U1703 ( .A(n780), .B(n781), .Z(n776) );
  ANDN U1704 ( .A(n779), .B(n782), .Z(n781) );
  XNOR U1705 ( .A(n785), .B(n763), .Z(n774) );
  XOR U1706 ( .A(n784), .B(n782), .Z(n785) );
  XNOR U1707 ( .A(n740), .B(n739), .Z(n765) );
  XOR U1708 ( .A(n789), .B(n748), .Z(n739) );
  XNOR U1709 ( .A(n736), .B(n737), .Z(n748) );
  NANDN U1710 ( .B(n651), .A(n631), .Z(n737) );
  XNOR U1711 ( .A(n735), .B(n790), .Z(n736) );
  ANDN U1712 ( .A(n692), .B(n633), .Z(n790) );
  XNOR U1713 ( .A(n747), .B(n738), .Z(n789) );
  XOR U1714 ( .A(n797), .B(n743), .Z(n747) );
  XNOR U1715 ( .A(n742), .B(n798), .Z(n743) );
  ANDN U1716 ( .A(n799), .B(n559), .Z(n798) );
  XOR U1717 ( .A(n800), .B(n801), .Z(n742) );
  AND U1718 ( .A(n802), .B(n803), .Z(n801) );
  XNOR U1719 ( .A(n804), .B(n800), .Z(n803) );
  AND U1720 ( .A(n556), .B(n745), .Z(n744) );
  XNOR U1721 ( .A(n756), .B(n755), .Z(n740) );
  XOR U1722 ( .A(n808), .B(n752), .Z(n755) );
  XNOR U1723 ( .A(n751), .B(n809), .Z(n752) );
  ANDN U1724 ( .A(n624), .B(n717), .Z(n809) );
  AND U1725 ( .A(n715), .B(n583), .Z(n753) );
  XNOR U1726 ( .A(n761), .B(n762), .Z(n756) );
  NAND U1727 ( .A(n816), .B(n527), .Z(n762) );
  XNOR U1728 ( .A(n760), .B(n817), .Z(n761) );
  ANDN U1729 ( .A(n558), .B(n818), .Z(n817) );
  MUX U1730 ( .IN0(o[21]), .IN1(n447), .SEL(n479), .F(\_MxM/n334 ) );
  XOR U1731 ( .A(n828), .B(\_MxM/Y0[22] ), .Z(n447) );
  XNOR U1732 ( .A(n829), .B(n830), .Z(n828) );
  AND U1733 ( .A(n491), .B(n832), .Z(n831) );
  XNOR U1734 ( .A(n826), .B(n830), .Z(n832) );
  XNOR U1735 ( .A(n824), .B(n823), .Z(n830) );
  IV U1736 ( .A(n822), .Z(n823) );
  XNOR U1737 ( .A(n788), .B(n787), .Z(n824) );
  XOR U1738 ( .A(n836), .B(n779), .Z(n787) );
  XNOR U1739 ( .A(n782), .B(n837), .Z(n779) );
  NANDN U1740 ( .B(n838), .A(n526), .Z(n783) );
  XOR U1741 ( .A(n778), .B(n786), .Z(n836) );
  XNOR U1742 ( .A(n796), .B(n795), .Z(n788) );
  XOR U1743 ( .A(n850), .B(n807), .Z(n795) );
  XNOR U1744 ( .A(n792), .B(n793), .Z(n807) );
  NANDN U1745 ( .B(n651), .A(n671), .Z(n793) );
  XNOR U1746 ( .A(n791), .B(n851), .Z(n792) );
  ANDN U1747 ( .A(n692), .B(n673), .Z(n851) );
  XOR U1748 ( .A(n852), .B(n853), .Z(n791) );
  AND U1749 ( .A(n854), .B(n855), .Z(n853) );
  XOR U1750 ( .A(n856), .B(n852), .Z(n855) );
  XNOR U1751 ( .A(n806), .B(n794), .Z(n850) );
  XOR U1752 ( .A(n860), .B(n802), .Z(n806) );
  XNOR U1753 ( .A(n800), .B(n861), .Z(n802) );
  ANDN U1754 ( .A(n799), .B(n589), .Z(n861) );
  XOR U1755 ( .A(n862), .B(n863), .Z(n800) );
  AND U1756 ( .A(n864), .B(n865), .Z(n863) );
  XNOR U1757 ( .A(n866), .B(n862), .Z(n865) );
  AND U1758 ( .A(n587), .B(n745), .Z(n804) );
  XNOR U1759 ( .A(n815), .B(n814), .Z(n796) );
  XOR U1760 ( .A(n870), .B(n811), .Z(n814) );
  XNOR U1761 ( .A(n810), .B(n871), .Z(n811) );
  ANDN U1762 ( .A(n624), .B(n759), .Z(n871) );
  XOR U1763 ( .A(n872), .B(n873), .Z(n810) );
  AND U1764 ( .A(n874), .B(n875), .Z(n873) );
  XNOR U1765 ( .A(n876), .B(n872), .Z(n875) );
  AND U1766 ( .A(n757), .B(n583), .Z(n812) );
  XNOR U1767 ( .A(n820), .B(n821), .Z(n815) );
  NAND U1768 ( .A(n880), .B(n527), .Z(n821) );
  XNOR U1769 ( .A(n819), .B(n881), .Z(n820) );
  ANDN U1770 ( .A(n558), .B(n882), .Z(n881) );
  XOR U1771 ( .A(n883), .B(n884), .Z(n819) );
  AND U1772 ( .A(n885), .B(n886), .Z(n884) );
  XOR U1773 ( .A(n887), .B(n883), .Z(n886) );
  MUX U1774 ( .IN0(o[20]), .IN1(n444), .SEL(n479), .F(\_MxM/n333 ) );
  XOR U1775 ( .A(n891), .B(\_MxM/Y0[21] ), .Z(n444) );
  XNOR U1776 ( .A(n892), .B(n893), .Z(n891) );
  AND U1777 ( .A(n491), .B(n895), .Z(n894) );
  XNOR U1778 ( .A(n889), .B(n893), .Z(n895) );
  XNOR U1779 ( .A(n835), .B(n834), .Z(n893) );
  IV U1780 ( .A(n833), .Z(n834) );
  XNOR U1781 ( .A(n847), .B(n846), .Z(n835) );
  XOR U1782 ( .A(n899), .B(n849), .Z(n846) );
  XNOR U1783 ( .A(n844), .B(n843), .Z(n849) );
  XNOR U1784 ( .A(n900), .B(n901), .Z(n843) );
  IV U1785 ( .A(n842), .Z(n901) );
  XNOR U1786 ( .A(n840), .B(n841), .Z(n844) );
  NANDN U1787 ( .B(n838), .A(n556), .Z(n841) );
  XNOR U1788 ( .A(n839), .B(n907), .Z(n840) );
  ANDN U1789 ( .A(n908), .B(n559), .Z(n907) );
  XNOR U1790 ( .A(n859), .B(n858), .Z(n847) );
  XOR U1791 ( .A(n918), .B(n869), .Z(n858) );
  XNOR U1792 ( .A(n854), .B(n856), .Z(n869) );
  NANDN U1793 ( .B(n651), .A(n715), .Z(n856) );
  XNOR U1794 ( .A(n852), .B(n919), .Z(n854) );
  ANDN U1795 ( .A(n692), .B(n717), .Z(n919) );
  XOR U1796 ( .A(n920), .B(n921), .Z(n852) );
  AND U1797 ( .A(n922), .B(n923), .Z(n921) );
  XOR U1798 ( .A(n924), .B(n920), .Z(n923) );
  XNOR U1799 ( .A(n868), .B(n857), .Z(n918) );
  XOR U1800 ( .A(n928), .B(n864), .Z(n868) );
  XNOR U1801 ( .A(n862), .B(n929), .Z(n864) );
  ANDN U1802 ( .A(n799), .B(n633), .Z(n929) );
  XOR U1803 ( .A(n930), .B(n931), .Z(n862) );
  AND U1804 ( .A(n932), .B(n933), .Z(n931) );
  XNOR U1805 ( .A(n934), .B(n930), .Z(n933) );
  AND U1806 ( .A(n631), .B(n745), .Z(n866) );
  XNOR U1807 ( .A(n879), .B(n878), .Z(n859) );
  XOR U1808 ( .A(n938), .B(n874), .Z(n878) );
  XNOR U1809 ( .A(n872), .B(n939), .Z(n874) );
  ANDN U1810 ( .A(n624), .B(n818), .Z(n939) );
  XOR U1811 ( .A(n940), .B(n941), .Z(n872) );
  AND U1812 ( .A(n942), .B(n943), .Z(n941) );
  XNOR U1813 ( .A(n944), .B(n940), .Z(n943) );
  AND U1814 ( .A(n816), .B(n583), .Z(n876) );
  XNOR U1815 ( .A(n885), .B(n887), .Z(n879) );
  NAND U1816 ( .A(n948), .B(n527), .Z(n887) );
  XNOR U1817 ( .A(n883), .B(n949), .Z(n885) );
  ANDN U1818 ( .A(n558), .B(n950), .Z(n949) );
  XOR U1819 ( .A(n951), .B(n952), .Z(n883) );
  AND U1820 ( .A(n953), .B(n954), .Z(n952) );
  XOR U1821 ( .A(n955), .B(n951), .Z(n954) );
  MUX U1822 ( .IN0(o[19]), .IN1(n441), .SEL(n479), .F(\_MxM/n332 ) );
  XOR U1823 ( .A(n959), .B(\_MxM/Y0[20] ), .Z(n441) );
  XNOR U1824 ( .A(n960), .B(n961), .Z(n959) );
  AND U1825 ( .A(n491), .B(n963), .Z(n962) );
  XNOR U1826 ( .A(n957), .B(n961), .Z(n963) );
  XNOR U1827 ( .A(n898), .B(n897), .Z(n961) );
  IV U1828 ( .A(n896), .Z(n897) );
  XNOR U1829 ( .A(n914), .B(n913), .Z(n898) );
  XOR U1830 ( .A(n967), .B(n917), .Z(n913) );
  XNOR U1831 ( .A(n904), .B(n903), .Z(n917) );
  XOR U1832 ( .A(n972), .B(n905), .Z(n968) );
  AND U1833 ( .A(n973), .B(n526), .Z(n905) );
  IV U1834 ( .A(n902), .Z(n972) );
  XNOR U1835 ( .A(n910), .B(n911), .Z(n904) );
  NANDN U1836 ( .B(n838), .A(n587), .Z(n911) );
  XNOR U1837 ( .A(n909), .B(n977), .Z(n910) );
  ANDN U1838 ( .A(n908), .B(n589), .Z(n977) );
  XNOR U1839 ( .A(n916), .B(n912), .Z(n967) );
  IV U1840 ( .A(n915), .Z(n916) );
  XNOR U1841 ( .A(n927), .B(n926), .Z(n914) );
  XOR U1842 ( .A(n987), .B(n937), .Z(n926) );
  XNOR U1843 ( .A(n922), .B(n924), .Z(n937) );
  NANDN U1844 ( .B(n651), .A(n757), .Z(n924) );
  XNOR U1845 ( .A(n920), .B(n988), .Z(n922) );
  ANDN U1846 ( .A(n692), .B(n759), .Z(n988) );
  XOR U1847 ( .A(n989), .B(n990), .Z(n920) );
  AND U1848 ( .A(n991), .B(n992), .Z(n990) );
  XOR U1849 ( .A(n993), .B(n989), .Z(n992) );
  XNOR U1850 ( .A(n936), .B(n925), .Z(n987) );
  XOR U1851 ( .A(n997), .B(n932), .Z(n936) );
  XNOR U1852 ( .A(n930), .B(n998), .Z(n932) );
  ANDN U1853 ( .A(n799), .B(n673), .Z(n998) );
  XOR U1854 ( .A(n999), .B(n1000), .Z(n930) );
  AND U1855 ( .A(n1001), .B(n1002), .Z(n1000) );
  XNOR U1856 ( .A(n1003), .B(n999), .Z(n1002) );
  AND U1857 ( .A(n671), .B(n745), .Z(n934) );
  XNOR U1858 ( .A(n947), .B(n946), .Z(n927) );
  XOR U1859 ( .A(n1007), .B(n942), .Z(n946) );
  XNOR U1860 ( .A(n940), .B(n1008), .Z(n942) );
  ANDN U1861 ( .A(n624), .B(n882), .Z(n1008) );
  AND U1862 ( .A(n880), .B(n583), .Z(n944) );
  XNOR U1863 ( .A(n953), .B(n955), .Z(n947) );
  NAND U1864 ( .A(n1015), .B(n527), .Z(n955) );
  XNOR U1865 ( .A(n951), .B(n1016), .Z(n953) );
  ANDN U1866 ( .A(n558), .B(n1017), .Z(n1016) );
  XOR U1867 ( .A(n1018), .B(n1019), .Z(n951) );
  AND U1868 ( .A(n1020), .B(n1021), .Z(n1019) );
  XOR U1869 ( .A(n1022), .B(n1018), .Z(n1021) );
  MUX U1870 ( .IN0(o[18]), .IN1(n438), .SEL(n479), .F(\_MxM/n331 ) );
  XOR U1871 ( .A(n1026), .B(\_MxM/Y0[19] ), .Z(n438) );
  XNOR U1872 ( .A(n1027), .B(n1028), .Z(n1026) );
  AND U1873 ( .A(n491), .B(n1030), .Z(n1029) );
  XOR U1874 ( .A(n1024), .B(n1028), .Z(n1030) );
  XOR U1875 ( .A(n1023), .B(n1028), .Z(n1024) );
  XNOR U1876 ( .A(n966), .B(n965), .Z(n1028) );
  IV U1877 ( .A(n964), .Z(n965) );
  XNOR U1878 ( .A(n983), .B(n982), .Z(n966) );
  XOR U1879 ( .A(n1033), .B(n986), .Z(n982) );
  XNOR U1880 ( .A(n976), .B(n975), .Z(n986) );
  XOR U1881 ( .A(n1034), .B(n970), .Z(n975) );
  XNOR U1882 ( .A(n969), .B(n1035), .Z(n970) );
  ANDN U1883 ( .A(n1036), .B(n559), .Z(n1035) );
  XOR U1884 ( .A(n1037), .B(n1038), .Z(n969) );
  AND U1885 ( .A(n1039), .B(n1040), .Z(n1038) );
  XNOR U1886 ( .A(n1041), .B(n1037), .Z(n1040) );
  AND U1887 ( .A(n556), .B(n973), .Z(n971) );
  XNOR U1888 ( .A(n979), .B(n980), .Z(n976) );
  NANDN U1889 ( .B(n838), .A(n631), .Z(n980) );
  XNOR U1890 ( .A(n978), .B(n1045), .Z(n979) );
  ANDN U1891 ( .A(n908), .B(n633), .Z(n1045) );
  XNOR U1892 ( .A(n985), .B(n981), .Z(n1033) );
  XNOR U1893 ( .A(n1052), .B(n1053), .Z(n985) );
  IV U1894 ( .A(n984), .Z(n1053) );
  XNOR U1895 ( .A(n996), .B(n995), .Z(n983) );
  XOR U1896 ( .A(n1059), .B(n1006), .Z(n995) );
  XNOR U1897 ( .A(n991), .B(n993), .Z(n1006) );
  NANDN U1898 ( .B(n651), .A(n816), .Z(n993) );
  XNOR U1899 ( .A(n989), .B(n1060), .Z(n991) );
  ANDN U1900 ( .A(n692), .B(n818), .Z(n1060) );
  XOR U1901 ( .A(n1061), .B(n1062), .Z(n989) );
  AND U1902 ( .A(n1063), .B(n1064), .Z(n1062) );
  XOR U1903 ( .A(n1065), .B(n1061), .Z(n1064) );
  XNOR U1904 ( .A(n1005), .B(n994), .Z(n1059) );
  XOR U1905 ( .A(n1069), .B(n1001), .Z(n1005) );
  XNOR U1906 ( .A(n999), .B(n1070), .Z(n1001) );
  ANDN U1907 ( .A(n799), .B(n717), .Z(n1070) );
  XOR U1908 ( .A(n1071), .B(n1072), .Z(n999) );
  AND U1909 ( .A(n1073), .B(n1074), .Z(n1072) );
  XNOR U1910 ( .A(n1075), .B(n1071), .Z(n1074) );
  AND U1911 ( .A(n715), .B(n745), .Z(n1003) );
  XNOR U1912 ( .A(n1014), .B(n1013), .Z(n996) );
  XOR U1913 ( .A(n1079), .B(n1010), .Z(n1013) );
  XNOR U1914 ( .A(n1009), .B(n1080), .Z(n1010) );
  ANDN U1915 ( .A(n624), .B(n950), .Z(n1080) );
  XOR U1916 ( .A(n1081), .B(n1082), .Z(n1009) );
  AND U1917 ( .A(n1083), .B(n1084), .Z(n1082) );
  XNOR U1918 ( .A(n1085), .B(n1081), .Z(n1084) );
  AND U1919 ( .A(n948), .B(n583), .Z(n1011) );
  XNOR U1920 ( .A(n1020), .B(n1022), .Z(n1014) );
  NAND U1921 ( .A(n1089), .B(n527), .Z(n1022) );
  XNOR U1922 ( .A(n1018), .B(n1090), .Z(n1020) );
  ANDN U1923 ( .A(n558), .B(n1091), .Z(n1090) );
  NANDN U1924 ( .B(n1092), .A(n1093), .Z(n1018) );
  NAND U1925 ( .A(n1094), .B(n1095), .Z(n1093) );
  MUX U1926 ( .IN0(o[17]), .IN1(n435), .SEL(n479), .F(\_MxM/n330 ) );
  XOR U1927 ( .A(n1100), .B(\_MxM/Y0[18] ), .Z(n435) );
  XOR U1928 ( .A(n1101), .B(n1102), .Z(n1100) );
  AND U1929 ( .A(n491), .B(n1104), .Z(n1103) );
  XOR U1930 ( .A(n1098), .B(n1102), .Z(n1104) );
  XOR U1931 ( .A(n1097), .B(n1102), .Z(n1098) );
  XOR U1932 ( .A(n1032), .B(n1031), .Z(n1102) );
  XNOR U1933 ( .A(n1107), .B(n1056), .Z(n1050) );
  XNOR U1934 ( .A(n1044), .B(n1043), .Z(n1056) );
  XOR U1935 ( .A(n1108), .B(n1039), .Z(n1043) );
  XNOR U1936 ( .A(n1037), .B(n1109), .Z(n1039) );
  ANDN U1937 ( .A(n1036), .B(n589), .Z(n1109) );
  XOR U1938 ( .A(n1110), .B(n1111), .Z(n1037) );
  AND U1939 ( .A(n1112), .B(n1113), .Z(n1111) );
  XNOR U1940 ( .A(n1114), .B(n1110), .Z(n1113) );
  AND U1941 ( .A(n587), .B(n973), .Z(n1041) );
  XNOR U1942 ( .A(n1047), .B(n1048), .Z(n1044) );
  NANDN U1943 ( .B(n838), .A(n671), .Z(n1048) );
  XNOR U1944 ( .A(n1046), .B(n1118), .Z(n1047) );
  ANDN U1945 ( .A(n908), .B(n673), .Z(n1118) );
  XOR U1946 ( .A(n1119), .B(n1120), .Z(n1046) );
  AND U1947 ( .A(n1121), .B(n1122), .Z(n1120) );
  XOR U1948 ( .A(n1123), .B(n1119), .Z(n1122) );
  XNOR U1949 ( .A(n1055), .B(n1049), .Z(n1107) );
  XOR U1950 ( .A(n1127), .B(n1057), .Z(n1055) );
  NAND U1951 ( .A(n1131), .B(n1132), .Z(n1058) );
  NANDN U1952 ( .B(n1133), .A(n526), .Z(n1132) );
  NANDN U1953 ( .B(n1134), .A(n1135), .Z(n1131) );
  XNOR U1954 ( .A(n1068), .B(n1067), .Z(n1051) );
  XOR U1955 ( .A(n1139), .B(n1078), .Z(n1067) );
  XNOR U1956 ( .A(n1063), .B(n1065), .Z(n1078) );
  NANDN U1957 ( .B(n651), .A(n880), .Z(n1065) );
  XNOR U1958 ( .A(n1061), .B(n1140), .Z(n1063) );
  ANDN U1959 ( .A(n692), .B(n882), .Z(n1140) );
  XOR U1960 ( .A(n1141), .B(n1142), .Z(n1061) );
  AND U1961 ( .A(n1143), .B(n1144), .Z(n1142) );
  XOR U1962 ( .A(n1145), .B(n1141), .Z(n1144) );
  XNOR U1963 ( .A(n1077), .B(n1066), .Z(n1139) );
  XOR U1964 ( .A(n1149), .B(n1073), .Z(n1077) );
  XNOR U1965 ( .A(n1071), .B(n1150), .Z(n1073) );
  ANDN U1966 ( .A(n799), .B(n759), .Z(n1150) );
  XOR U1967 ( .A(n1151), .B(n1152), .Z(n1071) );
  AND U1968 ( .A(n1153), .B(n1154), .Z(n1152) );
  XNOR U1969 ( .A(n1155), .B(n1151), .Z(n1154) );
  AND U1970 ( .A(n757), .B(n745), .Z(n1075) );
  XOR U1971 ( .A(n1088), .B(n1087), .Z(n1068) );
  XOR U1972 ( .A(n1159), .B(n1083), .Z(n1087) );
  XNOR U1973 ( .A(n1081), .B(n1160), .Z(n1083) );
  ANDN U1974 ( .A(n624), .B(n1017), .Z(n1160) );
  AND U1975 ( .A(n1015), .B(n583), .Z(n1085) );
  XOR U1976 ( .A(n1095), .B(n1094), .Z(n1088) );
  NAND U1977 ( .A(n1167), .B(n527), .Z(n1094) );
  XNOR U1978 ( .A(n1092), .B(n1168), .Z(n1095) );
  ANDN U1979 ( .A(n558), .B(n1169), .Z(n1168) );
  NANDN U1980 ( .B(n1170), .A(n1171), .Z(n1092) );
  NAND U1981 ( .A(n1172), .B(n1173), .Z(n1171) );
  IV U1982 ( .A(n1096), .Z(n1097) );
  MUX U1983 ( .IN0(o[16]), .IN1(n432), .SEL(n479), .F(\_MxM/n329 ) );
  XOR U1984 ( .A(n1178), .B(\_MxM/Y0[17] ), .Z(n432) );
  XOR U1985 ( .A(n1179), .B(n1180), .Z(n1178) );
  AND U1986 ( .A(n491), .B(n1182), .Z(n1181) );
  XOR U1987 ( .A(n1176), .B(n1180), .Z(n1182) );
  XOR U1988 ( .A(n1175), .B(n1180), .Z(n1176) );
  XOR U1989 ( .A(n1106), .B(n1105), .Z(n1180) );
  XNOR U1990 ( .A(n1185), .B(n1138), .Z(n1125) );
  XNOR U1991 ( .A(n1117), .B(n1116), .Z(n1138) );
  XOR U1992 ( .A(n1186), .B(n1112), .Z(n1116) );
  XNOR U1993 ( .A(n1110), .B(n1187), .Z(n1112) );
  ANDN U1994 ( .A(n1036), .B(n633), .Z(n1187) );
  XOR U1995 ( .A(n1188), .B(n1189), .Z(n1110) );
  AND U1996 ( .A(n1190), .B(n1191), .Z(n1189) );
  XNOR U1997 ( .A(n1192), .B(n1188), .Z(n1191) );
  AND U1998 ( .A(n631), .B(n973), .Z(n1114) );
  XNOR U1999 ( .A(n1121), .B(n1123), .Z(n1117) );
  NANDN U2000 ( .B(n838), .A(n715), .Z(n1123) );
  XNOR U2001 ( .A(n1119), .B(n1196), .Z(n1121) );
  ANDN U2002 ( .A(n908), .B(n717), .Z(n1196) );
  XOR U2003 ( .A(n1197), .B(n1198), .Z(n1119) );
  AND U2004 ( .A(n1199), .B(n1200), .Z(n1198) );
  XOR U2005 ( .A(n1201), .B(n1197), .Z(n1200) );
  XOR U2006 ( .A(n1137), .B(n1124), .Z(n1185) );
  XNOR U2007 ( .A(n1205), .B(n1129), .Z(n1137) );
  XNOR U2008 ( .A(n1206), .B(n1135), .Z(n1129) );
  AND U2009 ( .A(n556), .B(n1207), .Z(n1135) );
  NAND U2010 ( .A(n1208), .B(n1134), .Z(n1206) );
  XOR U2011 ( .A(n1209), .B(n1210), .Z(n1134) );
  AND U2012 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR U2013 ( .A(n1213), .B(n1209), .Z(n1212) );
  NANDN U2014 ( .B(n559), .A(n1214), .Z(n1208) );
  XNOR U2015 ( .A(n1128), .B(n1136), .Z(n1205) );
  IV U2016 ( .A(n1130), .Z(n1128) );
  XNOR U2017 ( .A(n1148), .B(n1147), .Z(n1126) );
  XOR U2018 ( .A(n1220), .B(n1158), .Z(n1147) );
  XNOR U2019 ( .A(n1143), .B(n1145), .Z(n1158) );
  NANDN U2020 ( .B(n651), .A(n948), .Z(n1145) );
  XNOR U2021 ( .A(n1141), .B(n1221), .Z(n1143) );
  ANDN U2022 ( .A(n692), .B(n950), .Z(n1221) );
  XNOR U2023 ( .A(n1157), .B(n1146), .Z(n1220) );
  XOR U2024 ( .A(n1228), .B(n1153), .Z(n1157) );
  XNOR U2025 ( .A(n1151), .B(n1229), .Z(n1153) );
  ANDN U2026 ( .A(n799), .B(n818), .Z(n1229) );
  XOR U2027 ( .A(n1230), .B(n1231), .Z(n1151) );
  AND U2028 ( .A(n1232), .B(n1233), .Z(n1231) );
  XNOR U2029 ( .A(n1234), .B(n1230), .Z(n1233) );
  AND U2030 ( .A(n816), .B(n745), .Z(n1155) );
  XOR U2031 ( .A(n1166), .B(n1165), .Z(n1148) );
  XOR U2032 ( .A(n1238), .B(n1162), .Z(n1165) );
  XNOR U2033 ( .A(n1161), .B(n1239), .Z(n1162) );
  ANDN U2034 ( .A(n624), .B(n1091), .Z(n1239) );
  XOR U2035 ( .A(n1240), .B(n1241), .Z(n1161) );
  AND U2036 ( .A(n1242), .B(n1243), .Z(n1241) );
  XNOR U2037 ( .A(n1244), .B(n1240), .Z(n1243) );
  AND U2038 ( .A(n1089), .B(n583), .Z(n1163) );
  XOR U2039 ( .A(n1173), .B(n1172), .Z(n1166) );
  NAND U2040 ( .A(n1248), .B(n527), .Z(n1172) );
  XNOR U2041 ( .A(n1170), .B(n1249), .Z(n1173) );
  ANDN U2042 ( .A(n558), .B(n1250), .Z(n1249) );
  NAND U2043 ( .A(n1251), .B(n1252), .Z(n1170) );
  NAND U2044 ( .A(n1253), .B(n1254), .Z(n1251) );
  IV U2045 ( .A(n1174), .Z(n1175) );
  MUX U2046 ( .IN0(o[15]), .IN1(n429), .SEL(n479), .F(\_MxM/n328 ) );
  XOR U2047 ( .A(n1259), .B(\_MxM/Y0[16] ), .Z(n429) );
  XOR U2048 ( .A(n1260), .B(n1261), .Z(n1259) );
  AND U2049 ( .A(n491), .B(n1263), .Z(n1262) );
  XOR U2050 ( .A(n1257), .B(n1261), .Z(n1263) );
  XOR U2051 ( .A(n1256), .B(n1261), .Z(n1257) );
  XOR U2052 ( .A(n1184), .B(n1183), .Z(n1261) );
  XNOR U2053 ( .A(n1267), .B(n1217), .Z(n1203) );
  XNOR U2054 ( .A(n1195), .B(n1194), .Z(n1217) );
  XOR U2055 ( .A(n1268), .B(n1190), .Z(n1194) );
  XNOR U2056 ( .A(n1188), .B(n1269), .Z(n1190) );
  ANDN U2057 ( .A(n1036), .B(n673), .Z(n1269) );
  XOR U2058 ( .A(n1270), .B(n1271), .Z(n1188) );
  AND U2059 ( .A(n1272), .B(n1273), .Z(n1271) );
  XNOR U2060 ( .A(n1274), .B(n1270), .Z(n1273) );
  AND U2061 ( .A(n671), .B(n973), .Z(n1192) );
  XNOR U2062 ( .A(n1199), .B(n1201), .Z(n1195) );
  NANDN U2063 ( .B(n838), .A(n757), .Z(n1201) );
  XNOR U2064 ( .A(n1197), .B(n1278), .Z(n1199) );
  ANDN U2065 ( .A(n908), .B(n759), .Z(n1278) );
  XNOR U2066 ( .A(n1216), .B(n1202), .Z(n1267) );
  XOR U2067 ( .A(n1285), .B(n1219), .Z(n1216) );
  XNOR U2068 ( .A(n1211), .B(n1213), .Z(n1219) );
  NAND U2069 ( .A(n587), .B(n1207), .Z(n1213) );
  XNOR U2070 ( .A(n1209), .B(n1286), .Z(n1211) );
  ANDN U2071 ( .A(n1214), .B(n589), .Z(n1286) );
  XOR U2072 ( .A(n1287), .B(n1288), .Z(n1209) );
  AND U2073 ( .A(n1289), .B(n1290), .Z(n1288) );
  XOR U2074 ( .A(n1291), .B(n1287), .Z(n1290) );
  XNOR U2075 ( .A(n1218), .B(n1215), .Z(n1285) );
  AND U2076 ( .A(n1296), .B(n1297), .Z(n1295) );
  NANDN U2077 ( .B(n1298), .A(n526), .Z(n1297) );
  NANDN U2078 ( .B(n1299), .A(n1300), .Z(n1296) );
  XNOR U2079 ( .A(n1227), .B(n1226), .Z(n1204) );
  XOR U2080 ( .A(n1304), .B(n1237), .Z(n1226) );
  XNOR U2081 ( .A(n1223), .B(n1224), .Z(n1237) );
  NANDN U2082 ( .B(n651), .A(n1015), .Z(n1224) );
  XNOR U2083 ( .A(n1222), .B(n1305), .Z(n1223) );
  ANDN U2084 ( .A(n692), .B(n1017), .Z(n1305) );
  XNOR U2085 ( .A(n1236), .B(n1225), .Z(n1304) );
  XOR U2086 ( .A(n1312), .B(n1232), .Z(n1236) );
  XNOR U2087 ( .A(n1230), .B(n1313), .Z(n1232) );
  ANDN U2088 ( .A(n799), .B(n882), .Z(n1313) );
  XOR U2089 ( .A(n1314), .B(n1315), .Z(n1230) );
  AND U2090 ( .A(n1316), .B(n1317), .Z(n1315) );
  XNOR U2091 ( .A(n1318), .B(n1314), .Z(n1317) );
  AND U2092 ( .A(n880), .B(n745), .Z(n1234) );
  XOR U2093 ( .A(n1247), .B(n1246), .Z(n1227) );
  XOR U2094 ( .A(n1322), .B(n1242), .Z(n1246) );
  XNOR U2095 ( .A(n1240), .B(n1323), .Z(n1242) );
  ANDN U2096 ( .A(n624), .B(n1169), .Z(n1323) );
  XOR U2097 ( .A(n1324), .B(n1325), .Z(n1240) );
  AND U2098 ( .A(n1326), .B(n1327), .Z(n1325) );
  XNOR U2099 ( .A(n1328), .B(n1324), .Z(n1327) );
  AND U2100 ( .A(n1167), .B(n583), .Z(n1244) );
  XOR U2101 ( .A(n1254), .B(n1253), .Z(n1247) );
  NAND U2102 ( .A(n1332), .B(n527), .Z(n1253) );
  XOR U2103 ( .A(n1252), .B(n1333), .Z(n1254) );
  ANDN U2104 ( .A(n558), .B(n1334), .Z(n1333) );
  ANDN U2105 ( .A(n1335), .B(n1336), .Z(n1252) );
  NAND U2106 ( .A(n1337), .B(n1338), .Z(n1335) );
  IV U2107 ( .A(n1255), .Z(n1256) );
  MUX U2108 ( .IN0(o[14]), .IN1(n426), .SEL(n479), .F(\_MxM/n327 ) );
  XOR U2109 ( .A(n1343), .B(\_MxM/Y0[15] ), .Z(n426) );
  XOR U2110 ( .A(n1344), .B(n1345), .Z(n1343) );
  AND U2111 ( .A(n491), .B(n1347), .Z(n1346) );
  XOR U2112 ( .A(n1341), .B(n1345), .Z(n1347) );
  XOR U2113 ( .A(n1340), .B(n1345), .Z(n1341) );
  XNOR U2114 ( .A(n1266), .B(n1265), .Z(n1345) );
  XOR U2115 ( .A(n1348), .B(n1349), .Z(n1265) );
  XOR U2116 ( .A(n1350), .B(n1351), .Z(n1349) );
  XOR U2117 ( .A(n1352), .B(n1350), .Z(n1351) );
  XNOR U2118 ( .A(n1358), .B(n1294), .Z(n1283) );
  XNOR U2119 ( .A(n1277), .B(n1276), .Z(n1294) );
  XOR U2120 ( .A(n1359), .B(n1272), .Z(n1276) );
  XNOR U2121 ( .A(n1270), .B(n1360), .Z(n1272) );
  ANDN U2122 ( .A(n1036), .B(n717), .Z(n1360) );
  AND U2123 ( .A(n715), .B(n973), .Z(n1274) );
  XNOR U2124 ( .A(n1280), .B(n1281), .Z(n1277) );
  NANDN U2125 ( .B(n838), .A(n816), .Z(n1281) );
  XNOR U2126 ( .A(n1279), .B(n1367), .Z(n1280) );
  ANDN U2127 ( .A(n908), .B(n818), .Z(n1367) );
  XOR U2128 ( .A(n1368), .B(n1369), .Z(n1279) );
  AND U2129 ( .A(n1370), .B(n1371), .Z(n1369) );
  XOR U2130 ( .A(n1372), .B(n1368), .Z(n1371) );
  XNOR U2131 ( .A(n1293), .B(n1282), .Z(n1358) );
  XOR U2132 ( .A(n1376), .B(n1303), .Z(n1293) );
  XNOR U2133 ( .A(n1289), .B(n1291), .Z(n1303) );
  NAND U2134 ( .A(n631), .B(n1207), .Z(n1291) );
  XNOR U2135 ( .A(n1287), .B(n1377), .Z(n1289) );
  ANDN U2136 ( .A(n1214), .B(n633), .Z(n1377) );
  XOR U2137 ( .A(n1378), .B(n1379), .Z(n1287) );
  AND U2138 ( .A(n1380), .B(n1381), .Z(n1379) );
  XOR U2139 ( .A(n1382), .B(n1378), .Z(n1381) );
  XNOR U2140 ( .A(n1302), .B(n1292), .Z(n1376) );
  XOR U2141 ( .A(n1390), .B(n1300), .Z(n1386) );
  AND U2142 ( .A(n556), .B(n1391), .Z(n1300) );
  NAND U2143 ( .A(n1392), .B(n1299), .Z(n1390) );
  XOR U2144 ( .A(n1393), .B(n1394), .Z(n1299) );
  AND U2145 ( .A(n1395), .B(n1396), .Z(n1394) );
  XNOR U2146 ( .A(n1397), .B(n1393), .Z(n1396) );
  NANDN U2147 ( .B(n559), .A(n1398), .Z(n1392) );
  XNOR U2148 ( .A(n1311), .B(n1310), .Z(n1284) );
  XOR U2149 ( .A(n1399), .B(n1321), .Z(n1310) );
  XNOR U2150 ( .A(n1307), .B(n1308), .Z(n1321) );
  NANDN U2151 ( .B(n651), .A(n1089), .Z(n1308) );
  XNOR U2152 ( .A(n1306), .B(n1400), .Z(n1307) );
  ANDN U2153 ( .A(n692), .B(n1091), .Z(n1400) );
  XNOR U2154 ( .A(n1320), .B(n1309), .Z(n1399) );
  XOR U2155 ( .A(n1407), .B(n1316), .Z(n1320) );
  XNOR U2156 ( .A(n1314), .B(n1408), .Z(n1316) );
  ANDN U2157 ( .A(n799), .B(n950), .Z(n1408) );
  AND U2158 ( .A(n948), .B(n745), .Z(n1318) );
  XOR U2159 ( .A(n1331), .B(n1330), .Z(n1311) );
  XOR U2160 ( .A(n1415), .B(n1326), .Z(n1330) );
  XNOR U2161 ( .A(n1324), .B(n1416), .Z(n1326) );
  ANDN U2162 ( .A(n624), .B(n1250), .Z(n1416) );
  AND U2163 ( .A(n1248), .B(n583), .Z(n1328) );
  XOR U2164 ( .A(n1338), .B(n1337), .Z(n1331) );
  NAND U2165 ( .A(n1423), .B(n527), .Z(n1337) );
  XNOR U2166 ( .A(n1336), .B(n1424), .Z(n1338) );
  ANDN U2167 ( .A(n558), .B(n1425), .Z(n1424) );
  NAND U2168 ( .A(n1426), .B(n1427), .Z(n1336) );
  NAND U2169 ( .A(n1428), .B(n1429), .Z(n1426) );
  IV U2170 ( .A(n1339), .Z(n1340) );
  MUX U2171 ( .IN0(o[13]), .IN1(n423), .SEL(n479), .F(\_MxM/n326 ) );
  XOR U2172 ( .A(n1434), .B(\_MxM/Y0[14] ), .Z(n423) );
  XOR U2173 ( .A(n1435), .B(n1436), .Z(n1434) );
  AND U2174 ( .A(n491), .B(n1438), .Z(n1437) );
  XOR U2175 ( .A(n1432), .B(n1436), .Z(n1438) );
  XOR U2176 ( .A(n1431), .B(n1436), .Z(n1432) );
  XOR U2177 ( .A(n1439), .B(n1353), .Z(n1356) );
  NAND U2178 ( .A(n1350), .B(n1443), .Z(n1354) );
  AND U2179 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U2180 ( .B(n1446), .A(n526), .Z(n1445) );
  NANDN U2181 ( .B(n1447), .A(n1448), .Z(n1444) );
  AND U2182 ( .A(n1449), .B(n1450), .Z(n1350) );
  NANDN U2183 ( .B(n1451), .A(n1452), .Z(n1450) );
  OR U2184 ( .A(n1453), .B(n1454), .Z(n1449) );
  XNOR U2185 ( .A(n1375), .B(n1374), .Z(n1357) );
  XOR U2186 ( .A(n1458), .B(n1385), .Z(n1374) );
  XNOR U2187 ( .A(n1366), .B(n1365), .Z(n1385) );
  XOR U2188 ( .A(n1459), .B(n1362), .Z(n1365) );
  XNOR U2189 ( .A(n1361), .B(n1460), .Z(n1362) );
  ANDN U2190 ( .A(n1036), .B(n759), .Z(n1460) );
  XOR U2191 ( .A(n1461), .B(n1462), .Z(n1361) );
  AND U2192 ( .A(n1463), .B(n1464), .Z(n1462) );
  XNOR U2193 ( .A(n1465), .B(n1461), .Z(n1464) );
  AND U2194 ( .A(n757), .B(n973), .Z(n1363) );
  XNOR U2195 ( .A(n1370), .B(n1372), .Z(n1366) );
  NANDN U2196 ( .B(n838), .A(n880), .Z(n1372) );
  XNOR U2197 ( .A(n1368), .B(n1469), .Z(n1370) );
  ANDN U2198 ( .A(n908), .B(n882), .Z(n1469) );
  XNOR U2199 ( .A(n1384), .B(n1373), .Z(n1458) );
  XOR U2200 ( .A(n1476), .B(n1389), .Z(n1384) );
  XNOR U2201 ( .A(n1380), .B(n1382), .Z(n1389) );
  NAND U2202 ( .A(n671), .B(n1207), .Z(n1382) );
  XNOR U2203 ( .A(n1378), .B(n1477), .Z(n1380) );
  ANDN U2204 ( .A(n1214), .B(n673), .Z(n1477) );
  XOR U2205 ( .A(n1478), .B(n1479), .Z(n1378) );
  AND U2206 ( .A(n1480), .B(n1481), .Z(n1479) );
  XOR U2207 ( .A(n1482), .B(n1478), .Z(n1481) );
  XNOR U2208 ( .A(n1388), .B(n1383), .Z(n1476) );
  XOR U2209 ( .A(n1486), .B(n1395), .Z(n1388) );
  XNOR U2210 ( .A(n1393), .B(n1487), .Z(n1395) );
  ANDN U2211 ( .A(n1398), .B(n589), .Z(n1487) );
  XOR U2212 ( .A(n1488), .B(n1489), .Z(n1393) );
  AND U2213 ( .A(n1490), .B(n1491), .Z(n1489) );
  XNOR U2214 ( .A(n1492), .B(n1488), .Z(n1491) );
  AND U2215 ( .A(n587), .B(n1391), .Z(n1397) );
  XNOR U2216 ( .A(n1406), .B(n1405), .Z(n1375) );
  XOR U2217 ( .A(n1496), .B(n1414), .Z(n1405) );
  XNOR U2218 ( .A(n1402), .B(n1403), .Z(n1414) );
  NANDN U2219 ( .B(n651), .A(n1167), .Z(n1403) );
  XNOR U2220 ( .A(n1401), .B(n1497), .Z(n1402) );
  ANDN U2221 ( .A(n692), .B(n1169), .Z(n1497) );
  XNOR U2222 ( .A(n1413), .B(n1404), .Z(n1496) );
  XOR U2223 ( .A(n1504), .B(n1410), .Z(n1413) );
  XNOR U2224 ( .A(n1409), .B(n1505), .Z(n1410) );
  ANDN U2225 ( .A(n799), .B(n1017), .Z(n1505) );
  AND U2226 ( .A(n1015), .B(n745), .Z(n1411) );
  XOR U2227 ( .A(n1422), .B(n1421), .Z(n1406) );
  XOR U2228 ( .A(n1512), .B(n1418), .Z(n1421) );
  XNOR U2229 ( .A(n1417), .B(n1513), .Z(n1418) );
  ANDN U2230 ( .A(n624), .B(n1334), .Z(n1513) );
  AND U2231 ( .A(n1332), .B(n583), .Z(n1419) );
  XOR U2232 ( .A(n1429), .B(n1428), .Z(n1422) );
  NAND U2233 ( .A(n1520), .B(n527), .Z(n1428) );
  XOR U2234 ( .A(n1427), .B(n1521), .Z(n1429) );
  ANDN U2235 ( .A(n558), .B(n1522), .Z(n1521) );
  ANDN U2236 ( .A(n1523), .B(n1524), .Z(n1427) );
  NAND U2237 ( .A(n1525), .B(n1526), .Z(n1523) );
  IV U2238 ( .A(n1430), .Z(n1431) );
  MUX U2239 ( .IN0(o[12]), .IN1(n420), .SEL(n479), .F(\_MxM/n325 ) );
  XOR U2240 ( .A(n1531), .B(\_MxM/Y0[13] ), .Z(n420) );
  XNOR U2241 ( .A(n1532), .B(n1533), .Z(n1531) );
  AND U2242 ( .A(n491), .B(n1535), .Z(n1534) );
  XNOR U2243 ( .A(n1529), .B(n1533), .Z(n1535) );
  XNOR U2244 ( .A(n1528), .B(n1533), .Z(n1529) );
  XNOR U2245 ( .A(n1457), .B(n1456), .Z(n1533) );
  XOR U2246 ( .A(n1536), .B(n1441), .Z(n1456) );
  NANDN U2247 ( .B(n1537), .A(n1538), .Z(n1447) );
  XOR U2248 ( .A(n1541), .B(n1454), .Z(n1451) );
  NAND U2249 ( .A(n1542), .B(n556), .Z(n1454) );
  NAND U2250 ( .A(n1543), .B(n1453), .Z(n1541) );
  NANDN U2251 ( .B(n559), .A(n1547), .Z(n1543) );
  XNOR U2252 ( .A(n1440), .B(n1455), .Z(n1536) );
  IV U2253 ( .A(n1442), .Z(n1440) );
  XNOR U2254 ( .A(n1475), .B(n1474), .Z(n1457) );
  XOR U2255 ( .A(n1554), .B(n1485), .Z(n1474) );
  XNOR U2256 ( .A(n1468), .B(n1467), .Z(n1485) );
  XOR U2257 ( .A(n1555), .B(n1463), .Z(n1467) );
  XNOR U2258 ( .A(n1461), .B(n1556), .Z(n1463) );
  ANDN U2259 ( .A(n1036), .B(n818), .Z(n1556) );
  XOR U2260 ( .A(n1557), .B(n1558), .Z(n1461) );
  AND U2261 ( .A(n1559), .B(n1560), .Z(n1558) );
  XNOR U2262 ( .A(n1561), .B(n1557), .Z(n1560) );
  AND U2263 ( .A(n816), .B(n973), .Z(n1465) );
  XNOR U2264 ( .A(n1471), .B(n1472), .Z(n1468) );
  NANDN U2265 ( .B(n838), .A(n948), .Z(n1472) );
  XNOR U2266 ( .A(n1470), .B(n1565), .Z(n1471) );
  ANDN U2267 ( .A(n908), .B(n950), .Z(n1565) );
  XNOR U2268 ( .A(n1484), .B(n1473), .Z(n1554) );
  XOR U2269 ( .A(n1572), .B(n1495), .Z(n1484) );
  XNOR U2270 ( .A(n1480), .B(n1482), .Z(n1495) );
  NAND U2271 ( .A(n715), .B(n1207), .Z(n1482) );
  XNOR U2272 ( .A(n1478), .B(n1573), .Z(n1480) );
  ANDN U2273 ( .A(n1214), .B(n717), .Z(n1573) );
  XOR U2274 ( .A(n1574), .B(n1575), .Z(n1478) );
  AND U2275 ( .A(n1576), .B(n1577), .Z(n1575) );
  XOR U2276 ( .A(n1578), .B(n1574), .Z(n1577) );
  XNOR U2277 ( .A(n1494), .B(n1483), .Z(n1572) );
  XOR U2278 ( .A(n1582), .B(n1490), .Z(n1494) );
  XNOR U2279 ( .A(n1488), .B(n1583), .Z(n1490) );
  ANDN U2280 ( .A(n1398), .B(n633), .Z(n1583) );
  XOR U2281 ( .A(n1584), .B(n1585), .Z(n1488) );
  AND U2282 ( .A(n1586), .B(n1587), .Z(n1585) );
  XNOR U2283 ( .A(n1588), .B(n1584), .Z(n1587) );
  AND U2284 ( .A(n631), .B(n1391), .Z(n1492) );
  XNOR U2285 ( .A(n1503), .B(n1502), .Z(n1475) );
  XOR U2286 ( .A(n1592), .B(n1511), .Z(n1502) );
  XNOR U2287 ( .A(n1499), .B(n1500), .Z(n1511) );
  NANDN U2288 ( .B(n651), .A(n1248), .Z(n1500) );
  XNOR U2289 ( .A(n1498), .B(n1593), .Z(n1499) );
  ANDN U2290 ( .A(n692), .B(n1250), .Z(n1593) );
  XNOR U2291 ( .A(n1510), .B(n1501), .Z(n1592) );
  XOR U2292 ( .A(n1600), .B(n1507), .Z(n1510) );
  XNOR U2293 ( .A(n1506), .B(n1601), .Z(n1507) );
  ANDN U2294 ( .A(n799), .B(n1091), .Z(n1601) );
  AND U2295 ( .A(n1089), .B(n745), .Z(n1508) );
  XOR U2296 ( .A(n1519), .B(n1518), .Z(n1503) );
  XOR U2297 ( .A(n1608), .B(n1515), .Z(n1518) );
  XNOR U2298 ( .A(n1514), .B(n1609), .Z(n1515) );
  ANDN U2299 ( .A(n624), .B(n1425), .Z(n1609) );
  AND U2300 ( .A(n1423), .B(n583), .Z(n1516) );
  XOR U2301 ( .A(n1526), .B(n1525), .Z(n1519) );
  NAND U2302 ( .A(n1616), .B(n527), .Z(n1525) );
  XNOR U2303 ( .A(n1524), .B(n1617), .Z(n1526) );
  ANDN U2304 ( .A(n558), .B(n1618), .Z(n1617) );
  NAND U2305 ( .A(n1619), .B(n1620), .Z(n1524) );
  NAND U2306 ( .A(n1621), .B(n1622), .Z(n1619) );
  IV U2307 ( .A(n1527), .Z(n1528) );
  MUX U2308 ( .IN0(o[11]), .IN1(n417), .SEL(n479), .F(\_MxM/n324 ) );
  XOR U2309 ( .A(n1627), .B(\_MxM/Y0[12] ), .Z(n417) );
  XOR U2310 ( .A(n1628), .B(n1629), .Z(n1627) );
  AND U2311 ( .A(n491), .B(n1631), .Z(n1630) );
  XOR U2312 ( .A(n1625), .B(n1629), .Z(n1631) );
  XOR U2313 ( .A(n1624), .B(n1629), .Z(n1625) );
  XNOR U2314 ( .A(n1632), .B(n1553), .Z(n1549) );
  XOR U2315 ( .A(n1538), .B(n1537), .Z(n1553) );
  NANDN U2316 ( .B(n1633), .A(n1634), .Z(n1537) );
  AND U2317 ( .A(n1636), .B(n1637), .Z(n1635) );
  NANDN U2318 ( .B(n1638), .A(n526), .Z(n1637) );
  NANDN U2319 ( .B(n1639), .A(n1640), .Z(n1636) );
  XNOR U2320 ( .A(n1545), .B(n1546), .Z(n1540) );
  NAND U2321 ( .A(n1542), .B(n587), .Z(n1546) );
  XNOR U2322 ( .A(n1544), .B(n1644), .Z(n1545) );
  ANDN U2323 ( .A(n1547), .B(n589), .Z(n1644) );
  XNOR U2324 ( .A(n1552), .B(n1548), .Z(n1632) );
  IV U2325 ( .A(n1551), .Z(n1552) );
  XNOR U2326 ( .A(n1571), .B(n1570), .Z(n1550) );
  XOR U2327 ( .A(n1654), .B(n1581), .Z(n1570) );
  XNOR U2328 ( .A(n1564), .B(n1563), .Z(n1581) );
  XOR U2329 ( .A(n1655), .B(n1559), .Z(n1563) );
  XNOR U2330 ( .A(n1557), .B(n1656), .Z(n1559) );
  ANDN U2331 ( .A(n1036), .B(n882), .Z(n1656) );
  AND U2332 ( .A(n880), .B(n973), .Z(n1561) );
  XNOR U2333 ( .A(n1567), .B(n1568), .Z(n1564) );
  NANDN U2334 ( .B(n838), .A(n1015), .Z(n1568) );
  XNOR U2335 ( .A(n1566), .B(n1663), .Z(n1567) );
  ANDN U2336 ( .A(n908), .B(n1017), .Z(n1663) );
  XNOR U2337 ( .A(n1580), .B(n1569), .Z(n1654) );
  XOR U2338 ( .A(n1670), .B(n1591), .Z(n1580) );
  XNOR U2339 ( .A(n1576), .B(n1578), .Z(n1591) );
  NAND U2340 ( .A(n757), .B(n1207), .Z(n1578) );
  XNOR U2341 ( .A(n1574), .B(n1671), .Z(n1576) );
  ANDN U2342 ( .A(n1214), .B(n759), .Z(n1671) );
  XNOR U2343 ( .A(n1590), .B(n1579), .Z(n1670) );
  XOR U2344 ( .A(n1678), .B(n1586), .Z(n1590) );
  XNOR U2345 ( .A(n1584), .B(n1679), .Z(n1586) );
  ANDN U2346 ( .A(n1398), .B(n673), .Z(n1679) );
  XOR U2347 ( .A(n1680), .B(n1681), .Z(n1584) );
  AND U2348 ( .A(n1682), .B(n1683), .Z(n1681) );
  XNOR U2349 ( .A(n1684), .B(n1680), .Z(n1683) );
  AND U2350 ( .A(n671), .B(n1391), .Z(n1588) );
  XNOR U2351 ( .A(n1599), .B(n1598), .Z(n1571) );
  XOR U2352 ( .A(n1688), .B(n1607), .Z(n1598) );
  XNOR U2353 ( .A(n1595), .B(n1596), .Z(n1607) );
  NANDN U2354 ( .B(n651), .A(n1332), .Z(n1596) );
  XNOR U2355 ( .A(n1594), .B(n1689), .Z(n1595) );
  ANDN U2356 ( .A(n692), .B(n1334), .Z(n1689) );
  XNOR U2357 ( .A(n1606), .B(n1597), .Z(n1688) );
  XOR U2358 ( .A(n1696), .B(n1603), .Z(n1606) );
  XNOR U2359 ( .A(n1602), .B(n1697), .Z(n1603) );
  ANDN U2360 ( .A(n799), .B(n1169), .Z(n1697) );
  AND U2361 ( .A(n1167), .B(n745), .Z(n1604) );
  XOR U2362 ( .A(n1615), .B(n1614), .Z(n1599) );
  XOR U2363 ( .A(n1704), .B(n1611), .Z(n1614) );
  XNOR U2364 ( .A(n1610), .B(n1705), .Z(n1611) );
  ANDN U2365 ( .A(n624), .B(n1522), .Z(n1705) );
  AND U2366 ( .A(n1520), .B(n583), .Z(n1612) );
  XOR U2367 ( .A(n1622), .B(n1621), .Z(n1615) );
  NAND U2368 ( .A(n1712), .B(n527), .Z(n1621) );
  XOR U2369 ( .A(n1620), .B(n1713), .Z(n1622) );
  ANDN U2370 ( .A(n558), .B(n1714), .Z(n1713) );
  ANDN U2371 ( .A(n1715), .B(n1716), .Z(n1620) );
  NAND U2372 ( .A(n1717), .B(n1718), .Z(n1715) );
  IV U2373 ( .A(n1623), .Z(n1624) );
  MUX U2374 ( .IN0(o[10]), .IN1(n414), .SEL(n479), .F(\_MxM/n323 ) );
  XOR U2375 ( .A(n1723), .B(\_MxM/Y0[11] ), .Z(n414) );
  XNOR U2376 ( .A(n1724), .B(n1725), .Z(n1723) );
  AND U2377 ( .A(n491), .B(n1727), .Z(n1726) );
  XNOR U2378 ( .A(n1721), .B(n1725), .Z(n1727) );
  XNOR U2379 ( .A(n1720), .B(n1725), .Z(n1721) );
  XNOR U2380 ( .A(n1650), .B(n1649), .Z(n1725) );
  XOR U2381 ( .A(n1728), .B(n1653), .Z(n1649) );
  XOR U2382 ( .A(n1643), .B(n1642), .Z(n1633) );
  XOR U2383 ( .A(n1736), .B(n1640), .Z(n1732) );
  AND U2384 ( .A(n1737), .B(n556), .Z(n1640) );
  NAND U2385 ( .A(n1738), .B(n1639), .Z(n1736) );
  XOR U2386 ( .A(n1739), .B(n1740), .Z(n1639) );
  AND U2387 ( .A(n1741), .B(n1742), .Z(n1740) );
  XNOR U2388 ( .A(n1743), .B(n1739), .Z(n1742) );
  NANDN U2389 ( .B(n559), .A(n1744), .Z(n1738) );
  XNOR U2390 ( .A(n1646), .B(n1647), .Z(n1643) );
  NAND U2391 ( .A(n1542), .B(n631), .Z(n1647) );
  XNOR U2392 ( .A(n1645), .B(n1745), .Z(n1646) );
  ANDN U2393 ( .A(n1547), .B(n633), .Z(n1745) );
  XNOR U2394 ( .A(n1652), .B(n1648), .Z(n1728) );
  IV U2395 ( .A(n1651), .Z(n1652) );
  XNOR U2396 ( .A(n1669), .B(n1668), .Z(n1650) );
  XOR U2397 ( .A(n1755), .B(n1677), .Z(n1668) );
  XNOR U2398 ( .A(n1662), .B(n1661), .Z(n1677) );
  XOR U2399 ( .A(n1756), .B(n1658), .Z(n1661) );
  XNOR U2400 ( .A(n1657), .B(n1757), .Z(n1658) );
  ANDN U2401 ( .A(n1036), .B(n950), .Z(n1757) );
  AND U2402 ( .A(n948), .B(n973), .Z(n1659) );
  XNOR U2403 ( .A(n1665), .B(n1666), .Z(n1662) );
  NANDN U2404 ( .B(n838), .A(n1089), .Z(n1666) );
  XNOR U2405 ( .A(n1664), .B(n1764), .Z(n1665) );
  ANDN U2406 ( .A(n908), .B(n1091), .Z(n1764) );
  XNOR U2407 ( .A(n1676), .B(n1667), .Z(n1755) );
  XOR U2408 ( .A(n1771), .B(n1687), .Z(n1676) );
  XNOR U2409 ( .A(n1673), .B(n1674), .Z(n1687) );
  NAND U2410 ( .A(n816), .B(n1207), .Z(n1674) );
  XNOR U2411 ( .A(n1672), .B(n1772), .Z(n1673) );
  ANDN U2412 ( .A(n1214), .B(n818), .Z(n1772) );
  XNOR U2413 ( .A(n1686), .B(n1675), .Z(n1771) );
  XOR U2414 ( .A(n1779), .B(n1682), .Z(n1686) );
  XNOR U2415 ( .A(n1680), .B(n1780), .Z(n1682) );
  ANDN U2416 ( .A(n1398), .B(n717), .Z(n1780) );
  XOR U2417 ( .A(n1781), .B(n1782), .Z(n1680) );
  AND U2418 ( .A(n1783), .B(n1784), .Z(n1782) );
  XNOR U2419 ( .A(n1785), .B(n1781), .Z(n1784) );
  AND U2420 ( .A(n715), .B(n1391), .Z(n1684) );
  XNOR U2421 ( .A(n1695), .B(n1694), .Z(n1669) );
  XOR U2422 ( .A(n1789), .B(n1703), .Z(n1694) );
  XNOR U2423 ( .A(n1691), .B(n1692), .Z(n1703) );
  NANDN U2424 ( .B(n651), .A(n1423), .Z(n1692) );
  XNOR U2425 ( .A(n1690), .B(n1790), .Z(n1691) );
  ANDN U2426 ( .A(n692), .B(n1425), .Z(n1790) );
  XNOR U2427 ( .A(n1702), .B(n1693), .Z(n1789) );
  XOR U2428 ( .A(n1797), .B(n1699), .Z(n1702) );
  XNOR U2429 ( .A(n1698), .B(n1798), .Z(n1699) );
  ANDN U2430 ( .A(n799), .B(n1250), .Z(n1798) );
  AND U2431 ( .A(n1248), .B(n745), .Z(n1700) );
  XOR U2432 ( .A(n1711), .B(n1710), .Z(n1695) );
  XOR U2433 ( .A(n1805), .B(n1707), .Z(n1710) );
  XNOR U2434 ( .A(n1706), .B(n1806), .Z(n1707) );
  ANDN U2435 ( .A(n624), .B(n1618), .Z(n1806) );
  AND U2436 ( .A(n1616), .B(n583), .Z(n1708) );
  XOR U2437 ( .A(n1718), .B(n1717), .Z(n1711) );
  NAND U2438 ( .A(n1813), .B(n527), .Z(n1717) );
  XNOR U2439 ( .A(n1716), .B(n1814), .Z(n1718) );
  ANDN U2440 ( .A(n558), .B(n1815), .Z(n1814) );
  NAND U2441 ( .A(n1816), .B(n1817), .Z(n1716) );
  NAND U2442 ( .A(n1818), .B(n1819), .Z(n1816) );
  IV U2443 ( .A(n1719), .Z(n1720) );
  MUX U2444 ( .IN0(o[9]), .IN1(n411), .SEL(n479), .F(\_MxM/n322 ) );
  XOR U2445 ( .A(n1824), .B(\_MxM/Y0[10] ), .Z(n411) );
  XOR U2446 ( .A(n1825), .B(n1826), .Z(n1824) );
  AND U2447 ( .A(n491), .B(n1828), .Z(n1827) );
  XOR U2448 ( .A(n1822), .B(n1826), .Z(n1828) );
  XOR U2449 ( .A(n1821), .B(n1826), .Z(n1822) );
  XNOR U2450 ( .A(n1829), .B(n1754), .Z(n1750) );
  XNOR U2451 ( .A(n1731), .B(n1730), .Z(n1754) );
  XOR U2452 ( .A(n1729), .B(n1830), .Z(n1730) );
  AND U2453 ( .A(n1831), .B(n1832), .Z(n1830) );
  NANDN U2454 ( .B(n1833), .A(n1834), .Z(n1832) );
  AND U2455 ( .A(n1835), .B(n1836), .Z(n1831) );
  NANDN U2456 ( .B(n1837), .A(n526), .Z(n1836) );
  OR U2457 ( .A(n1838), .B(n1839), .Z(n1835) );
  XNOR U2458 ( .A(n1735), .B(n1734), .Z(n1731) );
  XOR U2459 ( .A(n1843), .B(n1741), .Z(n1734) );
  XNOR U2460 ( .A(n1739), .B(n1844), .Z(n1741) );
  ANDN U2461 ( .A(n1744), .B(n589), .Z(n1844) );
  XOR U2462 ( .A(n1845), .B(n1846), .Z(n1739) );
  AND U2463 ( .A(n1847), .B(n1848), .Z(n1846) );
  XNOR U2464 ( .A(n1849), .B(n1845), .Z(n1848) );
  AND U2465 ( .A(n1737), .B(n587), .Z(n1743) );
  XNOR U2466 ( .A(n1747), .B(n1748), .Z(n1735) );
  NAND U2467 ( .A(n1542), .B(n671), .Z(n1748) );
  XNOR U2468 ( .A(n1746), .B(n1853), .Z(n1747) );
  ANDN U2469 ( .A(n1547), .B(n673), .Z(n1853) );
  XNOR U2470 ( .A(n1753), .B(n1749), .Z(n1829) );
  IV U2471 ( .A(n1752), .Z(n1753) );
  XNOR U2472 ( .A(n1770), .B(n1769), .Z(n1751) );
  XOR U2473 ( .A(n1863), .B(n1778), .Z(n1769) );
  XNOR U2474 ( .A(n1763), .B(n1762), .Z(n1778) );
  XOR U2475 ( .A(n1864), .B(n1759), .Z(n1762) );
  XNOR U2476 ( .A(n1758), .B(n1865), .Z(n1759) );
  ANDN U2477 ( .A(n1036), .B(n1017), .Z(n1865) );
  AND U2478 ( .A(n1015), .B(n973), .Z(n1760) );
  XNOR U2479 ( .A(n1766), .B(n1767), .Z(n1763) );
  NANDN U2480 ( .B(n838), .A(n1167), .Z(n1767) );
  XNOR U2481 ( .A(n1765), .B(n1872), .Z(n1766) );
  ANDN U2482 ( .A(n908), .B(n1169), .Z(n1872) );
  XNOR U2483 ( .A(n1777), .B(n1768), .Z(n1863) );
  XOR U2484 ( .A(n1879), .B(n1788), .Z(n1777) );
  XNOR U2485 ( .A(n1774), .B(n1775), .Z(n1788) );
  NAND U2486 ( .A(n880), .B(n1207), .Z(n1775) );
  XNOR U2487 ( .A(n1773), .B(n1880), .Z(n1774) );
  ANDN U2488 ( .A(n1214), .B(n882), .Z(n1880) );
  XNOR U2489 ( .A(n1787), .B(n1776), .Z(n1879) );
  XOR U2490 ( .A(n1887), .B(n1783), .Z(n1787) );
  XNOR U2491 ( .A(n1781), .B(n1888), .Z(n1783) );
  ANDN U2492 ( .A(n1398), .B(n759), .Z(n1888) );
  AND U2493 ( .A(n757), .B(n1391), .Z(n1785) );
  XNOR U2494 ( .A(n1796), .B(n1795), .Z(n1770) );
  XOR U2495 ( .A(n1895), .B(n1804), .Z(n1795) );
  XNOR U2496 ( .A(n1792), .B(n1793), .Z(n1804) );
  NANDN U2497 ( .B(n651), .A(n1520), .Z(n1793) );
  XNOR U2498 ( .A(n1791), .B(n1896), .Z(n1792) );
  ANDN U2499 ( .A(n692), .B(n1522), .Z(n1896) );
  XNOR U2500 ( .A(n1803), .B(n1794), .Z(n1895) );
  XOR U2501 ( .A(n1903), .B(n1800), .Z(n1803) );
  XNOR U2502 ( .A(n1799), .B(n1904), .Z(n1800) );
  ANDN U2503 ( .A(n799), .B(n1334), .Z(n1904) );
  AND U2504 ( .A(n1332), .B(n745), .Z(n1801) );
  XOR U2505 ( .A(n1812), .B(n1811), .Z(n1796) );
  XOR U2506 ( .A(n1911), .B(n1808), .Z(n1811) );
  XNOR U2507 ( .A(n1807), .B(n1912), .Z(n1808) );
  ANDN U2508 ( .A(n624), .B(n1714), .Z(n1912) );
  AND U2509 ( .A(n1712), .B(n583), .Z(n1809) );
  XOR U2510 ( .A(n1819), .B(n1818), .Z(n1812) );
  NAND U2511 ( .A(n1919), .B(n527), .Z(n1818) );
  XOR U2512 ( .A(n1817), .B(n1920), .Z(n1819) );
  ANDN U2513 ( .A(n558), .B(n1921), .Z(n1920) );
  ANDN U2514 ( .A(n1922), .B(n1923), .Z(n1817) );
  NAND U2515 ( .A(n1924), .B(n1925), .Z(n1922) );
  IV U2516 ( .A(n1820), .Z(n1821) );
  MUX U2517 ( .IN0(o[8]), .IN1(n408), .SEL(n479), .F(\_MxM/n321 ) );
  XOR U2518 ( .A(n1930), .B(\_MxM/Y0[9] ), .Z(n408) );
  XOR U2519 ( .A(n1931), .B(n1932), .Z(n1930) );
  AND U2520 ( .A(n491), .B(n1934), .Z(n1933) );
  XOR U2521 ( .A(n1928), .B(n1932), .Z(n1934) );
  XOR U2522 ( .A(n1927), .B(n1932), .Z(n1928) );
  XNOR U2523 ( .A(n1935), .B(n1862), .Z(n1858) );
  XNOR U2524 ( .A(n1842), .B(n1841), .Z(n1862) );
  XOR U2525 ( .A(n1936), .B(n1838), .Z(n1841) );
  XNOR U2526 ( .A(n1937), .B(n1834), .Z(n1838) );
  AND U2527 ( .A(n1938), .B(n556), .Z(n1834) );
  NAND U2528 ( .A(n1939), .B(n1833), .Z(n1937) );
  NANDN U2529 ( .B(n559), .A(n1943), .Z(n1939) );
  XNOR U2530 ( .A(n1839), .B(n1840), .Z(n1936) );
  XNOR U2531 ( .A(n1947), .B(n1950), .Z(n1949) );
  XNOR U2532 ( .A(n1852), .B(n1851), .Z(n1842) );
  XOR U2533 ( .A(n1951), .B(n1847), .Z(n1851) );
  XNOR U2534 ( .A(n1845), .B(n1952), .Z(n1847) );
  ANDN U2535 ( .A(n1744), .B(n633), .Z(n1952) );
  XOR U2536 ( .A(n1953), .B(n1954), .Z(n1845) );
  AND U2537 ( .A(n1955), .B(n1956), .Z(n1954) );
  XNOR U2538 ( .A(n1957), .B(n1953), .Z(n1956) );
  AND U2539 ( .A(n1737), .B(n631), .Z(n1849) );
  XNOR U2540 ( .A(n1855), .B(n1856), .Z(n1852) );
  NAND U2541 ( .A(n1542), .B(n715), .Z(n1856) );
  XNOR U2542 ( .A(n1854), .B(n1961), .Z(n1855) );
  ANDN U2543 ( .A(n1547), .B(n717), .Z(n1961) );
  XNOR U2544 ( .A(n1861), .B(n1857), .Z(n1935) );
  IV U2545 ( .A(n1860), .Z(n1861) );
  XNOR U2546 ( .A(n1878), .B(n1877), .Z(n1859) );
  XOR U2547 ( .A(n1970), .B(n1886), .Z(n1877) );
  XNOR U2548 ( .A(n1871), .B(n1870), .Z(n1886) );
  XOR U2549 ( .A(n1971), .B(n1867), .Z(n1870) );
  XNOR U2550 ( .A(n1866), .B(n1972), .Z(n1867) );
  ANDN U2551 ( .A(n1036), .B(n1091), .Z(n1972) );
  AND U2552 ( .A(n1089), .B(n973), .Z(n1868) );
  XNOR U2553 ( .A(n1874), .B(n1875), .Z(n1871) );
  NANDN U2554 ( .B(n838), .A(n1248), .Z(n1875) );
  XNOR U2555 ( .A(n1873), .B(n1979), .Z(n1874) );
  ANDN U2556 ( .A(n908), .B(n1250), .Z(n1979) );
  XNOR U2557 ( .A(n1885), .B(n1876), .Z(n1970) );
  XOR U2558 ( .A(n1986), .B(n1894), .Z(n1885) );
  XNOR U2559 ( .A(n1882), .B(n1883), .Z(n1894) );
  NAND U2560 ( .A(n948), .B(n1207), .Z(n1883) );
  XNOR U2561 ( .A(n1881), .B(n1987), .Z(n1882) );
  ANDN U2562 ( .A(n1214), .B(n950), .Z(n1987) );
  XNOR U2563 ( .A(n1893), .B(n1884), .Z(n1986) );
  XOR U2564 ( .A(n1994), .B(n1890), .Z(n1893) );
  XNOR U2565 ( .A(n1889), .B(n1995), .Z(n1890) );
  ANDN U2566 ( .A(n1398), .B(n818), .Z(n1995) );
  AND U2567 ( .A(n816), .B(n1391), .Z(n1891) );
  XNOR U2568 ( .A(n1902), .B(n1901), .Z(n1878) );
  XOR U2569 ( .A(n2002), .B(n1910), .Z(n1901) );
  XNOR U2570 ( .A(n1898), .B(n1899), .Z(n1910) );
  NANDN U2571 ( .B(n651), .A(n1616), .Z(n1899) );
  XNOR U2572 ( .A(n1897), .B(n2003), .Z(n1898) );
  ANDN U2573 ( .A(n692), .B(n1618), .Z(n2003) );
  XNOR U2574 ( .A(n1909), .B(n1900), .Z(n2002) );
  XOR U2575 ( .A(n2010), .B(n1906), .Z(n1909) );
  XNOR U2576 ( .A(n1905), .B(n2011), .Z(n1906) );
  ANDN U2577 ( .A(n799), .B(n1425), .Z(n2011) );
  AND U2578 ( .A(n1423), .B(n745), .Z(n1907) );
  XOR U2579 ( .A(n1918), .B(n1917), .Z(n1902) );
  XOR U2580 ( .A(n2018), .B(n1914), .Z(n1917) );
  XNOR U2581 ( .A(n1913), .B(n2019), .Z(n1914) );
  ANDN U2582 ( .A(n624), .B(n1815), .Z(n2019) );
  AND U2583 ( .A(n1813), .B(n583), .Z(n1915) );
  XOR U2584 ( .A(n1925), .B(n1924), .Z(n1918) );
  NAND U2585 ( .A(n2026), .B(n527), .Z(n1924) );
  XNOR U2586 ( .A(n1923), .B(n2027), .Z(n1925) );
  ANDN U2587 ( .A(n558), .B(n2028), .Z(n2027) );
  NAND U2588 ( .A(n2029), .B(n2030), .Z(n1923) );
  NAND U2589 ( .A(n2031), .B(n2032), .Z(n2029) );
  IV U2590 ( .A(n1926), .Z(n1927) );
  MUX U2591 ( .IN0(o[7]), .IN1(n405), .SEL(n479), .F(\_MxM/n320 ) );
  XOR U2592 ( .A(n2037), .B(\_MxM/Y0[8] ), .Z(n405) );
  XOR U2593 ( .A(n2038), .B(n2039), .Z(n2037) );
  AND U2594 ( .A(n491), .B(n2041), .Z(n2040) );
  XOR U2595 ( .A(n2035), .B(n2039), .Z(n2041) );
  XOR U2596 ( .A(n2034), .B(n2039), .Z(n2035) );
  XNOR U2597 ( .A(n2042), .B(n1969), .Z(n1966) );
  XNOR U2598 ( .A(n1946), .B(n1945), .Z(n1969) );
  XOR U2599 ( .A(n2043), .B(n1950), .Z(n1945) );
  XNOR U2600 ( .A(n1941), .B(n1942), .Z(n1950) );
  NAND U2601 ( .A(n1938), .B(n587), .Z(n1942) );
  XNOR U2602 ( .A(n1940), .B(n2044), .Z(n1941) );
  ANDN U2603 ( .A(n1943), .B(n589), .Z(n2044) );
  XNOR U2604 ( .A(n1948), .B(n1944), .Z(n2043) );
  XOR U2605 ( .A(n1947), .B(n2051), .Z(n1948) );
  AND U2606 ( .A(n2052), .B(n2053), .Z(n2051) );
  NANDN U2607 ( .B(n2054), .A(n526), .Z(n2053) );
  NANDN U2608 ( .B(n2055), .A(n2056), .Z(n2052) );
  XNOR U2609 ( .A(n1960), .B(n1959), .Z(n1946) );
  XOR U2610 ( .A(n2060), .B(n1955), .Z(n1959) );
  XNOR U2611 ( .A(n1953), .B(n2061), .Z(n1955) );
  ANDN U2612 ( .A(n1744), .B(n673), .Z(n2061) );
  AND U2613 ( .A(n1737), .B(n671), .Z(n1957) );
  XNOR U2614 ( .A(n1963), .B(n1964), .Z(n1960) );
  NAND U2615 ( .A(n1542), .B(n757), .Z(n1964) );
  XNOR U2616 ( .A(n1962), .B(n2068), .Z(n1963) );
  ANDN U2617 ( .A(n1547), .B(n759), .Z(n2068) );
  XNOR U2618 ( .A(n1985), .B(n1984), .Z(n1967) );
  XOR U2619 ( .A(n2078), .B(n1993), .Z(n1984) );
  XNOR U2620 ( .A(n1978), .B(n1977), .Z(n1993) );
  XOR U2621 ( .A(n2079), .B(n1974), .Z(n1977) );
  XNOR U2622 ( .A(n1973), .B(n2080), .Z(n1974) );
  ANDN U2623 ( .A(n1036), .B(n1169), .Z(n2080) );
  AND U2624 ( .A(n1167), .B(n973), .Z(n1975) );
  XNOR U2625 ( .A(n1981), .B(n1982), .Z(n1978) );
  NANDN U2626 ( .B(n838), .A(n1332), .Z(n1982) );
  XNOR U2627 ( .A(n1980), .B(n2087), .Z(n1981) );
  ANDN U2628 ( .A(n908), .B(n1334), .Z(n2087) );
  XNOR U2629 ( .A(n1992), .B(n1983), .Z(n2078) );
  XOR U2630 ( .A(n2094), .B(n2001), .Z(n1992) );
  XNOR U2631 ( .A(n1989), .B(n1990), .Z(n2001) );
  NAND U2632 ( .A(n1015), .B(n1207), .Z(n1990) );
  XNOR U2633 ( .A(n1988), .B(n2095), .Z(n1989) );
  ANDN U2634 ( .A(n1214), .B(n1017), .Z(n2095) );
  XNOR U2635 ( .A(n2000), .B(n1991), .Z(n2094) );
  XOR U2636 ( .A(n2102), .B(n1997), .Z(n2000) );
  XNOR U2637 ( .A(n1996), .B(n2103), .Z(n1997) );
  ANDN U2638 ( .A(n1398), .B(n882), .Z(n2103) );
  AND U2639 ( .A(n880), .B(n1391), .Z(n1998) );
  XNOR U2640 ( .A(n2009), .B(n2008), .Z(n1985) );
  XOR U2641 ( .A(n2110), .B(n2017), .Z(n2008) );
  XNOR U2642 ( .A(n2005), .B(n2006), .Z(n2017) );
  NANDN U2643 ( .B(n651), .A(n1712), .Z(n2006) );
  XNOR U2644 ( .A(n2004), .B(n2111), .Z(n2005) );
  ANDN U2645 ( .A(n692), .B(n1714), .Z(n2111) );
  XNOR U2646 ( .A(n2016), .B(n2007), .Z(n2110) );
  XOR U2647 ( .A(n2118), .B(n2013), .Z(n2016) );
  XNOR U2648 ( .A(n2012), .B(n2119), .Z(n2013) );
  ANDN U2649 ( .A(n799), .B(n1522), .Z(n2119) );
  AND U2650 ( .A(n1520), .B(n745), .Z(n2014) );
  XOR U2651 ( .A(n2025), .B(n2024), .Z(n2009) );
  XOR U2652 ( .A(n2126), .B(n2021), .Z(n2024) );
  XNOR U2653 ( .A(n2020), .B(n2127), .Z(n2021) );
  ANDN U2654 ( .A(n624), .B(n1921), .Z(n2127) );
  AND U2655 ( .A(n1919), .B(n583), .Z(n2022) );
  XOR U2656 ( .A(n2032), .B(n2031), .Z(n2025) );
  NAND U2657 ( .A(n2134), .B(n527), .Z(n2031) );
  XOR U2658 ( .A(n2030), .B(n2135), .Z(n2032) );
  ANDN U2659 ( .A(n558), .B(n2136), .Z(n2135) );
  ANDN U2660 ( .A(n2137), .B(n2138), .Z(n2030) );
  NAND U2661 ( .A(n2139), .B(n2140), .Z(n2137) );
  IV U2662 ( .A(n2033), .Z(n2034) );
  MUX U2663 ( .IN0(o[6]), .IN1(n402), .SEL(n479), .F(\_MxM/n319 ) );
  XOR U2664 ( .A(n2145), .B(\_MxM/Y0[7] ), .Z(n402) );
  XOR U2665 ( .A(n2146), .B(n2147), .Z(n2145) );
  AND U2666 ( .A(n491), .B(n2149), .Z(n2148) );
  XOR U2667 ( .A(n2143), .B(n2147), .Z(n2149) );
  XOR U2668 ( .A(n2142), .B(n2147), .Z(n2143) );
  XNOR U2669 ( .A(n2150), .B(n2077), .Z(n2073) );
  XNOR U2670 ( .A(n2050), .B(n2049), .Z(n2077) );
  XOR U2671 ( .A(n2151), .B(n2059), .Z(n2049) );
  XNOR U2672 ( .A(n2046), .B(n2047), .Z(n2059) );
  NAND U2673 ( .A(n1938), .B(n631), .Z(n2047) );
  XNOR U2674 ( .A(n2045), .B(n2152), .Z(n2046) );
  ANDN U2675 ( .A(n1943), .B(n633), .Z(n2152) );
  XOR U2676 ( .A(n2153), .B(n2154), .Z(n2045) );
  AND U2677 ( .A(n2155), .B(n2156), .Z(n2154) );
  XOR U2678 ( .A(n2157), .B(n2153), .Z(n2156) );
  XNOR U2679 ( .A(n2058), .B(n2048), .Z(n2151) );
  XOR U2680 ( .A(n2165), .B(n2056), .Z(n2161) );
  AND U2681 ( .A(n2166), .B(n556), .Z(n2056) );
  NAND U2682 ( .A(n2167), .B(n2055), .Z(n2165) );
  XOR U2683 ( .A(n2168), .B(n2169), .Z(n2055) );
  AND U2684 ( .A(n2170), .B(n2171), .Z(n2169) );
  XNOR U2685 ( .A(n2172), .B(n2168), .Z(n2171) );
  NANDN U2686 ( .B(n559), .A(n2173), .Z(n2167) );
  XNOR U2687 ( .A(n2067), .B(n2066), .Z(n2050) );
  XOR U2688 ( .A(n2174), .B(n2063), .Z(n2066) );
  XNOR U2689 ( .A(n2062), .B(n2175), .Z(n2063) );
  ANDN U2690 ( .A(n1744), .B(n717), .Z(n2175) );
  AND U2691 ( .A(n1737), .B(n715), .Z(n2064) );
  XNOR U2692 ( .A(n2070), .B(n2071), .Z(n2067) );
  NAND U2693 ( .A(n1542), .B(n816), .Z(n2071) );
  XNOR U2694 ( .A(n2069), .B(n2182), .Z(n2070) );
  ANDN U2695 ( .A(n1547), .B(n818), .Z(n2182) );
  XNOR U2696 ( .A(n2076), .B(n2072), .Z(n2150) );
  XOR U2697 ( .A(n2193), .B(n2194), .Z(n2189) );
  NANDN U2698 ( .B(n2195), .A(n2196), .Z(n2193) );
  XNOR U2699 ( .A(n2093), .B(n2092), .Z(n2074) );
  XOR U2700 ( .A(n2197), .B(n2101), .Z(n2092) );
  XNOR U2701 ( .A(n2086), .B(n2085), .Z(n2101) );
  XOR U2702 ( .A(n2198), .B(n2082), .Z(n2085) );
  XNOR U2703 ( .A(n2081), .B(n2199), .Z(n2082) );
  ANDN U2704 ( .A(n1036), .B(n1250), .Z(n2199) );
  AND U2705 ( .A(n1248), .B(n973), .Z(n2083) );
  XNOR U2706 ( .A(n2089), .B(n2090), .Z(n2086) );
  NANDN U2707 ( .B(n838), .A(n1423), .Z(n2090) );
  XNOR U2708 ( .A(n2088), .B(n2206), .Z(n2089) );
  ANDN U2709 ( .A(n908), .B(n1425), .Z(n2206) );
  XNOR U2710 ( .A(n2100), .B(n2091), .Z(n2197) );
  XOR U2711 ( .A(n2213), .B(n2109), .Z(n2100) );
  XNOR U2712 ( .A(n2097), .B(n2098), .Z(n2109) );
  NAND U2713 ( .A(n1089), .B(n1207), .Z(n2098) );
  XNOR U2714 ( .A(n2096), .B(n2214), .Z(n2097) );
  ANDN U2715 ( .A(n1214), .B(n1091), .Z(n2214) );
  XNOR U2716 ( .A(n2108), .B(n2099), .Z(n2213) );
  XOR U2717 ( .A(n2221), .B(n2105), .Z(n2108) );
  XNOR U2718 ( .A(n2104), .B(n2222), .Z(n2105) );
  ANDN U2719 ( .A(n1398), .B(n950), .Z(n2222) );
  AND U2720 ( .A(n948), .B(n1391), .Z(n2106) );
  XNOR U2721 ( .A(n2117), .B(n2116), .Z(n2093) );
  XOR U2722 ( .A(n2229), .B(n2125), .Z(n2116) );
  XNOR U2723 ( .A(n2113), .B(n2114), .Z(n2125) );
  NANDN U2724 ( .B(n651), .A(n1813), .Z(n2114) );
  XNOR U2725 ( .A(n2112), .B(n2230), .Z(n2113) );
  ANDN U2726 ( .A(n692), .B(n1815), .Z(n2230) );
  XNOR U2727 ( .A(n2124), .B(n2115), .Z(n2229) );
  XOR U2728 ( .A(n2237), .B(n2121), .Z(n2124) );
  XNOR U2729 ( .A(n2120), .B(n2238), .Z(n2121) );
  ANDN U2730 ( .A(n799), .B(n1618), .Z(n2238) );
  AND U2731 ( .A(n1616), .B(n745), .Z(n2122) );
  XOR U2732 ( .A(n2133), .B(n2132), .Z(n2117) );
  XOR U2733 ( .A(n2245), .B(n2129), .Z(n2132) );
  XNOR U2734 ( .A(n2128), .B(n2246), .Z(n2129) );
  ANDN U2735 ( .A(n624), .B(n2028), .Z(n2246) );
  AND U2736 ( .A(n2026), .B(n583), .Z(n2130) );
  XOR U2737 ( .A(n2140), .B(n2139), .Z(n2133) );
  NAND U2738 ( .A(n2253), .B(n527), .Z(n2139) );
  XNOR U2739 ( .A(n2138), .B(n2254), .Z(n2140) );
  ANDN U2740 ( .A(n558), .B(n2255), .Z(n2254) );
  NAND U2741 ( .A(n2256), .B(n2257), .Z(n2138) );
  NAND U2742 ( .A(n2258), .B(n2259), .Z(n2256) );
  IV U2743 ( .A(n2141), .Z(n2142) );
  MUX U2744 ( .IN0(o[5]), .IN1(n399), .SEL(n479), .F(\_MxM/n318 ) );
  XOR U2745 ( .A(n2264), .B(\_MxM/Y0[6] ), .Z(n399) );
  XOR U2746 ( .A(n2265), .B(n2266), .Z(n2264) );
  AND U2747 ( .A(n491), .B(n2268), .Z(n2267) );
  XOR U2748 ( .A(n2262), .B(n2266), .Z(n2268) );
  XOR U2749 ( .A(n2261), .B(n2266), .Z(n2262) );
  XNOR U2750 ( .A(n2269), .B(n2192), .Z(n2187) );
  XNOR U2751 ( .A(n2160), .B(n2159), .Z(n2192) );
  XOR U2752 ( .A(n2270), .B(n2164), .Z(n2159) );
  XNOR U2753 ( .A(n2155), .B(n2157), .Z(n2164) );
  NAND U2754 ( .A(n1938), .B(n671), .Z(n2157) );
  XNOR U2755 ( .A(n2153), .B(n2271), .Z(n2155) );
  ANDN U2756 ( .A(n1943), .B(n673), .Z(n2271) );
  XNOR U2757 ( .A(n2163), .B(n2158), .Z(n2270) );
  XOR U2758 ( .A(n2278), .B(n2170), .Z(n2163) );
  XNOR U2759 ( .A(n2168), .B(n2279), .Z(n2170) );
  ANDN U2760 ( .A(n2173), .B(n589), .Z(n2279) );
  XOR U2761 ( .A(n2280), .B(n2281), .Z(n2168) );
  AND U2762 ( .A(n2282), .B(n2283), .Z(n2281) );
  XNOR U2763 ( .A(n2284), .B(n2280), .Z(n2283) );
  AND U2764 ( .A(n2166), .B(n587), .Z(n2172) );
  XNOR U2765 ( .A(n2181), .B(n2180), .Z(n2160) );
  XOR U2766 ( .A(n2288), .B(n2177), .Z(n2180) );
  XNOR U2767 ( .A(n2176), .B(n2289), .Z(n2177) );
  ANDN U2768 ( .A(n1744), .B(n759), .Z(n2289) );
  AND U2769 ( .A(n1737), .B(n757), .Z(n2178) );
  XNOR U2770 ( .A(n2184), .B(n2185), .Z(n2181) );
  NAND U2771 ( .A(n1542), .B(n880), .Z(n2185) );
  XNOR U2772 ( .A(n2183), .B(n2296), .Z(n2184) );
  ANDN U2773 ( .A(n1547), .B(n882), .Z(n2296) );
  XNOR U2774 ( .A(n2191), .B(n2186), .Z(n2269) );
  XOR U2775 ( .A(n2190), .B(n2303), .Z(n2191) );
  AND U2776 ( .A(n2194), .B(n2304), .Z(n2303) );
  AND U2777 ( .A(n2305), .B(n2306), .Z(n2304) );
  NANDN U2778 ( .B(n2307), .A(n526), .Z(n2306) );
  NAND U2779 ( .A(n2308), .B(n2309), .Z(n2305) );
  ANDN U2780 ( .A(n2196), .B(n2195), .Z(n2194) );
  ANDN U2781 ( .A(n2310), .B(n2311), .Z(n2195) );
  OR U2782 ( .A(n2312), .B(n2313), .Z(n2196) );
  XNOR U2783 ( .A(n2212), .B(n2211), .Z(n2188) );
  XOR U2784 ( .A(n2317), .B(n2220), .Z(n2211) );
  XNOR U2785 ( .A(n2205), .B(n2204), .Z(n2220) );
  XOR U2786 ( .A(n2318), .B(n2201), .Z(n2204) );
  XNOR U2787 ( .A(n2200), .B(n2319), .Z(n2201) );
  ANDN U2788 ( .A(n1036), .B(n1334), .Z(n2319) );
  AND U2789 ( .A(n1332), .B(n973), .Z(n2202) );
  XNOR U2790 ( .A(n2208), .B(n2209), .Z(n2205) );
  NANDN U2791 ( .B(n838), .A(n1520), .Z(n2209) );
  XNOR U2792 ( .A(n2207), .B(n2326), .Z(n2208) );
  ANDN U2793 ( .A(n908), .B(n1522), .Z(n2326) );
  XNOR U2794 ( .A(n2219), .B(n2210), .Z(n2317) );
  XOR U2795 ( .A(n2333), .B(n2228), .Z(n2219) );
  XNOR U2796 ( .A(n2216), .B(n2217), .Z(n2228) );
  NAND U2797 ( .A(n1167), .B(n1207), .Z(n2217) );
  XNOR U2798 ( .A(n2215), .B(n2334), .Z(n2216) );
  ANDN U2799 ( .A(n1214), .B(n1169), .Z(n2334) );
  XNOR U2800 ( .A(n2227), .B(n2218), .Z(n2333) );
  XOR U2801 ( .A(n2341), .B(n2224), .Z(n2227) );
  XNOR U2802 ( .A(n2223), .B(n2342), .Z(n2224) );
  ANDN U2803 ( .A(n1398), .B(n1017), .Z(n2342) );
  AND U2804 ( .A(n1015), .B(n1391), .Z(n2225) );
  XNOR U2805 ( .A(n2236), .B(n2235), .Z(n2212) );
  XOR U2806 ( .A(n2349), .B(n2244), .Z(n2235) );
  XNOR U2807 ( .A(n2232), .B(n2233), .Z(n2244) );
  NANDN U2808 ( .B(n651), .A(n1919), .Z(n2233) );
  XNOR U2809 ( .A(n2231), .B(n2350), .Z(n2232) );
  ANDN U2810 ( .A(n692), .B(n1921), .Z(n2350) );
  XNOR U2811 ( .A(n2243), .B(n2234), .Z(n2349) );
  XOR U2812 ( .A(n2357), .B(n2240), .Z(n2243) );
  XNOR U2813 ( .A(n2239), .B(n2358), .Z(n2240) );
  ANDN U2814 ( .A(n799), .B(n1714), .Z(n2358) );
  AND U2815 ( .A(n1712), .B(n745), .Z(n2241) );
  XOR U2816 ( .A(n2252), .B(n2251), .Z(n2236) );
  XOR U2817 ( .A(n2365), .B(n2248), .Z(n2251) );
  XNOR U2818 ( .A(n2247), .B(n2366), .Z(n2248) );
  ANDN U2819 ( .A(n624), .B(n2136), .Z(n2366) );
  AND U2820 ( .A(n2134), .B(n583), .Z(n2249) );
  XOR U2821 ( .A(n2259), .B(n2258), .Z(n2252) );
  NAND U2822 ( .A(n2373), .B(n527), .Z(n2258) );
  XOR U2823 ( .A(n2257), .B(n2374), .Z(n2259) );
  ANDN U2824 ( .A(n558), .B(n2375), .Z(n2374) );
  ANDN U2825 ( .A(n2376), .B(n2377), .Z(n2257) );
  NAND U2826 ( .A(n2378), .B(n2379), .Z(n2376) );
  IV U2827 ( .A(n2260), .Z(n2261) );
  MUX U2828 ( .IN0(o[4]), .IN1(n396), .SEL(n479), .F(\_MxM/n317 ) );
  XOR U2829 ( .A(n2384), .B(\_MxM/Y0[5] ), .Z(n396) );
  XOR U2830 ( .A(n2385), .B(n2386), .Z(n2384) );
  AND U2831 ( .A(n491), .B(n2388), .Z(n2387) );
  XOR U2832 ( .A(n2382), .B(n2386), .Z(n2388) );
  XOR U2833 ( .A(n2381), .B(n2386), .Z(n2382) );
  XNOR U2834 ( .A(n2389), .B(n2316), .Z(n2301) );
  XNOR U2835 ( .A(n2277), .B(n2276), .Z(n2316) );
  XOR U2836 ( .A(n2390), .B(n2287), .Z(n2276) );
  XNOR U2837 ( .A(n2273), .B(n2274), .Z(n2287) );
  NAND U2838 ( .A(n1938), .B(n715), .Z(n2274) );
  XNOR U2839 ( .A(n2272), .B(n2391), .Z(n2273) );
  ANDN U2840 ( .A(n1943), .B(n717), .Z(n2391) );
  XNOR U2841 ( .A(n2286), .B(n2275), .Z(n2390) );
  XOR U2842 ( .A(n2398), .B(n2282), .Z(n2286) );
  XNOR U2843 ( .A(n2280), .B(n2399), .Z(n2282) );
  ANDN U2844 ( .A(n2173), .B(n633), .Z(n2399) );
  XOR U2845 ( .A(n2400), .B(n2401), .Z(n2280) );
  AND U2846 ( .A(n2402), .B(n2403), .Z(n2401) );
  XNOR U2847 ( .A(n2404), .B(n2400), .Z(n2403) );
  AND U2848 ( .A(n2166), .B(n631), .Z(n2284) );
  XNOR U2849 ( .A(n2295), .B(n2294), .Z(n2277) );
  XOR U2850 ( .A(n2408), .B(n2291), .Z(n2294) );
  XNOR U2851 ( .A(n2290), .B(n2409), .Z(n2291) );
  ANDN U2852 ( .A(n1744), .B(n818), .Z(n2409) );
  AND U2853 ( .A(n1737), .B(n816), .Z(n2292) );
  XNOR U2854 ( .A(n2298), .B(n2299), .Z(n2295) );
  NAND U2855 ( .A(n1542), .B(n948), .Z(n2299) );
  XNOR U2856 ( .A(n2297), .B(n2416), .Z(n2298) );
  ANDN U2857 ( .A(n1547), .B(n950), .Z(n2416) );
  XOR U2858 ( .A(n2315), .B(n2300), .Z(n2389) );
  XOR U2859 ( .A(n2423), .B(n2308), .Z(n2315) );
  XOR U2860 ( .A(n2427), .B(n2313), .Z(n2311) );
  NAND U2861 ( .A(n2428), .B(n556), .Z(n2313) );
  NAND U2862 ( .A(n2429), .B(n2312), .Z(n2427) );
  NANDN U2863 ( .B(n559), .A(n2433), .Z(n2429) );
  ANDN U2864 ( .A(n2434), .B(n2435), .Z(n2309) );
  XNOR U2865 ( .A(n2332), .B(n2331), .Z(n2302) );
  XOR U2866 ( .A(n2439), .B(n2340), .Z(n2331) );
  XNOR U2867 ( .A(n2325), .B(n2324), .Z(n2340) );
  XOR U2868 ( .A(n2440), .B(n2321), .Z(n2324) );
  XNOR U2869 ( .A(n2320), .B(n2441), .Z(n2321) );
  ANDN U2870 ( .A(n1036), .B(n1425), .Z(n2441) );
  AND U2871 ( .A(n1423), .B(n973), .Z(n2322) );
  XNOR U2872 ( .A(n2328), .B(n2329), .Z(n2325) );
  NANDN U2873 ( .B(n838), .A(n1616), .Z(n2329) );
  XNOR U2874 ( .A(n2327), .B(n2448), .Z(n2328) );
  ANDN U2875 ( .A(n908), .B(n1618), .Z(n2448) );
  XNOR U2876 ( .A(n2339), .B(n2330), .Z(n2439) );
  XOR U2877 ( .A(n2455), .B(n2348), .Z(n2339) );
  XNOR U2878 ( .A(n2336), .B(n2337), .Z(n2348) );
  NAND U2879 ( .A(n1248), .B(n1207), .Z(n2337) );
  XNOR U2880 ( .A(n2335), .B(n2456), .Z(n2336) );
  ANDN U2881 ( .A(n1214), .B(n1250), .Z(n2456) );
  XNOR U2882 ( .A(n2347), .B(n2338), .Z(n2455) );
  XOR U2883 ( .A(n2463), .B(n2344), .Z(n2347) );
  XNOR U2884 ( .A(n2343), .B(n2464), .Z(n2344) );
  ANDN U2885 ( .A(n1398), .B(n1091), .Z(n2464) );
  AND U2886 ( .A(n1089), .B(n1391), .Z(n2345) );
  XNOR U2887 ( .A(n2356), .B(n2355), .Z(n2332) );
  XOR U2888 ( .A(n2471), .B(n2364), .Z(n2355) );
  XNOR U2889 ( .A(n2352), .B(n2353), .Z(n2364) );
  NANDN U2890 ( .B(n651), .A(n2026), .Z(n2353) );
  XNOR U2891 ( .A(n2351), .B(n2472), .Z(n2352) );
  ANDN U2892 ( .A(n692), .B(n2028), .Z(n2472) );
  XNOR U2893 ( .A(n2363), .B(n2354), .Z(n2471) );
  XOR U2894 ( .A(n2479), .B(n2360), .Z(n2363) );
  XNOR U2895 ( .A(n2359), .B(n2480), .Z(n2360) );
  ANDN U2896 ( .A(n799), .B(n1815), .Z(n2480) );
  AND U2897 ( .A(n1813), .B(n745), .Z(n2361) );
  XOR U2898 ( .A(n2372), .B(n2371), .Z(n2356) );
  XOR U2899 ( .A(n2487), .B(n2368), .Z(n2371) );
  XNOR U2900 ( .A(n2367), .B(n2488), .Z(n2368) );
  ANDN U2901 ( .A(n624), .B(n2255), .Z(n2488) );
  AND U2902 ( .A(n2253), .B(n583), .Z(n2369) );
  XOR U2903 ( .A(n2379), .B(n2378), .Z(n2372) );
  NAND U2904 ( .A(n2495), .B(n527), .Z(n2378) );
  XNOR U2905 ( .A(n2377), .B(n2496), .Z(n2379) );
  ANDN U2906 ( .A(n558), .B(n2497), .Z(n2496) );
  NAND U2907 ( .A(n2498), .B(n2499), .Z(n2377) );
  NAND U2908 ( .A(n2500), .B(n2501), .Z(n2498) );
  IV U2909 ( .A(n2380), .Z(n2381) );
  MUX U2910 ( .IN0(o[3]), .IN1(n393), .SEL(n479), .F(\_MxM/n316 ) );
  XNOR U2911 ( .A(n2505), .B(\_MxM/Y0[4] ), .Z(n393) );
  XNOR U2912 ( .A(n2507), .B(n2508), .Z(n2505) );
  XOR U2913 ( .A(n2506), .B(n2509), .Z(n2507) );
  AND U2914 ( .A(n491), .B(n2510), .Z(n2509) );
  XNOR U2915 ( .A(n2503), .B(n2508), .Z(n2510) );
  XOR U2916 ( .A(n2508), .B(n2502), .Z(n2503) );
  NOR U2917 ( .A(n2511), .B(n2512), .Z(n2502) );
  XNOR U2918 ( .A(n2513), .B(n2438), .Z(n2421) );
  XNOR U2919 ( .A(n2397), .B(n2396), .Z(n2438) );
  XOR U2920 ( .A(n2514), .B(n2407), .Z(n2396) );
  XNOR U2921 ( .A(n2393), .B(n2394), .Z(n2407) );
  NAND U2922 ( .A(n1938), .B(n757), .Z(n2394) );
  XNOR U2923 ( .A(n2392), .B(n2515), .Z(n2393) );
  ANDN U2924 ( .A(n1943), .B(n759), .Z(n2515) );
  XNOR U2925 ( .A(n2406), .B(n2395), .Z(n2514) );
  XOR U2926 ( .A(n2522), .B(n2402), .Z(n2406) );
  XNOR U2927 ( .A(n2400), .B(n2523), .Z(n2402) );
  ANDN U2928 ( .A(n2173), .B(n673), .Z(n2523) );
  AND U2929 ( .A(n2166), .B(n671), .Z(n2404) );
  XNOR U2930 ( .A(n2415), .B(n2414), .Z(n2397) );
  XOR U2931 ( .A(n2530), .B(n2411), .Z(n2414) );
  XNOR U2932 ( .A(n2410), .B(n2531), .Z(n2411) );
  ANDN U2933 ( .A(n1744), .B(n882), .Z(n2531) );
  AND U2934 ( .A(n1737), .B(n880), .Z(n2412) );
  XNOR U2935 ( .A(n2418), .B(n2419), .Z(n2415) );
  NAND U2936 ( .A(n1542), .B(n1015), .Z(n2419) );
  XNOR U2937 ( .A(n2417), .B(n2538), .Z(n2418) );
  ANDN U2938 ( .A(n1547), .B(n1017), .Z(n2538) );
  XNOR U2939 ( .A(n2437), .B(n2420), .Z(n2513) );
  XOR U2940 ( .A(n2545), .B(n2435), .Z(n2437) );
  XOR U2941 ( .A(n2426), .B(n2425), .Z(n2435) );
  XNOR U2942 ( .A(n2424), .B(n2546), .Z(n2425) );
  AND U2943 ( .A(n2547), .B(n2548), .Z(n2546) );
  NANDN U2944 ( .B(n2549), .A(n526), .Z(n2548) );
  NANDN U2945 ( .B(n2550), .A(n2551), .Z(n2547) );
  XNOR U2946 ( .A(n2431), .B(n2432), .Z(n2426) );
  NAND U2947 ( .A(n2428), .B(n587), .Z(n2432) );
  XNOR U2948 ( .A(n2430), .B(n2555), .Z(n2431) );
  ANDN U2949 ( .A(n2433), .B(n589), .Z(n2555) );
  NOR U2950 ( .A(n2559), .B(n2560), .Z(n2434) );
  XNOR U2951 ( .A(n2454), .B(n2453), .Z(n2422) );
  XOR U2952 ( .A(n2564), .B(n2462), .Z(n2453) );
  XNOR U2953 ( .A(n2447), .B(n2446), .Z(n2462) );
  XOR U2954 ( .A(n2565), .B(n2443), .Z(n2446) );
  XNOR U2955 ( .A(n2442), .B(n2566), .Z(n2443) );
  ANDN U2956 ( .A(n1036), .B(n1522), .Z(n2566) );
  AND U2957 ( .A(n1520), .B(n973), .Z(n2444) );
  XNOR U2958 ( .A(n2450), .B(n2451), .Z(n2447) );
  NANDN U2959 ( .B(n838), .A(n1712), .Z(n2451) );
  XNOR U2960 ( .A(n2449), .B(n2573), .Z(n2450) );
  ANDN U2961 ( .A(n908), .B(n1714), .Z(n2573) );
  XNOR U2962 ( .A(n2461), .B(n2452), .Z(n2564) );
  XOR U2963 ( .A(n2580), .B(n2470), .Z(n2461) );
  XNOR U2964 ( .A(n2458), .B(n2459), .Z(n2470) );
  NAND U2965 ( .A(n1332), .B(n1207), .Z(n2459) );
  XNOR U2966 ( .A(n2457), .B(n2581), .Z(n2458) );
  ANDN U2967 ( .A(n1214), .B(n1334), .Z(n2581) );
  XNOR U2968 ( .A(n2469), .B(n2460), .Z(n2580) );
  XOR U2969 ( .A(n2588), .B(n2466), .Z(n2469) );
  XNOR U2970 ( .A(n2465), .B(n2589), .Z(n2466) );
  ANDN U2971 ( .A(n1398), .B(n1169), .Z(n2589) );
  AND U2972 ( .A(n1167), .B(n1391), .Z(n2467) );
  XNOR U2973 ( .A(n2478), .B(n2477), .Z(n2454) );
  XOR U2974 ( .A(n2596), .B(n2486), .Z(n2477) );
  XNOR U2975 ( .A(n2474), .B(n2475), .Z(n2486) );
  NANDN U2976 ( .B(n651), .A(n2134), .Z(n2475) );
  XNOR U2977 ( .A(n2473), .B(n2597), .Z(n2474) );
  ANDN U2978 ( .A(n692), .B(n2136), .Z(n2597) );
  XNOR U2979 ( .A(n2485), .B(n2476), .Z(n2596) );
  XOR U2980 ( .A(n2604), .B(n2482), .Z(n2485) );
  XNOR U2981 ( .A(n2481), .B(n2605), .Z(n2482) );
  ANDN U2982 ( .A(n799), .B(n1921), .Z(n2605) );
  AND U2983 ( .A(n1919), .B(n745), .Z(n2483) );
  XOR U2984 ( .A(n2494), .B(n2493), .Z(n2478) );
  XOR U2985 ( .A(n2612), .B(n2490), .Z(n2493) );
  XNOR U2986 ( .A(n2489), .B(n2613), .Z(n2490) );
  ANDN U2987 ( .A(n624), .B(n2375), .Z(n2613) );
  AND U2988 ( .A(n2373), .B(n583), .Z(n2491) );
  XOR U2989 ( .A(n2501), .B(n2500), .Z(n2494) );
  NAND U2990 ( .A(n2620), .B(n527), .Z(n2500) );
  XOR U2991 ( .A(n2499), .B(n2621), .Z(n2501) );
  ANDN U2992 ( .A(n558), .B(n2622), .Z(n2621) );
  ANDN U2993 ( .A(n2623), .B(n2624), .Z(n2499) );
  NAND U2994 ( .A(n2625), .B(n2626), .Z(n2623) );
  IV U2995 ( .A(n2504), .Z(n2506) );
  MUX U2996 ( .IN0(o[2]), .IN1(n390), .SEL(n479), .F(\_MxM/n315 ) );
  IV U2997 ( .A(n2630), .Z(n479) );
  XNOR U2998 ( .A(n2628), .B(\_MxM/Y0[3] ), .Z(n390) );
  XNOR U2999 ( .A(n2631), .B(n2632), .Z(n2628) );
  XOR U3000 ( .A(n2629), .B(n2633), .Z(n2631) );
  AND U3001 ( .A(n491), .B(n2634), .Z(n2633) );
  XNOR U3002 ( .A(n2512), .B(n2632), .Z(n2634) );
  NANDN U3003 ( .B(n2635), .A(n2636), .Z(n2511) );
  XNOR U3004 ( .A(n2637), .B(n2563), .Z(n2543) );
  XNOR U3005 ( .A(n2521), .B(n2520), .Z(n2563) );
  XOR U3006 ( .A(n2638), .B(n2529), .Z(n2520) );
  XNOR U3007 ( .A(n2517), .B(n2518), .Z(n2529) );
  NAND U3008 ( .A(n1938), .B(n816), .Z(n2518) );
  XNOR U3009 ( .A(n2516), .B(n2639), .Z(n2517) );
  ANDN U3010 ( .A(n1943), .B(n818), .Z(n2639) );
  XNOR U3011 ( .A(n2528), .B(n2519), .Z(n2638) );
  XOR U3012 ( .A(n2646), .B(n2525), .Z(n2528) );
  XNOR U3013 ( .A(n2524), .B(n2647), .Z(n2525) );
  ANDN U3014 ( .A(n2173), .B(n717), .Z(n2647) );
  AND U3015 ( .A(n2166), .B(n715), .Z(n2526) );
  XNOR U3016 ( .A(n2537), .B(n2536), .Z(n2521) );
  XOR U3017 ( .A(n2654), .B(n2533), .Z(n2536) );
  XNOR U3018 ( .A(n2532), .B(n2655), .Z(n2533) );
  ANDN U3019 ( .A(n1744), .B(n950), .Z(n2655) );
  AND U3020 ( .A(n1737), .B(n948), .Z(n2534) );
  XNOR U3021 ( .A(n2540), .B(n2541), .Z(n2537) );
  NAND U3022 ( .A(n1542), .B(n1089), .Z(n2541) );
  XNOR U3023 ( .A(n2539), .B(n2662), .Z(n2540) );
  ANDN U3024 ( .A(n1547), .B(n1091), .Z(n2662) );
  XNOR U3025 ( .A(n2562), .B(n2542), .Z(n2637) );
  XOR U3026 ( .A(n2669), .B(n2560), .Z(n2562) );
  XOR U3027 ( .A(n2554), .B(n2553), .Z(n2560) );
  XOR U3028 ( .A(n2674), .B(n2551), .Z(n2670) );
  AND U3029 ( .A(n2675), .B(n556), .Z(n2551) );
  NAND U3030 ( .A(n2676), .B(n2550), .Z(n2674) );
  XOR U3031 ( .A(n2677), .B(n2678), .Z(n2550) );
  AND U3032 ( .A(n2679), .B(n2680), .Z(n2678) );
  XNOR U3033 ( .A(n2681), .B(n2677), .Z(n2680) );
  NANDN U3034 ( .B(n559), .A(n2682), .Z(n2676) );
  XNOR U3035 ( .A(n2557), .B(n2558), .Z(n2554) );
  NAND U3036 ( .A(n2428), .B(n631), .Z(n2558) );
  XNOR U3037 ( .A(n2556), .B(n2683), .Z(n2557) );
  ANDN U3038 ( .A(n2433), .B(n633), .Z(n2683) );
  XOR U3039 ( .A(n2684), .B(n2685), .Z(n2556) );
  AND U3040 ( .A(n2686), .B(n2687), .Z(n2685) );
  XOR U3041 ( .A(n2688), .B(n2684), .Z(n2687) );
  XNOR U3042 ( .A(n2559), .B(n2561), .Z(n2669) );
  XNOR U3043 ( .A(n2692), .B(n2695), .Z(n2694) );
  XNOR U3044 ( .A(n2579), .B(n2578), .Z(n2544) );
  XOR U3045 ( .A(n2696), .B(n2587), .Z(n2578) );
  XNOR U3046 ( .A(n2572), .B(n2571), .Z(n2587) );
  XOR U3047 ( .A(n2697), .B(n2568), .Z(n2571) );
  XNOR U3048 ( .A(n2567), .B(n2698), .Z(n2568) );
  ANDN U3049 ( .A(n1036), .B(n1618), .Z(n2698) );
  AND U3050 ( .A(n1616), .B(n973), .Z(n2569) );
  XNOR U3051 ( .A(n2575), .B(n2576), .Z(n2572) );
  NANDN U3052 ( .B(n838), .A(n1813), .Z(n2576) );
  XNOR U3053 ( .A(n2574), .B(n2705), .Z(n2575) );
  ANDN U3054 ( .A(n908), .B(n1815), .Z(n2705) );
  XNOR U3055 ( .A(n2586), .B(n2577), .Z(n2696) );
  XOR U3056 ( .A(n2712), .B(n2595), .Z(n2586) );
  XNOR U3057 ( .A(n2583), .B(n2584), .Z(n2595) );
  NAND U3058 ( .A(n1423), .B(n1207), .Z(n2584) );
  XNOR U3059 ( .A(n2582), .B(n2713), .Z(n2583) );
  ANDN U3060 ( .A(n1214), .B(n1425), .Z(n2713) );
  XNOR U3061 ( .A(n2594), .B(n2585), .Z(n2712) );
  XOR U3062 ( .A(n2720), .B(n2591), .Z(n2594) );
  XNOR U3063 ( .A(n2590), .B(n2721), .Z(n2591) );
  ANDN U3064 ( .A(n1398), .B(n1250), .Z(n2721) );
  AND U3065 ( .A(n1248), .B(n1391), .Z(n2592) );
  XNOR U3066 ( .A(n2603), .B(n2602), .Z(n2579) );
  XOR U3067 ( .A(n2728), .B(n2611), .Z(n2602) );
  XNOR U3068 ( .A(n2599), .B(n2600), .Z(n2611) );
  NANDN U3069 ( .B(n651), .A(n2253), .Z(n2600) );
  XNOR U3070 ( .A(n2598), .B(n2729), .Z(n2599) );
  ANDN U3071 ( .A(n692), .B(n2255), .Z(n2729) );
  XNOR U3072 ( .A(n2610), .B(n2601), .Z(n2728) );
  XOR U3073 ( .A(n2736), .B(n2607), .Z(n2610) );
  XNOR U3074 ( .A(n2606), .B(n2737), .Z(n2607) );
  ANDN U3075 ( .A(n799), .B(n2028), .Z(n2737) );
  AND U3076 ( .A(n2026), .B(n745), .Z(n2608) );
  XOR U3077 ( .A(n2619), .B(n2618), .Z(n2603) );
  XOR U3078 ( .A(n2744), .B(n2615), .Z(n2618) );
  XNOR U3079 ( .A(n2614), .B(n2745), .Z(n2615) );
  ANDN U3080 ( .A(n624), .B(n2497), .Z(n2745) );
  AND U3081 ( .A(n2495), .B(n583), .Z(n2616) );
  XOR U3082 ( .A(n2626), .B(n2625), .Z(n2619) );
  NAND U3083 ( .A(n2752), .B(n527), .Z(n2625) );
  XNOR U3084 ( .A(n2624), .B(n2753), .Z(n2626) );
  ANDN U3085 ( .A(n558), .B(n2754), .Z(n2753) );
  NAND U3086 ( .A(n2755), .B(n2756), .Z(n2624) );
  NAND U3087 ( .A(n2757), .B(n2758), .Z(n2755) );
  IV U3088 ( .A(n2627), .Z(n2629) );
  MUX U3089 ( .IN0(n387), .IN1(o[1]), .SEL(n2630), .F(\_MxM/n314 ) );
  XNOR U3090 ( .A(n2760), .B(\_MxM/Y0[2] ), .Z(n387) );
  XNOR U3091 ( .A(n2761), .B(n2762), .Z(n2760) );
  XNOR U3092 ( .A(n2759), .B(n2763), .Z(n2761) );
  AND U3093 ( .A(n491), .B(n2764), .Z(n2763) );
  XNOR U3094 ( .A(n2635), .B(n2762), .Z(n2764) );
  XOR U3095 ( .A(n2762), .B(n2636), .Z(n2635) );
  ANDN U3096 ( .A(n2765), .B(n2766), .Z(n2636) );
  XNOR U3097 ( .A(n2767), .B(n2691), .Z(n2667) );
  XNOR U3098 ( .A(n2645), .B(n2644), .Z(n2691) );
  XOR U3099 ( .A(n2768), .B(n2653), .Z(n2644) );
  XNOR U3100 ( .A(n2641), .B(n2642), .Z(n2653) );
  NAND U3101 ( .A(n1938), .B(n880), .Z(n2642) );
  XNOR U3102 ( .A(n2640), .B(n2769), .Z(n2641) );
  ANDN U3103 ( .A(n1943), .B(n882), .Z(n2769) );
  XNOR U3104 ( .A(n2652), .B(n2643), .Z(n2768) );
  XOR U3105 ( .A(n2776), .B(n2649), .Z(n2652) );
  XNOR U3106 ( .A(n2648), .B(n2777), .Z(n2649) );
  ANDN U3107 ( .A(n2173), .B(n759), .Z(n2777) );
  AND U3108 ( .A(n2166), .B(n757), .Z(n2650) );
  XNOR U3109 ( .A(n2661), .B(n2660), .Z(n2645) );
  XOR U3110 ( .A(n2784), .B(n2657), .Z(n2660) );
  XNOR U3111 ( .A(n2656), .B(n2785), .Z(n2657) );
  ANDN U3112 ( .A(n1744), .B(n1017), .Z(n2785) );
  AND U3113 ( .A(n1737), .B(n1015), .Z(n2658) );
  XNOR U3114 ( .A(n2664), .B(n2665), .Z(n2661) );
  NAND U3115 ( .A(n1542), .B(n1167), .Z(n2665) );
  XNOR U3116 ( .A(n2663), .B(n2792), .Z(n2664) );
  ANDN U3117 ( .A(n1547), .B(n1169), .Z(n2792) );
  XOR U3118 ( .A(n2690), .B(n2666), .Z(n2767) );
  XNOR U3119 ( .A(n2799), .B(n2695), .Z(n2690) );
  XNOR U3120 ( .A(n2673), .B(n2672), .Z(n2695) );
  XOR U3121 ( .A(n2800), .B(n2679), .Z(n2672) );
  XNOR U3122 ( .A(n2677), .B(n2801), .Z(n2679) );
  ANDN U3123 ( .A(n2682), .B(n589), .Z(n2801) );
  AND U3124 ( .A(n2675), .B(n587), .Z(n2681) );
  XNOR U3125 ( .A(n2686), .B(n2688), .Z(n2673) );
  NAND U3126 ( .A(n2428), .B(n671), .Z(n2688) );
  XNOR U3127 ( .A(n2684), .B(n2808), .Z(n2686) );
  ANDN U3128 ( .A(n2433), .B(n673), .Z(n2808) );
  XNOR U3129 ( .A(n2693), .B(n2689), .Z(n2799) );
  XOR U3130 ( .A(n2692), .B(n2815), .Z(n2693) );
  AND U3131 ( .A(n2816), .B(n2817), .Z(n2815) );
  NANDN U3132 ( .B(n2818), .A(n2819), .Z(n2817) );
  AND U3133 ( .A(n2820), .B(n2821), .Z(n2816) );
  NANDN U3134 ( .B(n2822), .A(n526), .Z(n2821) );
  OR U3135 ( .A(n2823), .B(n2824), .Z(n2820) );
  XNOR U3136 ( .A(n2711), .B(n2710), .Z(n2668) );
  XOR U3137 ( .A(n2828), .B(n2719), .Z(n2710) );
  XNOR U3138 ( .A(n2704), .B(n2703), .Z(n2719) );
  XOR U3139 ( .A(n2829), .B(n2700), .Z(n2703) );
  XNOR U3140 ( .A(n2699), .B(n2830), .Z(n2700) );
  ANDN U3141 ( .A(n1036), .B(n1714), .Z(n2830) );
  AND U3142 ( .A(n1712), .B(n973), .Z(n2701) );
  XNOR U3143 ( .A(n2707), .B(n2708), .Z(n2704) );
  NANDN U3144 ( .B(n838), .A(n1919), .Z(n2708) );
  XNOR U3145 ( .A(n2706), .B(n2837), .Z(n2707) );
  ANDN U3146 ( .A(n908), .B(n1921), .Z(n2837) );
  XNOR U3147 ( .A(n2718), .B(n2709), .Z(n2828) );
  XOR U3148 ( .A(n2844), .B(n2727), .Z(n2718) );
  XNOR U3149 ( .A(n2715), .B(n2716), .Z(n2727) );
  NAND U3150 ( .A(n1520), .B(n1207), .Z(n2716) );
  XNOR U3151 ( .A(n2714), .B(n2845), .Z(n2715) );
  ANDN U3152 ( .A(n1214), .B(n1522), .Z(n2845) );
  XNOR U3153 ( .A(n2726), .B(n2717), .Z(n2844) );
  XOR U3154 ( .A(n2852), .B(n2723), .Z(n2726) );
  XNOR U3155 ( .A(n2722), .B(n2853), .Z(n2723) );
  ANDN U3156 ( .A(n1398), .B(n1334), .Z(n2853) );
  AND U3157 ( .A(n1332), .B(n1391), .Z(n2724) );
  XNOR U3158 ( .A(n2735), .B(n2734), .Z(n2711) );
  XOR U3159 ( .A(n2860), .B(n2743), .Z(n2734) );
  XNOR U3160 ( .A(n2731), .B(n2732), .Z(n2743) );
  NANDN U3161 ( .B(n651), .A(n2373), .Z(n2732) );
  XNOR U3162 ( .A(n2730), .B(n2861), .Z(n2731) );
  ANDN U3163 ( .A(n692), .B(n2375), .Z(n2861) );
  XNOR U3164 ( .A(n2742), .B(n2733), .Z(n2860) );
  XOR U3165 ( .A(n2868), .B(n2739), .Z(n2742) );
  XNOR U3166 ( .A(n2738), .B(n2869), .Z(n2739) );
  ANDN U3167 ( .A(n799), .B(n2136), .Z(n2869) );
  AND U3168 ( .A(n2134), .B(n745), .Z(n2740) );
  XOR U3169 ( .A(n2751), .B(n2750), .Z(n2735) );
  XOR U3170 ( .A(n2876), .B(n2747), .Z(n2750) );
  XNOR U3171 ( .A(n2746), .B(n2877), .Z(n2747) );
  ANDN U3172 ( .A(n624), .B(n2622), .Z(n2877) );
  AND U3173 ( .A(n2620), .B(n583), .Z(n2748) );
  XOR U3174 ( .A(n2758), .B(n2757), .Z(n2751) );
  NAND U3175 ( .A(n2884), .B(n527), .Z(n2757) );
  XOR U3176 ( .A(n2756), .B(n2885), .Z(n2758) );
  ANDN U3177 ( .A(n558), .B(n2886), .Z(n2885) );
  ANDN U3178 ( .A(n2887), .B(n2888), .Z(n2756) );
  NAND U3179 ( .A(n2889), .B(n2890), .Z(n2887) );
  MUX U3180 ( .IN0(n383), .IN1(o[0]), .SEL(n2630), .F(\_MxM/n313 ) );
  NANDN U3181 ( .B(rst), .A(n478), .Z(n2630) );
  AND U3182 ( .A(n2893), .B(n2894), .Z(n478) );
  AND U3183 ( .A(n2895), .B(n2896), .Z(n2894) );
  ANDN U3184 ( .A(n2897), .B(\_MxM/n[3] ), .Z(n2896) );
  NOR U3185 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n2897) );
  ANDN U3186 ( .A(n2898), .B(\_MxM/n[13] ), .Z(n2895) );
  NOR U3187 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n2898) );
  AND U3188 ( .A(n2899), .B(n2900), .Z(n2893) );
  AND U3189 ( .A(n375), .B(n2901), .Z(n2900) );
  NOR U3190 ( .A(\_MxM/n[0] ), .B(\_MxM/n[10] ), .Z(n2901) );
  NOR U3191 ( .A(\_MxM/n[6] ), .B(\_MxM/n[7] ), .Z(n375) );
  AND U3192 ( .A(n373), .B(n376), .Z(n2899) );
  NOR U3193 ( .A(\_MxM/n[4] ), .B(\_MxM/n[5] ), .Z(n376) );
  NOR U3194 ( .A(\_MxM/n[12] ), .B(\_MxM/n[11] ), .Z(n373) );
  XOR U3195 ( .A(n2892), .B(\_MxM/Y0[1] ), .Z(n383) );
  XOR U3196 ( .A(n2902), .B(n2903), .Z(n2892) );
  XOR U3197 ( .A(n2904), .B(n2891), .Z(n2902) );
  NAND U3198 ( .A(n2905), .B(n491), .Z(n2904) );
  XOR U3199 ( .A(e_input[31]), .B(g_input[31]), .Z(n491) );
  XOR U3200 ( .A(n2765), .B(n2903), .Z(n2905) );
  XOR U3201 ( .A(n2766), .B(n2903), .Z(n2765) );
  XNOR U3202 ( .A(n2906), .B(n2814), .Z(n2797) );
  XNOR U3203 ( .A(n2775), .B(n2774), .Z(n2814) );
  XOR U3204 ( .A(n2907), .B(n2783), .Z(n2774) );
  XNOR U3205 ( .A(n2771), .B(n2772), .Z(n2783) );
  NAND U3206 ( .A(n1938), .B(n948), .Z(n2772) );
  XNOR U3207 ( .A(n2770), .B(n2908), .Z(n2771) );
  ANDN U3208 ( .A(n1943), .B(n950), .Z(n2908) );
  XNOR U3209 ( .A(n2782), .B(n2773), .Z(n2907) );
  XOR U3210 ( .A(n2915), .B(n2779), .Z(n2782) );
  XNOR U3211 ( .A(n2778), .B(n2916), .Z(n2779) );
  ANDN U3212 ( .A(n2173), .B(n818), .Z(n2916) );
  AND U3213 ( .A(n2166), .B(n816), .Z(n2780) );
  XNOR U3214 ( .A(n2791), .B(n2790), .Z(n2775) );
  XOR U3215 ( .A(n2923), .B(n2787), .Z(n2790) );
  XNOR U3216 ( .A(n2786), .B(n2924), .Z(n2787) );
  ANDN U3217 ( .A(n1744), .B(n1091), .Z(n2924) );
  AND U3218 ( .A(n1737), .B(n1089), .Z(n2788) );
  XNOR U3219 ( .A(n2794), .B(n2795), .Z(n2791) );
  NAND U3220 ( .A(n1542), .B(n1248), .Z(n2795) );
  XNOR U3221 ( .A(n2793), .B(n2931), .Z(n2794) );
  ANDN U3222 ( .A(n1547), .B(n1250), .Z(n2931) );
  XOR U3223 ( .A(n2813), .B(n2796), .Z(n2906) );
  XNOR U3224 ( .A(n2938), .B(n2827), .Z(n2813) );
  XNOR U3225 ( .A(n2807), .B(n2806), .Z(n2827) );
  XOR U3226 ( .A(n2939), .B(n2803), .Z(n2806) );
  XNOR U3227 ( .A(n2802), .B(n2940), .Z(n2803) );
  ANDN U3228 ( .A(n2682), .B(n633), .Z(n2940) );
  AND U3229 ( .A(n2675), .B(n631), .Z(n2804) );
  XNOR U3230 ( .A(n2810), .B(n2811), .Z(n2807) );
  NAND U3231 ( .A(n2428), .B(n715), .Z(n2811) );
  XNOR U3232 ( .A(n2809), .B(n2947), .Z(n2810) );
  ANDN U3233 ( .A(n2433), .B(n717), .Z(n2947) );
  XOR U3234 ( .A(n2826), .B(n2812), .Z(n2938) );
  XNOR U3235 ( .A(n2954), .B(n2823), .Z(n2826) );
  XNOR U3236 ( .A(n2955), .B(n2819), .Z(n2823) );
  AND U3237 ( .A(n2956), .B(n556), .Z(n2819) );
  NAND U3238 ( .A(n2957), .B(n2818), .Z(n2955) );
  NANDN U3239 ( .B(n559), .A(n2961), .Z(n2957) );
  XNOR U3240 ( .A(n2824), .B(n2825), .Z(n2954) );
  XNOR U3241 ( .A(n2965), .B(n2968), .Z(n2967) );
  XNOR U3242 ( .A(n2843), .B(n2842), .Z(n2798) );
  XOR U3243 ( .A(n2969), .B(n2851), .Z(n2842) );
  XNOR U3244 ( .A(n2836), .B(n2835), .Z(n2851) );
  XOR U3245 ( .A(n2970), .B(n2832), .Z(n2835) );
  XNOR U3246 ( .A(n2831), .B(n2971), .Z(n2832) );
  ANDN U3247 ( .A(n1036), .B(n1815), .Z(n2971) );
  AND U3248 ( .A(n1813), .B(n973), .Z(n2833) );
  XNOR U3249 ( .A(n2839), .B(n2840), .Z(n2836) );
  NANDN U3250 ( .B(n838), .A(n2026), .Z(n2840) );
  XNOR U3251 ( .A(n2838), .B(n2978), .Z(n2839) );
  ANDN U3252 ( .A(n908), .B(n2028), .Z(n2978) );
  XNOR U3253 ( .A(n2850), .B(n2841), .Z(n2969) );
  XOR U3254 ( .A(n2985), .B(n2859), .Z(n2850) );
  XNOR U3255 ( .A(n2847), .B(n2848), .Z(n2859) );
  NAND U3256 ( .A(n1616), .B(n1207), .Z(n2848) );
  XNOR U3257 ( .A(n2846), .B(n2986), .Z(n2847) );
  ANDN U3258 ( .A(n1214), .B(n1618), .Z(n2986) );
  XNOR U3259 ( .A(n2858), .B(n2849), .Z(n2985) );
  XOR U3260 ( .A(n2993), .B(n2855), .Z(n2858) );
  XNOR U3261 ( .A(n2854), .B(n2994), .Z(n2855) );
  ANDN U3262 ( .A(n1398), .B(n1425), .Z(n2994) );
  AND U3263 ( .A(n1423), .B(n1391), .Z(n2856) );
  XNOR U3264 ( .A(n2867), .B(n2866), .Z(n2843) );
  XOR U3265 ( .A(n3001), .B(n2875), .Z(n2866) );
  XNOR U3266 ( .A(n2863), .B(n2864), .Z(n2875) );
  NANDN U3267 ( .B(n651), .A(n2495), .Z(n2864) );
  XNOR U3268 ( .A(n2862), .B(n3002), .Z(n2863) );
  ANDN U3269 ( .A(n692), .B(n2497), .Z(n3002) );
  XNOR U3270 ( .A(n2874), .B(n2865), .Z(n3001) );
  XOR U3271 ( .A(n3009), .B(n2871), .Z(n2874) );
  XNOR U3272 ( .A(n2870), .B(n3010), .Z(n2871) );
  ANDN U3273 ( .A(n799), .B(n2255), .Z(n3010) );
  AND U3274 ( .A(n2253), .B(n745), .Z(n2872) );
  XOR U3275 ( .A(n2883), .B(n2882), .Z(n2867) );
  XOR U3276 ( .A(n3017), .B(n2879), .Z(n2882) );
  XNOR U3277 ( .A(n2878), .B(n3018), .Z(n2879) );
  ANDN U3278 ( .A(n624), .B(n2754), .Z(n3018) );
  AND U3279 ( .A(n2752), .B(n583), .Z(n2880) );
  XOR U3280 ( .A(n2890), .B(n2889), .Z(n2883) );
  NAND U3281 ( .A(n3025), .B(n527), .Z(n2889) );
  XNOR U3282 ( .A(n2888), .B(n3026), .Z(n2890) );
  ANDN U3283 ( .A(n558), .B(n3027), .Z(n3026) );
  NAND U3284 ( .A(n3028), .B(n3029), .Z(n2888) );
  NAND U3285 ( .A(n3030), .B(n3031), .Z(n3028) );
  XNOR U3286 ( .A(n3032), .B(n2953), .Z(n2936) );
  XNOR U3287 ( .A(n2914), .B(n2913), .Z(n2953) );
  XOR U3288 ( .A(n3033), .B(n2922), .Z(n2913) );
  XNOR U3289 ( .A(n2910), .B(n2911), .Z(n2922) );
  NAND U3290 ( .A(n1938), .B(n1015), .Z(n2911) );
  XNOR U3291 ( .A(n2909), .B(n3034), .Z(n2910) );
  ANDN U3292 ( .A(n1943), .B(n1017), .Z(n3034) );
  XOR U3293 ( .A(n3035), .B(n3036), .Z(n2909) );
  AND U3294 ( .A(n3037), .B(n3038), .Z(n3036) );
  XOR U3295 ( .A(n3039), .B(n3035), .Z(n3038) );
  XNOR U3296 ( .A(n2921), .B(n2912), .Z(n3033) );
  XOR U3297 ( .A(n3043), .B(n2918), .Z(n2921) );
  XNOR U3298 ( .A(n2917), .B(n3044), .Z(n2918) );
  ANDN U3299 ( .A(n2173), .B(n882), .Z(n3044) );
  XOR U3300 ( .A(n3045), .B(n3046), .Z(n2917) );
  AND U3301 ( .A(n3047), .B(n3048), .Z(n3046) );
  XNOR U3302 ( .A(n3049), .B(n3045), .Z(n3048) );
  AND U3303 ( .A(n2166), .B(n880), .Z(n2919) );
  XNOR U3304 ( .A(n2930), .B(n2929), .Z(n2914) );
  XOR U3305 ( .A(n3053), .B(n2926), .Z(n2929) );
  XNOR U3306 ( .A(n2925), .B(n3054), .Z(n2926) );
  ANDN U3307 ( .A(n1744), .B(n1169), .Z(n3054) );
  AND U3308 ( .A(n1737), .B(n1167), .Z(n2927) );
  XNOR U3309 ( .A(n2933), .B(n2934), .Z(n2930) );
  NAND U3310 ( .A(n1542), .B(n1332), .Z(n2934) );
  XNOR U3311 ( .A(n2932), .B(n3061), .Z(n2933) );
  ANDN U3312 ( .A(n1547), .B(n1334), .Z(n3061) );
  XNOR U3313 ( .A(n2952), .B(n2935), .Z(n3032) );
  XNOR U3314 ( .A(n3065), .B(n3066), .Z(n2935) );
  XNOR U3315 ( .A(n3067), .B(n2964), .Z(n2952) );
  XNOR U3316 ( .A(n2946), .B(n2945), .Z(n2964) );
  XOR U3317 ( .A(n3068), .B(n2942), .Z(n2945) );
  XNOR U3318 ( .A(n2941), .B(n3069), .Z(n2942) );
  ANDN U3319 ( .A(n2682), .B(n673), .Z(n3069) );
  XOR U3320 ( .A(n3070), .B(n3071), .Z(n2941) );
  AND U3321 ( .A(n3072), .B(n3073), .Z(n3071) );
  XNOR U3322 ( .A(n3074), .B(n3070), .Z(n3073) );
  AND U3323 ( .A(n2675), .B(n671), .Z(n2943) );
  XNOR U3324 ( .A(n2949), .B(n2950), .Z(n2946) );
  NAND U3325 ( .A(n2428), .B(n757), .Z(n2950) );
  XNOR U3326 ( .A(n2948), .B(n3078), .Z(n2949) );
  ANDN U3327 ( .A(n2433), .B(n759), .Z(n3078) );
  XOR U3328 ( .A(n3079), .B(n3080), .Z(n2948) );
  AND U3329 ( .A(n3081), .B(n3082), .Z(n3080) );
  XOR U3330 ( .A(n3083), .B(n3079), .Z(n3082) );
  XNOR U3331 ( .A(n2963), .B(n2951), .Z(n3067) );
  XOR U3332 ( .A(n3084), .B(n3085), .Z(n2951) );
  AND U3333 ( .A(n3086), .B(n3087), .Z(n3085) );
  XOR U3334 ( .A(n3088), .B(n3089), .Z(n3087) );
  XNOR U3335 ( .A(n3090), .B(n3084), .Z(n3088) );
  XNOR U3336 ( .A(n3041), .B(n3091), .Z(n3086) );
  XNOR U3337 ( .A(n3084), .B(n3042), .Z(n3091) );
  XNOR U3338 ( .A(n3060), .B(n3059), .Z(n3042) );
  XOR U3339 ( .A(n3092), .B(n3056), .Z(n3059) );
  XNOR U3340 ( .A(n3055), .B(n3093), .Z(n3056) );
  ANDN U3341 ( .A(n1744), .B(n1250), .Z(n3093) );
  AND U3342 ( .A(n1737), .B(n1248), .Z(n3057) );
  XNOR U3343 ( .A(n3063), .B(n3064), .Z(n3060) );
  NAND U3344 ( .A(n1423), .B(n1542), .Z(n3064) );
  XNOR U3345 ( .A(n3062), .B(n3100), .Z(n3063) );
  ANDN U3346 ( .A(n1547), .B(n1425), .Z(n3100) );
  XOR U3347 ( .A(n3104), .B(n3052), .Z(n3041) );
  XNOR U3348 ( .A(n3037), .B(n3039), .Z(n3052) );
  NAND U3349 ( .A(n1938), .B(n1089), .Z(n3039) );
  XNOR U3350 ( .A(n3035), .B(n3105), .Z(n3037) );
  ANDN U3351 ( .A(n1943), .B(n1091), .Z(n3105) );
  XNOR U3352 ( .A(n3051), .B(n3040), .Z(n3104) );
  XOR U3353 ( .A(n3112), .B(n3047), .Z(n3051) );
  XNOR U3354 ( .A(n3045), .B(n3113), .Z(n3047) );
  ANDN U3355 ( .A(n2173), .B(n950), .Z(n3113) );
  XOR U3356 ( .A(n3114), .B(n3115), .Z(n3045) );
  AND U3357 ( .A(n3116), .B(n3117), .Z(n3115) );
  XNOR U3358 ( .A(n3118), .B(n3114), .Z(n3117) );
  AND U3359 ( .A(n2166), .B(n948), .Z(n3049) );
  XOR U3360 ( .A(n3122), .B(n3123), .Z(n3084) );
  AND U3361 ( .A(n3124), .B(n3125), .Z(n3123) );
  XOR U3362 ( .A(n3126), .B(n3127), .Z(n3125) );
  XOR U3363 ( .A(n3122), .B(n3128), .Z(n3127) );
  XNOR U3364 ( .A(n3110), .B(n3129), .Z(n3124) );
  XNOR U3365 ( .A(n3122), .B(n3111), .Z(n3129) );
  XNOR U3366 ( .A(n3099), .B(n3098), .Z(n3111) );
  XOR U3367 ( .A(n3130), .B(n3095), .Z(n3098) );
  XNOR U3368 ( .A(n3094), .B(n3131), .Z(n3095) );
  ANDN U3369 ( .A(n1744), .B(n1334), .Z(n3131) );
  XOR U3370 ( .A(n3132), .B(n3133), .Z(n3094) );
  AND U3371 ( .A(n3134), .B(n3135), .Z(n3133) );
  XNOR U3372 ( .A(n3136), .B(n3132), .Z(n3135) );
  AND U3373 ( .A(n1737), .B(n1332), .Z(n3096) );
  XNOR U3374 ( .A(n3102), .B(n3103), .Z(n3099) );
  NAND U3375 ( .A(n1520), .B(n1542), .Z(n3103) );
  XNOR U3376 ( .A(n3101), .B(n3140), .Z(n3102) );
  ANDN U3377 ( .A(n1547), .B(n1522), .Z(n3140) );
  XOR U3378 ( .A(n3141), .B(n3142), .Z(n3101) );
  AND U3379 ( .A(n3143), .B(n3144), .Z(n3142) );
  XOR U3380 ( .A(n3145), .B(n3141), .Z(n3144) );
  XOR U3381 ( .A(n3146), .B(n3121), .Z(n3110) );
  XNOR U3382 ( .A(n3107), .B(n3108), .Z(n3121) );
  NAND U3383 ( .A(n1938), .B(n1167), .Z(n3108) );
  XNOR U3384 ( .A(n3106), .B(n3147), .Z(n3107) );
  ANDN U3385 ( .A(n1943), .B(n1169), .Z(n3147) );
  XOR U3386 ( .A(n3148), .B(n3149), .Z(n3106) );
  AND U3387 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U3388 ( .A(n3152), .B(n3148), .Z(n3151) );
  XNOR U3389 ( .A(n3120), .B(n3109), .Z(n3146) );
  XOR U3390 ( .A(n3156), .B(n3116), .Z(n3120) );
  XNOR U3391 ( .A(n3114), .B(n3157), .Z(n3116) );
  ANDN U3392 ( .A(n2173), .B(n1017), .Z(n3157) );
  XOR U3393 ( .A(n3158), .B(n3159), .Z(n3114) );
  AND U3394 ( .A(n3160), .B(n3161), .Z(n3159) );
  XNOR U3395 ( .A(n3162), .B(n3158), .Z(n3161) );
  XOR U3396 ( .A(n3163), .B(n3118), .Z(n3156) );
  AND U3397 ( .A(n2166), .B(n1015), .Z(n3118) );
  IV U3398 ( .A(n3119), .Z(n3163) );
  XOR U3399 ( .A(n3167), .B(n3168), .Z(n3122) );
  AND U3400 ( .A(n3169), .B(n3170), .Z(n3168) );
  XOR U3401 ( .A(n3171), .B(n3172), .Z(n3170) );
  XOR U3402 ( .A(n3167), .B(n3173), .Z(n3172) );
  XNOR U3403 ( .A(n3154), .B(n3174), .Z(n3169) );
  XNOR U3404 ( .A(n3167), .B(n3155), .Z(n3174) );
  XNOR U3405 ( .A(n3139), .B(n3138), .Z(n3155) );
  XOR U3406 ( .A(n3175), .B(n3134), .Z(n3138) );
  XNOR U3407 ( .A(n3132), .B(n3176), .Z(n3134) );
  ANDN U3408 ( .A(n1744), .B(n1425), .Z(n3176) );
  XOR U3409 ( .A(n3177), .B(n3178), .Z(n3132) );
  AND U3410 ( .A(n3179), .B(n3180), .Z(n3178) );
  XNOR U3411 ( .A(n3181), .B(n3177), .Z(n3180) );
  AND U3412 ( .A(n1423), .B(n1737), .Z(n3136) );
  XNOR U3413 ( .A(n3143), .B(n3145), .Z(n3139) );
  NAND U3414 ( .A(n1616), .B(n1542), .Z(n3145) );
  XNOR U3415 ( .A(n3141), .B(n3185), .Z(n3143) );
  ANDN U3416 ( .A(n1547), .B(n1618), .Z(n3185) );
  XOR U3417 ( .A(n3189), .B(n3166), .Z(n3154) );
  XNOR U3418 ( .A(n3150), .B(n3152), .Z(n3166) );
  NAND U3419 ( .A(n1938), .B(n1248), .Z(n3152) );
  XNOR U3420 ( .A(n3148), .B(n3190), .Z(n3150) );
  ANDN U3421 ( .A(n1943), .B(n1250), .Z(n3190) );
  XOR U3422 ( .A(n3191), .B(n3192), .Z(n3148) );
  AND U3423 ( .A(n3193), .B(n3194), .Z(n3192) );
  XOR U3424 ( .A(n3195), .B(n3191), .Z(n3194) );
  XNOR U3425 ( .A(n3165), .B(n3153), .Z(n3189) );
  XOR U3426 ( .A(n3199), .B(n3160), .Z(n3165) );
  XNOR U3427 ( .A(n3158), .B(n3200), .Z(n3160) );
  ANDN U3428 ( .A(n2173), .B(n1091), .Z(n3200) );
  XOR U3429 ( .A(n3201), .B(n3202), .Z(n3158) );
  AND U3430 ( .A(n3203), .B(n3204), .Z(n3202) );
  XNOR U3431 ( .A(n3205), .B(n3201), .Z(n3204) );
  AND U3432 ( .A(n2166), .B(n1089), .Z(n3162) );
  XOR U3433 ( .A(n3209), .B(n3210), .Z(n3167) );
  AND U3434 ( .A(n3211), .B(n3212), .Z(n3210) );
  XOR U3435 ( .A(n3213), .B(n3214), .Z(n3212) );
  XOR U3436 ( .A(n3209), .B(n3215), .Z(n3214) );
  XNOR U3437 ( .A(n3197), .B(n3216), .Z(n3211) );
  XNOR U3438 ( .A(n3209), .B(n3198), .Z(n3216) );
  XNOR U3439 ( .A(n3184), .B(n3183), .Z(n3198) );
  XOR U3440 ( .A(n3217), .B(n3179), .Z(n3183) );
  XNOR U3441 ( .A(n3177), .B(n3218), .Z(n3179) );
  ANDN U3442 ( .A(n1744), .B(n1522), .Z(n3218) );
  XOR U3443 ( .A(n3219), .B(n3220), .Z(n3177) );
  AND U3444 ( .A(n3221), .B(n3222), .Z(n3220) );
  XNOR U3445 ( .A(n3223), .B(n3219), .Z(n3222) );
  AND U3446 ( .A(n1520), .B(n1737), .Z(n3181) );
  XNOR U3447 ( .A(n3187), .B(n3188), .Z(n3184) );
  NAND U3448 ( .A(n1712), .B(n1542), .Z(n3188) );
  XNOR U3449 ( .A(n3186), .B(n3227), .Z(n3187) );
  ANDN U3450 ( .A(n1547), .B(n1714), .Z(n3227) );
  XOR U3451 ( .A(n3228), .B(n3229), .Z(n3186) );
  AND U3452 ( .A(n3230), .B(n3231), .Z(n3229) );
  XOR U3453 ( .A(n3232), .B(n3228), .Z(n3231) );
  XOR U3454 ( .A(n3233), .B(n3208), .Z(n3197) );
  XNOR U3455 ( .A(n3193), .B(n3195), .Z(n3208) );
  NAND U3456 ( .A(n1938), .B(n1332), .Z(n3195) );
  XNOR U3457 ( .A(n3191), .B(n3234), .Z(n3193) );
  ANDN U3458 ( .A(n1943), .B(n1334), .Z(n3234) );
  XNOR U3459 ( .A(n3207), .B(n3196), .Z(n3233) );
  XOR U3460 ( .A(n3241), .B(n3203), .Z(n3207) );
  XNOR U3461 ( .A(n3201), .B(n3242), .Z(n3203) );
  ANDN U3462 ( .A(n2173), .B(n1169), .Z(n3242) );
  XOR U3463 ( .A(n3243), .B(n3244), .Z(n3201) );
  AND U3464 ( .A(n3245), .B(n3246), .Z(n3244) );
  XNOR U3465 ( .A(n3247), .B(n3243), .Z(n3246) );
  XOR U3466 ( .A(n3248), .B(n3205), .Z(n3241) );
  AND U3467 ( .A(n2166), .B(n1167), .Z(n3205) );
  IV U3468 ( .A(n3206), .Z(n3248) );
  XOR U3469 ( .A(n3252), .B(n3253), .Z(n3209) );
  AND U3470 ( .A(n3254), .B(n3255), .Z(n3253) );
  XOR U3471 ( .A(n3256), .B(n3257), .Z(n3255) );
  XOR U3472 ( .A(n3252), .B(n3258), .Z(n3257) );
  XNOR U3473 ( .A(n3239), .B(n3259), .Z(n3254) );
  XNOR U3474 ( .A(n3252), .B(n3240), .Z(n3259) );
  XNOR U3475 ( .A(n3226), .B(n3225), .Z(n3240) );
  XOR U3476 ( .A(n3260), .B(n3221), .Z(n3225) );
  XNOR U3477 ( .A(n3219), .B(n3261), .Z(n3221) );
  ANDN U3478 ( .A(n1744), .B(n1618), .Z(n3261) );
  XOR U3479 ( .A(n3262), .B(n3263), .Z(n3219) );
  AND U3480 ( .A(n3264), .B(n3265), .Z(n3263) );
  XNOR U3481 ( .A(n3266), .B(n3262), .Z(n3265) );
  AND U3482 ( .A(n1616), .B(n1737), .Z(n3223) );
  XNOR U3483 ( .A(n3230), .B(n3232), .Z(n3226) );
  NAND U3484 ( .A(n1813), .B(n1542), .Z(n3232) );
  XNOR U3485 ( .A(n3228), .B(n3270), .Z(n3230) );
  ANDN U3486 ( .A(n1547), .B(n1815), .Z(n3270) );
  XOR U3487 ( .A(n3274), .B(n3251), .Z(n3239) );
  XNOR U3488 ( .A(n3236), .B(n3237), .Z(n3251) );
  NAND U3489 ( .A(n1423), .B(n1938), .Z(n3237) );
  XNOR U3490 ( .A(n3235), .B(n3275), .Z(n3236) );
  ANDN U3491 ( .A(n1943), .B(n1425), .Z(n3275) );
  XOR U3492 ( .A(n3276), .B(n3277), .Z(n3235) );
  AND U3493 ( .A(n3278), .B(n3279), .Z(n3277) );
  XOR U3494 ( .A(n3280), .B(n3276), .Z(n3279) );
  XNOR U3495 ( .A(n3250), .B(n3238), .Z(n3274) );
  XOR U3496 ( .A(n3284), .B(n3245), .Z(n3250) );
  XNOR U3497 ( .A(n3243), .B(n3285), .Z(n3245) );
  ANDN U3498 ( .A(n2173), .B(n1250), .Z(n3285) );
  XOR U3499 ( .A(n3286), .B(n3287), .Z(n3243) );
  AND U3500 ( .A(n3288), .B(n3289), .Z(n3287) );
  XNOR U3501 ( .A(n3290), .B(n3286), .Z(n3289) );
  AND U3502 ( .A(n2166), .B(n1248), .Z(n3247) );
  XOR U3503 ( .A(n3294), .B(n3295), .Z(n3252) );
  AND U3504 ( .A(n3296), .B(n3297), .Z(n3295) );
  XOR U3505 ( .A(n3298), .B(n3299), .Z(n3297) );
  XOR U3506 ( .A(n3294), .B(n3300), .Z(n3299) );
  XNOR U3507 ( .A(n3282), .B(n3301), .Z(n3296) );
  XNOR U3508 ( .A(n3294), .B(n3283), .Z(n3301) );
  XNOR U3509 ( .A(n3269), .B(n3268), .Z(n3283) );
  XOR U3510 ( .A(n3302), .B(n3264), .Z(n3268) );
  XNOR U3511 ( .A(n3262), .B(n3303), .Z(n3264) );
  ANDN U3512 ( .A(n1744), .B(n1714), .Z(n3303) );
  XOR U3513 ( .A(n3304), .B(n3305), .Z(n3262) );
  AND U3514 ( .A(n3306), .B(n3307), .Z(n3305) );
  XNOR U3515 ( .A(n3308), .B(n3304), .Z(n3307) );
  XOR U3516 ( .A(n3309), .B(n3266), .Z(n3302) );
  AND U3517 ( .A(n1712), .B(n1737), .Z(n3266) );
  IV U3518 ( .A(n3267), .Z(n3309) );
  XNOR U3519 ( .A(n3272), .B(n3273), .Z(n3269) );
  NAND U3520 ( .A(n1919), .B(n1542), .Z(n3273) );
  XNOR U3521 ( .A(n3271), .B(n3313), .Z(n3272) );
  ANDN U3522 ( .A(n1547), .B(n1921), .Z(n3313) );
  XOR U3523 ( .A(n3314), .B(n3315), .Z(n3271) );
  AND U3524 ( .A(n3316), .B(n3317), .Z(n3315) );
  XOR U3525 ( .A(n3318), .B(n3314), .Z(n3317) );
  XOR U3526 ( .A(n3319), .B(n3293), .Z(n3282) );
  XNOR U3527 ( .A(n3278), .B(n3280), .Z(n3293) );
  NAND U3528 ( .A(n1520), .B(n1938), .Z(n3280) );
  XNOR U3529 ( .A(n3276), .B(n3320), .Z(n3278) );
  ANDN U3530 ( .A(n1943), .B(n1522), .Z(n3320) );
  XOR U3531 ( .A(n3321), .B(n3322), .Z(n3276) );
  AND U3532 ( .A(n3323), .B(n3324), .Z(n3322) );
  XOR U3533 ( .A(n3325), .B(n3321), .Z(n3324) );
  XNOR U3534 ( .A(n3292), .B(n3281), .Z(n3319) );
  XOR U3535 ( .A(n3329), .B(n3288), .Z(n3292) );
  XNOR U3536 ( .A(n3286), .B(n3330), .Z(n3288) );
  ANDN U3537 ( .A(n2173), .B(n1334), .Z(n3330) );
  XOR U3538 ( .A(n3331), .B(n3332), .Z(n3286) );
  AND U3539 ( .A(n3333), .B(n3334), .Z(n3332) );
  XNOR U3540 ( .A(n3335), .B(n3331), .Z(n3334) );
  XOR U3541 ( .A(n3336), .B(n3290), .Z(n3329) );
  AND U3542 ( .A(n2166), .B(n1332), .Z(n3290) );
  IV U3543 ( .A(n3291), .Z(n3336) );
  XOR U3544 ( .A(n3340), .B(n3341), .Z(n3294) );
  AND U3545 ( .A(n3342), .B(n3343), .Z(n3341) );
  XOR U3546 ( .A(n3344), .B(n3345), .Z(n3343) );
  XOR U3547 ( .A(n3340), .B(n3346), .Z(n3345) );
  XNOR U3548 ( .A(n3327), .B(n3347), .Z(n3342) );
  XNOR U3549 ( .A(n3340), .B(n3328), .Z(n3347) );
  XNOR U3550 ( .A(n3312), .B(n3311), .Z(n3328) );
  XOR U3551 ( .A(n3348), .B(n3306), .Z(n3311) );
  XNOR U3552 ( .A(n3304), .B(n3349), .Z(n3306) );
  ANDN U3553 ( .A(n1744), .B(n1815), .Z(n3349) );
  XOR U3554 ( .A(n3350), .B(n3351), .Z(n3304) );
  AND U3555 ( .A(n3352), .B(n3353), .Z(n3351) );
  XNOR U3556 ( .A(n3354), .B(n3350), .Z(n3353) );
  XOR U3557 ( .A(n3355), .B(n3308), .Z(n3348) );
  AND U3558 ( .A(n1813), .B(n1737), .Z(n3308) );
  IV U3559 ( .A(n3310), .Z(n3355) );
  XNOR U3560 ( .A(n3316), .B(n3318), .Z(n3312) );
  NAND U3561 ( .A(n2026), .B(n1542), .Z(n3318) );
  XNOR U3562 ( .A(n3314), .B(n3359), .Z(n3316) );
  ANDN U3563 ( .A(n1547), .B(n2028), .Z(n3359) );
  XOR U3564 ( .A(n3360), .B(n3361), .Z(n3314) );
  AND U3565 ( .A(n3362), .B(n3363), .Z(n3361) );
  XOR U3566 ( .A(n3364), .B(n3360), .Z(n3363) );
  XOR U3567 ( .A(n3365), .B(n3339), .Z(n3327) );
  XNOR U3568 ( .A(n3323), .B(n3325), .Z(n3339) );
  NAND U3569 ( .A(n1616), .B(n1938), .Z(n3325) );
  XNOR U3570 ( .A(n3321), .B(n3366), .Z(n3323) );
  ANDN U3571 ( .A(n1943), .B(n1618), .Z(n3366) );
  XNOR U3572 ( .A(n3338), .B(n3326), .Z(n3365) );
  XOR U3573 ( .A(n3373), .B(n3333), .Z(n3338) );
  XNOR U3574 ( .A(n3331), .B(n3374), .Z(n3333) );
  ANDN U3575 ( .A(n2173), .B(n1425), .Z(n3374) );
  XOR U3576 ( .A(n3375), .B(n3376), .Z(n3331) );
  AND U3577 ( .A(n3377), .B(n3378), .Z(n3376) );
  XNOR U3578 ( .A(n3379), .B(n3375), .Z(n3378) );
  XOR U3579 ( .A(n3380), .B(n3335), .Z(n3373) );
  AND U3580 ( .A(n1423), .B(n2166), .Z(n3335) );
  IV U3581 ( .A(n3337), .Z(n3380) );
  XOR U3582 ( .A(n3384), .B(n3385), .Z(n3340) );
  AND U3583 ( .A(n3386), .B(n3387), .Z(n3385) );
  XOR U3584 ( .A(n3388), .B(n3389), .Z(n3387) );
  XOR U3585 ( .A(n3384), .B(n3390), .Z(n3389) );
  XNOR U3586 ( .A(n3371), .B(n3391), .Z(n3386) );
  XNOR U3587 ( .A(n3384), .B(n3372), .Z(n3391) );
  XNOR U3588 ( .A(n3358), .B(n3357), .Z(n3372) );
  XOR U3589 ( .A(n3392), .B(n3352), .Z(n3357) );
  XNOR U3590 ( .A(n3350), .B(n3393), .Z(n3352) );
  ANDN U3591 ( .A(n1744), .B(n1921), .Z(n3393) );
  XOR U3592 ( .A(n3394), .B(n3395), .Z(n3350) );
  AND U3593 ( .A(n3396), .B(n3397), .Z(n3395) );
  XNOR U3594 ( .A(n3398), .B(n3394), .Z(n3397) );
  XOR U3595 ( .A(n3399), .B(n3354), .Z(n3392) );
  AND U3596 ( .A(n1919), .B(n1737), .Z(n3354) );
  IV U3597 ( .A(n3356), .Z(n3399) );
  XNOR U3598 ( .A(n3362), .B(n3364), .Z(n3358) );
  NAND U3599 ( .A(n2134), .B(n1542), .Z(n3364) );
  XNOR U3600 ( .A(n3360), .B(n3403), .Z(n3362) );
  ANDN U3601 ( .A(n1547), .B(n2136), .Z(n3403) );
  XOR U3602 ( .A(n3404), .B(n3405), .Z(n3360) );
  AND U3603 ( .A(n3406), .B(n3407), .Z(n3405) );
  XOR U3604 ( .A(n3408), .B(n3404), .Z(n3407) );
  XOR U3605 ( .A(n3409), .B(n3383), .Z(n3371) );
  XNOR U3606 ( .A(n3368), .B(n3369), .Z(n3383) );
  NAND U3607 ( .A(n1712), .B(n1938), .Z(n3369) );
  XNOR U3608 ( .A(n3367), .B(n3410), .Z(n3368) );
  ANDN U3609 ( .A(n1943), .B(n1714), .Z(n3410) );
  XOR U3610 ( .A(n3411), .B(n3412), .Z(n3367) );
  AND U3611 ( .A(n3413), .B(n3414), .Z(n3412) );
  XOR U3612 ( .A(n3415), .B(n3411), .Z(n3414) );
  XNOR U3613 ( .A(n3382), .B(n3370), .Z(n3409) );
  XOR U3614 ( .A(n3419), .B(n3377), .Z(n3382) );
  XNOR U3615 ( .A(n3375), .B(n3420), .Z(n3377) );
  ANDN U3616 ( .A(n2173), .B(n1522), .Z(n3420) );
  XOR U3617 ( .A(n3421), .B(n3422), .Z(n3375) );
  AND U3618 ( .A(n3423), .B(n3424), .Z(n3422) );
  XNOR U3619 ( .A(n3425), .B(n3421), .Z(n3424) );
  XOR U3620 ( .A(n3426), .B(n3379), .Z(n3419) );
  AND U3621 ( .A(n1520), .B(n2166), .Z(n3379) );
  IV U3622 ( .A(n3381), .Z(n3426) );
  XOR U3623 ( .A(n3430), .B(n3431), .Z(n3384) );
  AND U3624 ( .A(n3432), .B(n3433), .Z(n3431) );
  XOR U3625 ( .A(n3434), .B(n3435), .Z(n3433) );
  XOR U3626 ( .A(n3430), .B(n3436), .Z(n3435) );
  XNOR U3627 ( .A(n3417), .B(n3437), .Z(n3432) );
  XNOR U3628 ( .A(n3430), .B(n3418), .Z(n3437) );
  XNOR U3629 ( .A(n3402), .B(n3401), .Z(n3418) );
  XOR U3630 ( .A(n3438), .B(n3396), .Z(n3401) );
  XNOR U3631 ( .A(n3394), .B(n3439), .Z(n3396) );
  ANDN U3632 ( .A(n1744), .B(n2028), .Z(n3439) );
  XOR U3633 ( .A(n3440), .B(n3441), .Z(n3394) );
  AND U3634 ( .A(n3442), .B(n3443), .Z(n3441) );
  XNOR U3635 ( .A(n3444), .B(n3440), .Z(n3443) );
  XOR U3636 ( .A(n3445), .B(n3398), .Z(n3438) );
  AND U3637 ( .A(n2026), .B(n1737), .Z(n3398) );
  IV U3638 ( .A(n3400), .Z(n3445) );
  XNOR U3639 ( .A(n3406), .B(n3408), .Z(n3402) );
  NAND U3640 ( .A(n2253), .B(n1542), .Z(n3408) );
  XNOR U3641 ( .A(n3404), .B(n3449), .Z(n3406) );
  ANDN U3642 ( .A(n1547), .B(n2255), .Z(n3449) );
  XOR U3643 ( .A(n3450), .B(n3451), .Z(n3404) );
  AND U3644 ( .A(n3452), .B(n3453), .Z(n3451) );
  XOR U3645 ( .A(n3454), .B(n3450), .Z(n3453) );
  XOR U3646 ( .A(n3455), .B(n3429), .Z(n3417) );
  XNOR U3647 ( .A(n3413), .B(n3415), .Z(n3429) );
  NAND U3648 ( .A(n1813), .B(n1938), .Z(n3415) );
  XNOR U3649 ( .A(n3411), .B(n3456), .Z(n3413) );
  ANDN U3650 ( .A(n1943), .B(n1815), .Z(n3456) );
  XOR U3651 ( .A(n3457), .B(n3458), .Z(n3411) );
  AND U3652 ( .A(n3459), .B(n3460), .Z(n3458) );
  XOR U3653 ( .A(n3461), .B(n3457), .Z(n3460) );
  XNOR U3654 ( .A(n3428), .B(n3416), .Z(n3455) );
  XOR U3655 ( .A(n3465), .B(n3423), .Z(n3428) );
  XNOR U3656 ( .A(n3421), .B(n3466), .Z(n3423) );
  ANDN U3657 ( .A(n2173), .B(n1618), .Z(n3466) );
  XOR U3658 ( .A(n3467), .B(n3468), .Z(n3421) );
  AND U3659 ( .A(n3469), .B(n3470), .Z(n3468) );
  XNOR U3660 ( .A(n3471), .B(n3467), .Z(n3470) );
  XOR U3661 ( .A(n3472), .B(n3425), .Z(n3465) );
  AND U3662 ( .A(n1616), .B(n2166), .Z(n3425) );
  IV U3663 ( .A(n3427), .Z(n3472) );
  XOR U3664 ( .A(n3476), .B(n3477), .Z(n3430) );
  AND U3665 ( .A(n3478), .B(n3479), .Z(n3477) );
  XOR U3666 ( .A(n3480), .B(n3481), .Z(n3479) );
  XOR U3667 ( .A(n3476), .B(n3482), .Z(n3481) );
  XNOR U3668 ( .A(n3463), .B(n3483), .Z(n3478) );
  XNOR U3669 ( .A(n3476), .B(n3464), .Z(n3483) );
  XNOR U3670 ( .A(n3448), .B(n3447), .Z(n3464) );
  XOR U3671 ( .A(n3484), .B(n3442), .Z(n3447) );
  XNOR U3672 ( .A(n3440), .B(n3485), .Z(n3442) );
  ANDN U3673 ( .A(n1744), .B(n2136), .Z(n3485) );
  XOR U3674 ( .A(n3486), .B(n3487), .Z(n3440) );
  AND U3675 ( .A(n3488), .B(n3489), .Z(n3487) );
  XNOR U3676 ( .A(n3490), .B(n3486), .Z(n3489) );
  XOR U3677 ( .A(n3491), .B(n3444), .Z(n3484) );
  AND U3678 ( .A(n2134), .B(n1737), .Z(n3444) );
  IV U3679 ( .A(n3446), .Z(n3491) );
  XNOR U3680 ( .A(n3452), .B(n3454), .Z(n3448) );
  NAND U3681 ( .A(n2373), .B(n1542), .Z(n3454) );
  XNOR U3682 ( .A(n3450), .B(n3495), .Z(n3452) );
  ANDN U3683 ( .A(n1547), .B(n2375), .Z(n3495) );
  XOR U3684 ( .A(n3496), .B(n3497), .Z(n3450) );
  AND U3685 ( .A(n3498), .B(n3499), .Z(n3497) );
  XOR U3686 ( .A(n3500), .B(n3496), .Z(n3499) );
  XOR U3687 ( .A(n3501), .B(n3475), .Z(n3463) );
  XNOR U3688 ( .A(n3459), .B(n3461), .Z(n3475) );
  NAND U3689 ( .A(n1919), .B(n1938), .Z(n3461) );
  XNOR U3690 ( .A(n3457), .B(n3502), .Z(n3459) );
  ANDN U3691 ( .A(n1943), .B(n1921), .Z(n3502) );
  XOR U3692 ( .A(n3503), .B(n3504), .Z(n3457) );
  AND U3693 ( .A(n3505), .B(n3506), .Z(n3504) );
  XOR U3694 ( .A(n3507), .B(n3503), .Z(n3506) );
  XNOR U3695 ( .A(n3474), .B(n3462), .Z(n3501) );
  XOR U3696 ( .A(n3511), .B(n3469), .Z(n3474) );
  XNOR U3697 ( .A(n3467), .B(n3512), .Z(n3469) );
  ANDN U3698 ( .A(n2173), .B(n1714), .Z(n3512) );
  XOR U3699 ( .A(n3513), .B(n3514), .Z(n3467) );
  AND U3700 ( .A(n3515), .B(n3516), .Z(n3514) );
  XNOR U3701 ( .A(n3517), .B(n3513), .Z(n3516) );
  XOR U3702 ( .A(n3518), .B(n3471), .Z(n3511) );
  AND U3703 ( .A(n1712), .B(n2166), .Z(n3471) );
  IV U3704 ( .A(n3473), .Z(n3518) );
  XOR U3705 ( .A(n3522), .B(n3523), .Z(n3476) );
  AND U3706 ( .A(n3524), .B(n3525), .Z(n3523) );
  XOR U3707 ( .A(n3526), .B(n3527), .Z(n3525) );
  XOR U3708 ( .A(n3522), .B(n3528), .Z(n3527) );
  XNOR U3709 ( .A(n3509), .B(n3529), .Z(n3524) );
  XNOR U3710 ( .A(n3522), .B(n3510), .Z(n3529) );
  XNOR U3711 ( .A(n3494), .B(n3493), .Z(n3510) );
  XOR U3712 ( .A(n3530), .B(n3488), .Z(n3493) );
  XNOR U3713 ( .A(n3486), .B(n3531), .Z(n3488) );
  ANDN U3714 ( .A(n1744), .B(n2255), .Z(n3531) );
  XOR U3715 ( .A(n3532), .B(n3533), .Z(n3486) );
  AND U3716 ( .A(n3534), .B(n3535), .Z(n3533) );
  XNOR U3717 ( .A(n3536), .B(n3532), .Z(n3535) );
  XOR U3718 ( .A(n3537), .B(n3490), .Z(n3530) );
  AND U3719 ( .A(n2253), .B(n1737), .Z(n3490) );
  IV U3720 ( .A(n3492), .Z(n3537) );
  XNOR U3721 ( .A(n3498), .B(n3500), .Z(n3494) );
  NAND U3722 ( .A(n2495), .B(n1542), .Z(n3500) );
  XNOR U3723 ( .A(n3496), .B(n3541), .Z(n3498) );
  ANDN U3724 ( .A(n1547), .B(n2497), .Z(n3541) );
  XOR U3725 ( .A(n3545), .B(n3521), .Z(n3509) );
  XNOR U3726 ( .A(n3505), .B(n3507), .Z(n3521) );
  NAND U3727 ( .A(n2026), .B(n1938), .Z(n3507) );
  XNOR U3728 ( .A(n3503), .B(n3546), .Z(n3505) );
  ANDN U3729 ( .A(n1943), .B(n2028), .Z(n3546) );
  XOR U3730 ( .A(n3547), .B(n3548), .Z(n3503) );
  AND U3731 ( .A(n3549), .B(n3550), .Z(n3548) );
  XOR U3732 ( .A(n3551), .B(n3547), .Z(n3550) );
  XNOR U3733 ( .A(n3520), .B(n3508), .Z(n3545) );
  XOR U3734 ( .A(n3555), .B(n3515), .Z(n3520) );
  XNOR U3735 ( .A(n3513), .B(n3556), .Z(n3515) );
  ANDN U3736 ( .A(n2173), .B(n1815), .Z(n3556) );
  XOR U3737 ( .A(n3557), .B(n3558), .Z(n3513) );
  AND U3738 ( .A(n3559), .B(n3560), .Z(n3558) );
  XNOR U3739 ( .A(n3561), .B(n3557), .Z(n3560) );
  XOR U3740 ( .A(n3562), .B(n3517), .Z(n3555) );
  AND U3741 ( .A(n1813), .B(n2166), .Z(n3517) );
  IV U3742 ( .A(n3519), .Z(n3562) );
  XOR U3743 ( .A(n3566), .B(n3567), .Z(n3522) );
  AND U3744 ( .A(n3568), .B(n3569), .Z(n3567) );
  XOR U3745 ( .A(n3570), .B(n3571), .Z(n3569) );
  XOR U3746 ( .A(n3566), .B(n3572), .Z(n3571) );
  XNOR U3747 ( .A(n3553), .B(n3573), .Z(n3568) );
  XNOR U3748 ( .A(n3566), .B(n3554), .Z(n3573) );
  XNOR U3749 ( .A(n3540), .B(n3539), .Z(n3554) );
  XOR U3750 ( .A(n3574), .B(n3534), .Z(n3539) );
  XNOR U3751 ( .A(n3532), .B(n3575), .Z(n3534) );
  ANDN U3752 ( .A(n1744), .B(n2375), .Z(n3575) );
  XOR U3753 ( .A(n3576), .B(n3577), .Z(n3532) );
  AND U3754 ( .A(n3578), .B(n3579), .Z(n3577) );
  XNOR U3755 ( .A(n3580), .B(n3576), .Z(n3579) );
  XOR U3756 ( .A(n3581), .B(n3536), .Z(n3574) );
  AND U3757 ( .A(n2373), .B(n1737), .Z(n3536) );
  IV U3758 ( .A(n3538), .Z(n3581) );
  XNOR U3759 ( .A(n3543), .B(n3544), .Z(n3540) );
  NAND U3760 ( .A(n2620), .B(n1542), .Z(n3544) );
  XNOR U3761 ( .A(n3542), .B(n3585), .Z(n3543) );
  ANDN U3762 ( .A(n1547), .B(n2622), .Z(n3585) );
  XOR U3763 ( .A(n3586), .B(n3587), .Z(n3542) );
  AND U3764 ( .A(n3588), .B(n3589), .Z(n3587) );
  XOR U3765 ( .A(n3590), .B(n3586), .Z(n3589) );
  XOR U3766 ( .A(n3591), .B(n3565), .Z(n3553) );
  XNOR U3767 ( .A(n3549), .B(n3551), .Z(n3565) );
  NAND U3768 ( .A(n2134), .B(n1938), .Z(n3551) );
  XNOR U3769 ( .A(n3547), .B(n3592), .Z(n3549) );
  ANDN U3770 ( .A(n1943), .B(n2136), .Z(n3592) );
  XOR U3771 ( .A(n3593), .B(n3594), .Z(n3547) );
  AND U3772 ( .A(n3595), .B(n3596), .Z(n3594) );
  XOR U3773 ( .A(n3597), .B(n3593), .Z(n3596) );
  XNOR U3774 ( .A(n3564), .B(n3552), .Z(n3591) );
  XOR U3775 ( .A(n3601), .B(n3559), .Z(n3564) );
  XNOR U3776 ( .A(n3557), .B(n3602), .Z(n3559) );
  ANDN U3777 ( .A(n2173), .B(n1921), .Z(n3602) );
  XOR U3778 ( .A(n3603), .B(n3604), .Z(n3557) );
  AND U3779 ( .A(n3605), .B(n3606), .Z(n3604) );
  XNOR U3780 ( .A(n3607), .B(n3603), .Z(n3606) );
  XOR U3781 ( .A(n3608), .B(n3561), .Z(n3601) );
  AND U3782 ( .A(n1919), .B(n2166), .Z(n3561) );
  IV U3783 ( .A(n3563), .Z(n3608) );
  XOR U3784 ( .A(n3612), .B(n3613), .Z(n3566) );
  AND U3785 ( .A(n3614), .B(n3615), .Z(n3613) );
  XOR U3786 ( .A(n3616), .B(n3617), .Z(n3615) );
  XOR U3787 ( .A(n3612), .B(n3618), .Z(n3617) );
  XNOR U3788 ( .A(n3599), .B(n3619), .Z(n3614) );
  XNOR U3789 ( .A(n3612), .B(n3600), .Z(n3619) );
  XNOR U3790 ( .A(n3584), .B(n3583), .Z(n3600) );
  XOR U3791 ( .A(n3620), .B(n3578), .Z(n3583) );
  XNOR U3792 ( .A(n3576), .B(n3621), .Z(n3578) );
  ANDN U3793 ( .A(n1744), .B(n2497), .Z(n3621) );
  XOR U3794 ( .A(n3622), .B(n3623), .Z(n3576) );
  AND U3795 ( .A(n3624), .B(n3625), .Z(n3623) );
  XNOR U3796 ( .A(n3626), .B(n3622), .Z(n3625) );
  XOR U3797 ( .A(n3627), .B(n3580), .Z(n3620) );
  AND U3798 ( .A(n2495), .B(n1737), .Z(n3580) );
  IV U3799 ( .A(n3582), .Z(n3627) );
  XNOR U3800 ( .A(n3588), .B(n3590), .Z(n3584) );
  NAND U3801 ( .A(n2752), .B(n1542), .Z(n3590) );
  XNOR U3802 ( .A(n3586), .B(n3631), .Z(n3588) );
  ANDN U3803 ( .A(n1547), .B(n2754), .Z(n3631) );
  XOR U3804 ( .A(n3632), .B(n3633), .Z(n3586) );
  AND U3805 ( .A(n3634), .B(n3635), .Z(n3633) );
  XOR U3806 ( .A(n3636), .B(n3632), .Z(n3635) );
  XOR U3807 ( .A(n3637), .B(n3611), .Z(n3599) );
  XNOR U3808 ( .A(n3595), .B(n3597), .Z(n3611) );
  NAND U3809 ( .A(n2253), .B(n1938), .Z(n3597) );
  XNOR U3810 ( .A(n3593), .B(n3638), .Z(n3595) );
  ANDN U3811 ( .A(n1943), .B(n2255), .Z(n3638) );
  XOR U3812 ( .A(n3639), .B(n3640), .Z(n3593) );
  AND U3813 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U3814 ( .A(n3643), .B(n3639), .Z(n3642) );
  XNOR U3815 ( .A(n3610), .B(n3598), .Z(n3637) );
  XOR U3816 ( .A(n3647), .B(n3605), .Z(n3610) );
  XNOR U3817 ( .A(n3603), .B(n3648), .Z(n3605) );
  ANDN U3818 ( .A(n2173), .B(n2028), .Z(n3648) );
  XOR U3819 ( .A(n3649), .B(n3650), .Z(n3603) );
  AND U3820 ( .A(n3651), .B(n3652), .Z(n3650) );
  XNOR U3821 ( .A(n3653), .B(n3649), .Z(n3652) );
  XOR U3822 ( .A(n3654), .B(n3607), .Z(n3647) );
  AND U3823 ( .A(n2026), .B(n2166), .Z(n3607) );
  IV U3824 ( .A(n3609), .Z(n3654) );
  XOR U3825 ( .A(n3658), .B(n3659), .Z(n3612) );
  AND U3826 ( .A(n3660), .B(n3661), .Z(n3659) );
  XOR U3827 ( .A(n3662), .B(n3663), .Z(n3661) );
  XOR U3828 ( .A(n3658), .B(n3664), .Z(n3663) );
  XNOR U3829 ( .A(n3645), .B(n3665), .Z(n3660) );
  XNOR U3830 ( .A(n3658), .B(n3646), .Z(n3665) );
  XNOR U3831 ( .A(n3630), .B(n3629), .Z(n3646) );
  XOR U3832 ( .A(n3666), .B(n3624), .Z(n3629) );
  XNOR U3833 ( .A(n3622), .B(n3667), .Z(n3624) );
  ANDN U3834 ( .A(n1744), .B(n2622), .Z(n3667) );
  XOR U3835 ( .A(n3668), .B(n3669), .Z(n3622) );
  AND U3836 ( .A(n3670), .B(n3671), .Z(n3669) );
  XNOR U3837 ( .A(n3672), .B(n3668), .Z(n3671) );
  XOR U3838 ( .A(n3673), .B(n3626), .Z(n3666) );
  AND U3839 ( .A(n2620), .B(n1737), .Z(n3626) );
  IV U3840 ( .A(n3628), .Z(n3673) );
  XNOR U3841 ( .A(n3634), .B(n3636), .Z(n3630) );
  NAND U3842 ( .A(n2884), .B(n1542), .Z(n3636) );
  XNOR U3843 ( .A(n3632), .B(n3677), .Z(n3634) );
  ANDN U3844 ( .A(n1547), .B(n2886), .Z(n3677) );
  XOR U3845 ( .A(n3678), .B(n3679), .Z(n3632) );
  AND U3846 ( .A(n3680), .B(n3681), .Z(n3679) );
  XOR U3847 ( .A(n3682), .B(n3678), .Z(n3681) );
  XOR U3848 ( .A(n3683), .B(n3657), .Z(n3645) );
  XNOR U3849 ( .A(n3641), .B(n3643), .Z(n3657) );
  NAND U3850 ( .A(n2373), .B(n1938), .Z(n3643) );
  XNOR U3851 ( .A(n3639), .B(n3684), .Z(n3641) );
  ANDN U3852 ( .A(n1943), .B(n2375), .Z(n3684) );
  XOR U3853 ( .A(n3685), .B(n3686), .Z(n3639) );
  AND U3854 ( .A(n3687), .B(n3688), .Z(n3686) );
  XOR U3855 ( .A(n3689), .B(n3685), .Z(n3688) );
  XNOR U3856 ( .A(n3656), .B(n3644), .Z(n3683) );
  XOR U3857 ( .A(n3693), .B(n3651), .Z(n3656) );
  XNOR U3858 ( .A(n3649), .B(n3694), .Z(n3651) );
  ANDN U3859 ( .A(n2173), .B(n2136), .Z(n3694) );
  XOR U3860 ( .A(n3695), .B(n3696), .Z(n3649) );
  AND U3861 ( .A(n3697), .B(n3698), .Z(n3696) );
  XNOR U3862 ( .A(n3699), .B(n3695), .Z(n3698) );
  XOR U3863 ( .A(n3700), .B(n3653), .Z(n3693) );
  AND U3864 ( .A(n2134), .B(n2166), .Z(n3653) );
  IV U3865 ( .A(n3655), .Z(n3700) );
  XOR U3866 ( .A(n3704), .B(n3705), .Z(n3658) );
  AND U3867 ( .A(n3706), .B(n3707), .Z(n3705) );
  XOR U3868 ( .A(n3708), .B(n3709), .Z(n3707) );
  XOR U3869 ( .A(n3704), .B(n3710), .Z(n3709) );
  XNOR U3870 ( .A(n3691), .B(n3711), .Z(n3706) );
  XNOR U3871 ( .A(n3704), .B(n3692), .Z(n3711) );
  XNOR U3872 ( .A(n3676), .B(n3675), .Z(n3692) );
  XOR U3873 ( .A(n3712), .B(n3670), .Z(n3675) );
  XNOR U3874 ( .A(n3668), .B(n3713), .Z(n3670) );
  ANDN U3875 ( .A(n1744), .B(n2754), .Z(n3713) );
  XOR U3876 ( .A(n3717), .B(n3672), .Z(n3712) );
  AND U3877 ( .A(n2752), .B(n1737), .Z(n3672) );
  IV U3878 ( .A(n3674), .Z(n3717) );
  XNOR U3879 ( .A(n3680), .B(n3682), .Z(n3676) );
  NAND U3880 ( .A(n3025), .B(n1542), .Z(n3682) );
  XNOR U3881 ( .A(n3678), .B(n3721), .Z(n3680) );
  ANDN U3882 ( .A(n1547), .B(n3027), .Z(n3721) );
  XOR U3883 ( .A(n3725), .B(n3703), .Z(n3691) );
  XNOR U3884 ( .A(n3687), .B(n3689), .Z(n3703) );
  NAND U3885 ( .A(n2495), .B(n1938), .Z(n3689) );
  XNOR U3886 ( .A(n3685), .B(n3726), .Z(n3687) );
  ANDN U3887 ( .A(n1943), .B(n2497), .Z(n3726) );
  XOR U3888 ( .A(n3727), .B(n3728), .Z(n3685) );
  AND U3889 ( .A(n3729), .B(n3730), .Z(n3728) );
  XOR U3890 ( .A(n3731), .B(n3727), .Z(n3730) );
  XNOR U3891 ( .A(n3702), .B(n3690), .Z(n3725) );
  XOR U3892 ( .A(n3735), .B(n3697), .Z(n3702) );
  XNOR U3893 ( .A(n3695), .B(n3736), .Z(n3697) );
  ANDN U3894 ( .A(n2173), .B(n2255), .Z(n3736) );
  XOR U3895 ( .A(n3737), .B(n3738), .Z(n3695) );
  AND U3896 ( .A(n3739), .B(n3740), .Z(n3738) );
  XNOR U3897 ( .A(n3741), .B(n3737), .Z(n3740) );
  XOR U3898 ( .A(n3742), .B(n3699), .Z(n3735) );
  AND U3899 ( .A(n2253), .B(n2166), .Z(n3699) );
  IV U3900 ( .A(n3701), .Z(n3742) );
  XOR U3901 ( .A(n3747), .B(n3748), .Z(n3066) );
  XOR U3902 ( .A(n3749), .B(n3746), .Z(n3747) );
  XNOR U3903 ( .A(n3734), .B(n3733), .Z(n3065) );
  XOR U3904 ( .A(n3750), .B(n3745), .Z(n3733) );
  XNOR U3905 ( .A(n3729), .B(n3731), .Z(n3745) );
  NAND U3906 ( .A(n2620), .B(n1938), .Z(n3731) );
  XNOR U3907 ( .A(n3727), .B(n3751), .Z(n3729) );
  ANDN U3908 ( .A(n1943), .B(n2622), .Z(n3751) );
  XOR U3909 ( .A(n3744), .B(n3732), .Z(n3750) );
  XOR U3910 ( .A(n3755), .B(n3756), .Z(n3732) );
  XOR U3911 ( .A(n3757), .B(n3739), .Z(n3744) );
  XNOR U3912 ( .A(n3737), .B(n3758), .Z(n3739) );
  ANDN U3913 ( .A(n2173), .B(n2375), .Z(n3758) );
  AND U3914 ( .A(n2373), .B(n2166), .Z(n3741) );
  XNOR U3915 ( .A(n3762), .B(n3763), .Z(n3743) );
  AND U3916 ( .A(n3764), .B(n3765), .Z(n3763) );
  XNOR U3917 ( .A(n3760), .B(n3766), .Z(n3765) );
  XNOR U3918 ( .A(n3761), .B(n3762), .Z(n3766) );
  AND U3919 ( .A(n2495), .B(n2166), .Z(n3761) );
  XOR U3920 ( .A(n3759), .B(n3767), .Z(n3760) );
  ANDN U3921 ( .A(n2173), .B(n2497), .Z(n3767) );
  XNOR U3922 ( .A(n3753), .B(n3771), .Z(n3764) );
  XNOR U3923 ( .A(n3754), .B(n3762), .Z(n3771) );
  AND U3924 ( .A(n2752), .B(n1938), .Z(n3754) );
  XOR U3925 ( .A(n3752), .B(n3772), .Z(n3753) );
  ANDN U3926 ( .A(n1943), .B(n2754), .Z(n3772) );
  XOR U3927 ( .A(n3776), .B(n3777), .Z(n3762) );
  AND U3928 ( .A(n3778), .B(n3779), .Z(n3777) );
  XNOR U3929 ( .A(n3769), .B(n3780), .Z(n3779) );
  XNOR U3930 ( .A(n3770), .B(n3776), .Z(n3780) );
  AND U3931 ( .A(n2620), .B(n2166), .Z(n3770) );
  XOR U3932 ( .A(n3768), .B(n3781), .Z(n3769) );
  ANDN U3933 ( .A(n2173), .B(n2622), .Z(n3781) );
  XNOR U3934 ( .A(n3774), .B(n3785), .Z(n3778) );
  XNOR U3935 ( .A(n3775), .B(n3776), .Z(n3785) );
  AND U3936 ( .A(n2884), .B(n1938), .Z(n3775) );
  XOR U3937 ( .A(n3773), .B(n3786), .Z(n3774) );
  ANDN U3938 ( .A(n1943), .B(n2886), .Z(n3786) );
  XOR U3939 ( .A(n3790), .B(n3791), .Z(n3776) );
  AND U3940 ( .A(n3792), .B(n3793), .Z(n3791) );
  XNOR U3941 ( .A(n3783), .B(n3794), .Z(n3793) );
  XNOR U3942 ( .A(n3784), .B(n3790), .Z(n3794) );
  AND U3943 ( .A(n2752), .B(n2166), .Z(n3784) );
  XOR U3944 ( .A(n3782), .B(n3795), .Z(n3783) );
  ANDN U3945 ( .A(n2173), .B(n2754), .Z(n3795) );
  XNOR U3946 ( .A(n3788), .B(n3799), .Z(n3792) );
  XNOR U3947 ( .A(n3789), .B(n3790), .Z(n3799) );
  AND U3948 ( .A(n3025), .B(n1938), .Z(n3789) );
  XOR U3949 ( .A(n3787), .B(n3800), .Z(n3788) );
  ANDN U3950 ( .A(n1943), .B(n3027), .Z(n3800) );
  XNOR U3951 ( .A(n3805), .B(n3797), .Z(n3756) );
  XNOR U3952 ( .A(n3796), .B(n3806), .Z(n3797) );
  ANDN U3953 ( .A(n2173), .B(n2886), .Z(n3806) );
  XNOR U3954 ( .A(n3809), .B(n3807), .Z(n3808) );
  ANDN U3955 ( .A(n2173), .B(n3027), .Z(n3809) );
  XNOR U3956 ( .A(n3804), .B(n3798), .Z(n3805) );
  AND U3957 ( .A(n2884), .B(n2166), .Z(n3798) );
  XNOR U3958 ( .A(n3802), .B(n3803), .Z(n3755) );
  NAND U3959 ( .A(n3813), .B(n1938), .Z(n3803) );
  XNOR U3960 ( .A(n3801), .B(n3814), .Z(n3802) );
  ANDN U3961 ( .A(n1943), .B(n3815), .Z(n3814) );
  NAND U3962 ( .A(g_input[0]), .B(n3816), .Z(n3801) );
  NANDN U3963 ( .B(n1938), .A(n3817), .Z(n3816) );
  NANDN U3964 ( .B(n3818), .A(n1943), .Z(n3817) );
  IV U3965 ( .A(n1837), .Z(n1938) );
  XNOR U3966 ( .A(n3811), .B(n3812), .Z(n3804) );
  NAND U3967 ( .A(n3813), .B(n2166), .Z(n3812) );
  XNOR U3968 ( .A(n3810), .B(n3821), .Z(n3811) );
  ANDN U3969 ( .A(n2173), .B(n3815), .Z(n3821) );
  NAND U3970 ( .A(g_input[0]), .B(n3822), .Z(n3810) );
  NANDN U3971 ( .B(n2166), .A(n3823), .Z(n3822) );
  NANDN U3972 ( .B(n3818), .A(n2173), .Z(n3823) );
  IV U3973 ( .A(n2054), .Z(n2166) );
  XNOR U3974 ( .A(n3720), .B(n3719), .Z(n3734) );
  XOR U3975 ( .A(n3826), .B(n3715), .Z(n3719) );
  XNOR U3976 ( .A(n3714), .B(n3827), .Z(n3715) );
  ANDN U3977 ( .A(n1744), .B(n2886), .Z(n3827) );
  XNOR U3978 ( .A(n3830), .B(n3828), .Z(n3829) );
  ANDN U3979 ( .A(n1744), .B(n3027), .Z(n3830) );
  XNOR U3980 ( .A(n3718), .B(n3716), .Z(n3826) );
  AND U3981 ( .A(n2884), .B(n1737), .Z(n3716) );
  XNOR U3982 ( .A(n3832), .B(n3833), .Z(n3718) );
  NAND U3983 ( .A(n3813), .B(n1737), .Z(n3833) );
  XNOR U3984 ( .A(n3831), .B(n3834), .Z(n3832) );
  ANDN U3985 ( .A(n1744), .B(n3815), .Z(n3834) );
  NAND U3986 ( .A(g_input[0]), .B(n3835), .Z(n3831) );
  NANDN U3987 ( .B(n1737), .A(n3836), .Z(n3835) );
  NANDN U3988 ( .B(n3818), .A(n1744), .Z(n3836) );
  IV U3989 ( .A(n1638), .Z(n1737) );
  XNOR U3990 ( .A(n3723), .B(n3724), .Z(n3720) );
  NAND U3991 ( .A(n3813), .B(n1542), .Z(n3724) );
  XNOR U3992 ( .A(n3722), .B(n3839), .Z(n3723) );
  ANDN U3993 ( .A(n1547), .B(n3815), .Z(n3839) );
  NAND U3994 ( .A(g_input[0]), .B(n3840), .Z(n3722) );
  NANDN U3995 ( .B(n1542), .A(n3841), .Z(n3840) );
  NANDN U3996 ( .B(n3818), .A(n1547), .Z(n3841) );
  IV U3997 ( .A(n1446), .Z(n1542) );
  XNOR U3998 ( .A(n3844), .B(n3845), .Z(n3746) );
  XOR U3999 ( .A(n3846), .B(n2968), .Z(n2963) );
  XNOR U4000 ( .A(n2959), .B(n2960), .Z(n2968) );
  NAND U4001 ( .A(n2956), .B(n587), .Z(n2960) );
  XNOR U4002 ( .A(n2958), .B(n3847), .Z(n2959) );
  ANDN U4003 ( .A(n2961), .B(n589), .Z(n3847) );
  XOR U4004 ( .A(n3848), .B(n3849), .Z(n2958) );
  AND U4005 ( .A(n3850), .B(n3851), .Z(n3849) );
  XOR U4006 ( .A(n3852), .B(n3848), .Z(n3851) );
  XNOR U4007 ( .A(n2966), .B(n2962), .Z(n3846) );
  XNOR U4008 ( .A(n3077), .B(n3076), .Z(n3089) );
  XOR U4009 ( .A(n3854), .B(n3072), .Z(n3076) );
  XNOR U4010 ( .A(n3070), .B(n3855), .Z(n3072) );
  ANDN U4011 ( .A(n2682), .B(n717), .Z(n3855) );
  XOR U4012 ( .A(n3856), .B(n3857), .Z(n3070) );
  AND U4013 ( .A(n3858), .B(n3859), .Z(n3857) );
  XNOR U4014 ( .A(n3860), .B(n3856), .Z(n3859) );
  AND U4015 ( .A(n2675), .B(n715), .Z(n3074) );
  XNOR U4016 ( .A(n3081), .B(n3083), .Z(n3077) );
  NAND U4017 ( .A(n2428), .B(n816), .Z(n3083) );
  XNOR U4018 ( .A(n3079), .B(n3864), .Z(n3081) );
  ANDN U4019 ( .A(n2433), .B(n818), .Z(n3864) );
  XOR U4020 ( .A(n3865), .B(n3866), .Z(n3079) );
  AND U4021 ( .A(n3867), .B(n3868), .Z(n3866) );
  XOR U4022 ( .A(n3869), .B(n3865), .Z(n3868) );
  XOR U4023 ( .A(n3870), .B(n3871), .Z(n3090) );
  XNOR U4024 ( .A(n3872), .B(n3853), .Z(n3870) );
  XOR U4025 ( .A(n3874), .B(n3875), .Z(n3128) );
  XOR U4026 ( .A(n3876), .B(n3873), .Z(n3874) );
  XNOR U4027 ( .A(n3863), .B(n3862), .Z(n3126) );
  XOR U4028 ( .A(n3877), .B(n3858), .Z(n3862) );
  XNOR U4029 ( .A(n3856), .B(n3878), .Z(n3858) );
  ANDN U4030 ( .A(n2682), .B(n759), .Z(n3878) );
  XOR U4031 ( .A(n3879), .B(n3880), .Z(n3856) );
  AND U4032 ( .A(n3881), .B(n3882), .Z(n3880) );
  XNOR U4033 ( .A(n3883), .B(n3879), .Z(n3882) );
  XOR U4034 ( .A(n3884), .B(n3860), .Z(n3877) );
  AND U4035 ( .A(n2675), .B(n757), .Z(n3860) );
  IV U4036 ( .A(n3861), .Z(n3884) );
  XNOR U4037 ( .A(n3867), .B(n3869), .Z(n3863) );
  NAND U4038 ( .A(n2428), .B(n880), .Z(n3869) );
  XNOR U4039 ( .A(n3865), .B(n3888), .Z(n3867) );
  ANDN U4040 ( .A(n2433), .B(n882), .Z(n3888) );
  XOR U4041 ( .A(n3889), .B(n3890), .Z(n3865) );
  AND U4042 ( .A(n3891), .B(n3892), .Z(n3890) );
  XOR U4043 ( .A(n3893), .B(n3889), .Z(n3892) );
  XOR U4044 ( .A(n3895), .B(n3896), .Z(n3173) );
  XOR U4045 ( .A(n3897), .B(n3894), .Z(n3895) );
  XNOR U4046 ( .A(n3887), .B(n3886), .Z(n3171) );
  XOR U4047 ( .A(n3898), .B(n3881), .Z(n3886) );
  XNOR U4048 ( .A(n3879), .B(n3899), .Z(n3881) );
  ANDN U4049 ( .A(n2682), .B(n818), .Z(n3899) );
  XOR U4050 ( .A(n3900), .B(n3901), .Z(n3879) );
  AND U4051 ( .A(n3902), .B(n3903), .Z(n3901) );
  XNOR U4052 ( .A(n3904), .B(n3900), .Z(n3903) );
  XOR U4053 ( .A(n3905), .B(n3883), .Z(n3898) );
  AND U4054 ( .A(n2675), .B(n816), .Z(n3883) );
  IV U4055 ( .A(n3885), .Z(n3905) );
  XNOR U4056 ( .A(n3891), .B(n3893), .Z(n3887) );
  NAND U4057 ( .A(n2428), .B(n948), .Z(n3893) );
  XNOR U4058 ( .A(n3889), .B(n3909), .Z(n3891) );
  ANDN U4059 ( .A(n2433), .B(n950), .Z(n3909) );
  XOR U4060 ( .A(n3910), .B(n3911), .Z(n3889) );
  AND U4061 ( .A(n3912), .B(n3913), .Z(n3911) );
  XOR U4062 ( .A(n3914), .B(n3910), .Z(n3913) );
  XOR U4063 ( .A(n3916), .B(n3917), .Z(n3215) );
  XOR U4064 ( .A(n3918), .B(n3915), .Z(n3916) );
  XNOR U4065 ( .A(n3908), .B(n3907), .Z(n3213) );
  XOR U4066 ( .A(n3919), .B(n3902), .Z(n3907) );
  XNOR U4067 ( .A(n3900), .B(n3920), .Z(n3902) );
  ANDN U4068 ( .A(n2682), .B(n882), .Z(n3920) );
  XOR U4069 ( .A(n3921), .B(n3922), .Z(n3900) );
  AND U4070 ( .A(n3923), .B(n3924), .Z(n3922) );
  XNOR U4071 ( .A(n3925), .B(n3921), .Z(n3924) );
  AND U4072 ( .A(n2675), .B(n880), .Z(n3904) );
  XNOR U4073 ( .A(n3912), .B(n3914), .Z(n3908) );
  NAND U4074 ( .A(n2428), .B(n1015), .Z(n3914) );
  XNOR U4075 ( .A(n3910), .B(n3929), .Z(n3912) );
  ANDN U4076 ( .A(n2433), .B(n1017), .Z(n3929) );
  XOR U4077 ( .A(n3930), .B(n3931), .Z(n3910) );
  AND U4078 ( .A(n3932), .B(n3933), .Z(n3931) );
  XOR U4079 ( .A(n3934), .B(n3930), .Z(n3933) );
  XOR U4080 ( .A(n3936), .B(n3937), .Z(n3258) );
  XOR U4081 ( .A(n3938), .B(n3935), .Z(n3936) );
  XNOR U4082 ( .A(n3928), .B(n3927), .Z(n3256) );
  XOR U4083 ( .A(n3939), .B(n3923), .Z(n3927) );
  XNOR U4084 ( .A(n3921), .B(n3940), .Z(n3923) );
  ANDN U4085 ( .A(n2682), .B(n950), .Z(n3940) );
  XOR U4086 ( .A(n3941), .B(n3942), .Z(n3921) );
  AND U4087 ( .A(n3943), .B(n3944), .Z(n3942) );
  XNOR U4088 ( .A(n3945), .B(n3941), .Z(n3944) );
  XOR U4089 ( .A(n3946), .B(n3925), .Z(n3939) );
  AND U4090 ( .A(n2675), .B(n948), .Z(n3925) );
  IV U4091 ( .A(n3926), .Z(n3946) );
  XNOR U4092 ( .A(n3932), .B(n3934), .Z(n3928) );
  NAND U4093 ( .A(n2428), .B(n1089), .Z(n3934) );
  XNOR U4094 ( .A(n3930), .B(n3950), .Z(n3932) );
  ANDN U4095 ( .A(n2433), .B(n1091), .Z(n3950) );
  XOR U4096 ( .A(n3951), .B(n3952), .Z(n3930) );
  AND U4097 ( .A(n3953), .B(n3954), .Z(n3952) );
  XOR U4098 ( .A(n3955), .B(n3951), .Z(n3954) );
  XOR U4099 ( .A(n3957), .B(n3958), .Z(n3300) );
  XOR U4100 ( .A(n3959), .B(n3956), .Z(n3957) );
  XNOR U4101 ( .A(n3949), .B(n3948), .Z(n3298) );
  XOR U4102 ( .A(n3960), .B(n3943), .Z(n3948) );
  XNOR U4103 ( .A(n3941), .B(n3961), .Z(n3943) );
  ANDN U4104 ( .A(n2682), .B(n1017), .Z(n3961) );
  XOR U4105 ( .A(n3962), .B(n3963), .Z(n3941) );
  AND U4106 ( .A(n3964), .B(n3965), .Z(n3963) );
  XNOR U4107 ( .A(n3966), .B(n3962), .Z(n3965) );
  XOR U4108 ( .A(n3967), .B(n3945), .Z(n3960) );
  AND U4109 ( .A(n2675), .B(n1015), .Z(n3945) );
  IV U4110 ( .A(n3947), .Z(n3967) );
  XNOR U4111 ( .A(n3953), .B(n3955), .Z(n3949) );
  NAND U4112 ( .A(n2428), .B(n1167), .Z(n3955) );
  XNOR U4113 ( .A(n3951), .B(n3971), .Z(n3953) );
  ANDN U4114 ( .A(n2433), .B(n1169), .Z(n3971) );
  XOR U4115 ( .A(n3972), .B(n3973), .Z(n3951) );
  AND U4116 ( .A(n3974), .B(n3975), .Z(n3973) );
  XOR U4117 ( .A(n3976), .B(n3972), .Z(n3975) );
  XOR U4118 ( .A(n3978), .B(n3979), .Z(n3346) );
  XOR U4119 ( .A(n3980), .B(n3977), .Z(n3978) );
  XNOR U4120 ( .A(n3970), .B(n3969), .Z(n3344) );
  XOR U4121 ( .A(n3981), .B(n3964), .Z(n3969) );
  XNOR U4122 ( .A(n3962), .B(n3982), .Z(n3964) );
  ANDN U4123 ( .A(n2682), .B(n1091), .Z(n3982) );
  XOR U4124 ( .A(n3983), .B(n3984), .Z(n3962) );
  AND U4125 ( .A(n3985), .B(n3986), .Z(n3984) );
  XNOR U4126 ( .A(n3987), .B(n3983), .Z(n3986) );
  XOR U4127 ( .A(n3988), .B(n3966), .Z(n3981) );
  AND U4128 ( .A(n2675), .B(n1089), .Z(n3966) );
  IV U4129 ( .A(n3968), .Z(n3988) );
  XNOR U4130 ( .A(n3974), .B(n3976), .Z(n3970) );
  NAND U4131 ( .A(n2428), .B(n1248), .Z(n3976) );
  XNOR U4132 ( .A(n3972), .B(n3992), .Z(n3974) );
  ANDN U4133 ( .A(n2433), .B(n1250), .Z(n3992) );
  XOR U4134 ( .A(n3993), .B(n3994), .Z(n3972) );
  AND U4135 ( .A(n3995), .B(n3996), .Z(n3994) );
  XOR U4136 ( .A(n3997), .B(n3993), .Z(n3996) );
  XOR U4137 ( .A(n3999), .B(n4000), .Z(n3390) );
  XOR U4138 ( .A(n4001), .B(n3998), .Z(n3999) );
  XNOR U4139 ( .A(n3991), .B(n3990), .Z(n3388) );
  XOR U4140 ( .A(n4002), .B(n3985), .Z(n3990) );
  XNOR U4141 ( .A(n3983), .B(n4003), .Z(n3985) );
  ANDN U4142 ( .A(n2682), .B(n1169), .Z(n4003) );
  XOR U4143 ( .A(n4004), .B(n4005), .Z(n3983) );
  AND U4144 ( .A(n4006), .B(n4007), .Z(n4005) );
  XNOR U4145 ( .A(n4008), .B(n4004), .Z(n4007) );
  XOR U4146 ( .A(n4009), .B(n3987), .Z(n4002) );
  AND U4147 ( .A(n2675), .B(n1167), .Z(n3987) );
  IV U4148 ( .A(n3989), .Z(n4009) );
  XNOR U4149 ( .A(n3995), .B(n3997), .Z(n3991) );
  NAND U4150 ( .A(n2428), .B(n1332), .Z(n3997) );
  XNOR U4151 ( .A(n3993), .B(n4013), .Z(n3995) );
  ANDN U4152 ( .A(n2433), .B(n1334), .Z(n4013) );
  XOR U4153 ( .A(n4014), .B(n4015), .Z(n3993) );
  AND U4154 ( .A(n4016), .B(n4017), .Z(n4015) );
  XOR U4155 ( .A(n4018), .B(n4014), .Z(n4017) );
  XOR U4156 ( .A(n4020), .B(n4021), .Z(n3436) );
  XOR U4157 ( .A(n4022), .B(n4019), .Z(n4020) );
  XNOR U4158 ( .A(n4012), .B(n4011), .Z(n3434) );
  XOR U4159 ( .A(n4023), .B(n4006), .Z(n4011) );
  XNOR U4160 ( .A(n4004), .B(n4024), .Z(n4006) );
  ANDN U4161 ( .A(n2682), .B(n1250), .Z(n4024) );
  XOR U4162 ( .A(n4025), .B(n4026), .Z(n4004) );
  AND U4163 ( .A(n4027), .B(n4028), .Z(n4026) );
  XNOR U4164 ( .A(n4029), .B(n4025), .Z(n4028) );
  XOR U4165 ( .A(n4030), .B(n4008), .Z(n4023) );
  AND U4166 ( .A(n2675), .B(n1248), .Z(n4008) );
  IV U4167 ( .A(n4010), .Z(n4030) );
  XNOR U4168 ( .A(n4016), .B(n4018), .Z(n4012) );
  NAND U4169 ( .A(n2428), .B(n1423), .Z(n4018) );
  XNOR U4170 ( .A(n4014), .B(n4034), .Z(n4016) );
  ANDN U4171 ( .A(n2433), .B(n1425), .Z(n4034) );
  XOR U4172 ( .A(n4035), .B(n4036), .Z(n4014) );
  AND U4173 ( .A(n4037), .B(n4038), .Z(n4036) );
  XOR U4174 ( .A(n4039), .B(n4035), .Z(n4038) );
  XOR U4175 ( .A(n4041), .B(n4042), .Z(n3482) );
  XOR U4176 ( .A(n4043), .B(n4040), .Z(n4041) );
  XNOR U4177 ( .A(n4033), .B(n4032), .Z(n3480) );
  XOR U4178 ( .A(n4044), .B(n4027), .Z(n4032) );
  XNOR U4179 ( .A(n4025), .B(n4045), .Z(n4027) );
  ANDN U4180 ( .A(n2682), .B(n1334), .Z(n4045) );
  XOR U4181 ( .A(n4046), .B(n4047), .Z(n4025) );
  AND U4182 ( .A(n4048), .B(n4049), .Z(n4047) );
  XNOR U4183 ( .A(n4050), .B(n4046), .Z(n4049) );
  XOR U4184 ( .A(n4051), .B(n4029), .Z(n4044) );
  AND U4185 ( .A(n2675), .B(n1332), .Z(n4029) );
  IV U4186 ( .A(n4031), .Z(n4051) );
  XNOR U4187 ( .A(n4037), .B(n4039), .Z(n4033) );
  NAND U4188 ( .A(n2428), .B(n1520), .Z(n4039) );
  XNOR U4189 ( .A(n4035), .B(n4055), .Z(n4037) );
  ANDN U4190 ( .A(n2433), .B(n1522), .Z(n4055) );
  XOR U4191 ( .A(n4056), .B(n4057), .Z(n4035) );
  AND U4192 ( .A(n4058), .B(n4059), .Z(n4057) );
  XOR U4193 ( .A(n4060), .B(n4056), .Z(n4059) );
  XOR U4194 ( .A(n4062), .B(n4063), .Z(n3528) );
  XOR U4195 ( .A(n4064), .B(n4061), .Z(n4062) );
  XNOR U4196 ( .A(n4054), .B(n4053), .Z(n3526) );
  XOR U4197 ( .A(n4065), .B(n4048), .Z(n4053) );
  XNOR U4198 ( .A(n4046), .B(n4066), .Z(n4048) );
  ANDN U4199 ( .A(n2682), .B(n1425), .Z(n4066) );
  XOR U4200 ( .A(n4067), .B(n4068), .Z(n4046) );
  AND U4201 ( .A(n4069), .B(n4070), .Z(n4068) );
  XNOR U4202 ( .A(n4071), .B(n4067), .Z(n4070) );
  XOR U4203 ( .A(n4072), .B(n4050), .Z(n4065) );
  AND U4204 ( .A(n2675), .B(n1423), .Z(n4050) );
  IV U4205 ( .A(n4052), .Z(n4072) );
  XNOR U4206 ( .A(n4058), .B(n4060), .Z(n4054) );
  NAND U4207 ( .A(n2428), .B(n1616), .Z(n4060) );
  XNOR U4208 ( .A(n4056), .B(n4076), .Z(n4058) );
  ANDN U4209 ( .A(n2433), .B(n1618), .Z(n4076) );
  XOR U4210 ( .A(n4077), .B(n4078), .Z(n4056) );
  AND U4211 ( .A(n4079), .B(n4080), .Z(n4078) );
  XOR U4212 ( .A(n4081), .B(n4077), .Z(n4080) );
  XOR U4213 ( .A(n4083), .B(n4084), .Z(n3572) );
  XOR U4214 ( .A(n4085), .B(n4082), .Z(n4083) );
  XNOR U4215 ( .A(n4075), .B(n4074), .Z(n3570) );
  XOR U4216 ( .A(n4086), .B(n4069), .Z(n4074) );
  XNOR U4217 ( .A(n4067), .B(n4087), .Z(n4069) );
  ANDN U4218 ( .A(n2682), .B(n1522), .Z(n4087) );
  XOR U4219 ( .A(n4088), .B(n4089), .Z(n4067) );
  AND U4220 ( .A(n4090), .B(n4091), .Z(n4089) );
  XNOR U4221 ( .A(n4092), .B(n4088), .Z(n4091) );
  XOR U4222 ( .A(n4093), .B(n4071), .Z(n4086) );
  AND U4223 ( .A(n2675), .B(n1520), .Z(n4071) );
  IV U4224 ( .A(n4073), .Z(n4093) );
  XNOR U4225 ( .A(n4079), .B(n4081), .Z(n4075) );
  NAND U4226 ( .A(n2428), .B(n1712), .Z(n4081) );
  XNOR U4227 ( .A(n4077), .B(n4097), .Z(n4079) );
  ANDN U4228 ( .A(n2433), .B(n1714), .Z(n4097) );
  XOR U4229 ( .A(n4098), .B(n4099), .Z(n4077) );
  AND U4230 ( .A(n4100), .B(n4101), .Z(n4099) );
  XOR U4231 ( .A(n4102), .B(n4098), .Z(n4101) );
  XOR U4232 ( .A(n4104), .B(n4105), .Z(n3618) );
  XOR U4233 ( .A(n4106), .B(n4103), .Z(n4104) );
  XNOR U4234 ( .A(n4096), .B(n4095), .Z(n3616) );
  XOR U4235 ( .A(n4107), .B(n4090), .Z(n4095) );
  XNOR U4236 ( .A(n4088), .B(n4108), .Z(n4090) );
  ANDN U4237 ( .A(n2682), .B(n1618), .Z(n4108) );
  XOR U4238 ( .A(n4109), .B(n4110), .Z(n4088) );
  AND U4239 ( .A(n4111), .B(n4112), .Z(n4110) );
  XNOR U4240 ( .A(n4113), .B(n4109), .Z(n4112) );
  XOR U4241 ( .A(n4114), .B(n4092), .Z(n4107) );
  AND U4242 ( .A(n2675), .B(n1616), .Z(n4092) );
  IV U4243 ( .A(n4094), .Z(n4114) );
  XNOR U4244 ( .A(n4100), .B(n4102), .Z(n4096) );
  NAND U4245 ( .A(n2428), .B(n1813), .Z(n4102) );
  XNOR U4246 ( .A(n4098), .B(n4118), .Z(n4100) );
  ANDN U4247 ( .A(n2433), .B(n1815), .Z(n4118) );
  XOR U4248 ( .A(n4119), .B(n4120), .Z(n4098) );
  AND U4249 ( .A(n4121), .B(n4122), .Z(n4120) );
  XOR U4250 ( .A(n4123), .B(n4119), .Z(n4122) );
  XOR U4251 ( .A(n4125), .B(n4126), .Z(n3664) );
  XOR U4252 ( .A(n4127), .B(n4124), .Z(n4125) );
  XNOR U4253 ( .A(n4117), .B(n4116), .Z(n3662) );
  XOR U4254 ( .A(n4128), .B(n4111), .Z(n4116) );
  XNOR U4255 ( .A(n4109), .B(n4129), .Z(n4111) );
  ANDN U4256 ( .A(n2682), .B(n1714), .Z(n4129) );
  XOR U4257 ( .A(n4130), .B(n4131), .Z(n4109) );
  AND U4258 ( .A(n4132), .B(n4133), .Z(n4131) );
  XNOR U4259 ( .A(n4134), .B(n4130), .Z(n4133) );
  XOR U4260 ( .A(n4135), .B(n4113), .Z(n4128) );
  AND U4261 ( .A(n2675), .B(n1712), .Z(n4113) );
  IV U4262 ( .A(n4115), .Z(n4135) );
  XNOR U4263 ( .A(n4121), .B(n4123), .Z(n4117) );
  NAND U4264 ( .A(n2428), .B(n1919), .Z(n4123) );
  XNOR U4265 ( .A(n4119), .B(n4139), .Z(n4121) );
  ANDN U4266 ( .A(n2433), .B(n1921), .Z(n4139) );
  XOR U4267 ( .A(n4140), .B(n4141), .Z(n4119) );
  AND U4268 ( .A(n4142), .B(n4143), .Z(n4141) );
  XOR U4269 ( .A(n4144), .B(n4140), .Z(n4143) );
  XOR U4270 ( .A(n4146), .B(n4147), .Z(n3710) );
  XOR U4271 ( .A(n4148), .B(n4145), .Z(n4146) );
  XNOR U4272 ( .A(n4138), .B(n4137), .Z(n3708) );
  XOR U4273 ( .A(n4149), .B(n4132), .Z(n4137) );
  XNOR U4274 ( .A(n4130), .B(n4150), .Z(n4132) );
  ANDN U4275 ( .A(n2682), .B(n1815), .Z(n4150) );
  XOR U4276 ( .A(n4151), .B(n4152), .Z(n4130) );
  AND U4277 ( .A(n4153), .B(n4154), .Z(n4152) );
  XNOR U4278 ( .A(n4155), .B(n4151), .Z(n4154) );
  XOR U4279 ( .A(n4156), .B(n4134), .Z(n4149) );
  AND U4280 ( .A(n2675), .B(n1813), .Z(n4134) );
  IV U4281 ( .A(n4136), .Z(n4156) );
  XNOR U4282 ( .A(n4142), .B(n4144), .Z(n4138) );
  NAND U4283 ( .A(n2428), .B(n2026), .Z(n4144) );
  XNOR U4284 ( .A(n4140), .B(n4160), .Z(n4142) );
  ANDN U4285 ( .A(n2433), .B(n2028), .Z(n4160) );
  XOR U4286 ( .A(n4161), .B(n4162), .Z(n4140) );
  AND U4287 ( .A(n4163), .B(n4164), .Z(n4162) );
  XOR U4288 ( .A(n4165), .B(n4161), .Z(n4164) );
  XOR U4289 ( .A(n4167), .B(n4168), .Z(n3749) );
  XOR U4290 ( .A(n4169), .B(n4166), .Z(n4167) );
  XNOR U4291 ( .A(n4159), .B(n4158), .Z(n3748) );
  XOR U4292 ( .A(n4170), .B(n4153), .Z(n4158) );
  XNOR U4293 ( .A(n4151), .B(n4171), .Z(n4153) );
  ANDN U4294 ( .A(n2682), .B(n1921), .Z(n4171) );
  AND U4295 ( .A(n2675), .B(n1919), .Z(n4155) );
  XNOR U4296 ( .A(n4163), .B(n4165), .Z(n4159) );
  NAND U4297 ( .A(n2428), .B(n2134), .Z(n4165) );
  XNOR U4298 ( .A(n4161), .B(n4178), .Z(n4163) );
  ANDN U4299 ( .A(n2433), .B(n2136), .Z(n4178) );
  XOR U4300 ( .A(n4182), .B(n4183), .Z(n4166) );
  AND U4301 ( .A(n4184), .B(n4185), .Z(n4183) );
  XOR U4302 ( .A(n4186), .B(n4187), .Z(n4185) );
  XNOR U4303 ( .A(n4182), .B(n4188), .Z(n4187) );
  XNOR U4304 ( .A(n4176), .B(n4189), .Z(n4184) );
  XNOR U4305 ( .A(n4182), .B(n4177), .Z(n4189) );
  XNOR U4306 ( .A(n4180), .B(n4181), .Z(n4177) );
  NAND U4307 ( .A(n2253), .B(n2428), .Z(n4181) );
  XNOR U4308 ( .A(n4179), .B(n4190), .Z(n4180) );
  ANDN U4309 ( .A(n2433), .B(n2255), .Z(n4190) );
  XOR U4310 ( .A(n4194), .B(n4173), .Z(n4176) );
  XNOR U4311 ( .A(n4172), .B(n4195), .Z(n4173) );
  ANDN U4312 ( .A(n2682), .B(n2028), .Z(n4195) );
  AND U4313 ( .A(n2675), .B(n2026), .Z(n4174) );
  XOR U4314 ( .A(n4202), .B(n4203), .Z(n4182) );
  AND U4315 ( .A(n4204), .B(n4205), .Z(n4203) );
  XOR U4316 ( .A(n4206), .B(n4207), .Z(n4205) );
  XNOR U4317 ( .A(n4202), .B(n4208), .Z(n4207) );
  XNOR U4318 ( .A(n4200), .B(n4209), .Z(n4204) );
  XNOR U4319 ( .A(n4202), .B(n4201), .Z(n4209) );
  XNOR U4320 ( .A(n4192), .B(n4193), .Z(n4201) );
  NAND U4321 ( .A(n2373), .B(n2428), .Z(n4193) );
  XNOR U4322 ( .A(n4191), .B(n4210), .Z(n4192) );
  ANDN U4323 ( .A(n2433), .B(n2375), .Z(n4210) );
  XOR U4324 ( .A(n4214), .B(n4197), .Z(n4200) );
  XNOR U4325 ( .A(n4196), .B(n4215), .Z(n4197) );
  ANDN U4326 ( .A(n2682), .B(n2136), .Z(n4215) );
  AND U4327 ( .A(n2675), .B(n2134), .Z(n4198) );
  XOR U4328 ( .A(n4222), .B(n4223), .Z(n4202) );
  AND U4329 ( .A(n4224), .B(n4225), .Z(n4223) );
  XOR U4330 ( .A(n4226), .B(n4227), .Z(n4225) );
  XNOR U4331 ( .A(n4222), .B(n4228), .Z(n4227) );
  XNOR U4332 ( .A(n4220), .B(n4229), .Z(n4224) );
  XNOR U4333 ( .A(n4222), .B(n4221), .Z(n4229) );
  XNOR U4334 ( .A(n4212), .B(n4213), .Z(n4221) );
  NAND U4335 ( .A(n2495), .B(n2428), .Z(n4213) );
  XNOR U4336 ( .A(n4211), .B(n4230), .Z(n4212) );
  ANDN U4337 ( .A(n2433), .B(n2497), .Z(n4230) );
  XOR U4338 ( .A(n4234), .B(n4217), .Z(n4220) );
  XNOR U4339 ( .A(n4216), .B(n4235), .Z(n4217) );
  ANDN U4340 ( .A(n2682), .B(n2255), .Z(n4235) );
  AND U4341 ( .A(n2253), .B(n2675), .Z(n4218) );
  XOR U4342 ( .A(n4242), .B(n4243), .Z(n4222) );
  AND U4343 ( .A(n4244), .B(n4245), .Z(n4243) );
  XOR U4344 ( .A(n4246), .B(n4247), .Z(n4245) );
  XNOR U4345 ( .A(n4242), .B(n4248), .Z(n4247) );
  XNOR U4346 ( .A(n4240), .B(n4249), .Z(n4244) );
  XNOR U4347 ( .A(n4242), .B(n4241), .Z(n4249) );
  XNOR U4348 ( .A(n4232), .B(n4233), .Z(n4241) );
  NAND U4349 ( .A(n2620), .B(n2428), .Z(n4233) );
  XNOR U4350 ( .A(n4231), .B(n4250), .Z(n4232) );
  ANDN U4351 ( .A(n2433), .B(n2622), .Z(n4250) );
  XOR U4352 ( .A(n4254), .B(n4237), .Z(n4240) );
  XNOR U4353 ( .A(n4236), .B(n4255), .Z(n4237) );
  ANDN U4354 ( .A(n2682), .B(n2375), .Z(n4255) );
  AND U4355 ( .A(n2373), .B(n2675), .Z(n4238) );
  XOR U4356 ( .A(n4262), .B(n4263), .Z(n4242) );
  AND U4357 ( .A(n4264), .B(n4265), .Z(n4263) );
  XOR U4358 ( .A(n4266), .B(n4267), .Z(n4265) );
  XNOR U4359 ( .A(n4262), .B(n4268), .Z(n4267) );
  XNOR U4360 ( .A(n4260), .B(n4269), .Z(n4264) );
  XNOR U4361 ( .A(n4262), .B(n4261), .Z(n4269) );
  XNOR U4362 ( .A(n4252), .B(n4253), .Z(n4261) );
  NAND U4363 ( .A(n2752), .B(n2428), .Z(n4253) );
  XNOR U4364 ( .A(n4251), .B(n4270), .Z(n4252) );
  ANDN U4365 ( .A(n2433), .B(n2754), .Z(n4270) );
  XOR U4366 ( .A(n4274), .B(n4257), .Z(n4260) );
  XNOR U4367 ( .A(n4256), .B(n4275), .Z(n4257) );
  ANDN U4368 ( .A(n2682), .B(n2497), .Z(n4275) );
  AND U4369 ( .A(n2495), .B(n2675), .Z(n4258) );
  XOR U4370 ( .A(n4282), .B(n4283), .Z(n4262) );
  AND U4371 ( .A(n4284), .B(n4285), .Z(n4283) );
  XOR U4372 ( .A(n4286), .B(n4287), .Z(n4285) );
  XNOR U4373 ( .A(n4282), .B(n4288), .Z(n4287) );
  XNOR U4374 ( .A(n4280), .B(n4289), .Z(n4284) );
  XNOR U4375 ( .A(n4282), .B(n4281), .Z(n4289) );
  XNOR U4376 ( .A(n4272), .B(n4273), .Z(n4281) );
  NAND U4377 ( .A(n2884), .B(n2428), .Z(n4273) );
  XNOR U4378 ( .A(n4271), .B(n4290), .Z(n4272) );
  ANDN U4379 ( .A(n2433), .B(n2886), .Z(n4290) );
  XOR U4380 ( .A(n4291), .B(n4292), .Z(n4271) );
  AND U4381 ( .A(n4293), .B(n4294), .Z(n4292) );
  XOR U4382 ( .A(n4295), .B(n4291), .Z(n4294) );
  XOR U4383 ( .A(n4296), .B(n4277), .Z(n4280) );
  XNOR U4384 ( .A(n4276), .B(n4297), .Z(n4277) );
  ANDN U4385 ( .A(n2682), .B(n2622), .Z(n4297) );
  XOR U4386 ( .A(n4298), .B(n4299), .Z(n4276) );
  AND U4387 ( .A(n4300), .B(n4301), .Z(n4299) );
  XNOR U4388 ( .A(n4302), .B(n4298), .Z(n4301) );
  AND U4389 ( .A(n2620), .B(n2675), .Z(n4278) );
  XOR U4390 ( .A(n4306), .B(n4307), .Z(n4282) );
  AND U4391 ( .A(n4308), .B(n4309), .Z(n4307) );
  XOR U4392 ( .A(n4310), .B(n4311), .Z(n4309) );
  XNOR U4393 ( .A(n4306), .B(n4312), .Z(n4311) );
  XNOR U4394 ( .A(n4304), .B(n4313), .Z(n4308) );
  XNOR U4395 ( .A(n4306), .B(n4305), .Z(n4313) );
  XNOR U4396 ( .A(n4293), .B(n4295), .Z(n4305) );
  NAND U4397 ( .A(n3025), .B(n2428), .Z(n4295) );
  XNOR U4398 ( .A(n4291), .B(n4314), .Z(n4293) );
  ANDN U4399 ( .A(n2433), .B(n3027), .Z(n4314) );
  XOR U4400 ( .A(n4318), .B(n4300), .Z(n4304) );
  XNOR U4401 ( .A(n4298), .B(n4319), .Z(n4300) );
  ANDN U4402 ( .A(n2682), .B(n2754), .Z(n4319) );
  XOR U4403 ( .A(n4320), .B(n4321), .Z(n4298) );
  AND U4404 ( .A(n4322), .B(n4323), .Z(n4321) );
  XNOR U4405 ( .A(n4324), .B(n4320), .Z(n4323) );
  AND U4406 ( .A(n2752), .B(n2675), .Z(n4302) );
  XOR U4407 ( .A(n4329), .B(n4330), .Z(n3845) );
  XNOR U4408 ( .A(n4327), .B(n4326), .Z(n3844) );
  XOR U4409 ( .A(n4332), .B(n4322), .Z(n4326) );
  XNOR U4410 ( .A(n4320), .B(n4333), .Z(n4322) );
  ANDN U4411 ( .A(n2682), .B(n2886), .Z(n4333) );
  XNOR U4412 ( .A(n4336), .B(n4334), .Z(n4335) );
  ANDN U4413 ( .A(n2682), .B(n3027), .Z(n4336) );
  XNOR U4414 ( .A(n4325), .B(n4324), .Z(n4332) );
  AND U4415 ( .A(n2884), .B(n2675), .Z(n4324) );
  XNOR U4416 ( .A(n4338), .B(n4339), .Z(n4325) );
  NAND U4417 ( .A(n3813), .B(n2675), .Z(n4339) );
  XNOR U4418 ( .A(n4337), .B(n4340), .Z(n4338) );
  ANDN U4419 ( .A(n2682), .B(n3815), .Z(n4340) );
  NAND U4420 ( .A(g_input[0]), .B(n4341), .Z(n4337) );
  NANDN U4421 ( .B(n2675), .A(n4342), .Z(n4341) );
  NANDN U4422 ( .B(n3818), .A(n2682), .Z(n4342) );
  IV U4423 ( .A(n2549), .Z(n2675) );
  XNOR U4424 ( .A(n4316), .B(n4317), .Z(n4327) );
  NAND U4425 ( .A(n3813), .B(n2428), .Z(n4317) );
  XNOR U4426 ( .A(n4315), .B(n4345), .Z(n4316) );
  ANDN U4427 ( .A(n2433), .B(n3815), .Z(n4345) );
  NAND U4428 ( .A(g_input[0]), .B(n4346), .Z(n4315) );
  NANDN U4429 ( .B(n2428), .A(n4347), .Z(n4346) );
  NANDN U4430 ( .B(n3818), .A(n2433), .Z(n4347) );
  IV U4431 ( .A(n2307), .Z(n2428) );
  XOR U4432 ( .A(n4350), .B(n4351), .Z(n4328) );
  XOR U4433 ( .A(n2965), .B(n4352), .Z(n2966) );
  AND U4434 ( .A(n4353), .B(n4354), .Z(n4352) );
  NANDN U4435 ( .B(n4355), .A(n526), .Z(n4354) );
  NANDN U4436 ( .B(n4356), .A(n4357), .Z(n4353) );
  XNOR U4437 ( .A(n3850), .B(n3852), .Z(n3871) );
  NAND U4438 ( .A(n2956), .B(n631), .Z(n3852) );
  XNOR U4439 ( .A(n3848), .B(n4359), .Z(n3850) );
  ANDN U4440 ( .A(n2961), .B(n633), .Z(n4359) );
  XOR U4441 ( .A(n4360), .B(n4361), .Z(n3848) );
  AND U4442 ( .A(n4362), .B(n4363), .Z(n4361) );
  XOR U4443 ( .A(n4364), .B(n4360), .Z(n4363) );
  XNOR U4444 ( .A(n4365), .B(n4366), .Z(n3872) );
  IV U4445 ( .A(n4358), .Z(n4366) );
  XOR U4446 ( .A(n4367), .B(n4357), .Z(n4365) );
  AND U4447 ( .A(n4368), .B(n556), .Z(n4357) );
  IV U4448 ( .A(n589), .Z(n556) );
  NAND U4449 ( .A(n4369), .B(n4356), .Z(n4367) );
  XOR U4450 ( .A(n4370), .B(n4371), .Z(n4356) );
  AND U4451 ( .A(n4372), .B(n4373), .Z(n4371) );
  XNOR U4452 ( .A(n4374), .B(n4370), .Z(n4373) );
  NANDN U4453 ( .B(n559), .A(e_input[0]), .Z(n4369) );
  IV U4454 ( .A(n526), .Z(n559) );
  AND U4455 ( .A(n4375), .B(n4376), .Z(n526) );
  ANDN U4456 ( .A(g_input[31]), .B(n4377), .Z(n4375) );
  XNOR U4457 ( .A(n4362), .B(n4364), .Z(n3875) );
  NAND U4458 ( .A(n2956), .B(n671), .Z(n4364) );
  XNOR U4459 ( .A(n4360), .B(n4379), .Z(n4362) );
  ANDN U4460 ( .A(n2961), .B(n673), .Z(n4379) );
  XOR U4461 ( .A(n4380), .B(n4381), .Z(n4360) );
  AND U4462 ( .A(n4382), .B(n4383), .Z(n4381) );
  XOR U4463 ( .A(n4384), .B(n4380), .Z(n4383) );
  XNOR U4464 ( .A(n4385), .B(n4372), .Z(n3876) );
  XNOR U4465 ( .A(n4370), .B(n4386), .Z(n4372) );
  ANDN U4466 ( .A(e_input[0]), .B(n589), .Z(n4386) );
  XNOR U4467 ( .A(n4377), .B(g_input[30]), .Z(n4376) );
  NANDN U4468 ( .B(n4387), .A(n4388), .Z(n4377) );
  XOR U4469 ( .A(n4389), .B(n4390), .Z(n4370) );
  AND U4470 ( .A(n4391), .B(n4392), .Z(n4390) );
  XNOR U4471 ( .A(n4393), .B(n4389), .Z(n4392) );
  XOR U4472 ( .A(n4394), .B(n4374), .Z(n4385) );
  AND U4473 ( .A(n4368), .B(n587), .Z(n4374) );
  IV U4474 ( .A(n633), .Z(n587) );
  IV U4475 ( .A(n4378), .Z(n4394) );
  XNOR U4476 ( .A(n4382), .B(n4384), .Z(n3896) );
  NAND U4477 ( .A(n2956), .B(n715), .Z(n4384) );
  XNOR U4478 ( .A(n4380), .B(n4396), .Z(n4382) );
  ANDN U4479 ( .A(n2961), .B(n717), .Z(n4396) );
  XOR U4480 ( .A(n4397), .B(n4398), .Z(n4380) );
  AND U4481 ( .A(n4399), .B(n4400), .Z(n4398) );
  XOR U4482 ( .A(n4401), .B(n4397), .Z(n4400) );
  XNOR U4483 ( .A(n4402), .B(n4391), .Z(n3897) );
  XNOR U4484 ( .A(n4389), .B(n4403), .Z(n4391) );
  ANDN U4485 ( .A(e_input[0]), .B(n633), .Z(n4403) );
  XNOR U4486 ( .A(n4388), .B(g_input[29]), .Z(n4387) );
  ANDN U4487 ( .A(n4404), .B(n4405), .Z(n4388) );
  XOR U4488 ( .A(n4406), .B(n4407), .Z(n4389) );
  AND U4489 ( .A(n4408), .B(n4409), .Z(n4407) );
  XNOR U4490 ( .A(n4410), .B(n4406), .Z(n4409) );
  XOR U4491 ( .A(n4411), .B(n4393), .Z(n4402) );
  AND U4492 ( .A(n4368), .B(n631), .Z(n4393) );
  IV U4493 ( .A(n673), .Z(n631) );
  IV U4494 ( .A(n4395), .Z(n4411) );
  XNOR U4495 ( .A(n4399), .B(n4401), .Z(n3917) );
  NAND U4496 ( .A(n2956), .B(n757), .Z(n4401) );
  XNOR U4497 ( .A(n4397), .B(n4413), .Z(n4399) );
  ANDN U4498 ( .A(n2961), .B(n759), .Z(n4413) );
  XOR U4499 ( .A(n4414), .B(n4415), .Z(n4397) );
  AND U4500 ( .A(n4416), .B(n4417), .Z(n4415) );
  XOR U4501 ( .A(n4418), .B(n4414), .Z(n4417) );
  XNOR U4502 ( .A(n4419), .B(n4408), .Z(n3918) );
  XNOR U4503 ( .A(n4406), .B(n4420), .Z(n4408) );
  ANDN U4504 ( .A(e_input[0]), .B(n673), .Z(n4420) );
  XNOR U4505 ( .A(n4404), .B(g_input[28]), .Z(n4405) );
  ANDN U4506 ( .A(n4421), .B(n4422), .Z(n4404) );
  XOR U4507 ( .A(n4423), .B(n4424), .Z(n4406) );
  AND U4508 ( .A(n4425), .B(n4426), .Z(n4424) );
  XNOR U4509 ( .A(n4427), .B(n4423), .Z(n4426) );
  AND U4510 ( .A(n4368), .B(n671), .Z(n4410) );
  IV U4511 ( .A(n717), .Z(n671) );
  XNOR U4512 ( .A(n4416), .B(n4418), .Z(n3937) );
  NAND U4513 ( .A(n2956), .B(n816), .Z(n4418) );
  XNOR U4514 ( .A(n4414), .B(n4429), .Z(n4416) );
  ANDN U4515 ( .A(n2961), .B(n818), .Z(n4429) );
  XOR U4516 ( .A(n4430), .B(n4431), .Z(n4414) );
  AND U4517 ( .A(n4432), .B(n4433), .Z(n4431) );
  XOR U4518 ( .A(n4434), .B(n4430), .Z(n4433) );
  XNOR U4519 ( .A(n4435), .B(n4425), .Z(n3938) );
  XNOR U4520 ( .A(n4423), .B(n4436), .Z(n4425) );
  ANDN U4521 ( .A(e_input[0]), .B(n717), .Z(n4436) );
  ANDN U4522 ( .A(n4437), .B(n4438), .Z(n4421) );
  XOR U4523 ( .A(n4439), .B(n4440), .Z(n4423) );
  AND U4524 ( .A(n4441), .B(n4442), .Z(n4440) );
  XNOR U4525 ( .A(n4443), .B(n4439), .Z(n4442) );
  AND U4526 ( .A(n4368), .B(n715), .Z(n4427) );
  IV U4527 ( .A(n759), .Z(n715) );
  XNOR U4528 ( .A(n4432), .B(n4434), .Z(n3958) );
  NAND U4529 ( .A(n2956), .B(n880), .Z(n4434) );
  XNOR U4530 ( .A(n4430), .B(n4445), .Z(n4432) );
  ANDN U4531 ( .A(n2961), .B(n882), .Z(n4445) );
  XOR U4532 ( .A(n4446), .B(n4447), .Z(n4430) );
  AND U4533 ( .A(n4448), .B(n4449), .Z(n4447) );
  XOR U4534 ( .A(n4450), .B(n4446), .Z(n4449) );
  XNOR U4535 ( .A(n4451), .B(n4441), .Z(n3959) );
  XNOR U4536 ( .A(n4439), .B(n4452), .Z(n4441) );
  ANDN U4537 ( .A(e_input[0]), .B(n759), .Z(n4452) );
  XNOR U4538 ( .A(n4437), .B(g_input[26]), .Z(n4438) );
  ANDN U4539 ( .A(n4453), .B(n4454), .Z(n4437) );
  XOR U4540 ( .A(n4455), .B(n4456), .Z(n4439) );
  AND U4541 ( .A(n4457), .B(n4458), .Z(n4456) );
  XNOR U4542 ( .A(n4459), .B(n4455), .Z(n4458) );
  XOR U4543 ( .A(n4460), .B(n4443), .Z(n4451) );
  AND U4544 ( .A(n4368), .B(n757), .Z(n4443) );
  IV U4545 ( .A(n818), .Z(n757) );
  IV U4546 ( .A(n4444), .Z(n4460) );
  XNOR U4547 ( .A(n4448), .B(n4450), .Z(n3979) );
  NAND U4548 ( .A(n2956), .B(n948), .Z(n4450) );
  XNOR U4549 ( .A(n4446), .B(n4462), .Z(n4448) );
  ANDN U4550 ( .A(n2961), .B(n950), .Z(n4462) );
  XOR U4551 ( .A(n4463), .B(n4464), .Z(n4446) );
  AND U4552 ( .A(n4465), .B(n4466), .Z(n4464) );
  XOR U4553 ( .A(n4467), .B(n4463), .Z(n4466) );
  XNOR U4554 ( .A(n4468), .B(n4457), .Z(n3980) );
  XNOR U4555 ( .A(n4455), .B(n4469), .Z(n4457) );
  ANDN U4556 ( .A(e_input[0]), .B(n818), .Z(n4469) );
  ANDN U4557 ( .A(n4470), .B(n4471), .Z(n4453) );
  XOR U4558 ( .A(n4472), .B(n4473), .Z(n4455) );
  AND U4559 ( .A(n4474), .B(n4475), .Z(n4473) );
  XNOR U4560 ( .A(n4476), .B(n4472), .Z(n4475) );
  XOR U4561 ( .A(n4477), .B(n4459), .Z(n4468) );
  AND U4562 ( .A(n4368), .B(n816), .Z(n4459) );
  IV U4563 ( .A(n882), .Z(n816) );
  IV U4564 ( .A(n4461), .Z(n4477) );
  XNOR U4565 ( .A(n4465), .B(n4467), .Z(n4000) );
  NAND U4566 ( .A(n2956), .B(n1015), .Z(n4467) );
  XNOR U4567 ( .A(n4463), .B(n4479), .Z(n4465) );
  ANDN U4568 ( .A(n2961), .B(n1017), .Z(n4479) );
  XOR U4569 ( .A(n4480), .B(n4481), .Z(n4463) );
  AND U4570 ( .A(n4482), .B(n4483), .Z(n4481) );
  XOR U4571 ( .A(n4484), .B(n4480), .Z(n4483) );
  XNOR U4572 ( .A(n4485), .B(n4474), .Z(n4001) );
  XNOR U4573 ( .A(n4472), .B(n4486), .Z(n4474) );
  ANDN U4574 ( .A(e_input[0]), .B(n882), .Z(n4486) );
  XNOR U4575 ( .A(n4470), .B(g_input[24]), .Z(n4471) );
  ANDN U4576 ( .A(n4487), .B(n4488), .Z(n4470) );
  XOR U4577 ( .A(n4489), .B(n4490), .Z(n4472) );
  AND U4578 ( .A(n4491), .B(n4492), .Z(n4490) );
  XNOR U4579 ( .A(n4493), .B(n4489), .Z(n4492) );
  XOR U4580 ( .A(n4494), .B(n4476), .Z(n4485) );
  AND U4581 ( .A(n4368), .B(n880), .Z(n4476) );
  IV U4582 ( .A(n950), .Z(n880) );
  IV U4583 ( .A(n4478), .Z(n4494) );
  XNOR U4584 ( .A(n4482), .B(n4484), .Z(n4021) );
  NAND U4585 ( .A(n2956), .B(n1089), .Z(n4484) );
  XNOR U4586 ( .A(n4480), .B(n4496), .Z(n4482) );
  ANDN U4587 ( .A(n2961), .B(n1091), .Z(n4496) );
  XOR U4588 ( .A(n4497), .B(n4498), .Z(n4480) );
  AND U4589 ( .A(n4499), .B(n4500), .Z(n4498) );
  XOR U4590 ( .A(n4501), .B(n4497), .Z(n4500) );
  XNOR U4591 ( .A(n4502), .B(n4491), .Z(n4022) );
  XNOR U4592 ( .A(n4489), .B(n4503), .Z(n4491) );
  ANDN U4593 ( .A(e_input[0]), .B(n950), .Z(n4503) );
  ANDN U4594 ( .A(n4504), .B(n4505), .Z(n4487) );
  XOR U4595 ( .A(n4506), .B(n4507), .Z(n4489) );
  AND U4596 ( .A(n4508), .B(n4509), .Z(n4507) );
  XNOR U4597 ( .A(n4510), .B(n4506), .Z(n4509) );
  XOR U4598 ( .A(n4511), .B(n4493), .Z(n4502) );
  AND U4599 ( .A(n4368), .B(n948), .Z(n4493) );
  IV U4600 ( .A(n1017), .Z(n948) );
  IV U4601 ( .A(n4495), .Z(n4511) );
  XNOR U4602 ( .A(n4499), .B(n4501), .Z(n4042) );
  NAND U4603 ( .A(n2956), .B(n1167), .Z(n4501) );
  XNOR U4604 ( .A(n4497), .B(n4513), .Z(n4499) );
  ANDN U4605 ( .A(n2961), .B(n1169), .Z(n4513) );
  XOR U4606 ( .A(n4514), .B(n4515), .Z(n4497) );
  AND U4607 ( .A(n4516), .B(n4517), .Z(n4515) );
  XOR U4608 ( .A(n4518), .B(n4514), .Z(n4517) );
  XNOR U4609 ( .A(n4519), .B(n4508), .Z(n4043) );
  XNOR U4610 ( .A(n4506), .B(n4520), .Z(n4508) );
  ANDN U4611 ( .A(e_input[0]), .B(n1017), .Z(n4520) );
  XNOR U4612 ( .A(n4504), .B(g_input[22]), .Z(n4505) );
  ANDN U4613 ( .A(n4521), .B(n4522), .Z(n4504) );
  XOR U4614 ( .A(n4523), .B(n4524), .Z(n4506) );
  AND U4615 ( .A(n4525), .B(n4526), .Z(n4524) );
  XNOR U4616 ( .A(n4527), .B(n4523), .Z(n4526) );
  XOR U4617 ( .A(n4528), .B(n4510), .Z(n4519) );
  AND U4618 ( .A(n4368), .B(n1015), .Z(n4510) );
  IV U4619 ( .A(n1091), .Z(n1015) );
  IV U4620 ( .A(n4512), .Z(n4528) );
  XNOR U4621 ( .A(n4516), .B(n4518), .Z(n4063) );
  NAND U4622 ( .A(n2956), .B(n1248), .Z(n4518) );
  XNOR U4623 ( .A(n4514), .B(n4530), .Z(n4516) );
  ANDN U4624 ( .A(n2961), .B(n1250), .Z(n4530) );
  XOR U4625 ( .A(n4531), .B(n4532), .Z(n4514) );
  AND U4626 ( .A(n4533), .B(n4534), .Z(n4532) );
  XOR U4627 ( .A(n4535), .B(n4531), .Z(n4534) );
  XNOR U4628 ( .A(n4536), .B(n4525), .Z(n4064) );
  XNOR U4629 ( .A(n4523), .B(n4537), .Z(n4525) );
  ANDN U4630 ( .A(e_input[0]), .B(n1091), .Z(n4537) );
  ANDN U4631 ( .A(n4538), .B(n4539), .Z(n4521) );
  XOR U4632 ( .A(n4540), .B(n4541), .Z(n4523) );
  AND U4633 ( .A(n4542), .B(n4543), .Z(n4541) );
  XNOR U4634 ( .A(n4544), .B(n4540), .Z(n4543) );
  XOR U4635 ( .A(n4545), .B(n4527), .Z(n4536) );
  AND U4636 ( .A(n4368), .B(n1089), .Z(n4527) );
  IV U4637 ( .A(n1169), .Z(n1089) );
  IV U4638 ( .A(n4529), .Z(n4545) );
  XNOR U4639 ( .A(n4533), .B(n4535), .Z(n4084) );
  NAND U4640 ( .A(n2956), .B(n1332), .Z(n4535) );
  XNOR U4641 ( .A(n4531), .B(n4547), .Z(n4533) );
  ANDN U4642 ( .A(n2961), .B(n1334), .Z(n4547) );
  XOR U4643 ( .A(n4548), .B(n4549), .Z(n4531) );
  AND U4644 ( .A(n4550), .B(n4551), .Z(n4549) );
  XOR U4645 ( .A(n4552), .B(n4548), .Z(n4551) );
  XNOR U4646 ( .A(n4553), .B(n4542), .Z(n4085) );
  XNOR U4647 ( .A(n4540), .B(n4554), .Z(n4542) );
  ANDN U4648 ( .A(e_input[0]), .B(n1169), .Z(n4554) );
  XNOR U4649 ( .A(n4538), .B(g_input[20]), .Z(n4539) );
  ANDN U4650 ( .A(n4555), .B(n4556), .Z(n4538) );
  XOR U4651 ( .A(n4557), .B(n4558), .Z(n4540) );
  AND U4652 ( .A(n4559), .B(n4560), .Z(n4558) );
  XNOR U4653 ( .A(n4561), .B(n4557), .Z(n4560) );
  XOR U4654 ( .A(n4562), .B(n4544), .Z(n4553) );
  AND U4655 ( .A(n4368), .B(n1167), .Z(n4544) );
  IV U4656 ( .A(n1250), .Z(n1167) );
  IV U4657 ( .A(n4546), .Z(n4562) );
  XNOR U4658 ( .A(n4550), .B(n4552), .Z(n4105) );
  NAND U4659 ( .A(n2956), .B(n1423), .Z(n4552) );
  XNOR U4660 ( .A(n4548), .B(n4564), .Z(n4550) );
  ANDN U4661 ( .A(n2961), .B(n1425), .Z(n4564) );
  XOR U4662 ( .A(n4565), .B(n4566), .Z(n4548) );
  AND U4663 ( .A(n4567), .B(n4568), .Z(n4566) );
  XOR U4664 ( .A(n4569), .B(n4565), .Z(n4568) );
  XNOR U4665 ( .A(n4570), .B(n4559), .Z(n4106) );
  XNOR U4666 ( .A(n4557), .B(n4571), .Z(n4559) );
  ANDN U4667 ( .A(e_input[0]), .B(n1250), .Z(n4571) );
  ANDN U4668 ( .A(n4572), .B(n4573), .Z(n4555) );
  XOR U4669 ( .A(n4574), .B(n4575), .Z(n4557) );
  AND U4670 ( .A(n4576), .B(n4577), .Z(n4575) );
  XNOR U4671 ( .A(n4578), .B(n4574), .Z(n4577) );
  XOR U4672 ( .A(n4579), .B(n4561), .Z(n4570) );
  AND U4673 ( .A(n4368), .B(n1248), .Z(n4561) );
  IV U4674 ( .A(n1334), .Z(n1248) );
  IV U4675 ( .A(n4563), .Z(n4579) );
  XNOR U4676 ( .A(n4567), .B(n4569), .Z(n4126) );
  NAND U4677 ( .A(n2956), .B(n1520), .Z(n4569) );
  XNOR U4678 ( .A(n4565), .B(n4581), .Z(n4567) );
  ANDN U4679 ( .A(n2961), .B(n1522), .Z(n4581) );
  XOR U4680 ( .A(n4582), .B(n4583), .Z(n4565) );
  AND U4681 ( .A(n4584), .B(n4585), .Z(n4583) );
  XOR U4682 ( .A(n4586), .B(n4582), .Z(n4585) );
  XNOR U4683 ( .A(n4587), .B(n4576), .Z(n4127) );
  XNOR U4684 ( .A(n4574), .B(n4588), .Z(n4576) );
  ANDN U4685 ( .A(e_input[0]), .B(n1334), .Z(n4588) );
  XNOR U4686 ( .A(n4572), .B(g_input[18]), .Z(n4573) );
  ANDN U4687 ( .A(n4589), .B(n4590), .Z(n4572) );
  XOR U4688 ( .A(n4591), .B(n4592), .Z(n4574) );
  AND U4689 ( .A(n4593), .B(n4594), .Z(n4592) );
  XNOR U4690 ( .A(n4595), .B(n4591), .Z(n4594) );
  XOR U4691 ( .A(n4596), .B(n4578), .Z(n4587) );
  AND U4692 ( .A(n4368), .B(n1332), .Z(n4578) );
  IV U4693 ( .A(n1425), .Z(n1332) );
  IV U4694 ( .A(n4580), .Z(n4596) );
  XNOR U4695 ( .A(n4584), .B(n4586), .Z(n4147) );
  NAND U4696 ( .A(n2956), .B(n1616), .Z(n4586) );
  XNOR U4697 ( .A(n4582), .B(n4598), .Z(n4584) );
  ANDN U4698 ( .A(n2961), .B(n1618), .Z(n4598) );
  XOR U4699 ( .A(n4599), .B(n4600), .Z(n4582) );
  AND U4700 ( .A(n4601), .B(n4602), .Z(n4600) );
  XOR U4701 ( .A(n4603), .B(n4599), .Z(n4602) );
  XNOR U4702 ( .A(n4604), .B(n4593), .Z(n4148) );
  XNOR U4703 ( .A(n4591), .B(n4605), .Z(n4593) );
  ANDN U4704 ( .A(e_input[0]), .B(n1425), .Z(n4605) );
  ANDN U4705 ( .A(n4606), .B(n4607), .Z(n4589) );
  XOR U4706 ( .A(n4608), .B(n4609), .Z(n4591) );
  AND U4707 ( .A(n4610), .B(n4611), .Z(n4609) );
  XNOR U4708 ( .A(n4612), .B(n4608), .Z(n4611) );
  XOR U4709 ( .A(n4613), .B(n4595), .Z(n4604) );
  AND U4710 ( .A(n4368), .B(n1423), .Z(n4595) );
  IV U4711 ( .A(n1522), .Z(n1423) );
  IV U4712 ( .A(n4597), .Z(n4613) );
  XNOR U4713 ( .A(n4601), .B(n4603), .Z(n4168) );
  NAND U4714 ( .A(n2956), .B(n1712), .Z(n4603) );
  XNOR U4715 ( .A(n4599), .B(n4615), .Z(n4601) );
  ANDN U4716 ( .A(n2961), .B(n1714), .Z(n4615) );
  XNOR U4717 ( .A(n4619), .B(n4610), .Z(n4169) );
  XNOR U4718 ( .A(n4608), .B(n4620), .Z(n4610) );
  ANDN U4719 ( .A(e_input[0]), .B(n1522), .Z(n4620) );
  AND U4720 ( .A(n4368), .B(n1520), .Z(n4612) );
  XNOR U4721 ( .A(n4617), .B(n4618), .Z(n4186) );
  NAND U4722 ( .A(n2956), .B(n1813), .Z(n4618) );
  XNOR U4723 ( .A(n4616), .B(n4625), .Z(n4617) );
  ANDN U4724 ( .A(n2961), .B(n1815), .Z(n4625) );
  XNOR U4725 ( .A(n4629), .B(n4622), .Z(n4188) );
  XNOR U4726 ( .A(n4621), .B(n4630), .Z(n4622) );
  ANDN U4727 ( .A(e_input[0]), .B(n1618), .Z(n4630) );
  AND U4728 ( .A(n4368), .B(n1616), .Z(n4623) );
  XNOR U4729 ( .A(n4627), .B(n4628), .Z(n4206) );
  NAND U4730 ( .A(n2956), .B(n1919), .Z(n4628) );
  XNOR U4731 ( .A(n4626), .B(n4635), .Z(n4627) );
  ANDN U4732 ( .A(n2961), .B(n1921), .Z(n4635) );
  XNOR U4733 ( .A(n4639), .B(n4632), .Z(n4208) );
  XNOR U4734 ( .A(n4631), .B(n4640), .Z(n4632) );
  ANDN U4735 ( .A(e_input[0]), .B(n1714), .Z(n4640) );
  AND U4736 ( .A(n4368), .B(n1712), .Z(n4633) );
  XNOR U4737 ( .A(n4637), .B(n4638), .Z(n4226) );
  NAND U4738 ( .A(n2956), .B(n2026), .Z(n4638) );
  XNOR U4739 ( .A(n4636), .B(n4645), .Z(n4637) );
  ANDN U4740 ( .A(n2961), .B(n2028), .Z(n4645) );
  XNOR U4741 ( .A(n4649), .B(n4642), .Z(n4228) );
  XNOR U4742 ( .A(n4641), .B(n4650), .Z(n4642) );
  ANDN U4743 ( .A(e_input[0]), .B(n1815), .Z(n4650) );
  XOR U4744 ( .A(n4651), .B(n4652), .Z(n4641) );
  AND U4745 ( .A(n4653), .B(n4654), .Z(n4652) );
  XNOR U4746 ( .A(n4655), .B(n4651), .Z(n4654) );
  AND U4747 ( .A(n4368), .B(n1813), .Z(n4643) );
  XNOR U4748 ( .A(n4647), .B(n4648), .Z(n4246) );
  NAND U4749 ( .A(n2956), .B(n2134), .Z(n4648) );
  XNOR U4750 ( .A(n4646), .B(n4657), .Z(n4647) );
  ANDN U4751 ( .A(n2961), .B(n2136), .Z(n4657) );
  XOR U4752 ( .A(n4658), .B(n4659), .Z(n4646) );
  AND U4753 ( .A(n4660), .B(n4661), .Z(n4659) );
  XOR U4754 ( .A(n4662), .B(n4658), .Z(n4661) );
  XNOR U4755 ( .A(n4663), .B(n4653), .Z(n4248) );
  XNOR U4756 ( .A(n4651), .B(n4664), .Z(n4653) );
  ANDN U4757 ( .A(e_input[0]), .B(n1921), .Z(n4664) );
  XOR U4758 ( .A(n4665), .B(n4666), .Z(n4651) );
  AND U4759 ( .A(n4667), .B(n4668), .Z(n4666) );
  XNOR U4760 ( .A(n4669), .B(n4665), .Z(n4668) );
  XOR U4761 ( .A(n4670), .B(n4655), .Z(n4663) );
  AND U4762 ( .A(n4368), .B(n1919), .Z(n4655) );
  IV U4763 ( .A(n4656), .Z(n4670) );
  XNOR U4764 ( .A(n4660), .B(n4662), .Z(n4266) );
  NAND U4765 ( .A(n2956), .B(n2253), .Z(n4662) );
  XNOR U4766 ( .A(n4658), .B(n4672), .Z(n4660) );
  ANDN U4767 ( .A(n2961), .B(n2255), .Z(n4672) );
  XOR U4768 ( .A(n4673), .B(n4674), .Z(n4658) );
  AND U4769 ( .A(n4675), .B(n4676), .Z(n4674) );
  XOR U4770 ( .A(n4677), .B(n4673), .Z(n4676) );
  XNOR U4771 ( .A(n4678), .B(n4667), .Z(n4268) );
  XNOR U4772 ( .A(n4665), .B(n4679), .Z(n4667) );
  ANDN U4773 ( .A(e_input[0]), .B(n2028), .Z(n4679) );
  XOR U4774 ( .A(n4680), .B(n4681), .Z(n4665) );
  AND U4775 ( .A(n4682), .B(n4683), .Z(n4681) );
  XNOR U4776 ( .A(n4684), .B(n4680), .Z(n4683) );
  XOR U4777 ( .A(n4685), .B(n4669), .Z(n4678) );
  AND U4778 ( .A(n4368), .B(n2026), .Z(n4669) );
  IV U4779 ( .A(n4671), .Z(n4685) );
  XNOR U4780 ( .A(n4675), .B(n4677), .Z(n4286) );
  NAND U4781 ( .A(n2956), .B(n2373), .Z(n4677) );
  XNOR U4782 ( .A(n4673), .B(n4687), .Z(n4675) );
  ANDN U4783 ( .A(n2961), .B(n2375), .Z(n4687) );
  XNOR U4784 ( .A(n4691), .B(n4682), .Z(n4288) );
  XNOR U4785 ( .A(n4680), .B(n4692), .Z(n4682) );
  ANDN U4786 ( .A(e_input[0]), .B(n2136), .Z(n4692) );
  XOR U4787 ( .A(n4693), .B(n4694), .Z(n4680) );
  AND U4788 ( .A(n4695), .B(n4696), .Z(n4694) );
  XNOR U4789 ( .A(n4697), .B(n4693), .Z(n4696) );
  AND U4790 ( .A(n4368), .B(n2134), .Z(n4684) );
  XNOR U4791 ( .A(n4689), .B(n4690), .Z(n4310) );
  NAND U4792 ( .A(n2956), .B(n2495), .Z(n4690) );
  XNOR U4793 ( .A(n4688), .B(n4699), .Z(n4689) );
  ANDN U4794 ( .A(n2961), .B(n2497), .Z(n4699) );
  XNOR U4795 ( .A(n4703), .B(n4695), .Z(n4312) );
  XNOR U4796 ( .A(n4693), .B(n4704), .Z(n4695) );
  ANDN U4797 ( .A(e_input[0]), .B(n2255), .Z(n4704) );
  XOR U4798 ( .A(n4705), .B(n4706), .Z(n4693) );
  AND U4799 ( .A(n4707), .B(n4708), .Z(n4706) );
  XNOR U4800 ( .A(n4709), .B(n4705), .Z(n4708) );
  AND U4801 ( .A(n4368), .B(n2253), .Z(n4697) );
  XNOR U4802 ( .A(n4701), .B(n4702), .Z(n4330) );
  NAND U4803 ( .A(n2956), .B(n2620), .Z(n4702) );
  XNOR U4804 ( .A(n4700), .B(n4711), .Z(n4701) );
  ANDN U4805 ( .A(n2961), .B(n2622), .Z(n4711) );
  XNOR U4806 ( .A(n4715), .B(n4707), .Z(n4331) );
  XNOR U4807 ( .A(n4705), .B(n4716), .Z(n4707) );
  ANDN U4808 ( .A(e_input[0]), .B(n2375), .Z(n4716) );
  AND U4809 ( .A(n4368), .B(n2373), .Z(n4709) );
  XNOR U4810 ( .A(n4720), .B(n4721), .Z(n4710) );
  AND U4811 ( .A(n4722), .B(n4723), .Z(n4721) );
  XNOR U4812 ( .A(n4718), .B(n4724), .Z(n4723) );
  XNOR U4813 ( .A(n4719), .B(n4720), .Z(n4724) );
  AND U4814 ( .A(n4368), .B(n2495), .Z(n4719) );
  XOR U4815 ( .A(n4717), .B(n4725), .Z(n4718) );
  ANDN U4816 ( .A(e_input[0]), .B(n2497), .Z(n4725) );
  XNOR U4817 ( .A(n4713), .B(n4729), .Z(n4722) );
  XNOR U4818 ( .A(n4714), .B(n4720), .Z(n4729) );
  AND U4819 ( .A(n2752), .B(n2956), .Z(n4714) );
  XOR U4820 ( .A(n4712), .B(n4730), .Z(n4713) );
  ANDN U4821 ( .A(n2961), .B(n2754), .Z(n4730) );
  XOR U4822 ( .A(n4734), .B(n4735), .Z(n4720) );
  AND U4823 ( .A(n4736), .B(n4737), .Z(n4735) );
  XNOR U4824 ( .A(n4727), .B(n4738), .Z(n4737) );
  XNOR U4825 ( .A(n4728), .B(n4734), .Z(n4738) );
  AND U4826 ( .A(n4368), .B(n2620), .Z(n4728) );
  XOR U4827 ( .A(n4726), .B(n4739), .Z(n4727) );
  ANDN U4828 ( .A(e_input[0]), .B(n2622), .Z(n4739) );
  XNOR U4829 ( .A(n4732), .B(n4743), .Z(n4736) );
  XNOR U4830 ( .A(n4733), .B(n4734), .Z(n4743) );
  AND U4831 ( .A(n2884), .B(n2956), .Z(n4733) );
  XOR U4832 ( .A(n4731), .B(n4744), .Z(n4732) );
  ANDN U4833 ( .A(n2961), .B(n2886), .Z(n4744) );
  XOR U4834 ( .A(n4745), .B(n4746), .Z(n4731) );
  ANDN U4835 ( .A(n4747), .B(n4748), .Z(n4746) );
  XNOR U4836 ( .A(n4749), .B(n4745), .Z(n4747) );
  XOR U4837 ( .A(n4750), .B(n4751), .Z(n4734) );
  AND U4838 ( .A(n4752), .B(n4753), .Z(n4751) );
  XNOR U4839 ( .A(n4741), .B(n4754), .Z(n4753) );
  XNOR U4840 ( .A(n4742), .B(n4750), .Z(n4754) );
  AND U4841 ( .A(n4368), .B(n2752), .Z(n4742) );
  XOR U4842 ( .A(n4740), .B(n4755), .Z(n4741) );
  ANDN U4843 ( .A(e_input[0]), .B(n2754), .Z(n4755) );
  XNOR U4844 ( .A(n4748), .B(n4759), .Z(n4752) );
  XNOR U4845 ( .A(n4749), .B(n4750), .Z(n4759) );
  AND U4846 ( .A(n3025), .B(n2956), .Z(n4749) );
  XOR U4847 ( .A(n4745), .B(n4760), .Z(n4748) );
  ANDN U4848 ( .A(n2961), .B(n3027), .Z(n4760) );
  XNOR U4849 ( .A(n4765), .B(n4757), .Z(n4351) );
  XNOR U4850 ( .A(n4756), .B(n4766), .Z(n4757) );
  ANDN U4851 ( .A(e_input[0]), .B(n2886), .Z(n4766) );
  XNOR U4852 ( .A(n4769), .B(n4767), .Z(n4768) );
  ANDN U4853 ( .A(e_input[0]), .B(n3027), .Z(n4769) );
  ANDN U4854 ( .A(n4368), .B(n3815), .Z(n4770) );
  XNOR U4855 ( .A(n4764), .B(n4758), .Z(n4765) );
  AND U4856 ( .A(n4368), .B(n2884), .Z(n4758) );
  XNOR U4857 ( .A(n4762), .B(n4763), .Z(n4350) );
  NAND U4858 ( .A(n3813), .B(n2956), .Z(n4763) );
  XNOR U4859 ( .A(n4761), .B(n4774), .Z(n4762) );
  ANDN U4860 ( .A(n2961), .B(n3815), .Z(n4774) );
  NAND U4861 ( .A(g_input[0]), .B(n4775), .Z(n4761) );
  NANDN U4862 ( .B(n2956), .A(n4776), .Z(n4775) );
  NANDN U4863 ( .B(n3818), .A(n2961), .Z(n4776) );
  IV U4864 ( .A(n2822), .Z(n2956) );
  XNOR U4865 ( .A(n4772), .B(n4773), .Z(n4764) );
  NAND U4866 ( .A(n3813), .B(n4368), .Z(n4773) );
  XNOR U4867 ( .A(n4771), .B(n4779), .Z(n4772) );
  ANDN U4868 ( .A(e_input[0]), .B(n3815), .Z(n4779) );
  NAND U4869 ( .A(g_input[0]), .B(n4780), .Z(n4771) );
  NANDN U4870 ( .B(n4368), .A(n4781), .Z(n4780) );
  NANDN U4871 ( .B(n3818), .A(e_input[0]), .Z(n4781) );
  IV U4872 ( .A(n4355), .Z(n4368) );
  XNOR U4873 ( .A(n2984), .B(n2983), .Z(n2937) );
  XOR U4874 ( .A(n4783), .B(n2992), .Z(n2983) );
  XNOR U4875 ( .A(n2977), .B(n2976), .Z(n2992) );
  XOR U4876 ( .A(n4784), .B(n2973), .Z(n2976) );
  XNOR U4877 ( .A(n2972), .B(n4785), .Z(n2973) );
  ANDN U4878 ( .A(n1036), .B(n1921), .Z(n4785) );
  AND U4879 ( .A(n1919), .B(n973), .Z(n2974) );
  XNOR U4880 ( .A(n2980), .B(n2981), .Z(n2977) );
  NANDN U4881 ( .B(n838), .A(n2134), .Z(n2981) );
  XNOR U4882 ( .A(n2979), .B(n4792), .Z(n2980) );
  ANDN U4883 ( .A(n908), .B(n2136), .Z(n4792) );
  XOR U4884 ( .A(n2991), .B(n2982), .Z(n4783) );
  XNOR U4885 ( .A(n4796), .B(n4797), .Z(n2982) );
  XOR U4886 ( .A(n4798), .B(n3000), .Z(n2991) );
  XNOR U4887 ( .A(n2988), .B(n2989), .Z(n3000) );
  NAND U4888 ( .A(n1712), .B(n1207), .Z(n2989) );
  XNOR U4889 ( .A(n2987), .B(n4799), .Z(n2988) );
  ANDN U4890 ( .A(n1214), .B(n1714), .Z(n4799) );
  XNOR U4891 ( .A(n2999), .B(n2990), .Z(n4798) );
  XOR U4892 ( .A(n4803), .B(n4804), .Z(n2990) );
  AND U4893 ( .A(n4805), .B(n4806), .Z(n4804) );
  XOR U4894 ( .A(n4807), .B(n4808), .Z(n4806) );
  XNOR U4895 ( .A(n4803), .B(n4809), .Z(n4808) );
  XNOR U4896 ( .A(n4790), .B(n4810), .Z(n4805) );
  XNOR U4897 ( .A(n4803), .B(n4791), .Z(n4810) );
  XNOR U4898 ( .A(n4794), .B(n4795), .Z(n4791) );
  NANDN U4899 ( .B(n838), .A(n2253), .Z(n4795) );
  XNOR U4900 ( .A(n4793), .B(n4811), .Z(n4794) );
  ANDN U4901 ( .A(n908), .B(n2255), .Z(n4811) );
  XOR U4902 ( .A(n4815), .B(n4787), .Z(n4790) );
  XNOR U4903 ( .A(n4786), .B(n4816), .Z(n4787) );
  ANDN U4904 ( .A(n1036), .B(n2028), .Z(n4816) );
  AND U4905 ( .A(n2026), .B(n973), .Z(n4788) );
  XOR U4906 ( .A(n4823), .B(n4824), .Z(n4803) );
  AND U4907 ( .A(n4825), .B(n4826), .Z(n4824) );
  XOR U4908 ( .A(n4827), .B(n4828), .Z(n4826) );
  XNOR U4909 ( .A(n4823), .B(n4829), .Z(n4828) );
  XNOR U4910 ( .A(n4821), .B(n4830), .Z(n4825) );
  XNOR U4911 ( .A(n4823), .B(n4822), .Z(n4830) );
  XNOR U4912 ( .A(n4813), .B(n4814), .Z(n4822) );
  NANDN U4913 ( .B(n838), .A(n2373), .Z(n4814) );
  XNOR U4914 ( .A(n4812), .B(n4831), .Z(n4813) );
  ANDN U4915 ( .A(n908), .B(n2375), .Z(n4831) );
  XOR U4916 ( .A(n4835), .B(n4818), .Z(n4821) );
  XNOR U4917 ( .A(n4817), .B(n4836), .Z(n4818) );
  ANDN U4918 ( .A(n1036), .B(n2136), .Z(n4836) );
  AND U4919 ( .A(n2134), .B(n973), .Z(n4819) );
  XOR U4920 ( .A(n4843), .B(n4844), .Z(n4823) );
  AND U4921 ( .A(n4845), .B(n4846), .Z(n4844) );
  XOR U4922 ( .A(n4847), .B(n4848), .Z(n4846) );
  XNOR U4923 ( .A(n4843), .B(n4849), .Z(n4848) );
  XNOR U4924 ( .A(n4841), .B(n4850), .Z(n4845) );
  XNOR U4925 ( .A(n4843), .B(n4842), .Z(n4850) );
  XNOR U4926 ( .A(n4833), .B(n4834), .Z(n4842) );
  NANDN U4927 ( .B(n838), .A(n2495), .Z(n4834) );
  XNOR U4928 ( .A(n4832), .B(n4851), .Z(n4833) );
  ANDN U4929 ( .A(n908), .B(n2497), .Z(n4851) );
  XOR U4930 ( .A(n4855), .B(n4838), .Z(n4841) );
  XNOR U4931 ( .A(n4837), .B(n4856), .Z(n4838) );
  ANDN U4932 ( .A(n1036), .B(n2255), .Z(n4856) );
  AND U4933 ( .A(n2253), .B(n973), .Z(n4839) );
  XOR U4934 ( .A(n4863), .B(n4864), .Z(n4843) );
  AND U4935 ( .A(n4865), .B(n4866), .Z(n4864) );
  XOR U4936 ( .A(n4867), .B(n4868), .Z(n4866) );
  XNOR U4937 ( .A(n4863), .B(n4869), .Z(n4868) );
  XNOR U4938 ( .A(n4861), .B(n4870), .Z(n4865) );
  XNOR U4939 ( .A(n4863), .B(n4862), .Z(n4870) );
  XNOR U4940 ( .A(n4853), .B(n4854), .Z(n4862) );
  NANDN U4941 ( .B(n838), .A(n2620), .Z(n4854) );
  XNOR U4942 ( .A(n4852), .B(n4871), .Z(n4853) );
  ANDN U4943 ( .A(n908), .B(n2622), .Z(n4871) );
  XOR U4944 ( .A(n4875), .B(n4858), .Z(n4861) );
  XNOR U4945 ( .A(n4857), .B(n4876), .Z(n4858) );
  ANDN U4946 ( .A(n1036), .B(n2375), .Z(n4876) );
  AND U4947 ( .A(n2373), .B(n973), .Z(n4859) );
  XOR U4948 ( .A(n4883), .B(n4884), .Z(n4863) );
  AND U4949 ( .A(n4885), .B(n4886), .Z(n4884) );
  XOR U4950 ( .A(n4887), .B(n4888), .Z(n4886) );
  XNOR U4951 ( .A(n4883), .B(n4889), .Z(n4888) );
  XNOR U4952 ( .A(n4881), .B(n4890), .Z(n4885) );
  XNOR U4953 ( .A(n4883), .B(n4882), .Z(n4890) );
  XNOR U4954 ( .A(n4873), .B(n4874), .Z(n4882) );
  NANDN U4955 ( .B(n838), .A(n2752), .Z(n4874) );
  XNOR U4956 ( .A(n4872), .B(n4891), .Z(n4873) );
  ANDN U4957 ( .A(n908), .B(n2754), .Z(n4891) );
  XOR U4958 ( .A(n4895), .B(n4878), .Z(n4881) );
  XNOR U4959 ( .A(n4877), .B(n4896), .Z(n4878) );
  ANDN U4960 ( .A(n1036), .B(n2497), .Z(n4896) );
  XOR U4961 ( .A(n4897), .B(n4898), .Z(n4877) );
  AND U4962 ( .A(n4899), .B(n4900), .Z(n4898) );
  XNOR U4963 ( .A(n4901), .B(n4897), .Z(n4900) );
  AND U4964 ( .A(n2495), .B(n973), .Z(n4879) );
  XOR U4965 ( .A(n4905), .B(n4906), .Z(n4883) );
  AND U4966 ( .A(n4907), .B(n4908), .Z(n4906) );
  XOR U4967 ( .A(n4909), .B(n4910), .Z(n4908) );
  XNOR U4968 ( .A(n4905), .B(n4911), .Z(n4910) );
  XNOR U4969 ( .A(n4903), .B(n4912), .Z(n4907) );
  XNOR U4970 ( .A(n4905), .B(n4904), .Z(n4912) );
  XNOR U4971 ( .A(n4893), .B(n4894), .Z(n4904) );
  NANDN U4972 ( .B(n838), .A(n2884), .Z(n4894) );
  XNOR U4973 ( .A(n4892), .B(n4913), .Z(n4893) );
  ANDN U4974 ( .A(n908), .B(n2886), .Z(n4913) );
  XOR U4975 ( .A(n4914), .B(n4915), .Z(n4892) );
  AND U4976 ( .A(n4916), .B(n4917), .Z(n4915) );
  XOR U4977 ( .A(n4918), .B(n4914), .Z(n4917) );
  XOR U4978 ( .A(n4919), .B(n4899), .Z(n4903) );
  XNOR U4979 ( .A(n4897), .B(n4920), .Z(n4899) );
  ANDN U4980 ( .A(n1036), .B(n2622), .Z(n4920) );
  XOR U4981 ( .A(n4921), .B(n4922), .Z(n4897) );
  AND U4982 ( .A(n4923), .B(n4924), .Z(n4922) );
  XNOR U4983 ( .A(n4925), .B(n4921), .Z(n4924) );
  AND U4984 ( .A(n2620), .B(n973), .Z(n4901) );
  XOR U4985 ( .A(n4929), .B(n4930), .Z(n4905) );
  AND U4986 ( .A(n4931), .B(n4932), .Z(n4930) );
  XOR U4987 ( .A(n4933), .B(n4934), .Z(n4932) );
  XNOR U4988 ( .A(n4929), .B(n4935), .Z(n4934) );
  XNOR U4989 ( .A(n4927), .B(n4936), .Z(n4931) );
  XNOR U4990 ( .A(n4929), .B(n4928), .Z(n4936) );
  XNOR U4991 ( .A(n4916), .B(n4918), .Z(n4928) );
  NANDN U4992 ( .B(n838), .A(n3025), .Z(n4918) );
  XNOR U4993 ( .A(n4914), .B(n4937), .Z(n4916) );
  ANDN U4994 ( .A(n908), .B(n3027), .Z(n4937) );
  XOR U4995 ( .A(n4941), .B(n4923), .Z(n4927) );
  XNOR U4996 ( .A(n4921), .B(n4942), .Z(n4923) );
  ANDN U4997 ( .A(n1036), .B(n2754), .Z(n4942) );
  AND U4998 ( .A(n2752), .B(n973), .Z(n4925) );
  XOR U4999 ( .A(n4950), .B(n4951), .Z(n4797) );
  XNOR U5000 ( .A(n4948), .B(n4947), .Z(n4796) );
  XOR U5001 ( .A(n4953), .B(n4944), .Z(n4947) );
  XNOR U5002 ( .A(n4943), .B(n4954), .Z(n4944) );
  ANDN U5003 ( .A(n1036), .B(n2886), .Z(n4954) );
  XNOR U5004 ( .A(n4957), .B(n4955), .Z(n4956) );
  ANDN U5005 ( .A(n1036), .B(n3027), .Z(n4957) );
  XNOR U5006 ( .A(n4946), .B(n4945), .Z(n4953) );
  AND U5007 ( .A(n2884), .B(n973), .Z(n4945) );
  XNOR U5008 ( .A(n4960), .B(n4961), .Z(n4946) );
  NAND U5009 ( .A(n3813), .B(n973), .Z(n4961) );
  XNOR U5010 ( .A(n4959), .B(n4962), .Z(n4960) );
  ANDN U5011 ( .A(n1036), .B(n3815), .Z(n4962) );
  NAND U5012 ( .A(g_input[0]), .B(n4963), .Z(n4959) );
  NANDN U5013 ( .B(n973), .A(n4964), .Z(n4963) );
  NANDN U5014 ( .B(n3818), .A(n1036), .Z(n4964) );
  IV U5015 ( .A(n4958), .Z(n973) );
  XNOR U5016 ( .A(n4939), .B(n4940), .Z(n4948) );
  NANDN U5017 ( .B(n838), .A(n3813), .Z(n4940) );
  XNOR U5018 ( .A(n4938), .B(n4967), .Z(n4939) );
  ANDN U5019 ( .A(n908), .B(n3815), .Z(n4967) );
  NAND U5020 ( .A(g_input[0]), .B(n4968), .Z(n4938) );
  NAND U5021 ( .A(n4969), .B(n838), .Z(n4968) );
  NANDN U5022 ( .B(n3818), .A(n908), .Z(n4969) );
  XOR U5023 ( .A(n4972), .B(n4973), .Z(n4949) );
  XOR U5024 ( .A(n4974), .B(n2996), .Z(n2999) );
  XNOR U5025 ( .A(n2995), .B(n4975), .Z(n2996) );
  ANDN U5026 ( .A(n1398), .B(n1522), .Z(n4975) );
  XNOR U5027 ( .A(n4606), .B(g_input[16]), .Z(n4607) );
  ANDN U5028 ( .A(n4976), .B(n4977), .Z(n4606) );
  AND U5029 ( .A(n1520), .B(n1391), .Z(n2997) );
  IV U5030 ( .A(n1618), .Z(n1520) );
  XNOR U5031 ( .A(n4801), .B(n4802), .Z(n4807) );
  NAND U5032 ( .A(n1813), .B(n1207), .Z(n4802) );
  XNOR U5033 ( .A(n4800), .B(n4982), .Z(n4801) );
  ANDN U5034 ( .A(n1214), .B(n1815), .Z(n4982) );
  XNOR U5035 ( .A(n4986), .B(n4979), .Z(n4809) );
  XNOR U5036 ( .A(n4978), .B(n4987), .Z(n4979) );
  ANDN U5037 ( .A(n1398), .B(n1618), .Z(n4987) );
  ANDN U5038 ( .A(n4988), .B(n4989), .Z(n4976) );
  AND U5039 ( .A(n1616), .B(n1391), .Z(n4980) );
  IV U5040 ( .A(n1714), .Z(n1616) );
  XNOR U5041 ( .A(n4984), .B(n4985), .Z(n4827) );
  NAND U5042 ( .A(n1919), .B(n1207), .Z(n4985) );
  XNOR U5043 ( .A(n4983), .B(n4994), .Z(n4984) );
  ANDN U5044 ( .A(n1214), .B(n1921), .Z(n4994) );
  XNOR U5045 ( .A(n4998), .B(n4991), .Z(n4829) );
  XNOR U5046 ( .A(n4990), .B(n4999), .Z(n4991) );
  ANDN U5047 ( .A(n1398), .B(n1714), .Z(n4999) );
  XNOR U5048 ( .A(n4988), .B(g_input[14]), .Z(n4989) );
  ANDN U5049 ( .A(n5000), .B(n5001), .Z(n4988) );
  AND U5050 ( .A(n1712), .B(n1391), .Z(n4992) );
  IV U5051 ( .A(n1815), .Z(n1712) );
  XNOR U5052 ( .A(n4996), .B(n4997), .Z(n4847) );
  NAND U5053 ( .A(n2026), .B(n1207), .Z(n4997) );
  XNOR U5054 ( .A(n4995), .B(n5006), .Z(n4996) );
  ANDN U5055 ( .A(n1214), .B(n2028), .Z(n5006) );
  XNOR U5056 ( .A(n5010), .B(n5003), .Z(n4849) );
  XNOR U5057 ( .A(n5002), .B(n5011), .Z(n5003) );
  ANDN U5058 ( .A(n1398), .B(n1815), .Z(n5011) );
  ANDN U5059 ( .A(n5012), .B(n5013), .Z(n5000) );
  AND U5060 ( .A(n1813), .B(n1391), .Z(n5004) );
  IV U5061 ( .A(n1921), .Z(n1813) );
  XNOR U5062 ( .A(n5008), .B(n5009), .Z(n4867) );
  NAND U5063 ( .A(n2134), .B(n1207), .Z(n5009) );
  XNOR U5064 ( .A(n5007), .B(n5018), .Z(n5008) );
  ANDN U5065 ( .A(n1214), .B(n2136), .Z(n5018) );
  XNOR U5066 ( .A(n5022), .B(n5015), .Z(n4869) );
  XNOR U5067 ( .A(n5014), .B(n5023), .Z(n5015) );
  ANDN U5068 ( .A(n1398), .B(n1921), .Z(n5023) );
  XNOR U5069 ( .A(n5012), .B(g_input[12]), .Z(n5013) );
  ANDN U5070 ( .A(n5024), .B(n5025), .Z(n5012) );
  AND U5071 ( .A(n1919), .B(n1391), .Z(n5016) );
  IV U5072 ( .A(n2028), .Z(n1919) );
  XNOR U5073 ( .A(n5020), .B(n5021), .Z(n4887) );
  NAND U5074 ( .A(n2253), .B(n1207), .Z(n5021) );
  XNOR U5075 ( .A(n5019), .B(n5030), .Z(n5020) );
  ANDN U5076 ( .A(n1214), .B(n2255), .Z(n5030) );
  XOR U5077 ( .A(n5031), .B(n5032), .Z(n5019) );
  AND U5078 ( .A(n5033), .B(n5034), .Z(n5032) );
  XOR U5079 ( .A(n5035), .B(n5031), .Z(n5034) );
  XNOR U5080 ( .A(n5036), .B(n5027), .Z(n4889) );
  XNOR U5081 ( .A(n5026), .B(n5037), .Z(n5027) );
  ANDN U5082 ( .A(n1398), .B(n2028), .Z(n5037) );
  ANDN U5083 ( .A(n5038), .B(n5039), .Z(n5024) );
  AND U5084 ( .A(n2026), .B(n1391), .Z(n5028) );
  IV U5085 ( .A(n2136), .Z(n2026) );
  XNOR U5086 ( .A(n5033), .B(n5035), .Z(n4909) );
  NAND U5087 ( .A(n2373), .B(n1207), .Z(n5035) );
  XNOR U5088 ( .A(n5031), .B(n5044), .Z(n5033) );
  ANDN U5089 ( .A(n1214), .B(n2375), .Z(n5044) );
  XOR U5090 ( .A(n5045), .B(n5046), .Z(n5031) );
  AND U5091 ( .A(n5047), .B(n5048), .Z(n5046) );
  XOR U5092 ( .A(n5049), .B(n5045), .Z(n5048) );
  XNOR U5093 ( .A(n5050), .B(n5041), .Z(n4911) );
  XNOR U5094 ( .A(n5040), .B(n5051), .Z(n5041) );
  ANDN U5095 ( .A(n1398), .B(n2136), .Z(n5051) );
  XNOR U5096 ( .A(n5038), .B(g_input[10]), .Z(n5039) );
  ANDN U5097 ( .A(n5052), .B(n5053), .Z(n5038) );
  XOR U5098 ( .A(n5054), .B(n5055), .Z(n5040) );
  AND U5099 ( .A(n5056), .B(n5057), .Z(n5055) );
  XNOR U5100 ( .A(n5058), .B(n5054), .Z(n5057) );
  XOR U5101 ( .A(n5059), .B(n5042), .Z(n5050) );
  AND U5102 ( .A(n2134), .B(n1391), .Z(n5042) );
  IV U5103 ( .A(n2255), .Z(n2134) );
  IV U5104 ( .A(n5043), .Z(n5059) );
  XNOR U5105 ( .A(n5047), .B(n5049), .Z(n4933) );
  NAND U5106 ( .A(n2495), .B(n1207), .Z(n5049) );
  XNOR U5107 ( .A(n5045), .B(n5061), .Z(n5047) );
  ANDN U5108 ( .A(n1214), .B(n2497), .Z(n5061) );
  XNOR U5109 ( .A(n5065), .B(n5056), .Z(n4935) );
  XNOR U5110 ( .A(n5054), .B(n5066), .Z(n5056) );
  ANDN U5111 ( .A(n1398), .B(n2255), .Z(n5066) );
  ANDN U5112 ( .A(n5067), .B(n5068), .Z(n5052) );
  XOR U5113 ( .A(n5069), .B(n5070), .Z(n5054) );
  AND U5114 ( .A(n5071), .B(n5072), .Z(n5070) );
  XNOR U5115 ( .A(n5073), .B(n5069), .Z(n5072) );
  AND U5116 ( .A(n2253), .B(n1391), .Z(n5058) );
  IV U5117 ( .A(n2375), .Z(n2253) );
  XNOR U5118 ( .A(n5063), .B(n5064), .Z(n4951) );
  NAND U5119 ( .A(n2620), .B(n1207), .Z(n5064) );
  XNOR U5120 ( .A(n5062), .B(n5075), .Z(n5063) );
  ANDN U5121 ( .A(n1214), .B(n2622), .Z(n5075) );
  XNOR U5122 ( .A(n5079), .B(n5071), .Z(n4952) );
  XNOR U5123 ( .A(n5069), .B(n5080), .Z(n5071) );
  ANDN U5124 ( .A(n1398), .B(n2375), .Z(n5080) );
  AND U5125 ( .A(n2373), .B(n1391), .Z(n5073) );
  XNOR U5126 ( .A(n5084), .B(n5085), .Z(n5074) );
  AND U5127 ( .A(n5086), .B(n5087), .Z(n5085) );
  XNOR U5128 ( .A(n5082), .B(n5088), .Z(n5087) );
  XNOR U5129 ( .A(n5083), .B(n5084), .Z(n5088) );
  AND U5130 ( .A(n2495), .B(n1391), .Z(n5083) );
  XOR U5131 ( .A(n5081), .B(n5089), .Z(n5082) );
  ANDN U5132 ( .A(n1398), .B(n2497), .Z(n5089) );
  XNOR U5133 ( .A(n5077), .B(n5093), .Z(n5086) );
  XNOR U5134 ( .A(n5078), .B(n5084), .Z(n5093) );
  AND U5135 ( .A(n2752), .B(n1207), .Z(n5078) );
  XOR U5136 ( .A(n5076), .B(n5094), .Z(n5077) );
  ANDN U5137 ( .A(n1214), .B(n2754), .Z(n5094) );
  XOR U5138 ( .A(n5098), .B(n5099), .Z(n5084) );
  AND U5139 ( .A(n5100), .B(n5101), .Z(n5099) );
  XNOR U5140 ( .A(n5091), .B(n5102), .Z(n5101) );
  XNOR U5141 ( .A(n5092), .B(n5098), .Z(n5102) );
  AND U5142 ( .A(n2620), .B(n1391), .Z(n5092) );
  XOR U5143 ( .A(n5090), .B(n5103), .Z(n5091) );
  ANDN U5144 ( .A(n1398), .B(n2622), .Z(n5103) );
  XNOR U5145 ( .A(n5096), .B(n5107), .Z(n5100) );
  XNOR U5146 ( .A(n5097), .B(n5098), .Z(n5107) );
  AND U5147 ( .A(n2884), .B(n1207), .Z(n5097) );
  XOR U5148 ( .A(n5095), .B(n5108), .Z(n5096) );
  ANDN U5149 ( .A(n1214), .B(n2886), .Z(n5108) );
  XOR U5150 ( .A(n5109), .B(n5110), .Z(n5095) );
  ANDN U5151 ( .A(n5111), .B(n5112), .Z(n5110) );
  XNOR U5152 ( .A(n5113), .B(n5109), .Z(n5111) );
  XOR U5153 ( .A(n5114), .B(n5115), .Z(n5098) );
  AND U5154 ( .A(n5116), .B(n5117), .Z(n5115) );
  XNOR U5155 ( .A(n5105), .B(n5118), .Z(n5117) );
  XNOR U5156 ( .A(n5106), .B(n5114), .Z(n5118) );
  AND U5157 ( .A(n2752), .B(n1391), .Z(n5106) );
  XOR U5158 ( .A(n5104), .B(n5119), .Z(n5105) );
  ANDN U5159 ( .A(n1398), .B(n2754), .Z(n5119) );
  XNOR U5160 ( .A(n5112), .B(n5123), .Z(n5116) );
  XNOR U5161 ( .A(n5113), .B(n5114), .Z(n5123) );
  AND U5162 ( .A(n3025), .B(n1207), .Z(n5113) );
  XOR U5163 ( .A(n5109), .B(n5124), .Z(n5112) );
  ANDN U5164 ( .A(n1214), .B(n3027), .Z(n5124) );
  XNOR U5165 ( .A(n5129), .B(n5121), .Z(n4973) );
  XNOR U5166 ( .A(n5120), .B(n5130), .Z(n5121) );
  ANDN U5167 ( .A(n1398), .B(n2886), .Z(n5130) );
  XNOR U5168 ( .A(n5133), .B(n5131), .Z(n5132) );
  ANDN U5169 ( .A(n1398), .B(n3027), .Z(n5133) );
  XNOR U5170 ( .A(n5128), .B(n5122), .Z(n5129) );
  AND U5171 ( .A(n2884), .B(n1391), .Z(n5122) );
  XNOR U5172 ( .A(n5126), .B(n5127), .Z(n4972) );
  NAND U5173 ( .A(n3813), .B(n1207), .Z(n5127) );
  XNOR U5174 ( .A(n5125), .B(n5137), .Z(n5126) );
  ANDN U5175 ( .A(n1214), .B(n3815), .Z(n5137) );
  NAND U5176 ( .A(g_input[0]), .B(n5138), .Z(n5125) );
  NANDN U5177 ( .B(n1207), .A(n5139), .Z(n5138) );
  NANDN U5178 ( .B(n3818), .A(n1214), .Z(n5139) );
  IV U5179 ( .A(n1133), .Z(n1207) );
  XNOR U5180 ( .A(n5135), .B(n5136), .Z(n5128) );
  NAND U5181 ( .A(n3813), .B(n1391), .Z(n5136) );
  XNOR U5182 ( .A(n5134), .B(n5142), .Z(n5135) );
  ANDN U5183 ( .A(n1398), .B(n3815), .Z(n5142) );
  NAND U5184 ( .A(g_input[0]), .B(n5143), .Z(n5134) );
  NANDN U5185 ( .B(n1391), .A(n5144), .Z(n5143) );
  NANDN U5186 ( .B(n3818), .A(n1398), .Z(n5144) );
  IV U5187 ( .A(n1298), .Z(n1391) );
  XNOR U5188 ( .A(n3008), .B(n3007), .Z(n2984) );
  XOR U5189 ( .A(n5147), .B(n3016), .Z(n3007) );
  XNOR U5190 ( .A(n3004), .B(n3005), .Z(n3016) );
  NANDN U5191 ( .B(n651), .A(n2620), .Z(n3005) );
  XNOR U5192 ( .A(n3003), .B(n5148), .Z(n3004) );
  ANDN U5193 ( .A(n692), .B(n2622), .Z(n5148) );
  XOR U5194 ( .A(n3015), .B(n3006), .Z(n5147) );
  XOR U5195 ( .A(n5152), .B(n5153), .Z(n3006) );
  XOR U5196 ( .A(n5154), .B(n3012), .Z(n3015) );
  XNOR U5197 ( .A(n3011), .B(n5155), .Z(n3012) );
  ANDN U5198 ( .A(n799), .B(n2375), .Z(n5155) );
  XNOR U5199 ( .A(n5067), .B(g_input[8]), .Z(n5068) );
  ANDN U5200 ( .A(n5156), .B(n5157), .Z(n5067) );
  AND U5201 ( .A(n2373), .B(n745), .Z(n3013) );
  IV U5202 ( .A(n2497), .Z(n2373) );
  XNOR U5203 ( .A(n5161), .B(n5162), .Z(n3014) );
  AND U5204 ( .A(n5163), .B(n5164), .Z(n5162) );
  XNOR U5205 ( .A(n5159), .B(n5165), .Z(n5164) );
  XNOR U5206 ( .A(n5160), .B(n5161), .Z(n5165) );
  AND U5207 ( .A(n2495), .B(n745), .Z(n5160) );
  IV U5208 ( .A(n2622), .Z(n2495) );
  XOR U5209 ( .A(n5158), .B(n5166), .Z(n5159) );
  ANDN U5210 ( .A(n799), .B(n2497), .Z(n5166) );
  ANDN U5211 ( .A(n5167), .B(n5168), .Z(n5156) );
  XNOR U5212 ( .A(n5150), .B(n5172), .Z(n5163) );
  XNOR U5213 ( .A(n5151), .B(n5161), .Z(n5172) );
  ANDN U5214 ( .A(n2752), .B(n651), .Z(n5151) );
  XOR U5215 ( .A(n5149), .B(n5173), .Z(n5150) );
  ANDN U5216 ( .A(n692), .B(n2754), .Z(n5173) );
  XOR U5217 ( .A(n5177), .B(n5178), .Z(n5161) );
  AND U5218 ( .A(n5179), .B(n5180), .Z(n5178) );
  XNOR U5219 ( .A(n5170), .B(n5181), .Z(n5180) );
  XNOR U5220 ( .A(n5171), .B(n5177), .Z(n5181) );
  AND U5221 ( .A(n2620), .B(n745), .Z(n5171) );
  IV U5222 ( .A(n2754), .Z(n2620) );
  XOR U5223 ( .A(n5169), .B(n5182), .Z(n5170) );
  ANDN U5224 ( .A(n799), .B(n2622), .Z(n5182) );
  XNOR U5225 ( .A(n5167), .B(g_input[6]), .Z(n5168) );
  ANDN U5226 ( .A(n5183), .B(n5184), .Z(n5167) );
  XNOR U5227 ( .A(n5175), .B(n5188), .Z(n5179) );
  XNOR U5228 ( .A(n5176), .B(n5177), .Z(n5188) );
  ANDN U5229 ( .A(n2884), .B(n651), .Z(n5176) );
  XOR U5230 ( .A(n5174), .B(n5189), .Z(n5175) );
  ANDN U5231 ( .A(n692), .B(n2886), .Z(n5189) );
  XOR U5232 ( .A(n5190), .B(n5191), .Z(n5174) );
  ANDN U5233 ( .A(n5192), .B(n5193), .Z(n5191) );
  XNOR U5234 ( .A(n5194), .B(n5190), .Z(n5192) );
  XOR U5235 ( .A(n5195), .B(n5196), .Z(n5177) );
  AND U5236 ( .A(n5197), .B(n5198), .Z(n5196) );
  XNOR U5237 ( .A(n5186), .B(n5199), .Z(n5198) );
  XNOR U5238 ( .A(n5187), .B(n5195), .Z(n5199) );
  AND U5239 ( .A(n2752), .B(n745), .Z(n5187) );
  XOR U5240 ( .A(n5185), .B(n5200), .Z(n5186) );
  ANDN U5241 ( .A(n799), .B(n2754), .Z(n5200) );
  ANDN U5242 ( .A(n5201), .B(n5202), .Z(n5183) );
  XNOR U5243 ( .A(n5193), .B(n5206), .Z(n5197) );
  XNOR U5244 ( .A(n5194), .B(n5195), .Z(n5206) );
  ANDN U5245 ( .A(n3025), .B(n651), .Z(n5194) );
  XOR U5246 ( .A(n5190), .B(n5207), .Z(n5193) );
  ANDN U5247 ( .A(n692), .B(n3027), .Z(n5207) );
  XNOR U5248 ( .A(n5212), .B(n5204), .Z(n5153) );
  XNOR U5249 ( .A(n5203), .B(n5213), .Z(n5204) );
  ANDN U5250 ( .A(n799), .B(n2886), .Z(n5213) );
  XNOR U5251 ( .A(n5216), .B(n5214), .Z(n5215) );
  ANDN U5252 ( .A(n799), .B(n3027), .Z(n5216) );
  XNOR U5253 ( .A(n5211), .B(n5205), .Z(n5212) );
  AND U5254 ( .A(n2884), .B(n745), .Z(n5205) );
  XNOR U5255 ( .A(n5209), .B(n5210), .Z(n5152) );
  NANDN U5256 ( .B(n651), .A(n3813), .Z(n5210) );
  XNOR U5257 ( .A(n5208), .B(n5221), .Z(n5209) );
  ANDN U5258 ( .A(n692), .B(n3815), .Z(n5221) );
  NAND U5259 ( .A(g_input[0]), .B(n5222), .Z(n5208) );
  NAND U5260 ( .A(n5223), .B(n651), .Z(n5222) );
  NANDN U5261 ( .B(n3818), .A(n692), .Z(n5223) );
  XNOR U5262 ( .A(n5219), .B(n5220), .Z(n5211) );
  NAND U5263 ( .A(n3813), .B(n745), .Z(n5220) );
  XNOR U5264 ( .A(n5218), .B(n5226), .Z(n5219) );
  ANDN U5265 ( .A(n799), .B(n3815), .Z(n5226) );
  NAND U5266 ( .A(g_input[0]), .B(n5227), .Z(n5218) );
  NANDN U5267 ( .B(n745), .A(n5228), .Z(n5227) );
  NANDN U5268 ( .B(n3818), .A(n799), .Z(n5228) );
  IV U5269 ( .A(n5217), .Z(n745) );
  XOR U5270 ( .A(n3024), .B(n3023), .Z(n3008) );
  XOR U5271 ( .A(n5231), .B(n3020), .Z(n3023) );
  XNOR U5272 ( .A(n3019), .B(n5232), .Z(n3020) );
  ANDN U5273 ( .A(n624), .B(n2886), .Z(n5232) );
  IV U5274 ( .A(n2752), .Z(n2886) );
  XNOR U5275 ( .A(n5201), .B(g_input[4]), .Z(n5202) );
  ANDN U5276 ( .A(n5233), .B(n5234), .Z(n5201) );
  XNOR U5277 ( .A(n5237), .B(n5235), .Z(n5236) );
  ANDN U5278 ( .A(n624), .B(n3027), .Z(n5237) );
  IV U5279 ( .A(n2884), .Z(n3027) );
  IV U5280 ( .A(n3815), .Z(n3025) );
  XNOR U5281 ( .A(n3022), .B(n3021), .Z(n5231) );
  AND U5282 ( .A(n2884), .B(n583), .Z(n3021) );
  ANDN U5283 ( .A(n5242), .B(n5243), .Z(n5233) );
  XNOR U5284 ( .A(n5240), .B(n5241), .Z(n3022) );
  NAND U5285 ( .A(n3813), .B(n583), .Z(n5241) );
  XNOR U5286 ( .A(n5239), .B(n5244), .Z(n5240) );
  ANDN U5287 ( .A(n624), .B(n3815), .Z(n5244) );
  NAND U5288 ( .A(g_input[0]), .B(n5245), .Z(n5239) );
  NANDN U5289 ( .B(n583), .A(n5246), .Z(n5245) );
  NANDN U5290 ( .B(n3818), .A(n624), .Z(n5246) );
  IV U5291 ( .A(n5238), .Z(n583) );
  XOR U5292 ( .A(n3031), .B(n3030), .Z(n3024) );
  NAND U5293 ( .A(n3813), .B(n527), .Z(n3030) );
  IV U5294 ( .A(n3818), .Z(n3813) );
  XOR U5295 ( .A(n3029), .B(n5249), .Z(n3031) );
  ANDN U5296 ( .A(n558), .B(n3815), .Z(n5249) );
  XNOR U5297 ( .A(n5242), .B(g_input[2]), .Z(n5243) );
  NOR U5298 ( .A(g_input[0]), .B(n5250), .Z(n5242) );
  NANDN U5299 ( .B(n527), .A(n5252), .Z(n5251) );
  NANDN U5300 ( .B(n3818), .A(n558), .Z(n5252) );
  XOR U5301 ( .A(g_input[0]), .B(g_input[1]), .Z(n5250) );
  AND U5302 ( .A(n5254), .B(n5253), .Z(n527) );
  ANDN U5303 ( .A(e_input[31]), .B(n5255), .Z(n5254) );
  NANDN U5304 ( .B(n5256), .A(n5248), .Z(n5255) );
  XNOR U5305 ( .A(n5256), .B(e_input[29]), .Z(n5248) );
  NAND U5306 ( .A(n5247), .B(n5257), .Z(n5256) );
  XOR U5307 ( .A(n5257), .B(e_input[28]), .Z(n5247) );
  ANDN U5308 ( .A(n5224), .B(n5258), .Z(n5257) );
  XNOR U5309 ( .A(n5258), .B(e_input[27]), .Z(n5224) );
  NAND U5310 ( .A(n5225), .B(n5259), .Z(n5258) );
  XOR U5311 ( .A(n5259), .B(e_input[26]), .Z(n5225) );
  ANDN U5312 ( .A(n5230), .B(n5260), .Z(n5259) );
  XNOR U5313 ( .A(n5260), .B(e_input[25]), .Z(n5230) );
  NAND U5314 ( .A(n5229), .B(n5261), .Z(n5260) );
  XOR U5315 ( .A(n5261), .B(e_input[24]), .Z(n5229) );
  ANDN U5316 ( .A(n4970), .B(n5262), .Z(n5261) );
  XNOR U5317 ( .A(n5262), .B(e_input[23]), .Z(n4970) );
  NAND U5318 ( .A(n4971), .B(n5263), .Z(n5262) );
  XOR U5319 ( .A(n5263), .B(e_input[22]), .Z(n4971) );
  ANDN U5320 ( .A(n4966), .B(n5264), .Z(n5263) );
  XNOR U5321 ( .A(n5264), .B(e_input[21]), .Z(n4966) );
  NAND U5322 ( .A(n4965), .B(n5265), .Z(n5264) );
  XOR U5323 ( .A(n5265), .B(e_input[20]), .Z(n4965) );
  ANDN U5324 ( .A(n5141), .B(n5266), .Z(n5265) );
  XNOR U5325 ( .A(n5266), .B(e_input[19]), .Z(n5141) );
  NAND U5326 ( .A(n5140), .B(n5267), .Z(n5266) );
  XOR U5327 ( .A(n5267), .B(e_input[18]), .Z(n5140) );
  ANDN U5328 ( .A(n5146), .B(n5268), .Z(n5267) );
  XNOR U5329 ( .A(n5268), .B(e_input[17]), .Z(n5146) );
  NAND U5330 ( .A(n5145), .B(n5269), .Z(n5268) );
  XOR U5331 ( .A(n5269), .B(e_input[16]), .Z(n5145) );
  ANDN U5332 ( .A(n3843), .B(n5270), .Z(n5269) );
  XNOR U5333 ( .A(n5270), .B(e_input[15]), .Z(n3843) );
  NAND U5334 ( .A(n3842), .B(n5271), .Z(n5270) );
  XOR U5335 ( .A(n5271), .B(e_input[14]), .Z(n3842) );
  ANDN U5336 ( .A(n3838), .B(n5272), .Z(n5271) );
  XNOR U5337 ( .A(n5272), .B(e_input[13]), .Z(n3838) );
  NAND U5338 ( .A(n3837), .B(n5273), .Z(n5272) );
  XOR U5339 ( .A(n5273), .B(e_input[12]), .Z(n3837) );
  ANDN U5340 ( .A(n3820), .B(n5274), .Z(n5273) );
  XNOR U5341 ( .A(n5274), .B(e_input[11]), .Z(n3820) );
  NAND U5342 ( .A(n3819), .B(n5275), .Z(n5274) );
  XOR U5343 ( .A(n5275), .B(e_input[10]), .Z(n3819) );
  ANDN U5344 ( .A(n3825), .B(n5276), .Z(n5275) );
  XNOR U5345 ( .A(n5276), .B(e_input[9]), .Z(n3825) );
  NAND U5346 ( .A(n3824), .B(n5277), .Z(n5276) );
  XOR U5347 ( .A(n5277), .B(e_input[8]), .Z(n3824) );
  ANDN U5348 ( .A(n4349), .B(n5278), .Z(n5277) );
  XNOR U5349 ( .A(n5278), .B(e_input[7]), .Z(n4349) );
  NAND U5350 ( .A(n4348), .B(n5279), .Z(n5278) );
  XOR U5351 ( .A(n5279), .B(e_input[6]), .Z(n4348) );
  ANDN U5352 ( .A(n4344), .B(n5280), .Z(n5279) );
  XNOR U5353 ( .A(n5280), .B(e_input[5]), .Z(n4344) );
  NAND U5354 ( .A(n4343), .B(n5281), .Z(n5280) );
  XOR U5355 ( .A(n5281), .B(e_input[4]), .Z(n4343) );
  ANDN U5356 ( .A(n4778), .B(n5282), .Z(n5281) );
  XNOR U5357 ( .A(n5282), .B(e_input[3]), .Z(n4778) );
  NAND U5358 ( .A(n4777), .B(n5283), .Z(n5282) );
  XOR U5359 ( .A(n5283), .B(e_input[2]), .Z(n4777) );
  NOR U5360 ( .A(n4782), .B(e_input[0]), .Z(n5283) );
  XOR U5361 ( .A(e_input[0]), .B(e_input[1]), .Z(n4782) );
endmodule

