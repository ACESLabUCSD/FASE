
module MxM_W8_N100 ( clk, rst, A, X, Y );
  input [7:0] A;
  input [7:0] X;
  output [7:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, \add_25/carry[6] , \add_25/carry[5] ,
         \add_25/carry[4] , \add_25/carry[3] , \add_25/carry[2] , n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554;
  wire   [7:0] Y0;
  wire   [6:0] n;

  DFF \n_reg[0]  ( .D(n133), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n132), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n131), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n130), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n129), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n128), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n127), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \Y0_reg[0]  ( .D(n126), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n125), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n124), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n123), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n122), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n121), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n120), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n119), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y_reg[7]  ( .D(n118), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n117), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n116), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n115), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n114), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n113), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n112), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n111), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  MUX U136 ( .IN0(n452), .IN1(n468), .SEL(n454), .F(n433) );
  MUX U137 ( .IN0(A[3]), .IN1(n517), .SEL(A[7]), .F(n134) );
  IV U138 ( .A(n134), .Z(n362) );
  MUX U139 ( .IN0(n402), .IN1(n400), .SEL(n401), .F(n357) );
  NAND U140 ( .A(n275), .B(n309), .Z(n308) );
  MUX U141 ( .IN0(n385), .IN1(n135), .SEL(n384), .F(n340) );
  IV U142 ( .A(n383), .Z(n135) );
  MUX U143 ( .IN0(n136), .IN1(n285), .SEL(n286), .F(n253) );
  IV U144 ( .A(Y0[3]), .Z(n136) );
  XOR U145 ( .A(n516), .B(A[3]), .Z(n517) );
  XNOR U146 ( .A(n504), .B(n505), .Z(n483) );
  MUX U147 ( .IN0(X[6]), .IN1(n542), .SEL(X[7]), .F(n251) );
  MUX U148 ( .IN0(X[3]), .IN1(n492), .SEL(X[7]), .F(n343) );
  MUX U149 ( .IN0(n346), .IN1(n137), .SEL(n347), .F(n298) );
  IV U150 ( .A(n348), .Z(n137) );
  XNOR U151 ( .A(n349), .B(n314), .Z(n306) );
  MUX U152 ( .IN0(n138), .IN1(n368), .SEL(n369), .F(n323) );
  IV U153 ( .A(Y0[1]), .Z(n138) );
  XOR U154 ( .A(n221), .B(n231), .Z(n229) );
  MUX U155 ( .IN0(n139), .IN1(n522), .SEL(n523), .F(n518) );
  IV U156 ( .A(n524), .Z(n139) );
  MUX U157 ( .IN0(A[4]), .IN1(n469), .SEL(A[7]), .F(n140) );
  IV U158 ( .A(n140), .Z(n316) );
  MUX U159 ( .IN0(A[5]), .IN1(n451), .SEL(A[7]), .F(n279) );
  XOR U160 ( .A(n365), .B(n404), .Z(n366) );
  MUX U161 ( .IN0(A[6]), .IN1(n423), .SEL(A[7]), .F(n252) );
  MUX U162 ( .IN0(n386), .IN1(n141), .SEL(n387), .F(n346) );
  IV U163 ( .A(n388), .Z(n141) );
  XNOR U164 ( .A(n268), .B(n269), .Z(n292) );
  XOR U165 ( .A(n253), .B(n263), .Z(n261) );
  NOR U166 ( .A(A[0]), .B(n539), .Z(n527) );
  MUX U167 ( .IN0(n142), .IN1(n416), .SEL(n417), .F(n463) );
  IV U168 ( .A(n483), .Z(n142) );
  MUX U169 ( .IN0(n518), .IN1(n521), .SEL(n519), .F(n394) );
  MUX U170 ( .IN0(n433), .IN1(n449), .SEL(n435), .F(n427) );
  MUX U171 ( .IN0(n278), .IN1(n302), .SEL(n277), .F(n240) );
  NAND U172 ( .A(n340), .B(n381), .Z(n380) );
  XNOR U173 ( .A(n402), .B(n401), .Z(n388) );
  XNOR U174 ( .A(n307), .B(n306), .Z(n300) );
  XNOR U175 ( .A(n361), .B(n360), .Z(n348) );
  MUX U176 ( .IN0(Y0[6]), .IN1(n203), .SEL(n198), .F(n191) );
  XOR U177 ( .A(n285), .B(n293), .Z(n291) );
  MUX U178 ( .IN0(A[2]), .IN1(n526), .SEL(A[7]), .F(n403) );
  XOR U179 ( .A(n493), .B(n474), .Z(n417) );
  XNOR U180 ( .A(n392), .B(n354), .Z(n360) );
  MUX U181 ( .IN0(n391), .IN1(n389), .SEL(n390), .F(n143) );
  IV U182 ( .A(n143), .Z(n345) );
  AND U183 ( .A(n246), .B(n212), .Z(n245) );
  MUX U184 ( .IN0(n144), .IN1(n300), .SEL(n299), .F(n269) );
  IV U185 ( .A(n298), .Z(n144) );
  MUX U186 ( .IN0(n145), .IN1(n323), .SEL(n324), .F(n285) );
  IV U187 ( .A(Y0[2]), .Z(n145) );
  MUX U188 ( .IN0(Y0[7]), .IN1(n191), .SEL(n192), .F(n146) );
  IV U189 ( .A(n146), .Z(n188) );
  XOR U190 ( .A(n369), .B(Y0[1]), .Z(n157) );
  ANDN U191 ( .A(n147), .B(n[0]), .Z(n133) );
  AND U192 ( .A(N8), .B(n147), .Z(n132) );
  AND U193 ( .A(N9), .B(n147), .Z(n131) );
  AND U194 ( .A(N10), .B(n147), .Z(n130) );
  AND U195 ( .A(N11), .B(n147), .Z(n129) );
  AND U196 ( .A(N12), .B(n147), .Z(n128) );
  AND U197 ( .A(n147), .B(n148), .Z(n127) );
  XOR U198 ( .A(n[6]), .B(\add_25/carry[6] ), .Z(n148) );
  ANDN U199 ( .A(n149), .B(rst), .Z(n147) );
  NAND U200 ( .A(n150), .B(n151), .Z(n149) );
  AND U201 ( .A(n[0]), .B(n152), .Z(n151) );
  NOR U202 ( .A(n153), .B(n[2]), .Z(n152) );
  AND U203 ( .A(n154), .B(n[6]), .Z(n150) );
  AND U204 ( .A(n[5]), .B(n[1]), .Z(n154) );
  NAND U205 ( .A(n155), .B(n156), .Z(n126) );
  OR U206 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U207 ( .B(n159), .A(Y0[0]), .Z(n155) );
  NAND U208 ( .A(n160), .B(n161), .Z(n125) );
  NANDN U209 ( .B(n158), .A(n162), .Z(n161) );
  NANDN U210 ( .B(n163), .A(rst), .Z(n160) );
  NAND U211 ( .A(n164), .B(n165), .Z(n124) );
  NANDN U212 ( .B(n158), .A(n166), .Z(n165) );
  NANDN U213 ( .B(n159), .A(Y0[2]), .Z(n164) );
  NAND U214 ( .A(n167), .B(n168), .Z(n123) );
  NANDN U215 ( .B(n158), .A(n169), .Z(n168) );
  NANDN U216 ( .B(n159), .A(Y0[3]), .Z(n167) );
  NAND U217 ( .A(n170), .B(n171), .Z(n122) );
  NANDN U218 ( .B(n158), .A(n172), .Z(n171) );
  NANDN U219 ( .B(n159), .A(Y0[4]), .Z(n170) );
  NAND U220 ( .A(n173), .B(n174), .Z(n121) );
  NANDN U221 ( .B(n158), .A(n175), .Z(n174) );
  NANDN U222 ( .B(n159), .A(Y0[5]), .Z(n173) );
  NAND U223 ( .A(n176), .B(n177), .Z(n120) );
  OR U224 ( .A(n178), .B(n158), .Z(n177) );
  NANDN U225 ( .B(n159), .A(Y0[6]), .Z(n176) );
  NAND U226 ( .A(n179), .B(n180), .Z(n119) );
  OR U227 ( .A(n158), .B(n181), .Z(n180) );
  NANDN U228 ( .B(n182), .A(n159), .Z(n158) );
  NANDN U229 ( .B(n159), .A(Y0[7]), .Z(n179) );
  NAND U230 ( .A(n183), .B(n184), .Z(n118) );
  NANDN U231 ( .B(n159), .A(Y[7]), .Z(n184) );
  AND U232 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U233 ( .B(n182), .A(Y[7]), .Z(n186) );
  OR U234 ( .A(n181), .B(n187), .Z(n185) );
  XOR U235 ( .A(n188), .B(n189), .Z(n181) );
  XNOR U236 ( .A(Y0[7]), .B(n190), .Z(n189) );
  NAND U237 ( .A(n193), .B(n194), .Z(n117) );
  NANDN U238 ( .B(n159), .A(Y[6]), .Z(n194) );
  AND U239 ( .A(n195), .B(n196), .Z(n193) );
  NANDN U240 ( .B(n182), .A(Y[6]), .Z(n196) );
  OR U241 ( .A(n178), .B(n187), .Z(n195) );
  XOR U242 ( .A(n192), .B(Y0[7]), .Z(n178) );
  XOR U243 ( .A(n191), .B(n190), .Z(n192) );
  NAND U244 ( .A(n199), .B(n200), .Z(n116) );
  NANDN U245 ( .B(n159), .A(Y[5]), .Z(n200) );
  AND U246 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U247 ( .B(n182), .A(Y[5]), .Z(n202) );
  NANDN U248 ( .B(n187), .A(n175), .Z(n201) );
  XNOR U249 ( .A(n198), .B(Y0[6]), .Z(n175) );
  XOR U250 ( .A(n203), .B(n204), .Z(n198) );
  ANDN U251 ( .A(n190), .B(n205), .Z(n204) );
  NANDN U252 ( .B(n206), .A(n207), .Z(n190) );
  ANDN U253 ( .A(n208), .B(n205), .Z(n206) );
  NAND U254 ( .A(n209), .B(n210), .Z(n205) );
  OR U255 ( .A(n211), .B(n212), .Z(n210) );
  AND U256 ( .A(n213), .B(n214), .Z(n209) );
  OR U257 ( .A(n215), .B(n216), .Z(n214) );
  OR U258 ( .A(n217), .B(n218), .Z(n213) );
  NOR U259 ( .A(n219), .B(n220), .Z(n208) );
  IV U260 ( .A(n197), .Z(n203) );
  XOR U261 ( .A(n221), .B(n222), .Z(n197) );
  ANDN U262 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U263 ( .A(Y0[5]), .B(n221), .Z(n223) );
  NAND U264 ( .A(n225), .B(n226), .Z(n115) );
  NANDN U265 ( .B(n159), .A(Y[4]), .Z(n226) );
  AND U266 ( .A(n227), .B(n228), .Z(n225) );
  NANDN U267 ( .B(n182), .A(Y[4]), .Z(n228) );
  NANDN U268 ( .B(n187), .A(n172), .Z(n227) );
  XNOR U269 ( .A(n224), .B(Y0[5]), .Z(n172) );
  XNOR U270 ( .A(n229), .B(n230), .Z(n224) );
  AND U271 ( .A(n207), .B(n232), .Z(n231) );
  XOR U272 ( .A(n219), .B(n233), .Z(n232) );
  XOR U273 ( .A(n233), .B(n220), .Z(n219) );
  OR U274 ( .A(n234), .B(n235), .Z(n220) );
  IV U275 ( .A(n230), .Z(n233) );
  XNOR U276 ( .A(n218), .B(n217), .Z(n230) );
  OR U277 ( .A(n236), .B(n237), .Z(n217) );
  AND U278 ( .A(n238), .B(n239), .Z(n218) );
  XNOR U279 ( .A(n240), .B(n241), .Z(n239) );
  ANDN U280 ( .A(n242), .B(n243), .Z(n241) );
  XOR U281 ( .A(n240), .B(n244), .Z(n242) );
  XNOR U282 ( .A(n211), .B(n245), .Z(n238) );
  NAND U283 ( .A(n247), .B(n248), .Z(n212) );
  NANDN U284 ( .B(n249), .A(n250), .Z(n247) );
  NANDN U285 ( .B(n215), .A(n251), .Z(n246) );
  NANDN U286 ( .B(n216), .A(n252), .Z(n211) );
  XOR U287 ( .A(n253), .B(n254), .Z(n221) );
  ANDN U288 ( .A(n255), .B(n256), .Z(n254) );
  XNOR U289 ( .A(Y0[4]), .B(n253), .Z(n255) );
  NAND U290 ( .A(n257), .B(n258), .Z(n114) );
  NANDN U291 ( .B(n159), .A(Y[3]), .Z(n258) );
  AND U292 ( .A(n259), .B(n260), .Z(n257) );
  NANDN U293 ( .B(n182), .A(Y[3]), .Z(n260) );
  NANDN U294 ( .B(n187), .A(n169), .Z(n259) );
  XNOR U295 ( .A(n256), .B(Y0[4]), .Z(n169) );
  XNOR U296 ( .A(n261), .B(n262), .Z(n256) );
  AND U297 ( .A(n207), .B(n264), .Z(n263) );
  XOR U298 ( .A(n234), .B(n265), .Z(n264) );
  XOR U299 ( .A(n265), .B(n235), .Z(n234) );
  OR U300 ( .A(n266), .B(n267), .Z(n235) );
  IV U301 ( .A(n262), .Z(n265) );
  XNOR U302 ( .A(n237), .B(n236), .Z(n262) );
  OR U303 ( .A(n268), .B(n269), .Z(n236) );
  XOR U304 ( .A(n244), .B(n243), .Z(n237) );
  XOR U305 ( .A(n240), .B(n270), .Z(n243) );
  AND U306 ( .A(n271), .B(n272), .Z(n270) );
  NANDN U307 ( .B(n215), .A(n273), .Z(n272) );
  OR U308 ( .A(n274), .B(n275), .Z(n271) );
  XOR U309 ( .A(n249), .B(n250), .Z(n244) );
  NANDN U310 ( .B(n216), .A(n279), .Z(n250) );
  XNOR U311 ( .A(n248), .B(n280), .Z(n249) );
  AND U312 ( .A(n252), .B(n251), .Z(n280) );
  ANDN U313 ( .A(n281), .B(n282), .Z(n248) );
  NANDN U314 ( .B(n283), .A(n284), .Z(n281) );
  NAND U315 ( .A(n287), .B(n288), .Z(n113) );
  NANDN U316 ( .B(n159), .A(Y[2]), .Z(n288) );
  AND U317 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U318 ( .B(n182), .A(Y[2]), .Z(n290) );
  NANDN U319 ( .B(n187), .A(n166), .Z(n289) );
  XNOR U320 ( .A(n286), .B(Y0[3]), .Z(n166) );
  XNOR U321 ( .A(n291), .B(n292), .Z(n286) );
  AND U322 ( .A(n207), .B(n294), .Z(n293) );
  XOR U323 ( .A(n266), .B(n295), .Z(n294) );
  XOR U324 ( .A(n295), .B(n267), .Z(n266) );
  OR U325 ( .A(n296), .B(n297), .Z(n267) );
  IV U326 ( .A(n292), .Z(n295) );
  XOR U327 ( .A(n278), .B(n277), .Z(n268) );
  XNOR U328 ( .A(n301), .B(n302), .Z(n277) );
  IV U329 ( .A(n276), .Z(n302) );
  XOR U330 ( .A(n303), .B(n304), .Z(n276) );
  ANDN U331 ( .A(n305), .B(n306), .Z(n304) );
  XOR U332 ( .A(n303), .B(n307), .Z(n305) );
  XNOR U333 ( .A(n308), .B(n274), .Z(n301) );
  NAND U334 ( .A(n273), .B(n252), .Z(n274) );
  NANDN U335 ( .B(n215), .A(n310), .Z(n309) );
  XNOR U336 ( .A(n311), .B(n312), .Z(n275) );
  ANDN U337 ( .A(n313), .B(n314), .Z(n312) );
  XNOR U338 ( .A(n315), .B(n311), .Z(n313) );
  XOR U339 ( .A(n283), .B(n284), .Z(n278) );
  OR U340 ( .A(n316), .B(n216), .Z(n284) );
  XNOR U341 ( .A(n317), .B(n318), .Z(n283) );
  AND U342 ( .A(n279), .B(n251), .Z(n318) );
  IV U343 ( .A(n282), .Z(n317) );
  NAND U344 ( .A(n319), .B(n320), .Z(n282) );
  NANDN U345 ( .B(n321), .A(n322), .Z(n319) );
  NAND U346 ( .A(n325), .B(n326), .Z(n112) );
  NANDN U347 ( .B(n159), .A(Y[1]), .Z(n326) );
  AND U348 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U349 ( .B(n182), .A(Y[1]), .Z(n328) );
  NANDN U350 ( .B(n187), .A(n162), .Z(n327) );
  XNOR U351 ( .A(n324), .B(Y0[2]), .Z(n162) );
  XNOR U352 ( .A(n329), .B(n330), .Z(n324) );
  XOR U353 ( .A(n323), .B(n331), .Z(n329) );
  AND U354 ( .A(n207), .B(n332), .Z(n331) );
  XOR U355 ( .A(n296), .B(n333), .Z(n332) );
  XOR U356 ( .A(n333), .B(n297), .Z(n296) );
  NANDN U357 ( .B(n334), .A(n335), .Z(n297) );
  IV U358 ( .A(n330), .Z(n333) );
  XOR U359 ( .A(n300), .B(n299), .Z(n330) );
  XNOR U360 ( .A(n298), .B(n336), .Z(n299) );
  AND U361 ( .A(n337), .B(n338), .Z(n336) );
  OR U362 ( .A(n339), .B(n340), .Z(n338) );
  AND U363 ( .A(n341), .B(n342), .Z(n337) );
  NANDN U364 ( .B(n215), .A(n343), .Z(n342) );
  NAND U365 ( .A(n344), .B(n345), .Z(n341) );
  XNOR U366 ( .A(n311), .B(n350), .Z(n314) );
  AND U367 ( .A(n252), .B(n310), .Z(n350) );
  XOR U368 ( .A(n351), .B(n352), .Z(n311) );
  ANDN U369 ( .A(n353), .B(n354), .Z(n352) );
  XNOR U370 ( .A(n355), .B(n351), .Z(n353) );
  XOR U371 ( .A(n356), .B(n315), .Z(n349) );
  NAND U372 ( .A(n273), .B(n279), .Z(n315) );
  IV U373 ( .A(n303), .Z(n356) );
  XOR U374 ( .A(n357), .B(n358), .Z(n303) );
  ANDN U375 ( .A(n359), .B(n360), .Z(n358) );
  XOR U376 ( .A(n357), .B(n361), .Z(n359) );
  XNOR U377 ( .A(n321), .B(n322), .Z(n307) );
  OR U378 ( .A(n362), .B(n216), .Z(n322) );
  XNOR U379 ( .A(n320), .B(n363), .Z(n321) );
  ANDN U380 ( .A(n251), .B(n316), .Z(n363) );
  ANDN U381 ( .A(n364), .B(n365), .Z(n320) );
  NANDN U382 ( .B(n366), .A(n367), .Z(n364) );
  NAND U383 ( .A(n370), .B(n371), .Z(n111) );
  NANDN U384 ( .B(n159), .A(Y[0]), .Z(n371) );
  AND U385 ( .A(n372), .B(n373), .Z(n370) );
  NANDN U386 ( .B(n182), .A(Y[0]), .Z(n373) );
  IV U387 ( .A(n374), .Z(n182) );
  OR U388 ( .A(n187), .B(n157), .Z(n372) );
  IV U389 ( .A(Y0[1]), .Z(n163) );
  XOR U390 ( .A(n375), .B(n376), .Z(n369) );
  XNOR U391 ( .A(n377), .B(n368), .Z(n375) );
  NAND U392 ( .A(Y0[0]), .B(n334), .Z(n368) );
  NAND U393 ( .A(n378), .B(n207), .Z(n377) );
  XOR U394 ( .A(A[7]), .B(X[7]), .Z(n207) );
  XNOR U395 ( .A(n335), .B(n376), .Z(n378) );
  XNOR U396 ( .A(n334), .B(n376), .Z(n335) );
  XNOR U397 ( .A(n348), .B(n347), .Z(n376) );
  XNOR U398 ( .A(n379), .B(n344), .Z(n347) );
  XNOR U399 ( .A(n380), .B(n339), .Z(n344) );
  NAND U400 ( .A(n252), .B(n343), .Z(n339) );
  NANDN U401 ( .B(n215), .A(n382), .Z(n381) );
  XNOR U402 ( .A(n345), .B(n346), .Z(n379) );
  XNOR U403 ( .A(n351), .B(n393), .Z(n354) );
  AND U404 ( .A(n279), .B(n310), .Z(n393) );
  XOR U405 ( .A(n394), .B(n395), .Z(n351) );
  ANDN U406 ( .A(n396), .B(n397), .Z(n395) );
  XNOR U407 ( .A(n398), .B(n394), .Z(n396) );
  XOR U408 ( .A(n399), .B(n355), .Z(n392) );
  NANDN U409 ( .B(n316), .A(n273), .Z(n355) );
  IV U410 ( .A(n357), .Z(n399) );
  XNOR U411 ( .A(n366), .B(n367), .Z(n361) );
  NANDN U412 ( .B(n216), .A(n403), .Z(n367) );
  ANDN U413 ( .A(n251), .B(n362), .Z(n404) );
  NAND U414 ( .A(n405), .B(n406), .Z(n365) );
  NANDN U415 ( .B(n407), .A(n408), .Z(n405) );
  XNOR U416 ( .A(n388), .B(n387), .Z(n334) );
  XNOR U417 ( .A(n409), .B(n391), .Z(n387) );
  XNOR U418 ( .A(n384), .B(n385), .Z(n391) );
  NAND U419 ( .A(n279), .B(n343), .Z(n385) );
  XNOR U420 ( .A(n383), .B(n410), .Z(n384) );
  AND U421 ( .A(n382), .B(n252), .Z(n410) );
  XOR U422 ( .A(n411), .B(n412), .Z(n383) );
  AND U423 ( .A(n413), .B(n414), .Z(n412) );
  XNOR U424 ( .A(n415), .B(n411), .Z(n414) );
  XNOR U425 ( .A(n390), .B(n386), .Z(n409) );
  XOR U426 ( .A(n416), .B(n417), .Z(n386) );
  XOR U427 ( .A(n418), .B(n419), .Z(n390) );
  AND U428 ( .A(n420), .B(n421), .Z(n419) );
  NANDN U429 ( .B(n215), .A(n422), .Z(n421) );
  NANDN U430 ( .B(n423), .A(n424), .Z(n215) );
  AND U431 ( .A(n425), .B(A[7]), .Z(n424) );
  NANDN U432 ( .B(n426), .A(n427), .Z(n420) );
  IV U433 ( .A(n389), .Z(n418) );
  XNOR U434 ( .A(n428), .B(n429), .Z(n389) );
  AND U435 ( .A(n430), .B(n431), .Z(n429) );
  XOR U436 ( .A(n427), .B(n432), .Z(n431) );
  XNOR U437 ( .A(n426), .B(n428), .Z(n432) );
  NAND U438 ( .A(n252), .B(n422), .Z(n426) );
  XNOR U439 ( .A(n436), .B(n433), .Z(n435) );
  XOR U440 ( .A(n413), .B(n437), .Z(n430) );
  XNOR U441 ( .A(n415), .B(n428), .Z(n437) );
  NANDN U442 ( .B(n316), .A(n343), .Z(n415) );
  XOR U443 ( .A(n411), .B(n438), .Z(n413) );
  AND U444 ( .A(n382), .B(n279), .Z(n438) );
  XOR U445 ( .A(n439), .B(n440), .Z(n411) );
  AND U446 ( .A(n441), .B(n442), .Z(n440) );
  XNOR U447 ( .A(n443), .B(n439), .Z(n442) );
  XOR U448 ( .A(n444), .B(n445), .Z(n428) );
  AND U449 ( .A(n446), .B(n447), .Z(n445) );
  XOR U450 ( .A(n434), .B(n448), .Z(n447) );
  XNOR U451 ( .A(n436), .B(n444), .Z(n448) );
  NAND U452 ( .A(n279), .B(n422), .Z(n436) );
  XOR U453 ( .A(n433), .B(n449), .Z(n434) );
  AND U454 ( .A(n252), .B(X[0]), .Z(n449) );
  XNOR U455 ( .A(n425), .B(A[6]), .Z(n423) );
  NOR U456 ( .A(n450), .B(n451), .Z(n425) );
  XNOR U457 ( .A(n455), .B(n452), .Z(n454) );
  XOR U458 ( .A(n441), .B(n456), .Z(n446) );
  XNOR U459 ( .A(n443), .B(n444), .Z(n456) );
  NANDN U460 ( .B(n362), .A(n343), .Z(n443) );
  XOR U461 ( .A(n439), .B(n457), .Z(n441) );
  ANDN U462 ( .A(n382), .B(n316), .Z(n457) );
  XOR U463 ( .A(n458), .B(n459), .Z(n439) );
  AND U464 ( .A(n460), .B(n461), .Z(n459) );
  XNOR U465 ( .A(n462), .B(n458), .Z(n461) );
  XOR U466 ( .A(n463), .B(n464), .Z(n444) );
  AND U467 ( .A(n465), .B(n466), .Z(n464) );
  XOR U468 ( .A(n453), .B(n467), .Z(n466) );
  XNOR U469 ( .A(n455), .B(n463), .Z(n467) );
  NANDN U470 ( .B(n316), .A(n422), .Z(n455) );
  XOR U471 ( .A(n452), .B(n468), .Z(n453) );
  AND U472 ( .A(n279), .B(X[0]), .Z(n468) );
  XOR U473 ( .A(n450), .B(A[5]), .Z(n451) );
  NANDN U474 ( .B(n469), .A(n470), .Z(n450) );
  XOR U475 ( .A(n471), .B(n472), .Z(n452) );
  ANDN U476 ( .A(n473), .B(n474), .Z(n472) );
  XNOR U477 ( .A(n475), .B(n471), .Z(n473) );
  XOR U478 ( .A(n460), .B(n476), .Z(n465) );
  XNOR U479 ( .A(n462), .B(n463), .Z(n476) );
  NAND U480 ( .A(n343), .B(n403), .Z(n462) );
  XOR U481 ( .A(n458), .B(n477), .Z(n460) );
  ANDN U482 ( .A(n382), .B(n362), .Z(n477) );
  XOR U483 ( .A(n478), .B(n479), .Z(n458) );
  ANDN U484 ( .A(n480), .B(n481), .Z(n479) );
  XNOR U485 ( .A(n482), .B(n478), .Z(n480) );
  XNOR U486 ( .A(n484), .B(n482), .Z(n416) );
  NAND U487 ( .A(n343), .B(n485), .Z(n482) );
  IV U488 ( .A(n481), .Z(n484) );
  XNOR U489 ( .A(n478), .B(n486), .Z(n481) );
  AND U490 ( .A(n403), .B(n382), .Z(n486) );
  AND U491 ( .A(n487), .B(A[0]), .Z(n478) );
  NANDN U492 ( .B(n343), .A(n488), .Z(n487) );
  NAND U493 ( .A(n485), .B(n382), .Z(n488) );
  XNOR U494 ( .A(n489), .B(X[2]), .Z(n382) );
  NAND U495 ( .A(n490), .B(X[7]), .Z(n489) );
  XOR U496 ( .A(n491), .B(X[2]), .Z(n490) );
  XNOR U497 ( .A(n471), .B(n494), .Z(n474) );
  ANDN U498 ( .A(X[0]), .B(n316), .Z(n494) );
  XOR U499 ( .A(n495), .B(n496), .Z(n471) );
  AND U500 ( .A(n497), .B(n498), .Z(n496) );
  XOR U501 ( .A(n499), .B(n495), .Z(n498) );
  ANDN U502 ( .A(X[0]), .B(n362), .Z(n499) );
  XOR U503 ( .A(n500), .B(n495), .Z(n497) );
  AND U504 ( .A(n422), .B(n403), .Z(n500) );
  XOR U505 ( .A(n501), .B(n502), .Z(n495) );
  ANDN U506 ( .A(n503), .B(n504), .Z(n502) );
  XNOR U507 ( .A(n505), .B(n501), .Z(n503) );
  XOR U508 ( .A(n506), .B(n475), .Z(n493) );
  NANDN U509 ( .B(n362), .A(n422), .Z(n475) );
  IV U510 ( .A(n483), .Z(n506) );
  NAND U511 ( .A(n422), .B(n485), .Z(n505) );
  XNOR U512 ( .A(n501), .B(n507), .Z(n504) );
  AND U513 ( .A(n403), .B(X[0]), .Z(n507) );
  AND U514 ( .A(n508), .B(A[0]), .Z(n501) );
  NANDN U515 ( .B(n422), .A(n509), .Z(n508) );
  NAND U516 ( .A(n485), .B(X[0]), .Z(n509) );
  XNOR U517 ( .A(n510), .B(X[1]), .Z(n422) );
  NAND U518 ( .A(n511), .B(X[7]), .Z(n510) );
  XNOR U519 ( .A(X[1]), .B(n512), .Z(n511) );
  XOR U520 ( .A(n513), .B(n514), .Z(n401) );
  IV U521 ( .A(n397), .Z(n514) );
  XNOR U522 ( .A(n394), .B(n515), .Z(n397) );
  ANDN U523 ( .A(n310), .B(n316), .Z(n515) );
  XNOR U524 ( .A(n470), .B(A[4]), .Z(n469) );
  NOR U525 ( .A(n516), .B(n517), .Z(n470) );
  XOR U526 ( .A(n520), .B(n518), .Z(n519) );
  ANDN U527 ( .A(n310), .B(n362), .Z(n520) );
  AND U528 ( .A(n403), .B(n273), .Z(n521) );
  XOR U529 ( .A(n525), .B(n398), .Z(n513) );
  NANDN U530 ( .B(n362), .A(n273), .Z(n398) );
  NANDN U531 ( .B(n526), .A(n527), .Z(n516) );
  IV U532 ( .A(n400), .Z(n525) );
  XOR U533 ( .A(n528), .B(n524), .Z(n400) );
  NAND U534 ( .A(n273), .B(n485), .Z(n524) );
  IV U535 ( .A(n523), .Z(n528) );
  XNOR U536 ( .A(n522), .B(n529), .Z(n523) );
  AND U537 ( .A(n403), .B(n310), .Z(n529) );
  AND U538 ( .A(n530), .B(A[0]), .Z(n522) );
  NANDN U539 ( .B(n273), .A(n531), .Z(n530) );
  NAND U540 ( .A(n485), .B(n310), .Z(n531) );
  XNOR U541 ( .A(n532), .B(X[4]), .Z(n310) );
  NAND U542 ( .A(n533), .B(X[7]), .Z(n532) );
  XOR U543 ( .A(n534), .B(X[4]), .Z(n533) );
  XNOR U544 ( .A(n535), .B(X[5]), .Z(n273) );
  NAND U545 ( .A(n536), .B(X[7]), .Z(n535) );
  XOR U546 ( .A(n537), .B(X[5]), .Z(n536) );
  XNOR U547 ( .A(n407), .B(n408), .Z(n402) );
  NANDN U548 ( .B(n216), .A(n485), .Z(n408) );
  XNOR U549 ( .A(n406), .B(n538), .Z(n407) );
  AND U550 ( .A(n403), .B(n251), .Z(n538) );
  XNOR U551 ( .A(n527), .B(A[2]), .Z(n526) );
  AND U552 ( .A(n540), .B(A[0]), .Z(n406) );
  NAND U553 ( .A(n541), .B(n216), .Z(n540) );
  NANDN U554 ( .B(n542), .A(n543), .Z(n216) );
  ANDN U555 ( .A(X[7]), .B(n544), .Z(n543) );
  NAND U556 ( .A(n485), .B(n251), .Z(n541) );
  XOR U557 ( .A(n544), .B(X[6]), .Z(n542) );
  OR U558 ( .A(n537), .B(n545), .Z(n544) );
  XOR U559 ( .A(n545), .B(X[5]), .Z(n537) );
  OR U560 ( .A(n534), .B(n546), .Z(n545) );
  XOR U561 ( .A(n546), .B(X[4]), .Z(n534) );
  OR U562 ( .A(n492), .B(n547), .Z(n546) );
  XOR U563 ( .A(n547), .B(X[3]), .Z(n492) );
  OR U564 ( .A(n491), .B(n548), .Z(n547) );
  XOR U565 ( .A(n548), .B(X[2]), .Z(n491) );
  NANDN U566 ( .B(X[0]), .A(n512), .Z(n548) );
  XNOR U567 ( .A(X[0]), .B(X[1]), .Z(n512) );
  XNOR U568 ( .A(n549), .B(A[1]), .Z(n485) );
  NAND U569 ( .A(n550), .B(A[7]), .Z(n549) );
  XOR U570 ( .A(A[1]), .B(n539), .Z(n550) );
  XOR U571 ( .A(A[0]), .B(A[1]), .Z(n539) );
  NANDN U572 ( .B(n374), .A(n159), .Z(n187) );
  IV U573 ( .A(rst), .Z(n159) );
  NAND U574 ( .A(n551), .B(n552), .Z(n374) );
  ANDN U575 ( .A(n553), .B(n[2]), .Z(n552) );
  NOR U576 ( .A(n[6]), .B(n[5]), .Z(n553) );
  ANDN U577 ( .A(n554), .B(n153), .Z(n551) );
  OR U578 ( .A(n[4]), .B(n[3]), .Z(n153) );
  NOR U579 ( .A(n[0]), .B(n[1]), .Z(n554) );
endmodule

