
module MxM_TG_W32_N1000 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MxM/n177 , \_MxM/n174 , \_MxM/n171 , \_MxM/n168 , \_MxM/n165 ,
         \_MxM/n162 , \_MxM/n159 , \_MxM/n156 , \_MxM/n153 , \_MxM/n150 ,
         \_MxM/n147 , \_MxM/n144 , \_MxM/n141 , \_MxM/n138 , \_MxM/n135 ,
         \_MxM/n132 , \_MxM/n129 , \_MxM/n126 , \_MxM/n123 , \_MxM/n120 ,
         \_MxM/n117 , \_MxM/n114 , \_MxM/n111 , \_MxM/n108 , \_MxM/n105 ,
         \_MxM/n102 , \_MxM/n99 , \_MxM/n96 , \_MxM/n93 , \_MxM/n90 ,
         \_MxM/n87 , \_MxM/n84 , \_MxM/N23 , \_MxM/N22 , \_MxM/N21 ,
         \_MxM/N20 , \_MxM/N19 , \_MxM/N18 , \_MxM/N17 , \_MxM/N16 ,
         \_MxM/N15 , \_MxM/N14 , \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 ,
         \_MxM/N8 , \_MxM/N7 , \_MxM/N6 , \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/Y1[0] , \_MxM/Y1[1] ,
         \_MxM/Y1[2] , \_MxM/Y1[3] , \_MxM/Y1[4] , \_MxM/Y1[5] , \_MxM/Y1[6] ,
         \_MxM/Y1[7] , \_MxM/Y1[8] , \_MxM/Y1[9] , \_MxM/Y1[10] ,
         \_MxM/Y1[11] , \_MxM/Y1[12] , \_MxM/Y1[13] , \_MxM/Y1[14] ,
         \_MxM/Y1[15] , \_MxM/Y1[16] , \_MxM/Y1[17] , \_MxM/Y1[18] ,
         \_MxM/Y1[19] , \_MxM/Y1[20] , \_MxM/Y1[21] , \_MxM/Y1[22] ,
         \_MxM/Y1[23] , \_MxM/Y1[24] , \_MxM/Y1[25] , \_MxM/Y1[26] ,
         \_MxM/Y1[27] , \_MxM/Y1[28] , \_MxM/Y1[29] , \_MxM/Y1[30] ,
         \_MxM/Y1[31] , \_MxM/Y0[31] , \_MxM/Y0[30] , \_MxM/Y0[29] ,
         \_MxM/Y0[28] , \_MxM/Y0[27] , \_MxM/Y0[26] , \_MxM/Y0[25] ,
         \_MxM/Y0[24] , \_MxM/Y0[23] , \_MxM/Y0[22] , \_MxM/Y0[21] ,
         \_MxM/Y0[20] , \_MxM/Y0[19] , \_MxM/Y0[18] , \_MxM/Y0[17] ,
         \_MxM/Y0[16] , \_MxM/Y0[15] , \_MxM/Y0[14] , \_MxM/Y0[13] ,
         \_MxM/Y0[12] , \_MxM/Y0[11] , \_MxM/Y0[10] , \_MxM/Y0[9] ,
         \_MxM/Y0[8] , \_MxM/Y0[7] , \_MxM/Y0[6] , \_MxM/Y0[5] , \_MxM/Y0[4] ,
         \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] , \_MxM/Y0[0] ,
         \_MxM/add_43/carry[9] , \_MxM/add_43/carry[8] ,
         \_MxM/add_43/carry[7] , \_MxM/add_43/carry[6] ,
         \_MxM/add_43/carry[5] , \_MxM/add_43/carry[4] ,
         \_MxM/add_43/carry[3] , \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222;

  DFF \_MxM/Y_reg[31]  ( .D(\_MxM/n84 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[31]) );
  DFF \_MxM/Y0_reg[31]  ( .D(\_MxM/Y1[31] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[31] ) );
  DFF \_MxM/Y_reg[30]  ( .D(\_MxM/n87 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[30]) );
  DFF \_MxM/Y0_reg[30]  ( .D(\_MxM/Y1[30] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[30] ) );
  DFF \_MxM/Y_reg[29]  ( .D(\_MxM/n90 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[29]) );
  DFF \_MxM/Y0_reg[29]  ( .D(\_MxM/Y1[29] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[29] ) );
  DFF \_MxM/Y_reg[28]  ( .D(\_MxM/n93 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[28]) );
  DFF \_MxM/Y0_reg[28]  ( .D(\_MxM/Y1[28] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[28] ) );
  DFF \_MxM/Y_reg[27]  ( .D(\_MxM/n96 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[27]) );
  DFF \_MxM/Y0_reg[27]  ( .D(\_MxM/Y1[27] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[27] ) );
  DFF \_MxM/Y_reg[26]  ( .D(\_MxM/n99 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[26]) );
  DFF \_MxM/Y0_reg[26]  ( .D(\_MxM/Y1[26] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[26] ) );
  DFF \_MxM/Y_reg[25]  ( .D(\_MxM/n102 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[25]) );
  DFF \_MxM/Y0_reg[25]  ( .D(\_MxM/Y1[25] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[25] ) );
  DFF \_MxM/Y_reg[24]  ( .D(\_MxM/n105 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[24]) );
  DFF \_MxM/Y0_reg[24]  ( .D(\_MxM/Y1[24] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[24] ) );
  DFF \_MxM/Y_reg[23]  ( .D(\_MxM/n108 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[23]) );
  DFF \_MxM/Y0_reg[23]  ( .D(\_MxM/Y1[23] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[23] ) );
  DFF \_MxM/Y_reg[22]  ( .D(\_MxM/n111 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[22]) );
  DFF \_MxM/Y0_reg[22]  ( .D(\_MxM/Y1[22] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[22] ) );
  DFF \_MxM/Y_reg[21]  ( .D(\_MxM/n114 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[21]) );
  DFF \_MxM/Y0_reg[21]  ( .D(\_MxM/Y1[21] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[21] ) );
  DFF \_MxM/Y_reg[20]  ( .D(\_MxM/n117 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[20]) );
  DFF \_MxM/Y0_reg[20]  ( .D(\_MxM/Y1[20] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[20] ) );
  DFF \_MxM/Y_reg[19]  ( .D(\_MxM/n120 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[19]) );
  DFF \_MxM/Y0_reg[19]  ( .D(\_MxM/Y1[19] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[19] ) );
  DFF \_MxM/Y_reg[18]  ( .D(\_MxM/n123 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[18]) );
  DFF \_MxM/Y0_reg[18]  ( .D(\_MxM/Y1[18] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[18] ) );
  DFF \_MxM/Y_reg[17]  ( .D(\_MxM/n126 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[17]) );
  DFF \_MxM/Y0_reg[17]  ( .D(\_MxM/Y1[17] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[17] ) );
  DFF \_MxM/Y_reg[16]  ( .D(\_MxM/n129 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[16]) );
  DFF \_MxM/Y0_reg[16]  ( .D(\_MxM/Y1[16] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[16] ) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n132 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/Y1[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n135 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/Y1[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n138 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/Y1[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n141 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/Y1[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n144 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/Y1[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n147 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/Y1[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n150 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/Y1[9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n153 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/Y1[8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n156 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n159 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n162 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n165 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n168 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n171 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n174 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n177 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N14 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_43/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_43/carry[6] ), .COUT(\_MxM/add_43/carry[7] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_43/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_43/carry[7] ), .COUT(\_MxM/add_43/carry[8] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_43/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_43/carry[8] ), .COUT(\_MxM/add_43/carry[9] ), .SUM(\_MxM/N12 ) );
  XOR U1 ( .A(n4520), .B(n4512), .Z(n4122) );
  XOR U2 ( .A(n4453), .B(n4454), .Z(n4053) );
  MUX U3 ( .IN0(n4864), .IN1(n4862), .SEL(n4863), .F(n4841) );
  MUX U4 ( .IN0(n4424), .IN1(n1), .SEL(n4003), .F(n4411) );
  IV U5 ( .A(n4002), .Z(n1) );
  MUX U6 ( .IN0(n4585), .IN1(n2), .SEL(n4243), .F(n4574) );
  IV U7 ( .A(n4241), .Z(n2) );
  MUX U8 ( .IN0(n4359), .IN1(n3), .SEL(n3918), .F(n4346) );
  IV U9 ( .A(n3917), .Z(n3) );
  MUX U10 ( .IN0(n4), .IN1(n2837), .SEL(n2838), .F(n2708) );
  IV U11 ( .A(n2839), .Z(n4) );
  MUX U12 ( .IN0(n5), .IN1(n2734), .SEL(n2735), .F(n2606) );
  IV U13 ( .A(n2736), .Z(n5) );
  MUX U14 ( .IN0(n2562), .IN1(n2560), .SEL(n2561), .F(n2438) );
  MUX U15 ( .IN0(n2253), .IN1(n2251), .SEL(n2252), .F(n2138) );
  MUX U16 ( .IN0(n1591), .IN1(n1589), .SEL(n1590), .F(n1496) );
  MUX U17 ( .IN0(n1549), .IN1(n1547), .SEL(n1548), .F(n1462) );
  MUX U18 ( .IN0(n1143), .IN1(n1141), .SEL(n1142), .F(n1075) );
  MUX U19 ( .IN0(n854), .IN1(n852), .SEL(n853), .F(n815) );
  MUX U20 ( .IN0(n6), .IN1(n1356), .SEL(n1357), .F(n1287) );
  IV U21 ( .A(n1358), .Z(n6) );
  MUX U22 ( .IN0(n7), .IN1(n1225), .SEL(n1226), .F(n1159) );
  IV U23 ( .A(n1227), .Z(n7) );
  MUX U24 ( .IN0(n2552), .IN1(n2550), .SEL(n2551), .F(n2428) );
  MUX U25 ( .IN0(n8), .IN1(n1086), .SEL(n1087), .F(n1026) );
  IV U26 ( .A(n1088), .Z(n8) );
  XNOR U27 ( .A(n712), .B(n711), .Z(n709) );
  MUX U28 ( .IN0(n1668), .IN1(n9), .SEL(n1669), .F(n1579) );
  IV U29 ( .A(n1670), .Z(n9) );
  OR U30 ( .A(n833), .B(n834), .Z(n794) );
  XNOR U31 ( .A(n736), .B(n733), .Z(n732) );
  MUX U32 ( .IN0(n3764), .IN1(n3766), .SEL(n3765), .F(n3726) );
  MUX U33 ( .IN0(n4114), .IN1(n4112), .SEL(n4113), .F(n4095) );
  MUX U34 ( .IN0(n4515), .IN1(n10), .SEL(n4122), .F(n4502) );
  IV U35 ( .A(n4121), .Z(n10) );
  MUX U36 ( .IN0(n3593), .IN1(n3591), .SEL(n3592), .F(n3553) );
  XOR U37 ( .A(n4468), .B(n4460), .Z(n4054) );
  XOR U38 ( .A(n4440), .B(n4441), .Z(n4036) );
  XNOR U39 ( .A(n4038), .B(n4024), .Z(n4028) );
  MUX U40 ( .IN0(n4618), .IN1(n11), .SEL(n4303), .F(n4607) );
  IV U41 ( .A(n4302), .Z(n11) );
  MUX U42 ( .IN0(n4276), .IN1(n12), .SEL(n4277), .F(n4255) );
  IV U43 ( .A(n4278), .Z(n12) );
  MUX U44 ( .IN0(n4977), .IN1(n13), .SEL(n4850), .F(n4964) );
  IV U45 ( .A(n4848), .Z(n13) );
  MUX U46 ( .IN0(n4820), .IN1(n14), .SEL(n4821), .F(n4799) );
  IV U47 ( .A(n4822), .Z(n14) );
  MUX U48 ( .IN0(n3961), .IN1(n3959), .SEL(n3960), .F(n3942) );
  MUX U49 ( .IN0(n15), .IN1(n4570), .SEL(n4571), .F(n4559) );
  IV U50 ( .A(n4572), .Z(n15) );
  MUX U51 ( .IN0(n16), .IN1(n4209), .SEL(n4210), .F(n4188) );
  IV U52 ( .A(n4211), .Z(n16) );
  MUX U53 ( .IN0(n4398), .IN1(n17), .SEL(n3969), .F(n4385) );
  IV U54 ( .A(n3968), .Z(n17) );
  MUX U55 ( .IN0(n18), .IN1(n3921), .SEL(n3922), .F(n3904) );
  IV U56 ( .A(n3923), .Z(n18) );
  MUX U57 ( .IN0(n4925), .IN1(n19), .SEL(n4766), .F(n4912) );
  IV U58 ( .A(n4764), .Z(n19) );
  XOR U59 ( .A(n4351), .B(n4340), .Z(n3901) );
  MUX U60 ( .IN0(n20), .IN1(n2766), .SEL(n2767), .F(n2639) );
  IV U61 ( .A(n2768), .Z(n20) );
  MUX U62 ( .IN0(n21), .IN1(n2648), .SEL(n2649), .F(n2524) );
  IV U63 ( .A(n2650), .Z(n21) );
  MUX U64 ( .IN0(n22), .IN1(n2580), .SEL(n2581), .F(n2458) );
  IV U65 ( .A(n2582), .Z(n22) );
  MUX U66 ( .IN0(n23), .IN1(n1824), .SEL(n1825), .F(n1728) );
  IV U67 ( .A(n1826), .Z(n23) );
  MUX U68 ( .IN0(n24), .IN1(n1335), .SEL(n1336), .F(n1265) );
  IV U69 ( .A(n1337), .Z(n24) );
  MUX U70 ( .IN0(n25), .IN1(n1309), .SEL(n1310), .F(n1239) );
  IV U71 ( .A(n1311), .Z(n25) );
  MUX U72 ( .IN0(n3143), .IN1(n3141), .SEL(n3142), .F(n3005) );
  MUX U73 ( .IN0(n3035), .IN1(n3037), .SEL(n3036), .F(n2899) );
  MUX U74 ( .IN0(n2957), .IN1(n2955), .SEL(n2956), .F(n2817) );
  MUX U75 ( .IN0(n2910), .IN1(n2908), .SEL(n2909), .F(n2779) );
  MUX U76 ( .IN0(n2927), .IN1(n2925), .SEL(n2926), .F(n2791) );
  MUX U77 ( .IN0(n2612), .IN1(n2610), .SEL(n2611), .F(n2488) );
  MUX U78 ( .IN0(n2409), .IN1(n2407), .SEL(n2408), .F(n2292) );
  MUX U79 ( .IN0(n2201), .IN1(n2199), .SEL(n2200), .F(n2088) );
  MUX U80 ( .IN0(n2140), .IN1(n2138), .SEL(n2139), .F(n2033) );
  MUX U81 ( .IN0(n2007), .IN1(n2009), .SEL(n2008), .F(n1902) );
  MUX U82 ( .IN0(n1498), .IN1(n1496), .SEL(n1497), .F(n1412) );
  MUX U83 ( .IN0(n1515), .IN1(n1517), .SEL(n1516), .F(n26) );
  IV U84 ( .A(n26), .Z(n1436) );
  MUX U85 ( .IN0(n1538), .IN1(n1540), .SEL(n1539), .F(n1453) );
  MUX U86 ( .IN0(n1464), .IN1(n1462), .SEL(n1463), .F(n1385) );
  MUX U87 ( .IN0(n1355), .IN1(n27), .SEL(n1354), .F(n1286) );
  IV U88 ( .A(n1353), .Z(n27) );
  MUX U89 ( .IN0(n1056), .IN1(n1054), .SEL(n1055), .F(n1000) );
  MUX U90 ( .IN0(n28), .IN1(n1714), .SEL(n1715), .F(n1621) );
  IV U91 ( .A(n1716), .Z(n28) );
  MUX U92 ( .IN0(n1217), .IN1(n1215), .SEL(n1216), .F(n1151) );
  MUX U93 ( .IN0(n29), .IN1(n1159), .SEL(n1160), .F(n1098) );
  IV U94 ( .A(n1161), .Z(n29) );
  MUX U95 ( .IN0(n30), .IN1(n878), .SEL(n879), .F(n840) );
  IV U96 ( .A(n880), .Z(n30) );
  MUX U97 ( .IN0(n817), .IN1(n815), .SEL(n816), .F(n775) );
  MUX U98 ( .IN0(n2430), .IN1(n2428), .SEL(n2429), .F(n2303) );
  MUX U99 ( .IN0(n31), .IN1(n1346), .SEL(n1347), .F(n1276) );
  IV U100 ( .A(n1348), .Z(n31) );
  MUX U101 ( .IN0(n32), .IN1(n973), .SEL(n974), .F(n914) );
  IV U102 ( .A(n975), .Z(n32) );
  MUX U103 ( .IN0(n2076), .IN1(n33), .SEL(n2077), .F(n1971) );
  IV U104 ( .A(n2078), .Z(n33) );
  NANDN U105 ( .B(n1869), .A(n1870), .Z(n1769) );
  MUX U106 ( .IN0(n34), .IN1(n1581), .SEL(n1580), .F(n1486) );
  IV U107 ( .A(n1579), .Z(n34) );
  OR U108 ( .A(n708), .B(n709), .Z(n686) );
  OR U109 ( .A(n731), .B(n732), .Z(n706) );
  OR U110 ( .A(n1133), .B(n1134), .Z(n1070) );
  OR U111 ( .A(n831), .B(n832), .Z(n792) );
  MUX U112 ( .IN0(n3745), .IN1(n3743), .SEL(n3744), .F(n3705) );
  MUX U113 ( .IN0(n4131), .IN1(n4129), .SEL(n4130), .F(n4112) );
  XOR U114 ( .A(n4507), .B(n4499), .Z(n4105) );
  XOR U115 ( .A(n3720), .B(n3685), .Z(n3689) );
  XNOR U116 ( .A(n4072), .B(n4058), .Z(n4062) );
  XOR U117 ( .A(n4455), .B(n4447), .Z(n4037) );
  MUX U118 ( .IN0(n35), .IN1(n3494), .SEL(n3495), .F(n3456) );
  IV U119 ( .A(n3496), .Z(n35) );
  XNOR U120 ( .A(n3509), .B(n3474), .Z(n3478) );
  MUX U121 ( .IN0(n4012), .IN1(n4010), .SEL(n4011), .F(n3993) );
  MUX U122 ( .IN0(n36), .IN1(n4598), .SEL(n4599), .F(n4587) );
  IV U123 ( .A(n4600), .Z(n36) );
  MUX U124 ( .IN0(n4299), .IN1(n4297), .SEL(n4298), .F(n4276) );
  MUX U125 ( .IN0(n37), .IN1(n4837), .SEL(n4838), .F(n4816) );
  IV U126 ( .A(n4839), .Z(n37) );
  XNOR U127 ( .A(n3395), .B(n3360), .Z(n3364) );
  XOR U128 ( .A(n4403), .B(n4395), .Z(n3969) );
  MUX U129 ( .IN0(n4964), .IN1(n38), .SEL(n4829), .F(n4951) );
  IV U130 ( .A(n4827), .Z(n38) );
  XOR U131 ( .A(n3416), .B(n3381), .Z(n3385) );
  XOR U132 ( .A(n4375), .B(n4376), .Z(n3951) );
  MUX U133 ( .IN0(n4574), .IN1(n39), .SEL(n4222), .F(n4563) );
  IV U134 ( .A(n4220), .Z(n39) );
  MUX U135 ( .IN0(n4213), .IN1(n40), .SEL(n4214), .F(n4192) );
  IV U136 ( .A(n4215), .Z(n40) );
  MUX U137 ( .IN0(n3927), .IN1(n3925), .SEL(n3926), .F(n3908) );
  MUX U138 ( .IN0(n4757), .IN1(n41), .SEL(n4758), .F(n4736) );
  IV U139 ( .A(n4759), .Z(n41) );
  MUX U140 ( .IN0(n3251), .IN1(n3249), .SEL(n3250), .F(n3211) );
  XOR U141 ( .A(n4344), .B(n4345), .Z(n3900) );
  MUX U142 ( .IN0(n4912), .IN1(n42), .SEL(n4745), .F(n4899) );
  IV U143 ( .A(n4743), .Z(n42) );
  MUX U144 ( .IN0(n43), .IN1(n4708), .SEL(n4709), .F(n3095) );
  IV U145 ( .A(n4710), .Z(n43) );
  MUX U146 ( .IN0(n44), .IN1(n3170), .SEL(n3171), .F(n3040) );
  IV U147 ( .A(n3172), .Z(n44) );
  MUX U148 ( .IN0(n45), .IN1(n2639), .SEL(n2640), .F(n2515) );
  IV U149 ( .A(n2641), .Z(n45) );
  MUX U150 ( .IN0(n46), .IN1(n2597), .SEL(n2598), .F(n2475) );
  IV U151 ( .A(n2599), .Z(n46) );
  MUX U152 ( .IN0(n47), .IN1(n2288), .SEL(n2289), .F(n2174) );
  IV U153 ( .A(n2290), .Z(n47) );
  MUX U154 ( .IN0(n48), .IN1(n2337), .SEL(n2338), .F(n2219) );
  IV U155 ( .A(n2339), .Z(n48) );
  MUX U156 ( .IN0(n49), .IN1(n2125), .SEL(n2126), .F(n2020) );
  IV U157 ( .A(n2127), .Z(n49) );
  MUX U158 ( .IN0(n50), .IN1(n1798), .SEL(n1799), .F(n1702) );
  IV U159 ( .A(n1800), .Z(n50) );
  MUX U160 ( .IN0(n51), .IN1(n1300), .SEL(n1301), .F(n1230) );
  IV U161 ( .A(n1302), .Z(n51) );
  MUX U162 ( .IN0(n52), .IN1(n1041), .SEL(n1042), .F(n987) );
  IV U163 ( .A(n1043), .Z(n52) );
  MUX U164 ( .IN0(n53), .IN1(n996), .SEL(n997), .F(n938) );
  IV U165 ( .A(n998), .Z(n53) );
  MUX U166 ( .IN0(n3063), .IN1(n3061), .SEL(n3062), .F(n2925) );
  MUX U167 ( .IN0(n2899), .IN1(n2901), .SEL(n2900), .F(n2770) );
  MUX U168 ( .IN0(n2841), .IN1(n2843), .SEL(n2842), .F(n2712) );
  MUX U169 ( .IN0(n2819), .IN1(n2817), .SEL(n2818), .F(n2688) );
  MUX U170 ( .IN0(n2869), .IN1(n2867), .SEL(n2868), .F(n2738) );
  MUX U171 ( .IN0(n2858), .IN1(n2860), .SEL(n2859), .F(n2729) );
  MUX U172 ( .IN0(n2654), .IN1(n2652), .SEL(n2653), .F(n2528) );
  MUX U173 ( .IN0(n2799), .IN1(n54), .SEL(n2798), .F(n2668) );
  IV U174 ( .A(n2797), .Z(n54) );
  MUX U175 ( .IN0(n2398), .IN1(n2400), .SEL(n2399), .F(n2277) );
  MUX U176 ( .IN0(n2319), .IN1(n2317), .SEL(n2318), .F(n2199) );
  MUX U177 ( .IN0(n2369), .IN1(n2367), .SEL(n2368), .F(n2251) );
  MUX U178 ( .IN0(n2071), .IN1(n2069), .SEL(n2070), .F(n1964) );
  MUX U179 ( .IN0(n1880), .IN1(n1878), .SEL(n1879), .F(n1778) );
  MUX U180 ( .IN0(n1930), .IN1(n1928), .SEL(n1929), .F(n1828) );
  MUX U181 ( .IN0(n1819), .IN1(n1821), .SEL(n1820), .F(n1723) );
  MUX U182 ( .IN0(n1414), .IN1(n1412), .SEL(n1413), .F(n1339) );
  MUX U183 ( .IN0(n1453), .IN1(n1455), .SEL(n1454), .F(n1376) );
  MUX U184 ( .IN0(n1438), .IN1(n1436), .SEL(n1437), .F(n55) );
  IV U185 ( .A(n55), .Z(n1359) );
  MUX U186 ( .IN0(n1387), .IN1(n1385), .SEL(n1386), .F(n1313) );
  MUX U187 ( .IN0(n933), .IN1(n935), .SEL(n934), .F(n883) );
  MUX U188 ( .IN0(n56), .IN1(n3123), .SEL(n3124), .F(n2987) );
  IV U189 ( .A(n3125), .Z(n56) );
  MUX U190 ( .IN0(n57), .IN1(n3026), .SEL(n3027), .F(n2890) );
  IV U191 ( .A(n3028), .Z(n57) );
  MUX U192 ( .IN0(n58), .IN1(n2592), .SEL(n2593), .F(n2470) );
  IV U193 ( .A(n2594), .Z(n58) );
  MUX U194 ( .IN0(n2103), .IN1(n59), .SEL(n2104), .F(n1998) );
  IV U195 ( .A(n2105), .Z(n59) );
  MUX U196 ( .IN0(n60), .IN1(n1621), .SEL(n1622), .F(n1529) );
  IV U197 ( .A(n1623), .Z(n60) );
  MUX U198 ( .IN0(n1289), .IN1(n61), .SEL(n1288), .F(n1215) );
  IV U199 ( .A(n1287), .Z(n61) );
  MUX U200 ( .IN0(n62), .IN1(n1098), .SEL(n1099), .F(n1036) );
  IV U201 ( .A(n1100), .Z(n62) );
  MUX U202 ( .IN0(n1077), .IN1(n1075), .SEL(n1076), .F(n1019) );
  MUX U203 ( .IN0(n63), .IN1(n840), .SEL(n841), .F(n805) );
  IV U204 ( .A(n842), .Z(n63) );
  XNOR U205 ( .A(n808), .B(n771), .Z(n776) );
  MUX U206 ( .IN0(n64), .IN1(n2324), .SEL(n2325), .F(n2206) );
  IV U207 ( .A(n2326), .Z(n64) );
  MUX U208 ( .IN0(n2305), .IN1(n2303), .SEL(n2304), .F(n2188) );
  MUX U209 ( .IN0(n65), .IN1(n1785), .SEL(n1786), .F(n1689) );
  IV U210 ( .A(n1787), .Z(n65) );
  MUX U211 ( .IN0(n66), .IN1(n1210), .SEL(n1211), .F(n1148) );
  IV U212 ( .A(n1212), .Z(n66) );
  MUX U213 ( .IN0(n1971), .IN1(n67), .SEL(n1972), .F(n1866) );
  IV U214 ( .A(n1973), .Z(n67) );
  NANDN U215 ( .B(n1769), .A(n1770), .Z(n1671) );
  MUX U216 ( .IN0(n1486), .IN1(n1488), .SEL(n1487), .F(n1402) );
  ANDN U217 ( .A(n1322), .B(n1323), .Z(n1252) );
  AND U218 ( .A(n1062), .B(n1063), .Z(n1008) );
  XNOR U219 ( .A(n880), .B(n879), .Z(n871) );
  AND U220 ( .A(n860), .B(n861), .Z(n823) );
  OR U221 ( .A(n1016), .B(n1017), .Z(n958) );
  OR U222 ( .A(n792), .B(n793), .Z(n759) );
  XNOR U223 ( .A(n732), .B(n731), .Z(n730) );
  ANDN U224 ( .A(n685), .B(n684), .Z(n683) );
  MUX U225 ( .IN0(n68), .IN1(n4125), .SEL(n4126), .F(n4108) );
  IV U226 ( .A(n4127), .Z(n68) );
  MUX U227 ( .IN0(n69), .IN1(n3709), .SEL(n3710), .F(n3671) );
  IV U228 ( .A(n3711), .Z(n69) );
  MUX U229 ( .IN0(n70), .IN1(n3722), .SEL(n3723), .F(n3684) );
  IV U230 ( .A(n3724), .Z(n70) );
  MUX U231 ( .IN0(n71), .IN1(n4524), .SEL(n4525), .F(n4511) );
  IV U232 ( .A(n4526), .Z(n71) );
  MUX U233 ( .IN0(n72), .IN1(n3755), .SEL(n3756), .F(n3717) );
  IV U234 ( .A(n3757), .Z(n72) );
  XNOR U235 ( .A(n3699), .B(n3664), .Z(n3668) );
  MUX U236 ( .IN0(n73), .IN1(n4504), .SEL(n4505), .F(n4491) );
  IV U237 ( .A(n4506), .Z(n73) );
  MUX U238 ( .IN0(n74), .IN1(n4119), .SEL(n3735), .F(n4102) );
  IV U239 ( .A(n3733), .Z(n74) );
  XOR U240 ( .A(n4494), .B(n4486), .Z(n4088) );
  XNOR U241 ( .A(n4089), .B(n4075), .Z(n4079) );
  XOR U242 ( .A(n4466), .B(n4467), .Z(n4070) );
  XOR U243 ( .A(n3644), .B(n3609), .Z(n3613) );
  XNOR U244 ( .A(n3585), .B(n3550), .Z(n3554) );
  MUX U245 ( .IN0(n4029), .IN1(n4027), .SEL(n4028), .F(n4010) );
  XOR U246 ( .A(n4442), .B(n4434), .Z(n4020) );
  MUX U247 ( .IN0(n75), .IN1(n4979), .SEL(n4980), .F(n4966) );
  IV U248 ( .A(n4981), .Z(n75) );
  MUX U249 ( .IN0(n76), .IN1(n4986), .SEL(n4987), .F(n4973) );
  IV U250 ( .A(n4988), .Z(n76) );
  XOR U251 ( .A(n3530), .B(n3495), .Z(n3499) );
  MUX U252 ( .IN0(n77), .IN1(n3989), .SEL(n3990), .F(n3972) );
  IV U253 ( .A(n3991), .Z(n77) );
  XOR U254 ( .A(n4268), .B(n4269), .Z(n4278) );
  MUX U255 ( .IN0(n3441), .IN1(n3439), .SEL(n3440), .F(n3401) );
  MUX U256 ( .IN0(n4607), .IN1(n78), .SEL(n4285), .F(n4596) );
  IV U257 ( .A(n4283), .Z(n78) );
  MUX U258 ( .IN0(n79), .IN1(n4251), .SEL(n4252), .F(n4230) );
  IV U259 ( .A(n4253), .Z(n79) );
  XOR U260 ( .A(n4856), .B(n4838), .Z(n4842) );
  XOR U261 ( .A(n4956), .B(n4948), .Z(n4808) );
  XOR U262 ( .A(n4390), .B(n4382), .Z(n3952) );
  MUX U263 ( .IN0(n3944), .IN1(n3942), .SEL(n3943), .F(n3925) );
  XNOR U264 ( .A(n3319), .B(n3284), .Z(n3288) );
  MUX U265 ( .IN0(n4778), .IN1(n80), .SEL(n4779), .F(n4757) );
  IV U266 ( .A(n4780), .Z(n80) );
  MUX U267 ( .IN0(n81), .IN1(n3904), .SEL(n3905), .F(n3884) );
  IV U268 ( .A(n3906), .Z(n81) );
  MUX U269 ( .IN0(n3308), .IN1(n3310), .SEL(n3309), .F(n3270) );
  MUX U270 ( .IN0(n4563), .IN1(n82), .SEL(n4201), .F(n4552) );
  IV U271 ( .A(n4199), .Z(n82) );
  MUX U272 ( .IN0(n4192), .IN1(n83), .SEL(n4193), .F(n4171) );
  IV U273 ( .A(n4194), .Z(n83) );
  XOR U274 ( .A(n4728), .B(n4729), .Z(n4738) );
  MUX U275 ( .IN0(n84), .IN1(n4732), .SEL(n4733), .F(n4700) );
  IV U276 ( .A(n4734), .Z(n84) );
  MUX U277 ( .IN0(n85), .IN1(n3228), .SEL(n3229), .F(n3161) );
  IV U278 ( .A(n3230), .Z(n85) );
  XOR U279 ( .A(n4904), .B(n4896), .Z(n4724) );
  XOR U280 ( .A(n4709), .B(n4710), .Z(n4706) );
  MUX U281 ( .IN0(n86), .IN1(n3178), .SEL(n3179), .F(n3048) );
  IV U282 ( .A(n3180), .Z(n86) );
  XNOR U283 ( .A(n3205), .B(n3171), .Z(n3175) );
  XNOR U284 ( .A(n5169), .B(n5170), .Z(n3141) );
  MUX U285 ( .IN0(n3192), .IN1(n3190), .SEL(n3191), .F(n3061) );
  MUX U286 ( .IN0(n87), .IN1(n2992), .SEL(n2993), .F(n2854) );
  IV U287 ( .A(n2994), .Z(n87) );
  MUX U288 ( .IN0(n88), .IN1(n3001), .SEL(n3002), .F(n2863) );
  IV U289 ( .A(n3003), .Z(n88) );
  MUX U290 ( .IN0(n89), .IN1(n2813), .SEL(n2814), .F(n2684) );
  IV U291 ( .A(n2815), .Z(n89) );
  MUX U292 ( .IN0(n90), .IN1(n2921), .SEL(n2922), .F(n2797) );
  IV U293 ( .A(n2923), .Z(n90) );
  MUX U294 ( .IN0(n91), .IN1(n2524), .SEL(n2525), .F(n2403) );
  IV U295 ( .A(n2526), .Z(n91) );
  MUX U296 ( .IN0(n92), .IN1(n2515), .SEL(n2516), .F(n2394) );
  IV U297 ( .A(n2517), .Z(n92) );
  MUX U298 ( .IN0(n93), .IN1(n2450), .SEL(n2451), .F(n2329) );
  IV U299 ( .A(n2452), .Z(n93) );
  MUX U300 ( .IN0(n94), .IN1(n2203), .SEL(n2204), .F(n2092) );
  IV U301 ( .A(n2205), .Z(n94) );
  MUX U302 ( .IN0(n95), .IN1(n2065), .SEL(n2066), .F(n1960) );
  IV U303 ( .A(n2067), .Z(n95) );
  MUX U304 ( .IN0(n96), .IN1(n1774), .SEL(n1775), .F(n1676) );
  IV U305 ( .A(n1776), .Z(n96) );
  MUX U306 ( .IN0(n97), .IN1(n1265), .SEL(n1266), .F(n1199) );
  IV U307 ( .A(n1267), .Z(n97) );
  MUX U308 ( .IN0(n98), .IN1(n1173), .SEL(n1174), .F(n1112) );
  IV U309 ( .A(n1175), .Z(n98) );
  MUX U310 ( .IN0(n99), .IN1(n1182), .SEL(n1183), .F(n1121) );
  IV U311 ( .A(n1184), .Z(n99) );
  MUX U312 ( .IN0(n100), .IN1(n890), .SEL(n891), .F(n848) );
  IV U313 ( .A(n892), .Z(n100) );
  MUX U314 ( .IN0(n3896), .IN1(n4332), .SEL(n3897), .F(n101) );
  IV U315 ( .A(n101), .Z(n3081) );
  MUX U316 ( .IN0(n2781), .IN1(n2779), .SEL(n2780), .F(n2652) );
  MUX U317 ( .IN0(n2770), .IN1(n2772), .SEL(n2771), .F(n2643) );
  MUX U318 ( .IN0(n2729), .IN1(n2731), .SEL(n2730), .F(n2601) );
  MUX U319 ( .IN0(n2712), .IN1(n2714), .SEL(n2713), .F(n2584) );
  MUX U320 ( .IN0(n2671), .IN1(n102), .SEL(n2670), .F(n2539) );
  IV U321 ( .A(n2669), .Z(n102) );
  MUX U322 ( .IN0(n2440), .IN1(n2438), .SEL(n2439), .F(n2317) );
  MUX U323 ( .IN0(n2277), .IN1(n2279), .SEL(n2278), .F(n103) );
  IV U324 ( .A(n103), .Z(n2169) );
  MUX U325 ( .IN0(n2294), .IN1(n2292), .SEL(n2293), .F(n2178) );
  MUX U326 ( .IN0(n2240), .IN1(n2242), .SEL(n2241), .F(n2129) );
  MUX U327 ( .IN0(n2223), .IN1(n2225), .SEL(n2224), .F(n2112) );
  MUX U328 ( .IN0(n1802), .IN1(n1804), .SEL(n1803), .F(n1706) );
  MUX U329 ( .IN0(n1723), .IN1(n1725), .SEL(n1724), .F(n1630) );
  MUX U330 ( .IN0(n1341), .IN1(n1339), .SEL(n1340), .F(n1269) );
  MUX U331 ( .IN0(n1376), .IN1(n1378), .SEL(n1377), .F(n1304) );
  MUX U332 ( .IN0(n1315), .IN1(n1313), .SEL(n1314), .F(n1243) );
  MUX U333 ( .IN0(n1107), .IN1(n1109), .SEL(n1108), .F(n1045) );
  MUX U334 ( .IN0(n1002), .IN1(n1000), .SEL(n1001), .F(n942) );
  MUX U335 ( .IN0(n883), .IN1(n885), .SEL(n884), .F(n843) );
  MUX U336 ( .IN0(n3106), .IN1(n104), .SEL(n3107), .F(n2970) );
  IV U337 ( .A(n3108), .Z(n104) );
  MUX U338 ( .IN0(n105), .IN1(n2987), .SEL(n2988), .F(n2849) );
  IV U339 ( .A(n2989), .Z(n105) );
  MUX U340 ( .IN0(n106), .IN1(n2890), .SEL(n2891), .F(n2761) );
  IV U341 ( .A(n2892), .Z(n106) );
  XNOR U342 ( .A(n2732), .B(n2607), .Z(n2611) );
  MUX U343 ( .IN0(n2575), .IN1(n107), .SEL(n2576), .F(n2453) );
  IV U344 ( .A(n2577), .Z(n107) );
  MUX U345 ( .IN0(n108), .IN1(n2470), .SEL(n2471), .F(n2349) );
  IV U346 ( .A(n2472), .Z(n108) );
  XNOR U347 ( .A(n2243), .B(n2135), .Z(n2139) );
  MUX U348 ( .IN0(n2057), .IN1(n109), .SEL(n2058), .F(n1955) );
  IV U349 ( .A(n2059), .Z(n109) );
  XNOR U350 ( .A(n2082), .B(n1980), .Z(n1984) );
  MUX U351 ( .IN0(n110), .IN1(n2015), .SEL(n2016), .F(n1910) );
  IV U352 ( .A(n2017), .Z(n110) );
  XNOR U353 ( .A(n1726), .B(n1636), .Z(n1640) );
  MUX U354 ( .IN0(n1604), .IN1(n111), .SEL(n1605), .F(n1511) );
  IV U355 ( .A(n1606), .Z(n111) );
  MUX U356 ( .IN0(n112), .IN1(n1529), .SEL(n1530), .F(n1444) );
  IV U357 ( .A(n1531), .Z(n112) );
  MUX U358 ( .IN0(n113), .IN1(n1036), .SEL(n1037), .F(n981) );
  IV U359 ( .A(n1038), .Z(n113) );
  OR U360 ( .A(n1079), .B(n1080), .Z(n1073) );
  MUX U361 ( .IN0(n807), .IN1(n114), .SEL(n806), .F(n765) );
  IV U362 ( .A(n805), .Z(n114) );
  MUX U363 ( .IN0(n115), .IN1(n2695), .SEL(n2696), .F(n2567) );
  IV U364 ( .A(n2697), .Z(n115) );
  MUX U365 ( .IN0(n116), .IN1(n2206), .SEL(n2207), .F(n2095) );
  IV U366 ( .A(n2208), .Z(n116) );
  MUX U367 ( .IN0(n1661), .IN1(n1659), .SEL(n1660), .F(n1576) );
  NANDN U368 ( .B(n1218), .A(n1219), .Z(n1213) );
  MUX U369 ( .IN0(n777), .IN1(n775), .SEL(n776), .F(n739) );
  XNOR U370 ( .A(n2512), .B(n2511), .Z(n2552) );
  ANDN U371 ( .A(n2620), .B(n2619), .Z(n2497) );
  MUX U372 ( .IN0(n2299), .IN1(n117), .SEL(n2300), .F(n2185) );
  IV U373 ( .A(n2301), .Z(n117) );
  MUX U374 ( .IN0(n1866), .IN1(n118), .SEL(n1867), .F(n1766) );
  IV U375 ( .A(n1868), .Z(n118) );
  NANDN U376 ( .B(n1671), .A(n1672), .Z(n1565) );
  ANDN U377 ( .A(n1471), .B(n1472), .Z(n1394) );
  AND U378 ( .A(n1185), .B(n1186), .Z(n1124) );
  AND U379 ( .A(n950), .B(n951), .Z(n904) );
  OR U380 ( .A(n870), .B(n871), .Z(n833) );
  MUX U381 ( .IN0(n1404), .IN1(n1402), .SEL(n1403), .F(n1330) );
  XNOR U382 ( .A(n1088), .B(n1087), .Z(n1071) );
  OR U383 ( .A(n912), .B(n913), .Z(n868) );
  MUX U384 ( .IN0(n119), .IN1(n825), .SEL(n826), .F(n785) );
  IV U385 ( .A(\_MxM/Y0[26] ), .Z(n119) );
  OR U386 ( .A(n759), .B(n760), .Z(n729) );
  AND U387 ( .A(n783), .B(n784), .Z(n750) );
  OR U388 ( .A(n706), .B(n707), .Z(n684) );
  MUX U389 ( .IN0(n120), .IN1(n2876), .SEL(n1128), .F(n2747) );
  IV U390 ( .A(\_MxM/Y0[2] ), .Z(n120) );
  MUX U391 ( .IN0(n2378), .IN1(n121), .SEL(n659), .F(n2262) );
  IV U392 ( .A(\_MxM/Y0[6] ), .Z(n121) );
  MUX U393 ( .IN0(n1939), .IN1(n122), .SEL(n655), .F(n1839) );
  IV U394 ( .A(\_MxM/Y0[10] ), .Z(n122) );
  MUX U395 ( .IN0(n1558), .IN1(n123), .SEL(n1559), .F(n1473) );
  IV U396 ( .A(\_MxM/Y0[14] ), .Z(n123) );
  MUX U397 ( .IN0(n1254), .IN1(n124), .SEL(n1255), .F(n1187) );
  IV U398 ( .A(\_MxM/Y0[18] ), .Z(n124) );
  MUX U399 ( .IN0(n125), .IN1(n1010), .SEL(n1011), .F(n952) );
  IV U400 ( .A(\_MxM/Y0[22] ), .Z(n125) );
  MUX U401 ( .IN0(n126), .IN1(n3760), .SEL(n3761), .F(n3722) );
  IV U402 ( .A(n3762), .Z(n126) );
  MUX U403 ( .IN0(n127), .IN1(n4116), .SEL(n4117), .F(n4099) );
  IV U404 ( .A(n4118), .Z(n127) );
  MUX U405 ( .IN0(n128), .IN1(n3714), .SEL(n3715), .F(n3676) );
  IV U406 ( .A(n3716), .Z(n128) );
  MUX U407 ( .IN0(n129), .IN1(n3671), .SEL(n3672), .F(n3633) );
  IV U408 ( .A(n3673), .Z(n129) );
  XNOR U409 ( .A(n4123), .B(n4109), .Z(n4113) );
  MUX U410 ( .IN0(n130), .IN1(n4511), .SEL(n4512), .F(n4498) );
  IV U411 ( .A(n4513), .Z(n130) );
  MUX U412 ( .IN0(n3717), .IN1(n131), .SEL(n3718), .F(n3679) );
  IV U413 ( .A(n3719), .Z(n131) );
  XNOR U414 ( .A(n3661), .B(n3626), .Z(n3630) );
  MUX U415 ( .IN0(n132), .IN1(n4491), .SEL(n4492), .F(n4478) );
  IV U416 ( .A(n4493), .Z(n132) );
  MUX U417 ( .IN0(n133), .IN1(n4102), .SEL(n3697), .F(n4085) );
  IV U418 ( .A(n3695), .Z(n133) );
  XOR U419 ( .A(n3682), .B(n3647), .Z(n3651) );
  XOR U420 ( .A(n4481), .B(n4473), .Z(n4071) );
  MUX U421 ( .IN0(n4063), .IN1(n4061), .SEL(n4062), .F(n4044) );
  MUX U422 ( .IN0(n134), .IN1(n3519), .SEL(n3520), .F(n3481) );
  IV U423 ( .A(n3521), .Z(n134) );
  XNOR U424 ( .A(n3547), .B(n3512), .Z(n3516) );
  XOR U425 ( .A(n3568), .B(n3533), .Z(n3537) );
  MUX U426 ( .IN0(n135), .IN1(n4293), .SEL(n4294), .F(n4272) );
  IV U427 ( .A(n4295), .Z(n135) );
  MUX U428 ( .IN0(n4437), .IN1(n136), .SEL(n4020), .F(n4424) );
  IV U429 ( .A(n4019), .Z(n136) );
  XOR U430 ( .A(n4982), .B(n4974), .Z(n4850) );
  MUX U431 ( .IN0(n3995), .IN1(n3993), .SEL(n3994), .F(n3976) );
  MUX U432 ( .IN0(n137), .IN1(n3972), .SEL(n3973), .F(n3955) );
  IV U433 ( .A(n3974), .Z(n137) );
  XNOR U434 ( .A(n3433), .B(n3398), .Z(n3402) );
  XOR U435 ( .A(n4601), .B(n4593), .Z(n4264) );
  MUX U436 ( .IN0(n138), .IN1(n4587), .SEL(n4588), .F(n4576) );
  IV U437 ( .A(n4589), .Z(n138) );
  MUX U438 ( .IN0(n4841), .IN1(n139), .SEL(n4842), .F(n4820) );
  IV U439 ( .A(n4843), .Z(n139) );
  MUX U440 ( .IN0(n140), .IN1(n3367), .SEL(n3368), .F(n3329) );
  IV U441 ( .A(n3369), .Z(n140) );
  XOR U442 ( .A(n3454), .B(n3419), .Z(n3423) );
  MUX U443 ( .IN0(n141), .IN1(n4674), .SEL(n4675), .F(n4659) );
  IV U444 ( .A(n4676), .Z(n141) );
  MUX U445 ( .IN0(n142), .IN1(n4669), .SEL(n4670), .F(n4653) );
  IV U446 ( .A(n4671), .Z(n142) );
  MUX U447 ( .IN0(n4255), .IN1(n143), .SEL(n4256), .F(n4234) );
  IV U448 ( .A(n4257), .Z(n143) );
  MUX U449 ( .IN0(n144), .IN1(n4400), .SEL(n4401), .F(n4387) );
  IV U450 ( .A(n4402), .Z(n144) );
  MUX U451 ( .IN0(n145), .IN1(n5046), .SEL(n5047), .F(n5031) );
  IV U452 ( .A(n5048), .Z(n145) );
  MUX U453 ( .IN0(n146), .IN1(n5041), .SEL(n5042), .F(n5025) );
  IV U454 ( .A(n5043), .Z(n146) );
  XOR U455 ( .A(n4954), .B(n4955), .Z(n4827) );
  MUX U456 ( .IN0(n147), .IN1(n4947), .SEL(n4948), .F(n4934) );
  IV U457 ( .A(n4949), .Z(n147) );
  MUX U458 ( .IN0(n148), .IN1(n4790), .SEL(n4791), .F(n4769) );
  IV U459 ( .A(n4792), .Z(n148) );
  MUX U460 ( .IN0(n149), .IN1(n4795), .SEL(n4796), .F(n4774) );
  IV U461 ( .A(n4797), .Z(n149) );
  MUX U462 ( .IN0(n150), .IN1(n3342), .SEL(n3343), .F(n3304) );
  IV U463 ( .A(n3344), .Z(n150) );
  MUX U464 ( .IN0(n151), .IN1(n3824), .SEL(n3825), .F(n3808) );
  IV U465 ( .A(n3826), .Z(n151) );
  XOR U466 ( .A(n4205), .B(n4206), .Z(n4215) );
  MUX U467 ( .IN0(n152), .IN1(n4927), .SEL(n4928), .F(n4914) );
  IV U468 ( .A(n4929), .Z(n152) );
  XOR U469 ( .A(n4184), .B(n4185), .Z(n4194) );
  XOR U470 ( .A(n4377), .B(n4369), .Z(n3935) );
  MUX U471 ( .IN0(n153), .IN1(n5151), .SEL(n5152), .F(n5147) );
  IV U472 ( .A(n5153), .Z(n153) );
  MUX U473 ( .IN0(n3289), .IN1(n3287), .SEL(n3288), .F(n3249) );
  XOR U474 ( .A(n4557), .B(n4549), .Z(n4180) );
  MUX U475 ( .IN0(n154), .IN1(n4543), .SEL(n4544), .F(n4532) );
  IV U476 ( .A(n4545), .Z(n154) );
  XOR U477 ( .A(n4163), .B(n4164), .Z(n4173) );
  MUX U478 ( .IN0(n155), .IN1(n4167), .SEL(n4168), .F(n4142) );
  IV U479 ( .A(n4169), .Z(n155) );
  XOR U480 ( .A(n4917), .B(n4909), .Z(n4745) );
  MUX U481 ( .IN0(n156), .IN1(n3207), .SEL(n3208), .F(n3170) );
  IV U482 ( .A(n3209), .Z(n156) );
  MUX U483 ( .IN0(n3910), .IN1(n3908), .SEL(n3909), .F(n3888) );
  MUX U484 ( .IN0(n3270), .IN1(n3272), .SEL(n3271), .F(n3232) );
  MUX U485 ( .IN0(n4736), .IN1(n157), .SEL(n4737), .F(n4704) );
  IV U486 ( .A(n4738), .Z(n157) );
  MUX U487 ( .IN0(n158), .IN1(n4700), .SEL(n4701), .F(n3087) );
  IV U488 ( .A(n4702), .Z(n158) );
  MUX U489 ( .IN0(n159), .IN1(n3161), .SEL(n3162), .F(n3031) );
  IV U490 ( .A(n3163), .Z(n159) );
  MUX U491 ( .IN0(n160), .IN1(n4343), .SEL(n4344), .F(n3878) );
  IV U492 ( .A(n4345), .Z(n160) );
  MUX U493 ( .IN0(n161), .IN1(n2775), .SEL(n2776), .F(n2648) );
  IV U494 ( .A(n2777), .Z(n161) );
  MUX U495 ( .IN0(n162), .IN1(n2821), .SEL(n2822), .F(n2692) );
  IV U496 ( .A(n2823), .Z(n162) );
  MUX U497 ( .IN0(n163), .IN1(n2475), .SEL(n2476), .F(n2354) );
  IV U498 ( .A(n2477), .Z(n163) );
  MUX U499 ( .IN0(n164), .IN1(n2174), .SEL(n2175), .F(n2065) );
  IV U500 ( .A(n2176), .Z(n164) );
  MUX U501 ( .IN0(n165), .IN1(n2195), .SEL(n2196), .F(n2084) );
  IV U502 ( .A(n2197), .Z(n165) );
  MUX U503 ( .IN0(n166), .IN1(n2108), .SEL(n2109), .F(n2003) );
  IV U504 ( .A(n2110), .Z(n166) );
  MUX U505 ( .IN0(n167), .IN1(n2020), .SEL(n2021), .F(n1915) );
  IV U506 ( .A(n2022), .Z(n167) );
  MUX U507 ( .IN0(n168), .IN1(n1987), .SEL(n1988), .F(n1882) );
  IV U508 ( .A(n1989), .Z(n168) );
  MUX U509 ( .IN0(n169), .IN1(n1694), .SEL(n1695), .F(n1601) );
  IV U510 ( .A(n1696), .Z(n169) );
  MUX U511 ( .IN0(n170), .IN1(n1702), .SEL(n1703), .F(n1609) );
  IV U512 ( .A(n1704), .Z(n170) );
  MUX U513 ( .IN0(n171), .IN1(n1458), .SEL(n1459), .F(n1381) );
  IV U514 ( .A(n1460), .Z(n171) );
  MUX U515 ( .IN0(n172), .IN1(n1230), .SEL(n1231), .F(n1164) );
  IV U516 ( .A(n1232), .Z(n172) );
  MUX U517 ( .IN0(n173), .IN1(n1156), .SEL(n1157), .F(n1095) );
  IV U518 ( .A(n1158), .Z(n173) );
  MUX U519 ( .IN0(n174), .IN1(n1059), .SEL(n1060), .F(n1005) );
  IV U520 ( .A(n1061), .Z(n174) );
  MUX U521 ( .IN0(n175), .IN1(n1050), .SEL(n1051), .F(n996) );
  IV U522 ( .A(n1052), .Z(n175) );
  MUX U523 ( .IN0(n176), .IN1(n1199), .SEL(n1200), .F(n1137) );
  IV U524 ( .A(n1201), .Z(n176) );
  MUX U525 ( .IN0(n177), .IN1(n987), .SEL(n988), .F(n928) );
  IV U526 ( .A(n989), .Z(n177) );
  MUX U527 ( .IN0(n178), .IN1(n921), .SEL(n922), .F(n875) );
  IV U528 ( .A(n923), .Z(n178) );
  MUX U529 ( .IN0(n3132), .IN1(n3134), .SEL(n3133), .F(n2996) );
  MUX U530 ( .IN0(n3046), .IN1(n3044), .SEL(n3045), .F(n2908) );
  MUX U531 ( .IN0(n3881), .IN1(n179), .SEL(n3203), .F(n3078) );
  IV U532 ( .A(n3202), .Z(n179) );
  MUX U533 ( .IN0(n2979), .IN1(n2981), .SEL(n2980), .F(n2841) );
  MUX U534 ( .IN0(n2793), .IN1(n2791), .SEL(n2792), .F(n2669) );
  XOR U535 ( .A(n2744), .B(n2871), .Z(n2745) );
  MUX U536 ( .IN0(n2643), .IN1(n2645), .SEL(n2644), .F(n2519) );
  MUX U537 ( .IN0(n2530), .IN1(n2528), .SEL(n2529), .F(n2407) );
  MUX U538 ( .IN0(n2601), .IN1(n2603), .SEL(n2602), .F(n2479) );
  MUX U539 ( .IN0(n2462), .IN1(n2464), .SEL(n2463), .F(n2341) );
  MUX U540 ( .IN0(n2285), .IN1(n180), .SEL(n2284), .F(n2168) );
  IV U541 ( .A(n2283), .Z(n180) );
  XOR U542 ( .A(n2039), .B(n2142), .Z(n2040) );
  MUX U543 ( .IN0(n2129), .IN1(n2131), .SEL(n2130), .F(n2024) );
  MUX U544 ( .IN0(n1966), .IN1(n1964), .SEL(n1965), .F(n1851) );
  MUX U545 ( .IN0(n1902), .IN1(n1904), .SEL(n1903), .F(n1802) );
  MUX U546 ( .IN0(n1630), .IN1(n1632), .SEL(n1631), .F(n1538) );
  MUX U547 ( .IN0(n1271), .IN1(n1269), .SEL(n1270), .F(n1203) );
  MUX U548 ( .IN0(n1304), .IN1(n1306), .SEL(n1305), .F(n1234) );
  MUX U549 ( .IN0(n1245), .IN1(n1243), .SEL(n1244), .F(n1177) );
  MUX U550 ( .IN0(n1045), .IN1(n1047), .SEL(n1046), .F(n991) );
  MUX U551 ( .IN0(n181), .IN1(n1145), .SEL(n1146), .F(n1083) );
  IV U552 ( .A(n1147), .Z(n181) );
  MUX U553 ( .IN0(n944), .IN1(n942), .SEL(n943), .F(n894) );
  XNOR U554 ( .A(n3135), .B(n3002), .Z(n3006) );
  XNOR U555 ( .A(n2949), .B(n2814), .Z(n2818) );
  MUX U556 ( .IN0(n182), .IN1(n2761), .SEL(n2762), .F(n2634) );
  IV U557 ( .A(n2763), .Z(n182) );
  MUX U558 ( .IN0(n183), .IN1(n2849), .SEL(n2850), .F(n2720) );
  IV U559 ( .A(n2851), .Z(n183) );
  XNOR U560 ( .A(n2554), .B(n2435), .Z(n2439) );
  XNOR U561 ( .A(n2604), .B(n2485), .Z(n2489) );
  MUX U562 ( .IN0(n184), .IN1(n2273), .SEL(n2274), .F(n2160) );
  IV U563 ( .A(n2275), .Z(n184) );
  MUX U564 ( .IN0(n185), .IN1(n2349), .SEL(n2350), .F(n2231) );
  IV U565 ( .A(n2351), .Z(n185) );
  XNOR U566 ( .A(n2132), .B(n2030), .Z(n2034) );
  XNOR U567 ( .A(n1977), .B(n1875), .Z(n1879) );
  MUX U568 ( .IN0(n186), .IN1(n1910), .SEL(n1911), .F(n1810) );
  IV U569 ( .A(n1912), .Z(n186) );
  XNOR U570 ( .A(n1822), .B(n1729), .Z(n1735) );
  MUX U571 ( .IN0(n1793), .IN1(n187), .SEL(n1794), .F(n1697) );
  IV U572 ( .A(n1795), .Z(n187) );
  XNOR U573 ( .A(n1583), .B(n1493), .Z(n1497) );
  XOR U574 ( .A(n1425), .B(n1426), .Z(n1438) );
  XOR U575 ( .A(n1354), .B(n1355), .Z(n1361) );
  MUX U576 ( .IN0(n188), .IN1(n1444), .SEL(n1445), .F(n1367) );
  IV U577 ( .A(n1446), .Z(n188) );
  MUX U578 ( .IN0(n189), .IN1(n981), .SEL(n982), .F(n924) );
  IV U579 ( .A(n983), .Z(n189) );
  MUX U580 ( .IN0(n843), .IN1(n845), .SEL(n844), .F(n190) );
  IV U581 ( .A(n190), .Z(n798) );
  MUX U582 ( .IN0(n191), .IN1(n3098), .SEL(n3099), .F(n2962) );
  IV U583 ( .A(n3100), .Z(n191) );
  MUX U584 ( .IN0(n192), .IN1(n3068), .SEL(n3069), .F(n2932) );
  IV U585 ( .A(n3070), .Z(n192) );
  MUX U586 ( .IN0(n193), .IN1(n2567), .SEL(n2568), .F(n2445) );
  IV U587 ( .A(n2569), .Z(n193) );
  MUX U588 ( .IN0(n194), .IN1(n2095), .SEL(n2096), .F(n1990) );
  IV U589 ( .A(n2097), .Z(n194) );
  MUX U590 ( .IN0(n195), .IN1(n1596), .SEL(n1597), .F(n1503) );
  IV U591 ( .A(n1598), .Z(n195) );
  MUX U592 ( .IN0(n196), .IN1(n1276), .SEL(n1277), .F(n1210) );
  IV U593 ( .A(n1278), .Z(n196) );
  MUX U594 ( .IN0(n1151), .IN1(n1153), .SEL(n1152), .F(n1089) );
  MUX U595 ( .IN0(n197), .IN1(n1026), .SEL(n1027), .F(n973) );
  IV U596 ( .A(n1028), .Z(n197) );
  MUX U597 ( .IN0(n1021), .IN1(n1019), .SEL(n1020), .F(n968) );
  XNOR U598 ( .A(n854), .B(n853), .Z(n842) );
  XNOR U599 ( .A(n817), .B(n816), .Z(n807) );
  XNOR U600 ( .A(n769), .B(n742), .Z(n740) );
  MUX U601 ( .IN0(n2786), .IN1(n198), .SEL(n2787), .F(n2659) );
  IV U602 ( .A(n2788), .Z(n198) );
  XNOR U603 ( .A(n2550), .B(n2549), .Z(n2662) );
  ANDN U604 ( .A(n2376), .B(n2377), .Z(n2260) );
  ANDN U605 ( .A(n1648), .B(n1649), .Z(n1556) );
  NOR U606 ( .A(n1484), .B(n1485), .Z(n1483) );
  AND U607 ( .A(n1124), .B(n1125), .Z(n1062) );
  AND U608 ( .A(n904), .B(n905), .Z(n860) );
  XOR U609 ( .A(n2079), .B(n2076), .Z(n2154) );
  XOR U610 ( .A(n1671), .B(n1668), .Z(n1751) );
  OR U611 ( .A(n1330), .B(n1331), .Z(n1260) );
  OR U612 ( .A(n1070), .B(n1071), .Z(n1016) );
  OR U613 ( .A(n868), .B(n869), .Z(n831) );
  MUX U614 ( .IN0(n199), .IN1(n785), .SEL(n786), .F(n752) );
  IV U615 ( .A(\_MxM/Y0[27] ), .Z(n199) );
  OR U616 ( .A(n729), .B(n730), .Z(n704) );
  MUX U617 ( .IN0(n200), .IN1(n2747), .SEL(n699), .F(n2621) );
  IV U618 ( .A(\_MxM/Y0[3] ), .Z(n200) );
  MUX U619 ( .IN0(n2262), .IN1(n201), .SEL(n658), .F(n2149) );
  IV U620 ( .A(\_MxM/Y0[7] ), .Z(n201) );
  MUX U621 ( .IN0(n1839), .IN1(n202), .SEL(n1840), .F(n1745) );
  IV U622 ( .A(\_MxM/Y0[11] ), .Z(n202) );
  MUX U623 ( .IN0(n1473), .IN1(n203), .SEL(n1474), .F(n1396) );
  IV U624 ( .A(\_MxM/Y0[15] ), .Z(n203) );
  MUX U625 ( .IN0(n204), .IN1(n1187), .SEL(n1188), .F(n1126) );
  IV U626 ( .A(\_MxM/Y0[19] ), .Z(n204) );
  MUX U627 ( .IN0(n205), .IN1(n952), .SEL(n953), .F(n906) );
  IV U628 ( .A(\_MxM/Y0[23] ), .Z(n205) );
  AND U629 ( .A(n692), .B(n693), .Z(n688) );
  MUX U630 ( .IN0(n206), .IN1(n3739), .SEL(n3740), .F(n3701) );
  IV U631 ( .A(n3741), .Z(n206) );
  MUX U632 ( .IN0(n207), .IN1(n3752), .SEL(n3753), .F(n3714) );
  IV U633 ( .A(n3754), .Z(n207) );
  MUX U634 ( .IN0(n208), .IN1(n4517), .SEL(n4518), .F(n4504) );
  IV U635 ( .A(n4519), .Z(n208) );
  MUX U636 ( .IN0(n3669), .IN1(n3667), .SEL(n3668), .F(n3629) );
  MUX U637 ( .IN0(n209), .IN1(n3767), .SEL(n3182), .F(n3729) );
  IV U638 ( .A(n3181), .Z(n209) );
  MUX U639 ( .IN0(n210), .IN1(n4082), .SEL(n4083), .F(n4065) );
  IV U640 ( .A(n4084), .Z(n210) );
  MUX U641 ( .IN0(n211), .IN1(n4074), .SEL(n4075), .F(n4057) );
  IV U642 ( .A(n4076), .Z(n211) );
  MUX U643 ( .IN0(n3688), .IN1(n3690), .SEL(n3689), .F(n3650) );
  MUX U644 ( .IN0(n4502), .IN1(n212), .SEL(n4105), .F(n4489) );
  IV U645 ( .A(n4104), .Z(n212) );
  MUX U646 ( .IN0(n213), .IN1(n3587), .SEL(n3588), .F(n3549) );
  IV U647 ( .A(n3589), .Z(n213) );
  MUX U648 ( .IN0(n214), .IN1(n3600), .SEL(n3601), .F(n3562) );
  IV U649 ( .A(n3602), .Z(n214) );
  MUX U650 ( .IN0(n215), .IN1(n3608), .SEL(n3609), .F(n3570) );
  IV U651 ( .A(n3610), .Z(n215) );
  MUX U652 ( .IN0(n216), .IN1(n4085), .SEL(n3659), .F(n4068) );
  IV U653 ( .A(n3657), .Z(n216) );
  MUX U654 ( .IN0(n4046), .IN1(n4044), .SEL(n4045), .F(n4027) );
  MUX U655 ( .IN0(n3603), .IN1(n217), .SEL(n3604), .F(n3565) );
  IV U656 ( .A(n3605), .Z(n217) );
  MUX U657 ( .IN0(n218), .IN1(n4452), .SEL(n4453), .F(n4439) );
  IV U658 ( .A(n4454), .Z(n218) );
  MUX U659 ( .IN0(n3517), .IN1(n3515), .SEL(n3516), .F(n3477) );
  MUX U660 ( .IN0(n219), .IN1(n4014), .SEL(n4015), .F(n3997) );
  IV U661 ( .A(n4016), .Z(n219) );
  MUX U662 ( .IN0(n220), .IN1(n4006), .SEL(n4007), .F(n3989) );
  IV U663 ( .A(n4008), .Z(n220) );
  MUX U664 ( .IN0(n3536), .IN1(n3538), .SEL(n3537), .F(n3498) );
  MUX U665 ( .IN0(n221), .IN1(n4609), .SEL(n4610), .F(n4598) );
  IV U666 ( .A(n4611), .Z(n221) );
  MUX U667 ( .IN0(n222), .IN1(n3435), .SEL(n3436), .F(n3397) );
  IV U668 ( .A(n3437), .Z(n222) );
  MUX U669 ( .IN0(n223), .IN1(n4446), .SEL(n4447), .F(n4433) );
  IV U670 ( .A(n4448), .Z(n223) );
  MUX U671 ( .IN0(n224), .IN1(n3448), .SEL(n3449), .F(n3410) );
  IV U672 ( .A(n3450), .Z(n224) );
  MUX U673 ( .IN0(n225), .IN1(n3456), .SEL(n3457), .F(n3418) );
  IV U674 ( .A(n3458), .Z(n225) );
  MUX U675 ( .IN0(n226), .IN1(n4603), .SEL(n4604), .F(n4592) );
  IV U676 ( .A(n4605), .Z(n226) );
  MUX U677 ( .IN0(n227), .IN1(n4966), .SEL(n4967), .F(n4953) );
  IV U678 ( .A(n4968), .Z(n227) );
  MUX U679 ( .IN0(n228), .IN1(n4973), .SEL(n4974), .F(n4960) );
  IV U680 ( .A(n4975), .Z(n228) );
  MUX U681 ( .IN0(n229), .IN1(n4832), .SEL(n4833), .F(n4811) );
  IV U682 ( .A(n4834), .Z(n229) );
  MUX U683 ( .IN0(n230), .IN1(n4017), .SEL(n3507), .F(n4000) );
  IV U684 ( .A(n3505), .Z(n230) );
  XOR U685 ( .A(n4291), .B(n4273), .Z(n4277) );
  XOR U686 ( .A(n4247), .B(n4248), .Z(n4257) );
  XOR U687 ( .A(n4416), .B(n4408), .Z(n3986) );
  MUX U688 ( .IN0(n3978), .IN1(n3976), .SEL(n3977), .F(n3959) );
  MUX U689 ( .IN0(n3451), .IN1(n231), .SEL(n3452), .F(n3413) );
  IV U690 ( .A(n3453), .Z(n231) );
  MUX U691 ( .IN0(n4596), .IN1(n232), .SEL(n4264), .F(n4585) );
  IV U692 ( .A(n4262), .Z(n232) );
  XOR U693 ( .A(n4226), .B(n4227), .Z(n4236) );
  MUX U694 ( .IN0(n233), .IN1(n4230), .SEL(n4231), .F(n4209) );
  IV U695 ( .A(n4232), .Z(n233) );
  MUX U696 ( .IN0(n3365), .IN1(n3363), .SEL(n3364), .F(n3325) );
  MUX U697 ( .IN0(n234), .IN1(n3946), .SEL(n3947), .F(n3929) );
  IV U698 ( .A(n3948), .Z(n234) );
  MUX U699 ( .IN0(n235), .IN1(n3938), .SEL(n3939), .F(n3921) );
  IV U700 ( .A(n3940), .Z(n235) );
  MUX U701 ( .IN0(n3384), .IN1(n3386), .SEL(n3385), .F(n3346) );
  MUX U702 ( .IN0(n236), .IN1(n4324), .SEL(n4325), .F(n4663) );
  IV U703 ( .A(n4677), .Z(n236) );
  MUX U704 ( .IN0(n4653), .IN1(n4668), .SEL(n4655), .F(n4637) );
  MUX U705 ( .IN0(n237), .IN1(n5136), .SEL(n5137), .F(n5119) );
  IV U706 ( .A(n5138), .Z(n237) );
  MUX U707 ( .IN0(n238), .IN1(n4889), .SEL(n4890), .F(n5035) );
  IV U708 ( .A(n5049), .Z(n238) );
  MUX U709 ( .IN0(n5025), .IN1(n5040), .SEL(n5027), .F(n5009) );
  XOR U710 ( .A(n4943), .B(n4935), .Z(n4787) );
  MUX U711 ( .IN0(n4799), .IN1(n239), .SEL(n4800), .F(n4778) );
  IV U712 ( .A(n4801), .Z(n239) );
  MUX U713 ( .IN0(n240), .IN1(n4774), .SEL(n4775), .F(n4753) );
  IV U714 ( .A(n4776), .Z(n240) );
  MUX U715 ( .IN0(n241), .IN1(n3283), .SEL(n3284), .F(n3245) );
  IV U716 ( .A(n3285), .Z(n241) );
  MUX U717 ( .IN0(n242), .IN1(n3304), .SEL(n3305), .F(n3266) );
  IV U718 ( .A(n3306), .Z(n242) );
  MUX U719 ( .IN0(n243), .IN1(n3777), .SEL(n3778), .F(n3818) );
  IV U720 ( .A(n3832), .Z(n243) );
  MUX U721 ( .IN0(n3808), .IN1(n3823), .SEL(n3810), .F(n3792) );
  MUX U722 ( .IN0(n244), .IN1(n4374), .SEL(n4375), .F(n4361) );
  IV U723 ( .A(n4376), .Z(n244) );
  MUX U724 ( .IN0(n5113), .IN1(n5128), .SEL(n5115), .F(n5095) );
  MUX U725 ( .IN0(n245), .IN1(n4914), .SEL(n4915), .F(n4901) );
  IV U726 ( .A(n4916), .Z(n245) );
  MUX U727 ( .IN0(n246), .IN1(n4381), .SEL(n4382), .F(n4368) );
  IV U728 ( .A(n4383), .Z(n246) );
  MUX U729 ( .IN0(n247), .IN1(n3949), .SEL(n3355), .F(n3932) );
  IV U730 ( .A(n3353), .Z(n247) );
  MUX U731 ( .IN0(n248), .IN1(n4548), .SEL(n4549), .F(n4537) );
  IV U732 ( .A(n4550), .Z(n248) );
  MUX U733 ( .IN0(n3299), .IN1(n249), .SEL(n3300), .F(n3261) );
  IV U734 ( .A(n3301), .Z(n249) );
  MUX U735 ( .IN0(n4552), .IN1(n250), .SEL(n4180), .F(n4541) );
  IV U736 ( .A(n4178), .Z(n250) );
  XOR U737 ( .A(n4186), .B(n4168), .Z(n4172) );
  XOR U738 ( .A(n4151), .B(n4152), .Z(n4148) );
  MUX U739 ( .IN0(n5164), .IN1(n5167), .SEL(n5165), .F(n3137) );
  MUX U740 ( .IN0(n3213), .IN1(n3211), .SEL(n3212), .F(n3174) );
  MUX U741 ( .IN0(n251), .IN1(n3194), .SEL(n3195), .F(n3065) );
  IV U742 ( .A(n3196), .Z(n251) );
  XNOR U743 ( .A(n3902), .B(n3885), .Z(n3889) );
  MUX U744 ( .IN0(n3232), .IN1(n3234), .SEL(n3233), .F(n3165) );
  MUX U745 ( .IN0(n252), .IN1(n3111), .SEL(n3112), .F(n2975) );
  IV U746 ( .A(n3113), .Z(n252) );
  MUX U747 ( .IN0(n253), .IN1(n3040), .SEL(n3041), .F(n2904) );
  IV U748 ( .A(n3042), .Z(n253) );
  MUX U749 ( .IN0(n254), .IN1(n3023), .SEL(n3024), .F(n2887) );
  IV U750 ( .A(n3025), .Z(n254) );
  MUX U751 ( .IN0(n255), .IN1(n3031), .SEL(n3032), .F(n2895) );
  IV U752 ( .A(n3033), .Z(n255) );
  MUX U753 ( .IN0(n256), .IN1(n3057), .SEL(n3058), .F(n2921) );
  IV U754 ( .A(n3059), .Z(n256) );
  MUX U755 ( .IN0(n257), .IN1(n3900), .SEL(n3901), .F(n4332) );
  IV U756 ( .A(n4346), .Z(n257) );
  MUX U757 ( .IN0(n4899), .IN1(n258), .SEL(n4724), .F(n3115) );
  IV U758 ( .A(n4722), .Z(n258) );
  MUX U759 ( .IN0(n4704), .IN1(n259), .SEL(n4705), .F(n3091) );
  IV U760 ( .A(n4706), .Z(n259) );
  MUX U761 ( .IN0(n260), .IN1(n2967), .SEL(n2968), .F(n2829) );
  IV U762 ( .A(n2969), .Z(n260) );
  MUX U763 ( .IN0(n261), .IN1(n2854), .SEL(n2855), .F(n2725) );
  IV U764 ( .A(n2856), .Z(n261) );
  MUX U765 ( .IN0(n262), .IN1(n2692), .SEL(n2693), .F(n2564) );
  IV U766 ( .A(n2694), .Z(n262) );
  MUX U767 ( .IN0(n263), .IN1(n2532), .SEL(n2533), .F(n2411) );
  IV U768 ( .A(n2534), .Z(n263) );
  MUX U769 ( .IN0(n264), .IN1(n2386), .SEL(n2387), .F(n2270) );
  IV U770 ( .A(n2388), .Z(n264) );
  MUX U771 ( .IN0(n265), .IN1(n2458), .SEL(n2459), .F(n2337) );
  IV U772 ( .A(n2460), .Z(n265) );
  MUX U773 ( .IN0(n266), .IN1(n2313), .SEL(n2314), .F(n2195) );
  IV U774 ( .A(n2315), .Z(n266) );
  MUX U775 ( .IN0(n267), .IN1(n2354), .SEL(n2355), .F(n2236) );
  IV U776 ( .A(n2356), .Z(n267) );
  MUX U777 ( .IN0(n268), .IN1(n2673), .SEL(n2674), .F(n2545) );
  IV U778 ( .A(n2675), .Z(n268) );
  MUX U779 ( .IN0(n269), .IN1(n2228), .SEL(n2229), .F(n2117) );
  IV U780 ( .A(n2230), .Z(n269) );
  MUX U781 ( .IN0(n270), .IN1(n2003), .SEL(n2004), .F(n1898) );
  IV U782 ( .A(n2005), .Z(n270) );
  MUX U783 ( .IN0(n271), .IN1(n1915), .SEL(n1916), .F(n1815) );
  IV U784 ( .A(n1917), .Z(n271) );
  MUX U785 ( .IN0(n272), .IN1(n1807), .SEL(n1808), .F(n1711) );
  IV U786 ( .A(n1809), .Z(n272) );
  MUX U787 ( .IN0(n273), .IN1(n1782), .SEL(n1783), .F(n1686) );
  IV U788 ( .A(n1784), .Z(n273) );
  MUX U789 ( .IN0(n274), .IN1(n1968), .SEL(n1969), .F(n1863) );
  IV U790 ( .A(n1970), .Z(n274) );
  MUX U791 ( .IN0(n275), .IN1(n1960), .SEL(n1961), .F(n1859) );
  IV U792 ( .A(n1962), .Z(n275) );
  MUX U793 ( .IN0(n276), .IN1(n1609), .SEL(n1610), .F(n1521) );
  IV U794 ( .A(n1611), .Z(n276) );
  MUX U795 ( .IN0(n277), .IN1(n1416), .SEL(n1417), .F(n1343) );
  IV U796 ( .A(n1418), .Z(n277) );
  MUX U797 ( .IN0(n278), .IN1(n1449), .SEL(n1450), .F(n1372) );
  IV U798 ( .A(n1451), .Z(n278) );
  MUX U799 ( .IN0(n279), .IN1(n1239), .SEL(n1240), .F(n1173) );
  IV U800 ( .A(n1241), .Z(n279) );
  MUX U801 ( .IN0(n280), .IN1(n1164), .SEL(n1165), .F(n1103) );
  IV U802 ( .A(n1166), .Z(n280) );
  MUX U803 ( .IN0(n2996), .IN1(n2998), .SEL(n2997), .F(n2858) );
  MUX U804 ( .IN0(n3077), .IN1(n281), .SEL(n3076), .F(n2939) );
  IV U805 ( .A(n3075), .Z(n281) );
  MUX U806 ( .IN0(n2584), .IN1(n2586), .SEL(n2585), .F(n2462) );
  MUX U807 ( .IN0(n2479), .IN1(n2481), .SEL(n2480), .F(n2358) );
  MUX U808 ( .IN0(n2180), .IN1(n2178), .SEL(n2179), .F(n2069) );
  MUX U809 ( .IN0(n2171), .IN1(n282), .SEL(n2170), .F(n2060) );
  IV U810 ( .A(n2169), .Z(n282) );
  MUX U811 ( .IN0(n2112), .IN1(n2114), .SEL(n2113), .F(n2007) );
  MUX U812 ( .IN0(n2090), .IN1(n2088), .SEL(n2089), .F(n1983) );
  MUX U813 ( .IN0(n2024), .IN1(n2026), .SEL(n2025), .F(n1919) );
  XOR U814 ( .A(n1645), .B(n1738), .Z(n1646) );
  MUX U815 ( .IN0(n1706), .IN1(n1708), .SEL(n1707), .F(n1613) );
  XNOR U816 ( .A(n1851), .B(n1852), .Z(n1850) );
  MUX U817 ( .IN0(n1234), .IN1(n1236), .SEL(n1235), .F(n1168) );
  MUX U818 ( .IN0(n1118), .IN1(n1116), .SEL(n1117), .F(n1054) );
  MUX U819 ( .IN0(n991), .IN1(n993), .SEL(n992), .F(n933) );
  MUX U820 ( .IN0(n283), .IN1(n3078), .SEL(n3079), .F(n2945) );
  IV U821 ( .A(n3080), .Z(n283) );
  XNOR U822 ( .A(n2999), .B(n2864), .Z(n2868) );
  XNOR U823 ( .A(n2773), .B(n2649), .Z(n2653) );
  XOR U824 ( .A(n2764), .B(n2640), .Z(n2644) );
  NAND U825 ( .A(n2668), .B(n2795), .Z(n2794) );
  MUX U826 ( .IN0(n2832), .IN1(n284), .SEL(n2833), .F(n2703) );
  IV U827 ( .A(n2834), .Z(n284) );
  XNOR U828 ( .A(n2811), .B(n2685), .Z(n2689) );
  MUX U829 ( .IN0(n285), .IN1(n2720), .SEL(n2721), .F(n2592) );
  IV U830 ( .A(n2722), .Z(n285) );
  MUX U831 ( .IN0(n286), .IN1(n2389), .SEL(n2390), .F(n2273) );
  IV U832 ( .A(n2391), .Z(n286) );
  XNOR U833 ( .A(n2482), .B(n2364), .Z(n2368) );
  MUX U834 ( .IN0(n2332), .IN1(n287), .SEL(n2333), .F(n2214) );
  IV U835 ( .A(n2334), .Z(n287) );
  MUX U836 ( .IN0(n288), .IN1(n2231), .SEL(n2232), .F(n2120) );
  IV U837 ( .A(n2233), .Z(n288) );
  XNOR U838 ( .A(n2027), .B(n1925), .Z(n1929) );
  MUX U839 ( .IN0(n1955), .IN1(n289), .SEL(n1956), .F(n1846) );
  IV U840 ( .A(n1957), .Z(n289) );
  MUX U841 ( .IN0(n1893), .IN1(n290), .SEL(n1894), .F(n1793) );
  IV U842 ( .A(n1895), .Z(n290) );
  MUX U843 ( .IN0(n291), .IN1(n1810), .SEL(n1811), .F(n1714) );
  IV U844 ( .A(n1812), .Z(n291) );
  XNOR U845 ( .A(n1772), .B(n1677), .Z(n1683) );
  XOR U846 ( .A(n1717), .B(n1627), .Z(n1631) );
  XNOR U847 ( .A(n1541), .B(n1459), .Z(n1463) );
  MUX U848 ( .IN0(n292), .IN1(n1427), .SEL(n1428), .F(n1356) );
  IV U849 ( .A(n1429), .Z(n292) );
  MUX U850 ( .IN0(n293), .IN1(n1359), .SEL(n1360), .F(n1280) );
  IV U851 ( .A(n1361), .Z(n293) );
  MUX U852 ( .IN0(n294), .IN1(n1367), .SEL(n1368), .F(n1295) );
  IV U853 ( .A(n1369), .Z(n294) );
  XNOR U854 ( .A(n1075), .B(n1080), .Z(n1136) );
  XNOR U855 ( .A(n936), .B(n891), .Z(n897) );
  AND U856 ( .A(n798), .B(n802), .Z(n801) );
  MUX U857 ( .IN0(n295), .IN1(n820), .SEL(n821), .F(n780) );
  IV U858 ( .A(n822), .Z(n295) );
  MUX U859 ( .IN0(n296), .IN1(n2962), .SEL(n2963), .F(n2824) );
  IV U860 ( .A(n2964), .Z(n296) );
  MUX U861 ( .IN0(n297), .IN1(n2932), .SEL(n2933), .F(n2804) );
  IV U862 ( .A(n2934), .Z(n297) );
  MUX U863 ( .IN0(n298), .IN1(n2445), .SEL(n2446), .F(n2324) );
  IV U864 ( .A(n2447), .Z(n298) );
  MUX U865 ( .IN0(n299), .IN1(n1990), .SEL(n1991), .F(n1885) );
  IV U866 ( .A(n1992), .Z(n299) );
  MUX U867 ( .IN0(n300), .IN1(n1503), .SEL(n1504), .F(n1419) );
  IV U868 ( .A(n1505), .Z(n300) );
  XNOR U869 ( .A(n1271), .B(n1270), .Z(n1289) );
  MUX U870 ( .IN0(n301), .IN1(n1148), .SEL(n1149), .F(n1086) );
  IV U871 ( .A(n1150), .Z(n301) );
  MUX U872 ( .IN0(n302), .IN1(n1023), .SEL(n1024), .F(n970) );
  IV U873 ( .A(n1025), .Z(n302) );
  MUX U874 ( .IN0(n2659), .IN1(n303), .SEL(n2660), .F(n2535) );
  IV U875 ( .A(n2661), .Z(n303) );
  XNOR U876 ( .A(n2428), .B(n2422), .Z(n2538) );
  ANDN U877 ( .A(n2497), .B(n2498), .Z(n2376) );
  MUX U878 ( .IN0(n2185), .IN1(n304), .SEL(n2186), .F(n2076) );
  IV U879 ( .A(n2187), .Z(n304) );
  NANDN U880 ( .B(n2079), .A(n2080), .Z(n1974) );
  ANDN U881 ( .A(n2042), .B(n2043), .Z(n1937) );
  MUX U882 ( .IN0(n1766), .IN1(n305), .SEL(n1767), .F(n1668) );
  IV U883 ( .A(n1768), .Z(n305) );
  ANDN U884 ( .A(n1556), .B(n1557), .Z(n1471) );
  ANDN U885 ( .A(n1252), .B(n1253), .Z(n1185) );
  XNOR U886 ( .A(n691), .B(n690), .Z(n687) );
  XNOR U887 ( .A(n1402), .B(n1484), .Z(n1479) );
  OR U888 ( .A(n1193), .B(n1194), .Z(n1133) );
  XNOR U889 ( .A(n1028), .B(n1027), .Z(n1017) );
  XNOR U890 ( .A(n975), .B(n974), .Z(n959) );
  XNOR U891 ( .A(n834), .B(n833), .Z(n832) );
  XNOR U892 ( .A(n764), .B(n761), .Z(n760) );
  AND U893 ( .A(n823), .B(n824), .Z(n783) );
  MUX U894 ( .IN0(n306), .IN1(n752), .SEL(n753), .F(n720) );
  IV U895 ( .A(\_MxM/Y0[28] ), .Z(n306) );
  XNOR U896 ( .A(n707), .B(n706), .Z(n705) );
  MUX U897 ( .IN0(n307), .IN1(n2621), .SEL(n661), .F(n2499) );
  IV U898 ( .A(\_MxM/Y0[4] ), .Z(n307) );
  MUX U899 ( .IN0(n2149), .IN1(n308), .SEL(n657), .F(n2044) );
  IV U900 ( .A(\_MxM/Y0[8] ), .Z(n308) );
  MUX U901 ( .IN0(n1745), .IN1(n309), .SEL(n1746), .F(n1650) );
  IV U902 ( .A(\_MxM/Y0[12] ), .Z(n309) );
  MUX U903 ( .IN0(n1396), .IN1(n310), .SEL(n1397), .F(n1324) );
  IV U904 ( .A(\_MxM/Y0[16] ), .Z(n310) );
  MUX U905 ( .IN0(n311), .IN1(n1126), .SEL(n1127), .F(n1064) );
  IV U906 ( .A(\_MxM/Y0[20] ), .Z(n311) );
  MUX U907 ( .IN0(n312), .IN1(n906), .SEL(n907), .F(n862) );
  IV U908 ( .A(\_MxM/Y0[24] ), .Z(n312) );
  NAND U909 ( .A(n673), .B(n674), .Z(n672) );
  MUX U910 ( .IN0(n313), .IN1(n4133), .SEL(n4134), .F(n4116) );
  IV U911 ( .A(n4135), .Z(n313) );
  MUX U912 ( .IN0(n3707), .IN1(n3705), .SEL(n3706), .F(n3667) );
  MUX U913 ( .IN0(n314), .IN1(n4136), .SEL(n3770), .F(n4119) );
  IV U914 ( .A(n3769), .Z(n314) );
  MUX U915 ( .IN0(n3726), .IN1(n3728), .SEL(n3727), .F(n3688) );
  XOR U916 ( .A(n4492), .B(n4493), .Z(n4104) );
  MUX U917 ( .IN0(n315), .IN1(n3633), .SEL(n3634), .F(n3595) );
  IV U918 ( .A(n3635), .Z(n315) );
  MUX U919 ( .IN0(n316), .IN1(n3625), .SEL(n3626), .F(n3587) );
  IV U920 ( .A(n3627), .Z(n316) );
  MUX U921 ( .IN0(n4097), .IN1(n4095), .SEL(n4096), .F(n4078) );
  MUX U922 ( .IN0(n317), .IN1(n3646), .SEL(n3647), .F(n3608) );
  IV U923 ( .A(n3648), .Z(n317) );
  XOR U924 ( .A(n4479), .B(n4480), .Z(n4087) );
  MUX U925 ( .IN0(n318), .IN1(n4498), .SEL(n4499), .F(n4485) );
  IV U926 ( .A(n4500), .Z(n318) );
  MUX U927 ( .IN0(n319), .IN1(n4057), .SEL(n4058), .F(n4040) );
  IV U928 ( .A(n4059), .Z(n319) );
  MUX U929 ( .IN0(n320), .IN1(n4048), .SEL(n4049), .F(n4031) );
  IV U930 ( .A(n4050), .Z(n320) );
  MUX U931 ( .IN0(n3641), .IN1(n321), .SEL(n3642), .F(n3603) );
  IV U932 ( .A(n3643), .Z(n321) );
  MUX U933 ( .IN0(n3555), .IN1(n3553), .SEL(n3554), .F(n3515) );
  MUX U934 ( .IN0(n322), .IN1(n4068), .SEL(n3621), .F(n4051) );
  IV U935 ( .A(n3619), .Z(n322) );
  MUX U936 ( .IN0(n3574), .IN1(n3576), .SEL(n3575), .F(n3536) );
  MUX U937 ( .IN0(n323), .IN1(n3481), .SEL(n3482), .F(n3443) );
  IV U938 ( .A(n3483), .Z(n323) );
  MUX U939 ( .IN0(n324), .IN1(n3473), .SEL(n3474), .F(n3435) );
  IV U940 ( .A(n3475), .Z(n324) );
  MUX U941 ( .IN0(n325), .IN1(n4288), .SEL(n4289), .F(n4267) );
  IV U942 ( .A(n4290), .Z(n325) );
  MUX U943 ( .IN0(n326), .IN1(n4614), .SEL(n4615), .F(n4603) );
  IV U944 ( .A(n4616), .Z(n326) );
  MUX U945 ( .IN0(n4450), .IN1(n327), .SEL(n4037), .F(n4437) );
  IV U946 ( .A(n4036), .Z(n327) );
  XNOR U947 ( .A(n4021), .B(n4007), .Z(n4011) );
  MUX U948 ( .IN0(n328), .IN1(n4433), .SEL(n4434), .F(n4420) );
  IV U949 ( .A(n4435), .Z(n328) );
  MUX U950 ( .IN0(n329), .IN1(n3980), .SEL(n3981), .F(n3963) );
  IV U951 ( .A(n3982), .Z(n329) );
  MUX U952 ( .IN0(n3489), .IN1(n330), .SEL(n3490), .F(n3451) );
  IV U953 ( .A(n3491), .Z(n330) );
  MUX U954 ( .IN0(n331), .IN1(n4300), .SEL(n3875), .F(n4279) );
  IV U955 ( .A(n3874), .Z(n331) );
  MUX U956 ( .IN0(n332), .IN1(n4413), .SEL(n4414), .F(n4400) );
  IV U957 ( .A(n4415), .Z(n332) );
  MUX U958 ( .IN0(n333), .IN1(n4865), .SEL(n4712), .F(n4844) );
  IV U959 ( .A(n4711), .Z(n333) );
  XOR U960 ( .A(n4969), .B(n4961), .Z(n4829) );
  MUX U961 ( .IN0(n3403), .IN1(n3401), .SEL(n3402), .F(n3363) );
  MUX U962 ( .IN0(n334), .IN1(n4000), .SEL(n3469), .F(n3983) );
  IV U963 ( .A(n3467), .Z(n334) );
  MUX U964 ( .IN0(n3422), .IN1(n3424), .SEL(n3423), .F(n3384) );
  MUX U965 ( .IN0(n335), .IN1(n3380), .SEL(n3381), .F(n3342) );
  IV U966 ( .A(n3382), .Z(n335) );
  XOR U967 ( .A(n4590), .B(n4582), .Z(n4243) );
  XOR U968 ( .A(n4835), .B(n4817), .Z(n4821) );
  XOR U969 ( .A(n4791), .B(n4792), .Z(n4801) );
  MUX U970 ( .IN0(n336), .IN1(n3329), .SEL(n3330), .F(n3291) );
  IV U971 ( .A(n3331), .Z(n336) );
  MUX U972 ( .IN0(n337), .IN1(n3321), .SEL(n3322), .F(n3283) );
  IV U973 ( .A(n3323), .Z(n337) );
  XNOR U974 ( .A(n3970), .B(n3956), .Z(n3960) );
  MUX U975 ( .IN0(n338), .IN1(n3829), .SEL(n3830), .F(n3814) );
  IV U976 ( .A(n3831), .Z(n338) );
  MUX U977 ( .IN0(n339), .IN1(n4204), .SEL(n4205), .F(n4183) );
  IV U978 ( .A(n4206), .Z(n339) );
  MUX U979 ( .IN0(n4659), .IN1(n4673), .SEL(n4661), .F(n4643) );
  MUX U980 ( .IN0(n340), .IN1(n4689), .SEL(n4690), .F(n4685) );
  IV U981 ( .A(n4691), .Z(n340) );
  XOR U982 ( .A(n4249), .B(n4231), .Z(n4235) );
  MUX U983 ( .IN0(n341), .IN1(n4565), .SEL(n4566), .F(n4554) );
  IV U984 ( .A(n4567), .Z(n341) );
  MUX U985 ( .IN0(n5031), .IN1(n5045), .SEL(n5033), .F(n5015) );
  MUX U986 ( .IN0(n342), .IN1(n5061), .SEL(n5062), .F(n5057) );
  IV U987 ( .A(n5063), .Z(n342) );
  XOR U988 ( .A(n4941), .B(n4942), .Z(n4806) );
  MUX U989 ( .IN0(n343), .IN1(n4934), .SEL(n4935), .F(n4921) );
  IV U990 ( .A(n4936), .Z(n343) );
  XOR U991 ( .A(n4770), .B(n4771), .Z(n4780) );
  MUX U992 ( .IN0(n344), .IN1(n3296), .SEL(n3297), .F(n3258) );
  IV U993 ( .A(n3298), .Z(n344) );
  MUX U994 ( .IN0(n345), .IN1(n3845), .SEL(n3846), .F(n3841) );
  IV U995 ( .A(n3847), .Z(n345) );
  MUX U996 ( .IN0(n346), .IN1(n4310), .SEL(n4311), .F(n4306) );
  IV U997 ( .A(n4312), .Z(n346) );
  MUX U998 ( .IN0(n347), .IN1(n4559), .SEL(n4560), .F(n4548) );
  IV U999 ( .A(n4561), .Z(n347) );
  MUX U1000 ( .IN0(n4385), .IN1(n348), .SEL(n3952), .F(n4372) );
  IV U1001 ( .A(n3951), .Z(n348) );
  MUX U1002 ( .IN0(n349), .IN1(n5076), .SEL(n5077), .F(n5123) );
  IV U1003 ( .A(n5139), .Z(n349) );
  MUX U1004 ( .IN0(n350), .IN1(n4875), .SEL(n4876), .F(n4871) );
  IV U1005 ( .A(n4877), .Z(n350) );
  XOR U1006 ( .A(n4928), .B(n4929), .Z(n4785) );
  XOR U1007 ( .A(n4749), .B(n4750), .Z(n4759) );
  MUX U1008 ( .IN0(n351), .IN1(n4753), .SEL(n4754), .F(n4732) );
  IV U1009 ( .A(n4755), .Z(n351) );
  MUX U1010 ( .IN0(n352), .IN1(n3912), .SEL(n3913), .F(n3892) );
  IV U1011 ( .A(n3914), .Z(n352) );
  MUX U1012 ( .IN0(n3337), .IN1(n353), .SEL(n3338), .F(n3299) );
  IV U1013 ( .A(n3339), .Z(n353) );
  MUX U1014 ( .IN0(n354), .IN1(n4361), .SEL(n4362), .F(n4348) );
  IV U1015 ( .A(n4363), .Z(n354) );
  MUX U1016 ( .IN0(n5095), .IN1(n5110), .SEL(n5097), .F(n5082) );
  MUX U1017 ( .IN0(n355), .IN1(n4901), .SEL(n4902), .F(n4715) );
  IV U1018 ( .A(n4903), .Z(n355) );
  MUX U1019 ( .IN0(n356), .IN1(n4368), .SEL(n4369), .F(n4355) );
  IV U1020 ( .A(n4370), .Z(n356) );
  MUX U1021 ( .IN0(n357), .IN1(n3932), .SEL(n3317), .F(n3915) );
  IV U1022 ( .A(n3315), .Z(n357) );
  XNOR U1023 ( .A(n3919), .B(n3905), .Z(n3909) );
  XOR U1024 ( .A(n3302), .B(n3267), .Z(n3271) );
  XNOR U1025 ( .A(n3251), .B(n3250), .Z(n3263) );
  MUX U1026 ( .IN0(n3856), .IN1(n3859), .SEL(n3857), .F(n3739) );
  MUX U1027 ( .IN0(n358), .IN1(n4142), .SEL(n4143), .F(n4125) );
  IV U1028 ( .A(n4144), .Z(n358) );
  MUX U1029 ( .IN0(n4171), .IN1(n359), .SEL(n4172), .F(n4146) );
  IV U1030 ( .A(n4173), .Z(n359) );
  MUX U1031 ( .IN0(n5072), .IN1(n5100), .SEL(n5074), .F(n3120) );
  XNOR U1032 ( .A(n3213), .B(n3212), .Z(n3225) );
  MUX U1033 ( .IN0(n4541), .IN1(n360), .SEL(n4159), .F(n4528) );
  IV U1034 ( .A(n4157), .Z(n360) );
  MUX U1035 ( .IN0(n361), .IN1(n3137), .SEL(n3138), .F(n3001) );
  IV U1036 ( .A(n3139), .Z(n361) );
  MUX U1037 ( .IN0(n362), .IN1(n3095), .SEL(n3096), .F(n2959) );
  IV U1038 ( .A(n3097), .Z(n362) );
  NAND U1039 ( .A(n4331), .B(n4335), .Z(n4334) );
  MUX U1040 ( .IN0(n363), .IN1(n2975), .SEL(n2976), .F(n2837) );
  IV U1041 ( .A(n2977), .Z(n363) );
  MUX U1042 ( .IN0(n364), .IN1(n2912), .SEL(n2913), .F(n2783) );
  IV U1043 ( .A(n2914), .Z(n364) );
  MUX U1044 ( .IN0(n365), .IN1(n2887), .SEL(n2888), .F(n2758) );
  IV U1045 ( .A(n2889), .Z(n365) );
  MUX U1046 ( .IN0(n366), .IN1(n2929), .SEL(n2930), .F(n2801) );
  IV U1047 ( .A(n2931), .Z(n366) );
  MUX U1048 ( .IN0(n367), .IN1(n2717), .SEL(n2718), .F(n2589) );
  IV U1049 ( .A(n2719), .Z(n367) );
  MUX U1050 ( .IN0(n368), .IN1(n2725), .SEL(n2726), .F(n2597) );
  IV U1051 ( .A(n2727), .Z(n368) );
  MUX U1052 ( .IN0(n369), .IN1(n2564), .SEL(n2565), .F(n2442) );
  IV U1053 ( .A(n2566), .Z(n369) );
  MUX U1054 ( .IN0(n370), .IN1(n2411), .SEL(n2412), .F(n2296) );
  IV U1055 ( .A(n2413), .Z(n370) );
  MUX U1056 ( .IN0(n371), .IN1(n2394), .SEL(n2395), .F(n2283) );
  IV U1057 ( .A(n2396), .Z(n371) );
  MUX U1058 ( .IN0(n372), .IN1(n2236), .SEL(n2237), .F(n2125) );
  IV U1059 ( .A(n2238), .Z(n372) );
  MUX U1060 ( .IN0(n373), .IN1(n2100), .SEL(n2101), .F(n1995) );
  IV U1061 ( .A(n2102), .Z(n373) );
  MUX U1062 ( .IN0(n374), .IN1(n2092), .SEL(n2093), .F(n1987) );
  IV U1063 ( .A(n2094), .Z(n374) );
  MUX U1064 ( .IN0(n375), .IN1(n1898), .SEL(n1899), .F(n1798) );
  IV U1065 ( .A(n1900), .Z(n375) );
  MUX U1066 ( .IN0(n376), .IN1(n1874), .SEL(n1875), .F(n1774) );
  IV U1067 ( .A(n1876), .Z(n376) );
  MUX U1068 ( .IN0(n377), .IN1(n1815), .SEL(n1816), .F(n1719) );
  IV U1069 ( .A(n1817), .Z(n377) );
  MUX U1070 ( .IN0(n378), .IN1(n1686), .SEL(n1687), .F(n1593) );
  IV U1071 ( .A(n1688), .Z(n378) );
  MUX U1072 ( .IN0(n379), .IN1(n1601), .SEL(n1602), .F(n1508) );
  IV U1073 ( .A(n1603), .Z(n379) );
  MUX U1074 ( .IN0(n380), .IN1(n1408), .SEL(n1409), .F(n1335) );
  IV U1075 ( .A(n1410), .Z(n380) );
  MUX U1076 ( .IN0(n381), .IN1(n1441), .SEL(n1442), .F(n1364) );
  IV U1077 ( .A(n1443), .Z(n381) );
  MUX U1078 ( .IN0(n382), .IN1(n1343), .SEL(n1344), .F(n1273) );
  IV U1079 ( .A(n1345), .Z(n382) );
  MUX U1080 ( .IN0(n383), .IN1(n1372), .SEL(n1373), .F(n1300) );
  IV U1081 ( .A(n1374), .Z(n383) );
  MUX U1082 ( .IN0(n384), .IN1(n1381), .SEL(n1382), .F(n1309) );
  IV U1083 ( .A(n1383), .Z(n384) );
  MUX U1084 ( .IN0(n385), .IN1(n1103), .SEL(n1104), .F(n1041) );
  IV U1085 ( .A(n1105), .Z(n385) );
  MUX U1086 ( .IN0(n386), .IN1(n1112), .SEL(n1113), .F(n1050) );
  IV U1087 ( .A(n1114), .Z(n386) );
  MUX U1088 ( .IN0(n387), .IN1(n1005), .SEL(n1006), .F(n947) );
  IV U1089 ( .A(n1007), .Z(n387) );
  XOR U1090 ( .A(n3011), .B(n3145), .Z(n3012) );
  MUX U1091 ( .IN0(n3115), .IN1(n3117), .SEL(n3116), .F(n2979) );
  XNOR U1092 ( .A(n4698), .B(n3088), .Z(n3092) );
  XOR U1093 ( .A(n3159), .B(n3032), .Z(n3036) );
  XNOR U1094 ( .A(n3184), .B(n3058), .Z(n3062) );
  XOR U1095 ( .A(n3076), .B(n3077), .Z(n3083) );
  MUX U1096 ( .IN0(n2519), .IN1(n2521), .SEL(n2520), .F(n2398) );
  XOR U1097 ( .A(n2494), .B(n2614), .Z(n2495) );
  MUX U1098 ( .IN0(n2358), .IN1(n2360), .SEL(n2359), .F(n2240) );
  XOR U1099 ( .A(n1834), .B(n1932), .Z(n1835) );
  MUX U1100 ( .IN0(n1919), .IN1(n1921), .SEL(n1920), .F(n1819) );
  MUX U1101 ( .IN0(n388), .IN1(n1863), .SEL(n1864), .F(n1763) );
  IV U1102 ( .A(n1865), .Z(n388) );
  MUX U1103 ( .IN0(n1205), .IN1(n1203), .SEL(n1204), .F(n1141) );
  MUX U1104 ( .IN0(n1179), .IN1(n1177), .SEL(n1178), .F(n1116) );
  MUX U1105 ( .IN0(n1168), .IN1(n1170), .SEL(n1169), .F(n1107) );
  MUX U1106 ( .IN0(n1139), .IN1(n389), .SEL(n1138), .F(n1079) );
  IV U1107 ( .A(n1137), .Z(n389) );
  MUX U1108 ( .IN0(n390), .IN1(n848), .SEL(n849), .F(n811) );
  IV U1109 ( .A(n850), .Z(n390) );
  XOR U1110 ( .A(n3126), .B(n2993), .Z(n2997) );
  XNOR U1111 ( .A(n3038), .B(n2905), .Z(n2909) );
  MUX U1112 ( .IN0(n2970), .IN1(n391), .SEL(n2971), .F(n2832) );
  IV U1113 ( .A(n2972), .Z(n391) );
  MUX U1114 ( .IN0(n2947), .IN1(n392), .SEL(n2946), .F(n2807) );
  IV U1115 ( .A(n2945), .Z(n392) );
  XNOR U1116 ( .A(n2861), .B(n2735), .Z(n2739) );
  MUX U1117 ( .IN0(n393), .IN1(n2634), .SEL(n2635), .F(n2510) );
  IV U1118 ( .A(n2636), .Z(n393) );
  XNOR U1119 ( .A(n2682), .B(n2557), .Z(n2561) );
  XOR U1120 ( .A(n2706), .B(n2581), .Z(n2585) );
  MUX U1121 ( .IN0(n2541), .IN1(n2539), .SEL(n2540), .F(n2427) );
  XNOR U1122 ( .A(n2522), .B(n2404), .Z(n2408) );
  MUX U1123 ( .IN0(n2453), .IN1(n394), .SEL(n2454), .F(n2332) );
  IV U1124 ( .A(n2455), .Z(n394) );
  XOR U1125 ( .A(n2335), .B(n2220), .Z(n2224) );
  XNOR U1126 ( .A(n2311), .B(n2196), .Z(n2200) );
  XNOR U1127 ( .A(n2361), .B(n2248), .Z(n2252) );
  MUX U1128 ( .IN0(n2160), .IN1(n395), .SEL(n2161), .F(n2057) );
  IV U1129 ( .A(n2162), .Z(n395) );
  MUX U1130 ( .IN0(n2062), .IN1(n2060), .SEL(n2061), .F(n396) );
  IV U1131 ( .A(n396), .Z(n1954) );
  XNOR U1132 ( .A(n2063), .B(n1961), .Z(n1965) );
  MUX U1133 ( .IN0(n397), .IN1(n2120), .SEL(n2121), .F(n2015) );
  IV U1134 ( .A(n2122), .Z(n397) );
  MUX U1135 ( .IN0(n1998), .IN1(n398), .SEL(n1999), .F(n1893) );
  IV U1136 ( .A(n2000), .Z(n398) );
  NAND U1137 ( .A(n1759), .B(n1857), .Z(n1856) );
  XNOR U1138 ( .A(n1922), .B(n1825), .Z(n1829) );
  XNOR U1139 ( .A(n1674), .B(n1586), .Z(n1590) );
  XOR U1140 ( .A(n1700), .B(n1610), .Z(n1614) );
  XOR U1141 ( .A(n1624), .B(n1535), .Z(n1539) );
  XNOR U1142 ( .A(n1633), .B(n1544), .Z(n1548) );
  MUX U1143 ( .IN0(n1511), .IN1(n399), .SEL(n1512), .F(n1427) );
  IV U1144 ( .A(n1513), .Z(n399) );
  XNOR U1145 ( .A(n1359), .B(n1430), .Z(n1360) );
  NAND U1146 ( .A(n1286), .B(n1351), .Z(n1350) );
  MUX U1147 ( .IN0(n400), .IN1(n1295), .SEL(n1296), .F(n1225) );
  IV U1148 ( .A(n1297), .Z(n400) );
  MUX U1149 ( .IN0(n401), .IN1(n1083), .SEL(n1084), .F(n1023) );
  IV U1150 ( .A(n1085), .Z(n401) );
  XNOR U1151 ( .A(n994), .B(n939), .Z(n943) );
  XOR U1152 ( .A(n984), .B(n929), .Z(n934) );
  XNOR U1153 ( .A(n3125), .B(n3124), .Z(n3100) );
  XNOR U1154 ( .A(n2869), .B(n2868), .Z(n2851) );
  MUX U1155 ( .IN0(n402), .IN1(n2804), .SEL(n2805), .F(n2678) );
  IV U1156 ( .A(n2806), .Z(n402) );
  MUX U1157 ( .IN0(n403), .IN1(n1885), .SEL(n1886), .F(n1785) );
  IV U1158 ( .A(n1887), .Z(n403) );
  MUX U1159 ( .IN0(n404), .IN1(n1419), .SEL(n1420), .F(n1346) );
  IV U1160 ( .A(n1421), .Z(n404) );
  ANDN U1161 ( .A(n964), .B(n965), .Z(n963) );
  XOR U1162 ( .A(n765), .B(n803), .Z(n796) );
  MUX U1163 ( .IN0(n2915), .IN1(n405), .SEL(n2916), .F(n2786) );
  IV U1164 ( .A(n2917), .Z(n405) );
  XNOR U1165 ( .A(n2594), .B(n2593), .Z(n2569) );
  MUX U1166 ( .IN0(n2414), .IN1(n406), .SEL(n2415), .F(n2299) );
  IV U1167 ( .A(n2416), .Z(n406) );
  XOR U1168 ( .A(n2302), .B(n2188), .Z(n2189) );
  ANDN U1169 ( .A(n2260), .B(n2261), .Z(n2147) );
  ANDN U1170 ( .A(n1837), .B(n1838), .Z(n1743) );
  ANDN U1171 ( .A(n1394), .B(n1395), .Z(n1322) );
  XOR U1172 ( .A(n1089), .B(n1086), .Z(n1135) );
  XNOR U1173 ( .A(n1038), .B(n1037), .Z(n1028) );
  AND U1174 ( .A(n1008), .B(n1009), .Z(n950) );
  OR U1175 ( .A(n742), .B(n743), .Z(n737) );
  MUX U1176 ( .IN0(n407), .IN1(n747), .SEL(n748), .F(n715) );
  IV U1177 ( .A(n749), .Z(n407) );
  XOR U1178 ( .A(n1869), .B(n1866), .Z(n1944) );
  XNOR U1179 ( .A(n1691), .B(n1690), .Z(n1670) );
  OR U1180 ( .A(n1260), .B(n1261), .Z(n1193) );
  XNOR U1181 ( .A(n1150), .B(n1149), .Z(n1134) );
  OR U1182 ( .A(n958), .B(n959), .Z(n912) );
  XNOR U1183 ( .A(n871), .B(n870), .Z(n869) );
  XNOR U1184 ( .A(n795), .B(n794), .Z(n793) );
  AND U1185 ( .A(n750), .B(n751), .Z(n718) );
  ANDN U1186 ( .A(n687), .B(n686), .Z(n682) );
  MUX U1187 ( .IN0(n2499), .IN1(n408), .SEL(n660), .F(n2378) );
  IV U1188 ( .A(\_MxM/Y0[5] ), .Z(n408) );
  MUX U1189 ( .IN0(n2044), .IN1(n409), .SEL(n656), .F(n1939) );
  IV U1190 ( .A(\_MxM/Y0[9] ), .Z(n409) );
  MUX U1191 ( .IN0(n1650), .IN1(n410), .SEL(n1651), .F(n1558) );
  IV U1192 ( .A(\_MxM/Y0[13] ), .Z(n410) );
  MUX U1193 ( .IN0(n1324), .IN1(n411), .SEL(n1325), .F(n1254) );
  IV U1194 ( .A(\_MxM/Y0[17] ), .Z(n411) );
  MUX U1195 ( .IN0(n412), .IN1(n1064), .SEL(n1065), .F(n1010) );
  IV U1196 ( .A(\_MxM/Y0[21] ), .Z(n412) );
  MUX U1197 ( .IN0(n413), .IN1(n862), .SEL(n863), .F(n825) );
  IV U1198 ( .A(\_MxM/Y0[25] ), .Z(n413) );
  XNOR U1199 ( .A(n720), .B(n721), .Z(n698) );
  OR U1200 ( .A(n704), .B(n705), .Z(n675) );
  MUX U1201 ( .IN0(n414), .IN1(n4108), .SEL(n4109), .F(n4091) );
  IV U1202 ( .A(n4110), .Z(n414) );
  XNOR U1203 ( .A(n3737), .B(n3702), .Z(n3706) );
  XOR U1204 ( .A(n3758), .B(n3723), .Z(n3727) );
  MUX U1205 ( .IN0(n415), .IN1(n3676), .SEL(n3677), .F(n3638) );
  IV U1206 ( .A(n3678), .Z(n415) );
  MUX U1207 ( .IN0(n416), .IN1(n4065), .SEL(n4066), .F(n4048) );
  IV U1208 ( .A(n4067), .Z(n416) );
  MUX U1209 ( .IN0(n4080), .IN1(n4078), .SEL(n4079), .F(n4061) );
  XNOR U1210 ( .A(n3623), .B(n3588), .Z(n3592) );
  MUX U1211 ( .IN0(n4489), .IN1(n417), .SEL(n4088), .F(n4476) );
  IV U1212 ( .A(n4087), .Z(n417) );
  MUX U1213 ( .IN0(n418), .IN1(n3557), .SEL(n3558), .F(n3519) );
  IV U1214 ( .A(n3559), .Z(n418) );
  MUX U1215 ( .IN0(n419), .IN1(n4485), .SEL(n4486), .F(n4472) );
  IV U1216 ( .A(n4487), .Z(n419) );
  MUX U1217 ( .IN0(n420), .IN1(n4040), .SEL(n4041), .F(n4023) );
  IV U1218 ( .A(n4042), .Z(n420) );
  MUX U1219 ( .IN0(n3612), .IN1(n3614), .SEL(n3613), .F(n3574) );
  MUX U1220 ( .IN0(n421), .IN1(n4465), .SEL(n4466), .F(n4452) );
  IV U1221 ( .A(n4467), .Z(n421) );
  MUX U1222 ( .IN0(n422), .IN1(n3524), .SEL(n3525), .F(n3486) );
  IV U1223 ( .A(n3526), .Z(n422) );
  MUX U1224 ( .IN0(n423), .IN1(n3532), .SEL(n3533), .F(n3494) );
  IV U1225 ( .A(n3534), .Z(n423) );
  MUX U1226 ( .IN0(n424), .IN1(n4051), .SEL(n3583), .F(n4034) );
  IV U1227 ( .A(n3581), .Z(n424) );
  MUX U1228 ( .IN0(n3565), .IN1(n425), .SEL(n3566), .F(n3527) );
  IV U1229 ( .A(n3567), .Z(n425) );
  XOR U1230 ( .A(n4427), .B(n4428), .Z(n4019) );
  MUX U1231 ( .IN0(n426), .IN1(n4853), .SEL(n4854), .F(n4832) );
  IV U1232 ( .A(n4855), .Z(n426) );
  MUX U1233 ( .IN0(n427), .IN1(n4858), .SEL(n4859), .F(n4837) );
  IV U1234 ( .A(n4860), .Z(n427) );
  MUX U1235 ( .IN0(n428), .IN1(n3997), .SEL(n3998), .F(n3980) );
  IV U1236 ( .A(n3999), .Z(n428) );
  XNOR U1237 ( .A(n3471), .B(n3436), .Z(n3440) );
  MUX U1238 ( .IN0(n429), .IN1(n4267), .SEL(n4268), .F(n4246) );
  IV U1239 ( .A(n4269), .Z(n429) );
  XOR U1240 ( .A(n4612), .B(n4604), .Z(n4285) );
  MUX U1241 ( .IN0(n430), .IN1(n4272), .SEL(n4273), .F(n4251) );
  IV U1242 ( .A(n4274), .Z(n430) );
  XOR U1243 ( .A(n4414), .B(n4415), .Z(n4002) );
  MUX U1244 ( .IN0(n4990), .IN1(n431), .SEL(n4868), .F(n4977) );
  IV U1245 ( .A(n4867), .Z(n431) );
  MUX U1246 ( .IN0(n432), .IN1(n3405), .SEL(n3406), .F(n3367) );
  IV U1247 ( .A(n3407), .Z(n432) );
  XNOR U1248 ( .A(n4004), .B(n3990), .Z(n3994) );
  MUX U1249 ( .IN0(n3460), .IN1(n3462), .SEL(n3461), .F(n3422) );
  MUX U1250 ( .IN0(n433), .IN1(n4953), .SEL(n4954), .F(n4940) );
  IV U1251 ( .A(n4955), .Z(n433) );
  MUX U1252 ( .IN0(n434), .IN1(n4960), .SEL(n4961), .F(n4947) );
  IV U1253 ( .A(n4962), .Z(n434) );
  MUX U1254 ( .IN0(n435), .IN1(n4420), .SEL(n4421), .F(n4407) );
  IV U1255 ( .A(n4422), .Z(n435) );
  MUX U1256 ( .IN0(n436), .IN1(n3372), .SEL(n3373), .F(n3334) );
  IV U1257 ( .A(n3374), .Z(n436) );
  MUX U1258 ( .IN0(n437), .IN1(n4581), .SEL(n4582), .F(n4570) );
  IV U1259 ( .A(n4583), .Z(n437) );
  XOR U1260 ( .A(n4588), .B(n4589), .Z(n4262) );
  MUX U1261 ( .IN0(n438), .IN1(n3983), .SEL(n3431), .F(n3966) );
  IV U1262 ( .A(n3429), .Z(n438) );
  MUX U1263 ( .IN0(n3413), .IN1(n439), .SEL(n3414), .F(n3375) );
  IV U1264 ( .A(n3415), .Z(n439) );
  XNOR U1265 ( .A(n3357), .B(n3322), .Z(n3326) );
  XOR U1266 ( .A(n4577), .B(n4578), .Z(n4241) );
  MUX U1267 ( .IN0(n4234), .IN1(n440), .SEL(n4235), .F(n4213) );
  IV U1268 ( .A(n4236), .Z(n440) );
  MUX U1269 ( .IN0(n441), .IN1(n4387), .SEL(n4388), .F(n4374) );
  IV U1270 ( .A(n4389), .Z(n441) );
  MUX U1271 ( .IN0(n442), .IN1(n5131), .SEL(n5132), .F(n5113) );
  IV U1272 ( .A(n5133), .Z(n442) );
  XOR U1273 ( .A(n4814), .B(n4796), .Z(n4800) );
  MUX U1274 ( .IN0(n443), .IN1(n4769), .SEL(n4770), .F(n4748) );
  IV U1275 ( .A(n4771), .Z(n443) );
  XNOR U1276 ( .A(n3953), .B(n3939), .Z(n3943) );
  MUX U1277 ( .IN0(n444), .IN1(n3929), .SEL(n3930), .F(n3912) );
  IV U1278 ( .A(n3931), .Z(n444) );
  MUX U1279 ( .IN0(n3814), .IN1(n3828), .SEL(n3816), .F(n3798) );
  MUX U1280 ( .IN0(n445), .IN1(n4183), .SEL(n4184), .F(n4162) );
  IV U1281 ( .A(n4185), .Z(n445) );
  MUX U1282 ( .IN0(n4643), .IN1(n4658), .SEL(n4645), .F(n4620) );
  MUX U1283 ( .IN0(n4637), .IN1(n4652), .SEL(n4639), .F(n4626) );
  XOR U1284 ( .A(n4566), .B(n4567), .Z(n4220) );
  MUX U1285 ( .IN0(n446), .IN1(n4188), .SEL(n4189), .F(n4167) );
  IV U1286 ( .A(n4190), .Z(n446) );
  MUX U1287 ( .IN0(n5015), .IN1(n5030), .SEL(n5017), .F(n4992) );
  MUX U1288 ( .IN0(n5009), .IN1(n5024), .SEL(n5011), .F(n4998) );
  MUX U1289 ( .IN0(n4938), .IN1(n447), .SEL(n4787), .F(n4925) );
  IV U1290 ( .A(n4785), .Z(n447) );
  MUX U1291 ( .IN0(n448), .IN1(n3253), .SEL(n3254), .F(n3215) );
  IV U1292 ( .A(n3255), .Z(n448) );
  XOR U1293 ( .A(n3340), .B(n3305), .Z(n3309) );
  MUX U1294 ( .IN0(n3792), .IN1(n3807), .SEL(n3794), .F(n3781) );
  MUX U1295 ( .IN0(n449), .IN1(n3860), .SEL(n3861), .F(n3856) );
  IV U1296 ( .A(n3862), .Z(n449) );
  XNOR U1297 ( .A(n4690), .B(n4691), .Z(n4677) );
  XOR U1298 ( .A(n4555), .B(n4556), .Z(n4199) );
  NOR U1299 ( .A(g_input[0]), .B(n5180), .Z(n5173) );
  MUX U1300 ( .IN0(n4372), .IN1(n450), .SEL(n3935), .F(n4359) );
  IV U1301 ( .A(n3934), .Z(n450) );
  MUX U1302 ( .IN0(n5101), .IN1(n5118), .SEL(n5103), .F(n5072) );
  XNOR U1303 ( .A(n5062), .B(n5063), .Z(n5049) );
  MUX U1304 ( .IN0(n451), .IN1(n4908), .SEL(n4909), .F(n4895) );
  IV U1305 ( .A(n4910), .Z(n451) );
  MUX U1306 ( .IN0(n452), .IN1(n3220), .SEL(n3221), .F(n3153) );
  IV U1307 ( .A(n3222), .Z(n452) );
  XNOR U1308 ( .A(n3243), .B(n3208), .Z(n3212) );
  XNOR U1309 ( .A(n3846), .B(n3847), .Z(n3832) );
  XNOR U1310 ( .A(n4311), .B(n4312), .Z(n4297) );
  MUX U1311 ( .IN0(n453), .IN1(n4537), .SEL(n4538), .F(n4524) );
  IV U1312 ( .A(n4539), .Z(n453) );
  XOR U1313 ( .A(n4544), .B(n4545), .Z(n4178) );
  XNOR U1314 ( .A(n5152), .B(n5153), .Z(n5139) );
  XNOR U1315 ( .A(n4876), .B(n4877), .Z(n4862) );
  XOR U1316 ( .A(n4751), .B(n4733), .Z(n4737) );
  MUX U1317 ( .IN0(n454), .IN1(n3186), .SEL(n3187), .F(n3057) );
  IV U1318 ( .A(n3188), .Z(n454) );
  MUX U1319 ( .IN0(n455), .IN1(n3915), .SEL(n3279), .F(n3898) );
  IV U1320 ( .A(n3277), .Z(n455) );
  MUX U1321 ( .IN0(n3890), .IN1(n3888), .SEL(n3889), .F(n3190) );
  MUX U1322 ( .IN0(n3261), .IN1(n456), .SEL(n3262), .F(n3223) );
  IV U1323 ( .A(n3263), .Z(n456) );
  MUX U1324 ( .IN0(n4146), .IN1(n457), .SEL(n4147), .F(n4129) );
  IV U1325 ( .A(n4148), .Z(n457) );
  XOR U1326 ( .A(n4533), .B(n4534), .Z(n4157) );
  MUX U1327 ( .IN0(n458), .IN1(n3128), .SEL(n3129), .F(n2992) );
  IV U1328 ( .A(n3130), .Z(n458) );
  MUX U1329 ( .IN0(n459), .IN1(n3103), .SEL(n3104), .F(n2967) );
  IV U1330 ( .A(n3105), .Z(n459) );
  XOR U1331 ( .A(n3879), .B(n3880), .Z(n3896) );
  MUX U1332 ( .IN0(n4341), .IN1(n460), .SEL(n4340), .F(n4331) );
  IV U1333 ( .A(n4339), .Z(n460) );
  XNOR U1334 ( .A(n3176), .B(n3175), .Z(n3158) );
  XOR U1335 ( .A(n3226), .B(n3162), .Z(n3166) );
  MUX U1336 ( .IN0(n461), .IN1(n2959), .SEL(n2960), .F(n2821) );
  IV U1337 ( .A(n2961), .Z(n461) );
  MUX U1338 ( .IN0(n462), .IN1(n2758), .SEL(n2759), .F(n2631) );
  IV U1339 ( .A(n2760), .Z(n462) );
  MUX U1340 ( .IN0(n463), .IN1(n2846), .SEL(n2847), .F(n2717) );
  IV U1341 ( .A(n2848), .Z(n463) );
  MUX U1342 ( .IN0(n464), .IN1(n2656), .SEL(n2657), .F(n2532) );
  IV U1343 ( .A(n2658), .Z(n464) );
  MUX U1344 ( .IN0(n465), .IN1(n2684), .SEL(n2685), .F(n2556) );
  IV U1345 ( .A(n2686), .Z(n465) );
  MUX U1346 ( .IN0(n466), .IN1(n2708), .SEL(n2709), .F(n2580) );
  IV U1347 ( .A(n2710), .Z(n466) );
  MUX U1348 ( .IN0(n467), .IN1(n2572), .SEL(n2573), .F(n2450) );
  IV U1349 ( .A(n2574), .Z(n467) );
  MUX U1350 ( .IN0(n468), .IN1(n2606), .SEL(n2607), .F(n2484) );
  IV U1351 ( .A(n2608), .Z(n468) );
  MUX U1352 ( .IN0(n469), .IN1(n2442), .SEL(n2443), .F(n2321) );
  IV U1353 ( .A(n2444), .Z(n469) );
  MUX U1354 ( .IN0(n470), .IN1(n2801), .SEL(n2802), .F(n2673) );
  IV U1355 ( .A(n2803), .Z(n470) );
  MUX U1356 ( .IN0(n471), .IN1(n2346), .SEL(n2347), .F(n2228) );
  IV U1357 ( .A(n2348), .Z(n471) );
  MUX U1358 ( .IN0(n472), .IN1(n2182), .SEL(n2183), .F(n2073) );
  IV U1359 ( .A(n2184), .Z(n472) );
  MUX U1360 ( .IN0(n473), .IN1(n2219), .SEL(n2220), .F(n2108) );
  IV U1361 ( .A(n2221), .Z(n473) );
  MUX U1362 ( .IN0(n474), .IN1(n2084), .SEL(n2085), .F(n1979) );
  IV U1363 ( .A(n2086), .Z(n474) );
  MUX U1364 ( .IN0(n475), .IN1(n2134), .SEL(n2135), .F(n2029) );
  IV U1365 ( .A(n2136), .Z(n475) );
  MUX U1366 ( .IN0(n476), .IN1(n2270), .SEL(n2271), .F(n2157) );
  IV U1367 ( .A(n2272), .Z(n476) );
  MUX U1368 ( .IN0(n477), .IN1(n1995), .SEL(n1996), .F(n1890) );
  IV U1369 ( .A(n1997), .Z(n477) );
  MUX U1370 ( .IN0(n478), .IN1(n1882), .SEL(n1883), .F(n1782) );
  IV U1371 ( .A(n1884), .Z(n478) );
  MUX U1372 ( .IN0(n479), .IN1(n1907), .SEL(n1908), .F(n1807) );
  IV U1373 ( .A(n1909), .Z(n479) );
  MUX U1374 ( .IN0(n480), .IN1(n1728), .SEL(n1729), .F(n1635) );
  IV U1375 ( .A(n1730), .Z(n480) );
  MUX U1376 ( .IN0(n481), .IN1(n1500), .SEL(n1501), .F(n1416) );
  IV U1377 ( .A(n1502), .Z(n481) );
  MUX U1378 ( .IN0(n482), .IN1(n1492), .SEL(n1493), .F(n1408) );
  IV U1379 ( .A(n1494), .Z(n482) );
  MUX U1380 ( .IN0(n483), .IN1(n1526), .SEL(n1527), .F(n1441) );
  IV U1381 ( .A(n1528), .Z(n483) );
  MUX U1382 ( .IN0(n484), .IN1(n1534), .SEL(n1535), .F(n1449) );
  IV U1383 ( .A(n1536), .Z(n484) );
  MUX U1384 ( .IN0(n485), .IN1(n1222), .SEL(n1223), .F(n1156) );
  IV U1385 ( .A(n1224), .Z(n485) );
  MUX U1386 ( .IN0(n486), .IN1(n1121), .SEL(n1122), .F(n1059) );
  IV U1387 ( .A(n1123), .Z(n486) );
  MUX U1388 ( .IN0(n487), .IN1(n978), .SEL(n979), .F(n921) );
  IV U1389 ( .A(n980), .Z(n487) );
  MUX U1390 ( .IN0(n488), .IN1(n938), .SEL(n939), .F(n890) );
  IV U1391 ( .A(n940), .Z(n488) );
  MUX U1392 ( .IN0(n489), .IN1(n901), .SEL(n902), .F(n857) );
  IV U1393 ( .A(n903), .Z(n489) );
  XNOR U1394 ( .A(n3745), .B(n3744), .Z(n3757) );
  MUX U1395 ( .IN0(n2341), .IN1(n2343), .SEL(n2342), .F(n2223) );
  MUX U1396 ( .IN0(n1613), .IN1(n1615), .SEL(n1614), .F(n1515) );
  MUX U1397 ( .IN0(n1641), .IN1(n1639), .SEL(n1640), .F(n1547) );
  XOR U1398 ( .A(n1468), .B(n1551), .Z(n1469) );
  MUX U1399 ( .IN0(n1523), .IN1(n490), .SEL(n1522), .F(n1435) );
  IV U1400 ( .A(n1521), .Z(n490) );
  MUX U1401 ( .IN0(n930), .IN1(n491), .SEL(n929), .F(n886) );
  IV U1402 ( .A(n928), .Z(n491) );
  XNOR U1403 ( .A(n3085), .B(n2952), .Z(n2956) );
  XOR U1404 ( .A(n3109), .B(n2976), .Z(n2980) );
  XNOR U1405 ( .A(n3143), .B(n3142), .Z(n3125) );
  XNOR U1406 ( .A(n3046), .B(n3045), .Z(n3028) );
  XNOR U1407 ( .A(n2902), .B(n2776), .Z(n2780) );
  XOR U1408 ( .A(n2893), .B(n2767), .Z(n2771) );
  XNOR U1409 ( .A(n2919), .B(n2798), .Z(n2792) );
  XOR U1410 ( .A(n2852), .B(n2726), .Z(n2730) );
  MUX U1411 ( .IN0(n2703), .IN1(n492), .SEL(n2704), .F(n2575) );
  IV U1412 ( .A(n2705), .Z(n492) );
  MUX U1413 ( .IN0(n493), .IN1(n2510), .SEL(n2511), .F(n2389) );
  IV U1414 ( .A(n2512), .Z(n493) );
  XOR U1415 ( .A(n2392), .B(n2284), .Z(n2278) );
  XNOR U1416 ( .A(n2401), .B(n2289), .Z(n2293) );
  XOR U1417 ( .A(n2473), .B(n2355), .Z(n2359) );
  XNOR U1418 ( .A(n2432), .B(n2314), .Z(n2318) );
  NAND U1419 ( .A(n2424), .B(n2543), .Z(n2542) );
  MUX U1420 ( .IN0(n2214), .IN1(n494), .SEL(n2215), .F(n2103) );
  IV U1421 ( .A(n2216), .Z(n494) );
  NAND U1422 ( .A(n1949), .B(n2052), .Z(n2051) );
  XOR U1423 ( .A(n2123), .B(n2021), .Z(n2025) );
  XNOR U1424 ( .A(n1958), .B(n1860), .Z(n1854) );
  XOR U1425 ( .A(n2001), .B(n1899), .Z(n1903) );
  XNOR U1426 ( .A(n1872), .B(n1775), .Z(n1779) );
  XOR U1427 ( .A(n1813), .B(n1720), .Z(n1724) );
  MUX U1428 ( .IN0(n1697), .IN1(n495), .SEL(n1698), .F(n1604) );
  IV U1429 ( .A(n1699), .Z(n495) );
  MUX U1430 ( .IN0(n496), .IN1(n1763), .SEL(n1764), .F(n1665) );
  IV U1431 ( .A(n1765), .Z(n496) );
  XNOR U1432 ( .A(n1333), .B(n1266), .Z(n1270) );
  XOR U1433 ( .A(n1370), .B(n1301), .Z(n1305) );
  XNOR U1434 ( .A(n1379), .B(n1310), .Z(n1314) );
  OR U1435 ( .A(n1280), .B(n1281), .Z(n1218) );
  XNOR U1436 ( .A(n1171), .B(n1113), .Z(n1117) );
  XOR U1437 ( .A(n1162), .B(n1104), .Z(n1108) );
  MUX U1438 ( .IN0(n497), .IN1(n924), .SEL(n925), .F(n878) );
  IV U1439 ( .A(n926), .Z(n497) );
  XNOR U1440 ( .A(n846), .B(n812), .Z(n816) );
  AND U1441 ( .A(n804), .B(n803), .Z(n800) );
  XNOR U1442 ( .A(n3007), .B(n3006), .Z(n2989) );
  XNOR U1443 ( .A(n2807), .B(n2935), .Z(n2808) );
  MUX U1444 ( .IN0(n498), .IN1(n2824), .SEL(n2825), .F(n2695) );
  IV U1445 ( .A(n2826), .Z(n498) );
  XNOR U1446 ( .A(n2740), .B(n2739), .Z(n2722) );
  MUX U1447 ( .IN0(n2680), .IN1(n499), .SEL(n2679), .F(n2550) );
  IV U1448 ( .A(n2678), .Z(n499) );
  XNOR U1449 ( .A(n2369), .B(n2368), .Z(n2351) );
  XNOR U1450 ( .A(n1966), .B(n1965), .Z(n1957) );
  XNOR U1451 ( .A(n2035), .B(n2034), .Z(n2017) );
  XNOR U1452 ( .A(n1736), .B(n1735), .Z(n1716) );
  XNOR U1453 ( .A(n1341), .B(n1340), .Z(n1358) );
  XNOR U1454 ( .A(n1205), .B(n1204), .Z(n1217) );
  XNOR U1455 ( .A(n1245), .B(n1244), .Z(n1227) );
  XNOR U1456 ( .A(n1143), .B(n1142), .Z(n1153) );
  XNOR U1457 ( .A(n1077), .B(n1076), .Z(n1092) );
  XNOR U1458 ( .A(n1021), .B(n1020), .Z(n1030) );
  XNOR U1459 ( .A(n969), .B(n968), .Z(n965) );
  XNOR U1460 ( .A(n777), .B(n776), .Z(n767) );
  MUX U1461 ( .IN0(n2535), .IN1(n500), .SEL(n2536), .F(n2414) );
  IV U1462 ( .A(n2537), .Z(n500) );
  XNOR U1463 ( .A(n2472), .B(n2471), .Z(n2447) );
  XNOR U1464 ( .A(n2233), .B(n2232), .Z(n2208) );
  MUX U1465 ( .IN0(n2188), .IN1(n2302), .SEL(n2190), .F(n2079) );
  XNOR U1466 ( .A(n1912), .B(n1911), .Z(n1887) );
  XNOR U1467 ( .A(n1812), .B(n1811), .Z(n1787) );
  ANDN U1468 ( .A(n1937), .B(n1938), .Z(n1837) );
  NANDN U1469 ( .B(n1565), .A(n1566), .Z(n1484) );
  XNOR U1470 ( .A(n1369), .B(n1368), .Z(n1348) );
  XNOR U1471 ( .A(n1161), .B(n1160), .Z(n1150) );
  XNOR U1472 ( .A(n983), .B(n982), .Z(n975) );
  XNOR U1473 ( .A(n842), .B(n841), .Z(n834) );
  XNOR U1474 ( .A(n2097), .B(n2096), .Z(n2078) );
  XOR U1475 ( .A(n1769), .B(n1766), .Z(n1845) );
  XNOR U1476 ( .A(n1598), .B(n1597), .Z(n1581) );
  XNOR U1477 ( .A(n1505), .B(n1504), .Z(n1488) );
  MUX U1478 ( .IN0(n712), .IN1(n710), .SEL(n711), .F(n690) );
  AND U1479 ( .A(n718), .B(n719), .Z(n673) );
  XOR U1480 ( .A(n1261), .B(n1260), .Z(n1327) );
  XNOR U1481 ( .A(n1071), .B(n1070), .Z(n1130) );
  XNOR U1482 ( .A(n913), .B(n912), .Z(n955) );
  XNOR U1483 ( .A(n793), .B(n792), .Z(n828) );
  ANDN U1484 ( .A(n676), .B(n675), .Z(n669) );
  MUX U1485 ( .IN0(\_MxM/Y0[30] ), .IN1(n698), .SEL(n697), .F(n665) );
  XOR U1486 ( .A(n2747), .B(n2750), .Z(n2748) );
  XOR U1487 ( .A(n2378), .B(n2381), .Z(n2379) );
  XOR U1488 ( .A(n2044), .B(n2047), .Z(n2045) );
  XOR U1489 ( .A(n1745), .B(n1749), .Z(n1747) );
  XOR U1490 ( .A(n1473), .B(n1477), .Z(n1475) );
  XOR U1491 ( .A(n1254), .B(n1258), .Z(n1256) );
  XOR U1492 ( .A(n1064), .B(n1068), .Z(n1066) );
  XOR U1493 ( .A(n906), .B(n910), .Z(n908) );
  MUX U1494 ( .IN0(n501), .IN1(n3747), .SEL(n3748), .F(n3709) );
  IV U1495 ( .A(n3749), .Z(n501) );
  MUX U1496 ( .IN0(n502), .IN1(n3701), .SEL(n3702), .F(n3663) );
  IV U1497 ( .A(n3703), .Z(n502) );
  XOR U1498 ( .A(n4505), .B(n4506), .Z(n4121) );
  MUX U1499 ( .IN0(n503), .IN1(n4099), .SEL(n4100), .F(n4082) );
  IV U1500 ( .A(n4101), .Z(n503) );
  XNOR U1501 ( .A(n4106), .B(n4092), .Z(n4096) );
  MUX U1502 ( .IN0(n504), .IN1(n3595), .SEL(n3596), .F(n3557) );
  IV U1503 ( .A(n3597), .Z(n504) );
  MUX U1504 ( .IN0(n3631), .IN1(n3629), .SEL(n3630), .F(n3591) );
  MUX U1505 ( .IN0(n3650), .IN1(n3652), .SEL(n3651), .F(n3612) );
  MUX U1506 ( .IN0(n3679), .IN1(n505), .SEL(n3680), .F(n3641) );
  IV U1507 ( .A(n3681), .Z(n505) );
  MUX U1508 ( .IN0(n506), .IN1(n4478), .SEL(n4479), .F(n4465) );
  IV U1509 ( .A(n4480), .Z(n506) );
  MUX U1510 ( .IN0(n507), .IN1(n3549), .SEL(n3550), .F(n3511) );
  IV U1511 ( .A(n3551), .Z(n507) );
  MUX U1512 ( .IN0(n508), .IN1(n3562), .SEL(n3563), .F(n3524) );
  IV U1513 ( .A(n3564), .Z(n508) );
  MUX U1514 ( .IN0(n509), .IN1(n3570), .SEL(n3571), .F(n3532) );
  IV U1515 ( .A(n3572), .Z(n509) );
  MUX U1516 ( .IN0(n510), .IN1(n4472), .SEL(n4473), .F(n4459) );
  IV U1517 ( .A(n4474), .Z(n510) );
  XNOR U1518 ( .A(n4055), .B(n4041), .Z(n4045) );
  MUX U1519 ( .IN0(n511), .IN1(n4031), .SEL(n4032), .F(n4014) );
  IV U1520 ( .A(n4033), .Z(n511) );
  MUX U1521 ( .IN0(n4463), .IN1(n512), .SEL(n4054), .F(n4450) );
  IV U1522 ( .A(n4053), .Z(n512) );
  MUX U1523 ( .IN0(n513), .IN1(n3443), .SEL(n3444), .F(n3405) );
  IV U1524 ( .A(n3445), .Z(n513) );
  MUX U1525 ( .IN0(n3479), .IN1(n3477), .SEL(n3478), .F(n3439) );
  MUX U1526 ( .IN0(n514), .IN1(n4034), .SEL(n3545), .F(n4017) );
  IV U1527 ( .A(n3543), .Z(n514) );
  MUX U1528 ( .IN0(n3498), .IN1(n3500), .SEL(n3499), .F(n3460) );
  MUX U1529 ( .IN0(n3527), .IN1(n515), .SEL(n3528), .F(n3489) );
  IV U1530 ( .A(n3529), .Z(n515) );
  MUX U1531 ( .IN0(n516), .IN1(n4426), .SEL(n4427), .F(n4413) );
  IV U1532 ( .A(n4428), .Z(n516) );
  XOR U1533 ( .A(n4833), .B(n4834), .Z(n4843) );
  MUX U1534 ( .IN0(n517), .IN1(n3397), .SEL(n3398), .F(n3359) );
  IV U1535 ( .A(n3399), .Z(n517) );
  MUX U1536 ( .IN0(n518), .IN1(n3410), .SEL(n3411), .F(n3372) );
  IV U1537 ( .A(n3412), .Z(n518) );
  MUX U1538 ( .IN0(n519), .IN1(n3418), .SEL(n3419), .F(n3380) );
  IV U1539 ( .A(n3420), .Z(n519) );
  MUX U1540 ( .IN0(n520), .IN1(n4246), .SEL(n4247), .F(n4225) );
  IV U1541 ( .A(n4248), .Z(n520) );
  XOR U1542 ( .A(n4599), .B(n4600), .Z(n4283) );
  XOR U1543 ( .A(n4967), .B(n4968), .Z(n4848) );
  XOR U1544 ( .A(n4812), .B(n4813), .Z(n4822) );
  MUX U1545 ( .IN0(n521), .IN1(n4816), .SEL(n4817), .F(n4795) );
  IV U1546 ( .A(n4818), .Z(n521) );
  XNOR U1547 ( .A(n3987), .B(n3973), .Z(n3977) );
  MUX U1548 ( .IN0(n522), .IN1(n3963), .SEL(n3964), .F(n3946) );
  IV U1549 ( .A(n3965), .Z(n522) );
  MUX U1550 ( .IN0(n4411), .IN1(n523), .SEL(n3986), .F(n4398) );
  IV U1551 ( .A(n3985), .Z(n523) );
  MUX U1552 ( .IN0(n524), .IN1(n4940), .SEL(n4941), .F(n4927) );
  IV U1553 ( .A(n4942), .Z(n524) );
  MUX U1554 ( .IN0(n525), .IN1(n4407), .SEL(n4408), .F(n4394) );
  IV U1555 ( .A(n4409), .Z(n525) );
  XOR U1556 ( .A(n4579), .B(n4571), .Z(n4222) );
  MUX U1557 ( .IN0(n526), .IN1(n3291), .SEL(n3292), .F(n3253) );
  IV U1558 ( .A(n3293), .Z(n526) );
  MUX U1559 ( .IN0(n3327), .IN1(n3325), .SEL(n3326), .F(n3287) );
  MUX U1560 ( .IN0(n527), .IN1(n3966), .SEL(n3393), .F(n3949) );
  IV U1561 ( .A(n3391), .Z(n527) );
  MUX U1562 ( .IN0(n3346), .IN1(n3348), .SEL(n3347), .F(n3308) );
  MUX U1563 ( .IN0(n3375), .IN1(n528), .SEL(n3376), .F(n3337) );
  IV U1564 ( .A(n3377), .Z(n528) );
  MUX U1565 ( .IN0(n4685), .IN1(n4688), .SEL(n4686), .F(n4669) );
  XOR U1566 ( .A(n4228), .B(n4210), .Z(n4214) );
  MUX U1567 ( .IN0(n529), .IN1(n4554), .SEL(n4555), .F(n4543) );
  IV U1568 ( .A(n4556), .Z(n529) );
  XOR U1569 ( .A(n4362), .B(n4363), .Z(n3934) );
  MUX U1570 ( .IN0(n5057), .IN1(n5060), .SEL(n5058), .F(n5041) );
  XOR U1571 ( .A(n4930), .B(n4922), .Z(n4766) );
  MUX U1572 ( .IN0(n530), .IN1(n4748), .SEL(n4749), .F(n4727) );
  IV U1573 ( .A(n4750), .Z(n530) );
  MUX U1574 ( .IN0(n531), .IN1(n3245), .SEL(n3246), .F(n3207) );
  IV U1575 ( .A(n3247), .Z(n531) );
  XNOR U1576 ( .A(n3936), .B(n3922), .Z(n3926) );
  MUX U1577 ( .IN0(n532), .IN1(n3258), .SEL(n3259), .F(n3220) );
  IV U1578 ( .A(n3260), .Z(n532) );
  MUX U1579 ( .IN0(n533), .IN1(n3266), .SEL(n3267), .F(n3228) );
  IV U1580 ( .A(n3268), .Z(n533) );
  MUX U1581 ( .IN0(n3798), .IN1(n3813), .SEL(n3800), .F(n3773) );
  MUX U1582 ( .IN0(n3841), .IN1(n3844), .SEL(n3842), .F(n3824) );
  MUX U1583 ( .IN0(n534), .IN1(n4162), .SEL(n4163), .F(n4150) );
  IV U1584 ( .A(n4164), .Z(n534) );
  MUX U1585 ( .IN0(n4626), .IN1(n4636), .SEL(n4628), .F(n4614) );
  XOR U1586 ( .A(n4349), .B(n4350), .Z(n3917) );
  MUX U1587 ( .IN0(n535), .IN1(n5168), .SEL(n5169), .F(n5164) );
  IV U1588 ( .A(n5170), .Z(n535) );
  MUX U1589 ( .IN0(n5147), .IN1(n5150), .SEL(n5148), .F(n5131) );
  MUX U1590 ( .IN0(n4998), .IN1(n5008), .SEL(n5000), .F(n4986) );
  XOR U1591 ( .A(n4772), .B(n4754), .Z(n4758) );
  MUX U1592 ( .IN0(n536), .IN1(n3892), .SEL(n3893), .F(n3194) );
  IV U1593 ( .A(n3894), .Z(n536) );
  MUX U1594 ( .IN0(n3781), .IN1(n3791), .SEL(n3783), .F(n3760) );
  XOR U1595 ( .A(n4675), .B(n4676), .Z(n4324) );
  XOR U1596 ( .A(n4546), .B(n4538), .Z(n4159) );
  XOR U1597 ( .A(n5047), .B(n5048), .Z(n4889) );
  XOR U1598 ( .A(n4902), .B(n4903), .Z(n4743) );
  MUX U1599 ( .IN0(n537), .IN1(n4895), .SEL(n4896), .F(n3111) );
  IV U1600 ( .A(n4897), .Z(n537) );
  MUX U1601 ( .IN0(n538), .IN1(n4355), .SEL(n4356), .F(n4339) );
  IV U1602 ( .A(n4357), .Z(n538) );
  XOR U1603 ( .A(n3830), .B(n3831), .Z(n3777) );
  XNOR U1604 ( .A(n3861), .B(n3862), .Z(n3743) );
  XNOR U1605 ( .A(n4304), .B(n4294), .Z(n4298) );
  XOR U1606 ( .A(n4610), .B(n4611), .Z(n4302) );
  XOR U1607 ( .A(n4165), .B(n4143), .Z(n4147) );
  XOR U1608 ( .A(n5162), .B(g_input[3]), .Z(n5163) );
  MUX U1609 ( .IN0(n539), .IN1(n3120), .SEL(n3121), .F(n2984) );
  IV U1610 ( .A(n3122), .Z(n539) );
  MUX U1611 ( .IN0(n540), .IN1(n3087), .SEL(n3088), .F(n2951) );
  IV U1612 ( .A(n3089), .Z(n540) );
  MUX U1613 ( .IN0(n541), .IN1(n3048), .SEL(n3049), .F(n2912) );
  IV U1614 ( .A(n3050), .Z(n541) );
  XOR U1615 ( .A(n5137), .B(n5138), .Z(n5076) );
  XNOR U1616 ( .A(n4869), .B(n4859), .Z(n4863) );
  XOR U1617 ( .A(n4980), .B(n4981), .Z(n4867) );
  XOR U1618 ( .A(n4716), .B(n4717), .Z(n4722) );
  MUX U1619 ( .IN0(n3176), .IN1(n3174), .SEL(n3175), .F(n3044) );
  MUX U1620 ( .IN0(n3165), .IN1(n3167), .SEL(n3166), .F(n3035) );
  MUX U1621 ( .IN0(n542), .IN1(n3898), .SEL(n3241), .F(n3881) );
  IV U1622 ( .A(n3239), .Z(n542) );
  XNOR U1623 ( .A(n3882), .B(n3187), .Z(n3191) );
  MUX U1624 ( .IN0(n3223), .IN1(n543), .SEL(n3224), .F(n3156) );
  IV U1625 ( .A(n3225), .Z(n543) );
  XOR U1626 ( .A(n4518), .B(n4519), .Z(n4138) );
  MUX U1627 ( .IN0(n544), .IN1(n2904), .SEL(n2905), .F(n2775) );
  IV U1628 ( .A(n2906), .Z(n544) );
  MUX U1629 ( .IN0(n545), .IN1(n2895), .SEL(n2896), .F(n2766) );
  IV U1630 ( .A(n2897), .Z(n545) );
  MUX U1631 ( .IN0(n546), .IN1(n3878), .SEL(n3879), .F(n3075) );
  IV U1632 ( .A(n3880), .Z(n546) );
  MUX U1633 ( .IN0(n547), .IN1(n2829), .SEL(n2830), .F(n2700) );
  IV U1634 ( .A(n2831), .Z(n547) );
  MUX U1635 ( .IN0(n548), .IN1(n2863), .SEL(n2864), .F(n2734) );
  IV U1636 ( .A(n2865), .Z(n548) );
  MUX U1637 ( .IN0(n549), .IN1(n2507), .SEL(n2508), .F(n2386) );
  IV U1638 ( .A(n2509), .Z(n549) );
  MUX U1639 ( .IN0(n550), .IN1(n2556), .SEL(n2557), .F(n2434) );
  IV U1640 ( .A(n2558), .Z(n550) );
  MUX U1641 ( .IN0(n551), .IN1(n2589), .SEL(n2590), .F(n2467) );
  IV U1642 ( .A(n2591), .Z(n551) );
  MUX U1643 ( .IN0(n552), .IN1(n2296), .SEL(n2297), .F(n2182) );
  IV U1644 ( .A(n2298), .Z(n552) );
  MUX U1645 ( .IN0(n553), .IN1(n2329), .SEL(n2330), .F(n2211) );
  IV U1646 ( .A(n2331), .Z(n553) );
  MUX U1647 ( .IN0(n554), .IN1(n2363), .SEL(n2364), .F(n2245) );
  IV U1648 ( .A(n2365), .Z(n554) );
  MUX U1649 ( .IN0(n555), .IN1(n2117), .SEL(n2118), .F(n2012) );
  IV U1650 ( .A(n2119), .Z(n555) );
  MUX U1651 ( .IN0(n556), .IN1(n1890), .SEL(n1891), .F(n1790) );
  IV U1652 ( .A(n1892), .Z(n556) );
  MUX U1653 ( .IN0(n557), .IN1(n1924), .SEL(n1925), .F(n1824) );
  IV U1654 ( .A(n1926), .Z(n557) );
  MUX U1655 ( .IN0(n558), .IN1(n1719), .SEL(n1720), .F(n1626) );
  IV U1656 ( .A(n1721), .Z(n558) );
  MUX U1657 ( .IN0(n559), .IN1(n1711), .SEL(n1712), .F(n1618) );
  IV U1658 ( .A(n1713), .Z(n559) );
  MUX U1659 ( .IN0(n560), .IN1(n1676), .SEL(n1677), .F(n1585) );
  IV U1660 ( .A(n1678), .Z(n560) );
  MUX U1661 ( .IN0(n561), .IN1(n1593), .SEL(n1594), .F(n1500) );
  IV U1662 ( .A(n1595), .Z(n561) );
  MUX U1663 ( .IN0(n562), .IN1(n1508), .SEL(n1509), .F(n1424) );
  IV U1664 ( .A(n1510), .Z(n562) );
  MUX U1665 ( .IN0(n563), .IN1(n1543), .SEL(n1544), .F(n1458) );
  IV U1666 ( .A(n1545), .Z(n563) );
  MUX U1667 ( .IN0(n564), .IN1(n1364), .SEL(n1365), .F(n1292) );
  IV U1668 ( .A(n1366), .Z(n564) );
  MUX U1669 ( .IN0(n565), .IN1(n1273), .SEL(n1274), .F(n1207) );
  IV U1670 ( .A(n1275), .Z(n565) );
  MUX U1671 ( .IN0(n566), .IN1(n1095), .SEL(n1096), .F(n1033) );
  IV U1672 ( .A(n1097), .Z(n566) );
  MUX U1673 ( .IN0(n567), .IN1(n947), .SEL(n948), .F(n901) );
  IV U1674 ( .A(n949), .Z(n567) );
  MUX U1675 ( .IN0(n3093), .IN1(n3091), .SEL(n3092), .F(n2955) );
  XOR U1676 ( .A(n5078), .B(n3129), .Z(n3133) );
  XNOR U1677 ( .A(n4131), .B(n4130), .Z(n3769) );
  MUX U1678 ( .IN0(n3007), .IN1(n3005), .SEL(n3006), .F(n2867) );
  MUX U1679 ( .IN0(n2490), .IN1(n2488), .SEL(n2489), .F(n2367) );
  MUX U1680 ( .IN0(n1830), .IN1(n1828), .SEL(n1829), .F(n1732) );
  MUX U1681 ( .IN0(n1780), .IN1(n1778), .SEL(n1779), .F(n1680) );
  MUX U1682 ( .IN0(n1861), .IN1(n568), .SEL(n1860), .F(n1759) );
  IV U1683 ( .A(n1859), .Z(n568) );
  MUX U1684 ( .IN0(n569), .IN1(n875), .SEL(n876), .F(n837) );
  IV U1685 ( .A(n877), .Z(n569) );
  MUX U1686 ( .IN0(n3083), .IN1(n570), .SEL(n3082), .F(n2944) );
  IV U1687 ( .A(n3081), .Z(n570) );
  XNOR U1688 ( .A(n3063), .B(n3062), .Z(n3080) );
  XNOR U1689 ( .A(n3757), .B(n3756), .Z(n3181) );
  XOR U1690 ( .A(n2973), .B(n2838), .Z(n2842) );
  XOR U1691 ( .A(n2790), .B(n2669), .Z(n2670) );
  XOR U1692 ( .A(n2637), .B(n2516), .Z(n2520) );
  XNOR U1693 ( .A(n2646), .B(n2525), .Z(n2529) );
  XOR U1694 ( .A(n2723), .B(n2598), .Z(n2602) );
  XOR U1695 ( .A(n2578), .B(n2459), .Z(n2463) );
  MUX U1696 ( .IN0(n2547), .IN1(n571), .SEL(n2546), .F(n2424) );
  IV U1697 ( .A(n2545), .Z(n571) );
  NAND U1698 ( .A(n2168), .B(n2281), .Z(n2280) );
  XNOR U1699 ( .A(n2286), .B(n2175), .Z(n2179) );
  XOR U1700 ( .A(n2352), .B(n2237), .Z(n2241) );
  XNOR U1701 ( .A(n2193), .B(n2085), .Z(n2089) );
  XOR U1702 ( .A(n2217), .B(n2109), .Z(n2113) );
  MUX U1703 ( .IN0(n2056), .IN1(n572), .SEL(n2055), .F(n1949) );
  IV U1704 ( .A(n2054), .Z(n572) );
  XOR U1705 ( .A(n2018), .B(n1916), .Z(n1920) );
  XOR U1706 ( .A(n1764), .B(n1765), .Z(n1761) );
  XOR U1707 ( .A(n1896), .B(n1799), .Z(n1803) );
  XOR U1708 ( .A(n1607), .B(n1522), .Z(n1516) );
  XOR U1709 ( .A(n1666), .B(n1667), .Z(n1661) );
  XNOR U1710 ( .A(n1490), .B(n1409), .Z(n1413) );
  XOR U1711 ( .A(n1532), .B(n1450), .Z(n1454) );
  XNOR U1712 ( .A(n1263), .B(n1200), .Z(n1204) );
  XNOR U1713 ( .A(n1307), .B(n1240), .Z(n1244) );
  XOR U1714 ( .A(n1298), .B(n1231), .Z(n1235) );
  XOR U1715 ( .A(n1101), .B(n1042), .Z(n1046) );
  XNOR U1716 ( .A(n1110), .B(n1051), .Z(n1055) );
  XOR U1717 ( .A(n927), .B(n886), .Z(n884) );
  XNOR U1718 ( .A(n888), .B(n849), .Z(n853) );
  XNOR U1719 ( .A(n2927), .B(n2926), .Z(n2947) );
  XNOR U1720 ( .A(n3028), .B(n3027), .Z(n3070) );
  XNOR U1721 ( .A(n2819), .B(n2818), .Z(n2834) );
  XNOR U1722 ( .A(n2781), .B(n2780), .Z(n2763) );
  XNOR U1723 ( .A(n2793), .B(n2792), .Z(n2809) );
  XNOR U1724 ( .A(n2654), .B(n2653), .Z(n2636) );
  XNOR U1725 ( .A(n2690), .B(n2689), .Z(n2705) );
  XNOR U1726 ( .A(n2612), .B(n2611), .Z(n2594) );
  XNOR U1727 ( .A(n2562), .B(n2561), .Z(n2577) );
  XNOR U1728 ( .A(n2319), .B(n2318), .Z(n2334) );
  XNOR U1729 ( .A(n2201), .B(n2200), .Z(n2216) );
  XNOR U1730 ( .A(n2253), .B(n2252), .Z(n2233) );
  XNOR U1731 ( .A(n2071), .B(n2070), .Z(n2059) );
  XNOR U1732 ( .A(n1985), .B(n1984), .Z(n2000) );
  XNOR U1733 ( .A(n1855), .B(n1854), .Z(n1848) );
  XNOR U1734 ( .A(n1930), .B(n1929), .Z(n1912) );
  XNOR U1735 ( .A(n1880), .B(n1879), .Z(n1895) );
  XNOR U1736 ( .A(n1641), .B(n1640), .Z(n1623) );
  MUX U1737 ( .IN0(n573), .IN1(n1689), .SEL(n1690), .F(n1596) );
  IV U1738 ( .A(n1691), .Z(n573) );
  XNOR U1739 ( .A(n1464), .B(n1463), .Z(n1446) );
  XNOR U1740 ( .A(n1387), .B(n1386), .Z(n1369) );
  XOR U1741 ( .A(n1280), .B(n1287), .Z(n1349) );
  XNOR U1742 ( .A(n1179), .B(n1178), .Z(n1161) );
  NOR U1743 ( .A(n1029), .B(n1030), .Z(n964) );
  XNOR U1744 ( .A(n1002), .B(n1001), .Z(n983) );
  ANDN U1745 ( .A(n969), .B(n968), .Z(n967) );
  MUX U1746 ( .IN0(n767), .IN1(n765), .SEL(n766), .F(n733) );
  MUX U1747 ( .IN0(n772), .IN1(n574), .SEL(n771), .F(n742) );
  IV U1748 ( .A(n770), .Z(n574) );
  MUX U1749 ( .IN0(n575), .IN1(n780), .SEL(n781), .F(n747) );
  IV U1750 ( .A(n782), .Z(n575) );
  XNOR U1751 ( .A(n2892), .B(n2891), .Z(n2934) );
  XNOR U1752 ( .A(n3100), .B(n3099), .Z(n3053) );
  XNOR U1753 ( .A(n2851), .B(n2850), .Z(n2826) );
  XNOR U1754 ( .A(n2722), .B(n2721), .Z(n2697) );
  XNOR U1755 ( .A(n2391), .B(n2390), .Z(n2430) );
  XNOR U1756 ( .A(n2275), .B(n2274), .Z(n2305) );
  XNOR U1757 ( .A(n2351), .B(n2350), .Z(n2326) );
  XNOR U1758 ( .A(n2122), .B(n2121), .Z(n2097) );
  XNOR U1759 ( .A(n2017), .B(n2016), .Z(n1992) );
  ANDN U1760 ( .A(n2147), .B(n2148), .Z(n2042) );
  XNOR U1761 ( .A(n1531), .B(n1530), .Z(n1505) );
  XNOR U1762 ( .A(n1297), .B(n1296), .Z(n1278) );
  XNOR U1763 ( .A(n1100), .B(n1099), .Z(n1088) );
  XNOR U1764 ( .A(n926), .B(n925), .Z(n918) );
  XNOR U1765 ( .A(n807), .B(n806), .Z(n795) );
  XNOR U1766 ( .A(n2964), .B(n2963), .Z(n2917) );
  XNOR U1767 ( .A(n2447), .B(n2446), .Z(n2416) );
  XOR U1768 ( .A(n1974), .B(n1971), .Z(n2049) );
  XNOR U1769 ( .A(n1787), .B(n1786), .Z(n1768) );
  XNOR U1770 ( .A(n1486), .B(n1485), .Z(n1564) );
  ANDN U1771 ( .A(n691), .B(n690), .Z(n689) );
  XNOR U1772 ( .A(n685), .B(n684), .Z(n676) );
  XOR U1773 ( .A(n1194), .B(n1193), .Z(n1257) );
  XNOR U1774 ( .A(n1017), .B(n1016), .Z(n1067) );
  XNOR U1775 ( .A(n869), .B(n868), .Z(n909) );
  XNOR U1776 ( .A(n760), .B(n759), .Z(n789) );
  XNOR U1777 ( .A(n705), .B(n704), .Z(n726) );
  XOR U1778 ( .A(n2621), .B(n2624), .Z(n2622) );
  XOR U1779 ( .A(n2262), .B(n2265), .Z(n2263) );
  XOR U1780 ( .A(n1939), .B(n1942), .Z(n1940) );
  XOR U1781 ( .A(n1650), .B(n1654), .Z(n1652) );
  XOR U1782 ( .A(n1396), .B(n1400), .Z(n1398) );
  XOR U1783 ( .A(n1187), .B(n1191), .Z(n1189) );
  XOR U1784 ( .A(n1010), .B(n1014), .Z(n1012) );
  XOR U1785 ( .A(n862), .B(n866), .Z(n864) );
  MUX U1786 ( .IN0(\_MxM/Y0[31] ), .IN1(n665), .SEL(n666), .F(n662) );
  MUX U1787 ( .IN0(n576), .IN1(n3663), .SEL(n3664), .F(n3625) );
  IV U1788 ( .A(n3665), .Z(n576) );
  MUX U1789 ( .IN0(n577), .IN1(n4091), .SEL(n4092), .F(n4074) );
  IV U1790 ( .A(n4093), .Z(n577) );
  MUX U1791 ( .IN0(n578), .IN1(n3684), .SEL(n3685), .F(n3646) );
  IV U1792 ( .A(n3686), .Z(n578) );
  XNOR U1793 ( .A(n3707), .B(n3706), .Z(n3719) );
  XNOR U1794 ( .A(n4114), .B(n4113), .Z(n3733) );
  MUX U1795 ( .IN0(n579), .IN1(n3638), .SEL(n3639), .F(n3600) );
  IV U1796 ( .A(n3640), .Z(n579) );
  XNOR U1797 ( .A(n3669), .B(n3668), .Z(n3681) );
  XNOR U1798 ( .A(n4097), .B(n4096), .Z(n3695) );
  XNOR U1799 ( .A(n3631), .B(n3630), .Z(n3643) );
  XNOR U1800 ( .A(n4080), .B(n4079), .Z(n3657) );
  XNOR U1801 ( .A(n3593), .B(n3592), .Z(n3605) );
  MUX U1802 ( .IN0(n4476), .IN1(n580), .SEL(n4071), .F(n4463) );
  IV U1803 ( .A(n4070), .Z(n580) );
  MUX U1804 ( .IN0(n581), .IN1(n3511), .SEL(n3512), .F(n3473) );
  IV U1805 ( .A(n3513), .Z(n581) );
  XNOR U1806 ( .A(n4063), .B(n4062), .Z(n3619) );
  XOR U1807 ( .A(n3606), .B(n3571), .Z(n3575) );
  MUX U1808 ( .IN0(n582), .IN1(n4023), .SEL(n4024), .F(n4006) );
  IV U1809 ( .A(n4025), .Z(n582) );
  XNOR U1810 ( .A(n3555), .B(n3554), .Z(n3567) );
  MUX U1811 ( .IN0(n583), .IN1(n4459), .SEL(n4460), .F(n4446) );
  IV U1812 ( .A(n4461), .Z(n583) );
  XNOR U1813 ( .A(n4046), .B(n4045), .Z(n3581) );
  MUX U1814 ( .IN0(n584), .IN1(n3486), .SEL(n3487), .F(n3448) );
  IV U1815 ( .A(n3488), .Z(n584) );
  XNOR U1816 ( .A(n3517), .B(n3516), .Z(n3529) );
  MUX U1817 ( .IN0(n585), .IN1(n4439), .SEL(n4440), .F(n4426) );
  IV U1818 ( .A(n4441), .Z(n585) );
  XNOR U1819 ( .A(n4029), .B(n4028), .Z(n3543) );
  XNOR U1820 ( .A(n3479), .B(n3478), .Z(n3491) );
  XOR U1821 ( .A(n4429), .B(n4421), .Z(n4003) );
  XNOR U1822 ( .A(n4012), .B(n4011), .Z(n3505) );
  XOR U1823 ( .A(n3492), .B(n3457), .Z(n3461) );
  XNOR U1824 ( .A(n3441), .B(n3440), .Z(n3453) );
  MUX U1825 ( .IN0(n586), .IN1(n4592), .SEL(n4593), .F(n4581) );
  IV U1826 ( .A(n4594), .Z(n586) );
  XOR U1827 ( .A(n4401), .B(n4402), .Z(n3985) );
  MUX U1828 ( .IN0(n587), .IN1(n4811), .SEL(n4812), .F(n4790) );
  IV U1829 ( .A(n4813), .Z(n587) );
  MUX U1830 ( .IN0(n588), .IN1(n3359), .SEL(n3360), .F(n3321) );
  IV U1831 ( .A(n3361), .Z(n588) );
  XNOR U1832 ( .A(n3995), .B(n3994), .Z(n3467) );
  MUX U1833 ( .IN0(n589), .IN1(n3955), .SEL(n3956), .F(n3938) );
  IV U1834 ( .A(n3957), .Z(n589) );
  XNOR U1835 ( .A(n3403), .B(n3402), .Z(n3415) );
  MUX U1836 ( .IN0(n590), .IN1(n4225), .SEL(n4226), .F(n4204) );
  IV U1837 ( .A(n4227), .Z(n590) );
  XOR U1838 ( .A(n4270), .B(n4252), .Z(n4256) );
  MUX U1839 ( .IN0(n591), .IN1(n4576), .SEL(n4577), .F(n4565) );
  IV U1840 ( .A(n4578), .Z(n591) );
  XOR U1841 ( .A(n4388), .B(n4389), .Z(n3968) );
  XNOR U1842 ( .A(n3978), .B(n3977), .Z(n3429) );
  MUX U1843 ( .IN0(n592), .IN1(n3334), .SEL(n3335), .F(n3296) );
  IV U1844 ( .A(n3336), .Z(n592) );
  XNOR U1845 ( .A(n3365), .B(n3364), .Z(n3377) );
  MUX U1846 ( .IN0(n4951), .IN1(n593), .SEL(n4808), .F(n4938) );
  IV U1847 ( .A(n4806), .Z(n593) );
  MUX U1848 ( .IN0(n594), .IN1(n4394), .SEL(n4395), .F(n4381) );
  IV U1849 ( .A(n4396), .Z(n594) );
  XNOR U1850 ( .A(n3961), .B(n3960), .Z(n3391) );
  XOR U1851 ( .A(n3378), .B(n3343), .Z(n3347) );
  XNOR U1852 ( .A(n3327), .B(n3326), .Z(n3339) );
  XOR U1853 ( .A(n4568), .B(n4560), .Z(n4201) );
  MUX U1854 ( .IN0(n5119), .IN1(n5135), .SEL(n5121), .F(n5101) );
  XOR U1855 ( .A(n4793), .B(n4775), .Z(n4779) );
  MUX U1856 ( .IN0(n595), .IN1(n4921), .SEL(n4922), .F(n4908) );
  IV U1857 ( .A(n4923), .Z(n595) );
  XNOR U1858 ( .A(n3944), .B(n3943), .Z(n3353) );
  XNOR U1859 ( .A(n3289), .B(n3288), .Z(n3301) );
  XNOR U1860 ( .A(n3281), .B(n3246), .Z(n3250) );
  MUX U1861 ( .IN0(n4306), .IN1(n4309), .SEL(n4307), .F(n4293) );
  MUX U1862 ( .IN0(n4620), .IN1(n4642), .SEL(n4622), .F(n4609) );
  XOR U1863 ( .A(n4207), .B(n4189), .Z(n4193) );
  XOR U1864 ( .A(n4364), .B(n4356), .Z(n3918) );
  MUX U1865 ( .IN0(n4871), .IN1(n4874), .SEL(n4872), .F(n4858) );
  MUX U1866 ( .IN0(n4992), .IN1(n5014), .SEL(n4994), .F(n4979) );
  XOR U1867 ( .A(n4915), .B(n4916), .Z(n4764) );
  MUX U1868 ( .IN0(n596), .IN1(n4727), .SEL(n4728), .F(n4708) );
  IV U1869 ( .A(n4729), .Z(n596) );
  MUX U1870 ( .IN0(n597), .IN1(n3215), .SEL(n3216), .F(n3178) );
  IV U1871 ( .A(n3217), .Z(n597) );
  XNOR U1872 ( .A(n3927), .B(n3926), .Z(n3315) );
  MUX U1873 ( .IN0(n598), .IN1(n3884), .SEL(n3885), .F(n3186) );
  IV U1874 ( .A(n3886), .Z(n598) );
  MUX U1875 ( .IN0(n3773), .IN1(n3797), .SEL(n3775), .F(n3752) );
  MUX U1876 ( .IN0(n599), .IN1(n4150), .SEL(n4151), .F(n4133) );
  IV U1877 ( .A(n4152), .Z(n599) );
  XOR U1878 ( .A(n4683), .B(n4670), .Z(n4325) );
  MUX U1879 ( .IN0(n600), .IN1(n4532), .SEL(n4533), .F(n4517) );
  IV U1880 ( .A(n4534), .Z(n600) );
  MUX U1881 ( .IN0(n601), .IN1(n4348), .SEL(n4349), .F(n4343) );
  IV U1882 ( .A(n4350), .Z(n601) );
  MUX U1883 ( .IN0(g_input[1]), .IN1(n5180), .SEL(g_input[31]), .F(n3833) );
  MUX U1884 ( .IN0(n5082), .IN1(n5092), .SEL(n5084), .F(n3128) );
  XOR U1885 ( .A(n5055), .B(n5042), .Z(n4890) );
  MUX U1886 ( .IN0(n602), .IN1(n4715), .SEL(n4716), .F(n3103) );
  IV U1887 ( .A(n4717), .Z(n602) );
  MUX U1888 ( .IN0(n603), .IN1(n3153), .SEL(n3154), .F(n3023) );
  IV U1889 ( .A(n3155), .Z(n603) );
  MUX U1890 ( .IN0(e_input[1]), .IN1(n604), .SEL(e_input[31]), .F(n4329) );
  IV U1891 ( .A(n4696), .Z(n604) );
  XNOR U1892 ( .A(n3910), .B(n3909), .Z(n3277) );
  XOR U1893 ( .A(n3264), .B(n3229), .Z(n3233) );
  XOR U1894 ( .A(n3839), .B(n3825), .Z(n3778) );
  XOR U1895 ( .A(n4624), .B(n4615), .Z(n4303) );
  MUX U1896 ( .IN0(g_input[2]), .IN1(n5172), .SEL(g_input[31]), .F(n3144) );
  MUX U1897 ( .IN0(n605), .IN1(n3065), .SEL(n3066), .F(n2929) );
  IV U1898 ( .A(n3067), .Z(n605) );
  XOR U1899 ( .A(n5145), .B(n5132), .Z(n5077) );
  XOR U1900 ( .A(n4996), .B(n4987), .Z(n4868) );
  XOR U1901 ( .A(n4730), .B(n4701), .Z(n4705) );
  XNOR U1902 ( .A(n3890), .B(n3889), .Z(n3239) );
  XOR U1903 ( .A(n3779), .B(n3761), .Z(n3765) );
  XNOR U1904 ( .A(n3854), .B(n3740), .Z(n3744) );
  XNOR U1905 ( .A(n4140), .B(n4126), .Z(n4130) );
  XNOR U1906 ( .A(n4299), .B(n4298), .Z(n3874) );
  XOR U1907 ( .A(n4535), .B(n4525), .Z(n4139) );
  MUX U1908 ( .IN0(n606), .IN1(n2951), .SEL(n2952), .F(n2813) );
  IV U1909 ( .A(n2953), .Z(n606) );
  MUX U1910 ( .IN0(n607), .IN1(n2984), .SEL(n2985), .F(n2846) );
  IV U1911 ( .A(n2986), .Z(n607) );
  MUX U1912 ( .IN0(g_input[3]), .IN1(n5163), .SEL(g_input[31]), .F(n608) );
  IV U1913 ( .A(n608), .Z(n3008) );
  MUX U1914 ( .IN0(n609), .IN1(n2783), .SEL(n2784), .F(n2656) );
  IV U1915 ( .A(n2785), .Z(n609) );
  MUX U1916 ( .IN0(e_input[4]), .IN1(n4317), .SEL(e_input[31]), .F(n2796) );
  MUX U1917 ( .IN0(g_input[4]), .IN1(n5129), .SEL(g_input[31]), .F(n610) );
  IV U1918 ( .A(n610), .Z(n2870) );
  MUX U1919 ( .IN0(n611), .IN1(n2631), .SEL(n2632), .F(n2507) );
  IV U1920 ( .A(n2633), .Z(n611) );
  MUX U1921 ( .IN0(g_input[5]), .IN1(n5112), .SEL(g_input[31]), .F(n2741) );
  MUX U1922 ( .IN0(n612), .IN1(n2700), .SEL(n2701), .F(n2572) );
  IV U1923 ( .A(n2702), .Z(n612) );
  MUX U1924 ( .IN0(g_input[6]), .IN1(n5093), .SEL(g_input[31]), .F(n2613) );
  MUX U1925 ( .IN0(n613), .IN1(n2403), .SEL(n2404), .F(n2288) );
  IV U1926 ( .A(n2405), .Z(n613) );
  MUX U1927 ( .IN0(n614), .IN1(n2467), .SEL(n2468), .F(n2346) );
  IV U1928 ( .A(n2469), .Z(n614) );
  MUX U1929 ( .IN0(g_input[7]), .IN1(n5081), .SEL(g_input[31]), .F(n2491) );
  MUX U1930 ( .IN0(n615), .IN1(n2484), .SEL(n2485), .F(n2363) );
  IV U1931 ( .A(n2486), .Z(n615) );
  MUX U1932 ( .IN0(n616), .IN1(n2434), .SEL(n2435), .F(n2313) );
  IV U1933 ( .A(n2436), .Z(n616) );
  MUX U1934 ( .IN0(e_input[8]), .IN1(n3852), .SEL(e_input[31]), .F(n2282) );
  MUX U1935 ( .IN0(n617), .IN1(n2321), .SEL(n2322), .F(n2203) );
  IV U1936 ( .A(n2323), .Z(n617) );
  MUX U1937 ( .IN0(g_input[8]), .IN1(n4984), .SEL(g_input[31]), .F(n2370) );
  MUX U1938 ( .IN0(e_input[9]), .IN1(n3853), .SEL(e_input[31]), .F(n2166) );
  MUX U1939 ( .IN0(g_input[9]), .IN1(n4972), .SEL(g_input[31]), .F(n2254) );
  MUX U1940 ( .IN0(n618), .IN1(n2211), .SEL(n2212), .F(n2100) );
  IV U1941 ( .A(n2213), .Z(n618) );
  MUX U1942 ( .IN0(n619), .IN1(n2073), .SEL(n2074), .F(n1968) );
  IV U1943 ( .A(n2075), .Z(n619) );
  MUX U1944 ( .IN0(g_input[10]), .IN1(n4958), .SEL(g_input[31]), .F(n2141) );
  MUX U1945 ( .IN0(n620), .IN1(n2012), .SEL(n2013), .F(n1907) );
  IV U1946 ( .A(n2014), .Z(n620) );
  MUX U1947 ( .IN0(g_input[11]), .IN1(n4946), .SEL(g_input[31]), .F(n2036) );
  MUX U1948 ( .IN0(n621), .IN1(n2029), .SEL(n2030), .F(n1924) );
  IV U1949 ( .A(n2031), .Z(n621) );
  MUX U1950 ( .IN0(n622), .IN1(n1979), .SEL(n1980), .F(n1874) );
  IV U1951 ( .A(n1981), .Z(n622) );
  MUX U1952 ( .IN0(e_input[12]), .IN1(n3867), .SEL(e_input[31]), .F(n1858) );
  MUX U1953 ( .IN0(g_input[12]), .IN1(n4932), .SEL(g_input[31]), .F(n1931) );
  MUX U1954 ( .IN0(g_input[13]), .IN1(n4920), .SEL(g_input[31]), .F(n1831) );
  MUX U1955 ( .IN0(n623), .IN1(n1790), .SEL(n1791), .F(n1694) );
  IV U1956 ( .A(n1792), .Z(n623) );
  MUX U1957 ( .IN0(g_input[14]), .IN1(n4906), .SEL(g_input[31]), .F(n1737) );
  MUX U1958 ( .IN0(n624), .IN1(n1585), .SEL(n1586), .F(n1492) );
  IV U1959 ( .A(n1587), .Z(n624) );
  MUX U1960 ( .IN0(n625), .IN1(n1618), .SEL(n1619), .F(n1526) );
  IV U1961 ( .A(n1620), .Z(n625) );
  MUX U1962 ( .IN0(n626), .IN1(n1626), .SEL(n1627), .F(n1534) );
  IV U1963 ( .A(n1628), .Z(n626) );
  MUX U1964 ( .IN0(g_input[15]), .IN1(n4894), .SEL(g_input[31]), .F(n1642) );
  MUX U1965 ( .IN0(n627), .IN1(n1635), .SEL(n1636), .F(n1543) );
  IV U1966 ( .A(n1637), .Z(n627) );
  MUX U1967 ( .IN0(e_input[16]), .IN1(n5068), .SEL(e_input[31]), .F(n1520) );
  MUX U1968 ( .IN0(g_input[16]), .IN1(n4522), .SEL(g_input[31]), .F(n1550) );
  MUX U1969 ( .IN0(e_input[17]), .IN1(n5069), .SEL(e_input[31]), .F(n1433) );
  MUX U1970 ( .IN0(g_input[17]), .IN1(n4510), .SEL(g_input[31]), .F(n1465) );
  MUX U1971 ( .IN0(g_input[18]), .IN1(n4496), .SEL(g_input[31]), .F(n1388) );
  MUX U1972 ( .IN0(n628), .IN1(n1424), .SEL(n1425), .F(n1353) );
  IV U1973 ( .A(n1426), .Z(n628) );
  MUX U1974 ( .IN0(g_input[19]), .IN1(n4484), .SEL(g_input[31]), .F(n1316) );
  MUX U1975 ( .IN0(n629), .IN1(n1292), .SEL(n1293), .F(n1222) );
  IV U1976 ( .A(n1294), .Z(n629) );
  MUX U1977 ( .IN0(g_input[20]), .IN1(n4470), .SEL(g_input[31]), .F(n1246) );
  MUX U1978 ( .IN0(e_input[20]), .IN1(n4882), .SEL(e_input[31]), .F(n1198) );
  MUX U1979 ( .IN0(e_input[21]), .IN1(n4883), .SEL(e_input[31]), .F(n1140) );
  MUX U1980 ( .IN0(g_input[21]), .IN1(n4458), .SEL(g_input[31]), .F(n1180) );
  MUX U1981 ( .IN0(g_input[22]), .IN1(n4444), .SEL(g_input[31]), .F(n1119) );
  MUX U1982 ( .IN0(n630), .IN1(n1033), .SEL(n1034), .F(n978) );
  IV U1983 ( .A(n1035), .Z(n630) );
  MUX U1984 ( .IN0(g_input[23]), .IN1(n4432), .SEL(g_input[31]), .F(n1057) );
  MUX U1985 ( .IN0(n631), .IN1(n1207), .SEL(n1208), .F(n1145) );
  IV U1986 ( .A(n1209), .Z(n631) );
  MUX U1987 ( .IN0(g_input[24]), .IN1(n4418), .SEL(g_input[31]), .F(n1003) );
  MUX U1988 ( .IN0(e_input[24]), .IN1(n5158), .SEL(e_input[31]), .F(n986) );
  MUX U1989 ( .IN0(e_input[25]), .IN1(n5159), .SEL(e_input[31]), .F(n932) );
  MUX U1990 ( .IN0(g_input[25]), .IN1(n4406), .SEL(g_input[31]), .F(n945) );
  MUX U1991 ( .IN0(g_input[26]), .IN1(n4392), .SEL(g_input[31]), .F(n899) );
  MUX U1992 ( .IN0(e_input[27]), .IN1(n5143), .SEL(e_input[31]), .F(n632) );
  IV U1993 ( .A(n632), .Z(n836) );
  MUX U1994 ( .IN0(e_input[26]), .IN1(n5144), .SEL(e_input[31]), .F(n874) );
  MUX U1995 ( .IN0(g_input[27]), .IN1(n4380), .SEL(g_input[31]), .F(n855) );
  MUX U1996 ( .IN0(e_input[2]), .IN1(n4681), .SEL(e_input[31]), .F(n3074) );
  XNOR U1997 ( .A(n5160), .B(n3138), .Z(n3142) );
  XNOR U1998 ( .A(n4864), .B(n4863), .Z(n4711) );
  XOR U1999 ( .A(n4891), .B(n3112), .Z(n3116) );
  XNOR U2000 ( .A(n3168), .B(n3041), .Z(n3045) );
  MUX U2001 ( .IN0(n3156), .IN1(n633), .SEL(n3157), .F(n3026) );
  IV U2002 ( .A(n3158), .Z(n633) );
  XNOR U2003 ( .A(n3081), .B(n4326), .Z(n3082) );
  XNOR U2004 ( .A(n3192), .B(n3191), .Z(n3202) );
  MUX U2005 ( .IN0(e_input[3]), .IN1(n4682), .SEL(e_input[31]), .F(n2942) );
  MUX U2006 ( .IN0(e_input[5]), .IN1(n4318), .SEL(e_input[31]), .F(n2666) );
  MUX U2007 ( .IN0(n2740), .IN1(n2738), .SEL(n2739), .F(n2610) );
  MUX U2008 ( .IN0(n2690), .IN1(n2688), .SEL(n2689), .F(n2560) );
  MUX U2009 ( .IN0(e_input[6]), .IN1(n4322), .SEL(e_input[31]), .F(n2544) );
  XOR U2010 ( .A(n2257), .B(n2371), .Z(n2258) );
  MUX U2011 ( .IN0(e_input[10]), .IN1(n3837), .SEL(e_input[31]), .F(n2053) );
  MUX U2012 ( .IN0(n634), .IN1(n2157), .SEL(n2158), .F(n2054) );
  IV U2013 ( .A(n2159), .Z(n634) );
  MUX U2014 ( .IN0(e_input[11]), .IN1(n3838), .SEL(e_input[31]), .F(n1952) );
  MUX U2015 ( .IN0(n2035), .IN1(n2033), .SEL(n2034), .F(n1928) );
  MUX U2016 ( .IN0(n1985), .IN1(n1983), .SEL(n1984), .F(n1878) );
  MUX U2017 ( .IN0(e_input[13]), .IN1(n3868), .SEL(e_input[31]), .F(n1757) );
  MUX U2018 ( .IN0(e_input[18]), .IN1(n5053), .SEL(e_input[31]), .F(n1352) );
  MUX U2019 ( .IN0(e_input[19]), .IN1(n5054), .SEL(e_input[31]), .F(n1284) );
  MUX U2020 ( .IN0(e_input[22]), .IN1(n4888), .SEL(e_input[31]), .F(n1082) );
  MUX U2021 ( .IN0(e_input[23]), .IN1(n4887), .SEL(e_input[31]), .F(n635) );
  IV U2022 ( .A(n635), .Z(n1022) );
  MUX U2023 ( .IN0(e_input[28]), .IN1(n5177), .SEL(e_input[31]), .F(n810) );
  MUX U2024 ( .IN0(e_input[29]), .IN1(n5178), .SEL(e_input[31]), .F(n774) );
  MUX U2025 ( .IN0(n636), .IN1(n857), .SEL(n858), .F(n820) );
  IV U2026 ( .A(n859), .Z(n636) );
  MUX U2027 ( .IN0(g_input[28]), .IN1(n4366), .SEL(g_input[31]), .F(n818) );
  XOR U2028 ( .A(n3029), .B(n2896), .Z(n2900) );
  XNOR U2029 ( .A(n3055), .B(n2922), .Z(n2926) );
  NAND U2030 ( .A(n2939), .B(n3073), .Z(n3072) );
  XNOR U2031 ( .A(n3093), .B(n3092), .Z(n3108) );
  XOR U2032 ( .A(n2990), .B(n2855), .Z(n2859) );
  XOR U2033 ( .A(n2674), .B(n2675), .Z(n2671) );
  XOR U2034 ( .A(n2835), .B(n2709), .Z(n2713) );
  XOR U2035 ( .A(n2546), .B(n2547), .Z(n2541) );
  XOR U2036 ( .A(n2513), .B(n2395), .Z(n2399) );
  XOR U2037 ( .A(n2595), .B(n2476), .Z(n2480) );
  MUX U2038 ( .IN0(e_input[7]), .IN1(n4323), .SEL(e_input[31]), .F(n2421) );
  XOR U2039 ( .A(n2456), .B(n2338), .Z(n2342) );
  XNOR U2040 ( .A(n2060), .B(n2163), .Z(n2061) );
  XNOR U2041 ( .A(n2172), .B(n2066), .Z(n2070) );
  XOR U2042 ( .A(n2234), .B(n2126), .Z(n2130) );
  XOR U2043 ( .A(n2106), .B(n2004), .Z(n2008) );
  XOR U2044 ( .A(n1913), .B(n1816), .Z(n1820) );
  XOR U2045 ( .A(n1796), .B(n1703), .Z(n1707) );
  MUX U2046 ( .IN0(n1761), .IN1(n1850), .SEL(n1760), .F(n1659) );
  MUX U2047 ( .IN0(e_input[14]), .IN1(n3872), .SEL(e_input[31]), .F(n1664) );
  NAND U2048 ( .A(n1435), .B(n1519), .Z(n1518) );
  XNOR U2049 ( .A(n1406), .B(n1336), .Z(n1340) );
  XNOR U2050 ( .A(n1456), .B(n1382), .Z(n1386) );
  XOR U2051 ( .A(n1447), .B(n1373), .Z(n1377) );
  XOR U2052 ( .A(n1228), .B(n1165), .Z(n1169) );
  XNOR U2053 ( .A(n1237), .B(n1174), .Z(n1178) );
  XNOR U2054 ( .A(n1196), .B(n1138), .Z(n1142) );
  XOR U2055 ( .A(n1039), .B(n988), .Z(n992) );
  XNOR U2056 ( .A(n1048), .B(n997), .Z(n1001) );
  OR U2057 ( .A(n886), .B(n887), .Z(n881) );
  MUX U2058 ( .IN0(n637), .IN1(n837), .SEL(n838), .F(n803) );
  IV U2059 ( .A(n839), .Z(n637) );
  MUX U2060 ( .IN0(n638), .IN1(n811), .SEL(n812), .F(n770) );
  IV U2061 ( .A(n813), .Z(n638) );
  MUX U2062 ( .IN0(g_input[29]), .IN1(n4354), .SEL(g_input[31]), .F(n778) );
  XNOR U2063 ( .A(n2957), .B(n2956), .Z(n2972) );
  XNOR U2064 ( .A(n2910), .B(n2909), .Z(n2892) );
  MUX U2065 ( .IN0(n2809), .IN1(n2807), .SEL(n2808), .F(n639) );
  IV U2066 ( .A(n639), .Z(n2677) );
  XNOR U2067 ( .A(n2530), .B(n2529), .Z(n2512) );
  XNOR U2068 ( .A(n2409), .B(n2408), .Z(n2391) );
  XNOR U2069 ( .A(n2440), .B(n2439), .Z(n2455) );
  XNOR U2070 ( .A(n2490), .B(n2489), .Z(n2472) );
  XNOR U2071 ( .A(n2294), .B(n2293), .Z(n2275) );
  XNOR U2072 ( .A(n2180), .B(n2179), .Z(n2162) );
  XNOR U2073 ( .A(n2140), .B(n2139), .Z(n2122) );
  XNOR U2074 ( .A(n2090), .B(n2089), .Z(n2105) );
  MUX U2075 ( .IN0(n1846), .IN1(n640), .SEL(n1847), .F(n1753) );
  IV U2076 ( .A(n1848), .Z(n640) );
  XNOR U2077 ( .A(n1780), .B(n1779), .Z(n1795) );
  XNOR U2078 ( .A(n1830), .B(n1829), .Z(n1812) );
  XNOR U2079 ( .A(n1684), .B(n1683), .Z(n1699) );
  XNOR U2080 ( .A(n1591), .B(n1590), .Z(n1606) );
  XNOR U2081 ( .A(n1498), .B(n1497), .Z(n1513) );
  XNOR U2082 ( .A(n1549), .B(n1548), .Z(n1531) );
  MUX U2083 ( .IN0(e_input[15]), .IN1(n3873), .SEL(e_input[31]), .F(n1570) );
  MUX U2084 ( .IN0(n641), .IN1(n1665), .SEL(n1666), .F(n1578) );
  IV U2085 ( .A(n1667), .Z(n641) );
  XNOR U2086 ( .A(n1414), .B(n1413), .Z(n1429) );
  XNOR U2087 ( .A(n1315), .B(n1314), .Z(n1297) );
  XNOR U2088 ( .A(n1215), .B(n1219), .Z(n1279) );
  XNOR U2089 ( .A(n1118), .B(n1117), .Z(n1100) );
  XNOR U2090 ( .A(n1056), .B(n1055), .Z(n1038) );
  AND U2091 ( .A(n970), .B(n971), .Z(n966) );
  XNOR U2092 ( .A(n944), .B(n943), .Z(n926) );
  XNOR U2093 ( .A(n898), .B(n897), .Z(n880) );
  MUX U2094 ( .IN0(g_input[30]), .IN1(n4336), .SEL(g_input[31]), .F(n744) );
  MUX U2095 ( .IN0(e_input[30]), .IN1(n5183), .SEL(e_input[31]), .F(n746) );
  XNOR U2096 ( .A(n2989), .B(n2988), .Z(n2964) );
  MUX U2097 ( .IN0(n3051), .IN1(n642), .SEL(n3052), .F(n2915) );
  IV U2098 ( .A(n3053), .Z(n642) );
  XNOR U2099 ( .A(n2763), .B(n2762), .Z(n2806) );
  XNOR U2100 ( .A(n2636), .B(n2635), .Z(n2680) );
  XNOR U2101 ( .A(n2303), .B(n2417), .Z(n2304) );
  NANDN U2102 ( .B(n1974), .A(n1975), .Z(n1869) );
  XNOR U2103 ( .A(n1716), .B(n1715), .Z(n1691) );
  XNOR U2104 ( .A(n1623), .B(n1622), .Z(n1598) );
  ANDN U2105 ( .A(n1743), .B(n1744), .Z(n1648) );
  XNOR U2106 ( .A(n1446), .B(n1445), .Z(n1421) );
  XNOR U2107 ( .A(n1227), .B(n1226), .Z(n1212) );
  XOR U2108 ( .A(n1029), .B(n1026), .Z(n1072) );
  OR U2109 ( .A(n794), .B(n795), .Z(n761) );
  MUX U2110 ( .IN0(n741), .IN1(n739), .SEL(n740), .F(n710) );
  XNOR U2111 ( .A(n709), .B(n708), .Z(n707) );
  XNOR U2112 ( .A(n2826), .B(n2825), .Z(n2788) );
  XNOR U2113 ( .A(n2697), .B(n2696), .Z(n2661) );
  XNOR U2114 ( .A(n2569), .B(n2568), .Z(n2537) );
  XNOR U2115 ( .A(n2326), .B(n2325), .Z(n2301) );
  XNOR U2116 ( .A(n2208), .B(n2207), .Z(n2187) );
  XNOR U2117 ( .A(n1992), .B(n1991), .Z(n1973) );
  XNOR U2118 ( .A(n1887), .B(n1886), .Z(n1868) );
  XOR U2119 ( .A(n1565), .B(n1579), .Z(n1656) );
  MUX U2120 ( .IN0(n643), .IN1(n715), .SEL(n716), .F(n692) );
  IV U2121 ( .A(n717), .Z(n643) );
  MUX U2122 ( .IN0(n3014), .IN1(n644), .SEL(n3015), .F(n2876) );
  IV U2123 ( .A(\_MxM/Y0[1] ), .Z(n644) );
  XOR U2124 ( .A(n1331), .B(n1330), .Z(n1399) );
  XNOR U2125 ( .A(n1134), .B(n1133), .Z(n1190) );
  XNOR U2126 ( .A(n959), .B(n958), .Z(n1013) );
  XNOR U2127 ( .A(n832), .B(n831), .Z(n865) );
  XNOR U2128 ( .A(n730), .B(n729), .Z(n756) );
  XNOR U2129 ( .A(n676), .B(n675), .Z(n701) );
  XOR U2130 ( .A(n2499), .B(n2502), .Z(n2500) );
  XOR U2131 ( .A(n2149), .B(n2152), .Z(n2150) );
  XOR U2132 ( .A(n1839), .B(n1843), .Z(n1841) );
  XOR U2133 ( .A(n1558), .B(n1562), .Z(n1560) );
  XOR U2134 ( .A(n1324), .B(n1328), .Z(n1326) );
  XOR U2135 ( .A(n1126), .B(n1131), .Z(n1129) );
  XOR U2136 ( .A(n952), .B(n956), .Z(n954) );
  XOR U2137 ( .A(n825), .B(n829), .Z(n827) );
  MUX U2138 ( .IN0(n662), .IN1(\_MxM/Y1[30] ), .SEL(n663), .F(\_MxM/Y1[31] )
         );
  MUX U2139 ( .IN0(\_MxM/Y1[26] ), .IN1(o[26]), .SEL(n645), .F(\_MxM/n99 ) );
  MUX U2140 ( .IN0(\_MxM/Y1[27] ), .IN1(o[27]), .SEL(n645), .F(\_MxM/n96 ) );
  MUX U2141 ( .IN0(\_MxM/Y1[28] ), .IN1(o[28]), .SEL(n645), .F(\_MxM/n93 ) );
  MUX U2142 ( .IN0(\_MxM/Y1[29] ), .IN1(o[29]), .SEL(n645), .F(\_MxM/n90 ) );
  MUX U2143 ( .IN0(\_MxM/Y1[30] ), .IN1(o[30]), .SEL(n645), .F(\_MxM/n87 ) );
  MUX U2144 ( .IN0(\_MxM/Y1[31] ), .IN1(o[31]), .SEL(n645), .F(\_MxM/n84 ) );
  MUX U2145 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n645), .F(\_MxM/n177 ) );
  MUX U2146 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n645), .F(\_MxM/n174 ) );
  MUX U2147 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n645), .F(\_MxM/n171 ) );
  MUX U2148 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n645), .F(\_MxM/n168 ) );
  MUX U2149 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n645), .F(\_MxM/n165 ) );
  MUX U2150 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n645), .F(\_MxM/n162 ) );
  MUX U2151 ( .IN0(\_MxM/Y1[6] ), .IN1(o[6]), .SEL(n645), .F(\_MxM/n159 ) );
  MUX U2152 ( .IN0(\_MxM/Y1[7] ), .IN1(o[7]), .SEL(n645), .F(\_MxM/n156 ) );
  MUX U2153 ( .IN0(\_MxM/Y1[8] ), .IN1(o[8]), .SEL(n645), .F(\_MxM/n153 ) );
  MUX U2154 ( .IN0(\_MxM/Y1[9] ), .IN1(o[9]), .SEL(n645), .F(\_MxM/n150 ) );
  MUX U2155 ( .IN0(\_MxM/Y1[10] ), .IN1(o[10]), .SEL(n645), .F(\_MxM/n147 ) );
  MUX U2156 ( .IN0(\_MxM/Y1[11] ), .IN1(o[11]), .SEL(n645), .F(\_MxM/n144 ) );
  MUX U2157 ( .IN0(\_MxM/Y1[12] ), .IN1(o[12]), .SEL(n645), .F(\_MxM/n141 ) );
  MUX U2158 ( .IN0(\_MxM/Y1[13] ), .IN1(o[13]), .SEL(n645), .F(\_MxM/n138 ) );
  MUX U2159 ( .IN0(\_MxM/Y1[14] ), .IN1(o[14]), .SEL(n645), .F(\_MxM/n135 ) );
  MUX U2160 ( .IN0(\_MxM/Y1[15] ), .IN1(o[15]), .SEL(n645), .F(\_MxM/n132 ) );
  MUX U2161 ( .IN0(\_MxM/Y1[16] ), .IN1(o[16]), .SEL(n645), .F(\_MxM/n129 ) );
  MUX U2162 ( .IN0(\_MxM/Y1[17] ), .IN1(o[17]), .SEL(n645), .F(\_MxM/n126 ) );
  MUX U2163 ( .IN0(\_MxM/Y1[18] ), .IN1(o[18]), .SEL(n645), .F(\_MxM/n123 ) );
  MUX U2164 ( .IN0(\_MxM/Y1[19] ), .IN1(o[19]), .SEL(n645), .F(\_MxM/n120 ) );
  MUX U2165 ( .IN0(\_MxM/Y1[20] ), .IN1(o[20]), .SEL(n645), .F(\_MxM/n117 ) );
  MUX U2166 ( .IN0(\_MxM/Y1[21] ), .IN1(o[21]), .SEL(n645), .F(\_MxM/n114 ) );
  MUX U2167 ( .IN0(\_MxM/Y1[22] ), .IN1(o[22]), .SEL(n645), .F(\_MxM/n111 ) );
  MUX U2168 ( .IN0(\_MxM/Y1[23] ), .IN1(o[23]), .SEL(n645), .F(\_MxM/n108 ) );
  IV U2169 ( .A(n646), .Z(n645) );
  MUX U2170 ( .IN0(o[24]), .IN1(\_MxM/Y1[24] ), .SEL(n646), .F(\_MxM/n105 ) );
  MUX U2171 ( .IN0(o[25]), .IN1(\_MxM/Y1[25] ), .SEL(n646), .F(\_MxM/n102 ) );
  AND U2172 ( .A(n647), .B(n648), .Z(n646) );
  AND U2173 ( .A(n649), .B(n650), .Z(n648) );
  ANDN U2174 ( .A(n651), .B(\_MxM/n[7] ), .Z(n650) );
  NOR U2175 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n651) );
  NOR U2176 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n649) );
  AND U2177 ( .A(n652), .B(n653), .Z(n647) );
  NOR U2178 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n653) );
  NOR U2179 ( .A(\_MxM/n[0] ), .B(n654), .Z(n652) );
  XOR U2180 ( .A(n655), .B(\_MxM/Y0[10] ), .Z(\_MxM/Y1[9] ) );
  XOR U2181 ( .A(n656), .B(\_MxM/Y0[9] ), .Z(\_MxM/Y1[8] ) );
  XOR U2182 ( .A(n657), .B(\_MxM/Y0[8] ), .Z(\_MxM/Y1[7] ) );
  XOR U2183 ( .A(n658), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XOR U2184 ( .A(n659), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XOR U2185 ( .A(n660), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U2186 ( .A(n661), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U2187 ( .A(\_MxM/Y0[31] ), .B(n664), .Z(n663) );
  XNOR U2188 ( .A(n666), .B(\_MxM/Y0[31] ), .Z(\_MxM/Y1[30] ) );
  XOR U2189 ( .A(n665), .B(n664), .Z(n666) );
  XOR U2190 ( .A(n667), .B(n668), .Z(n664) );
  XOR U2191 ( .A(n669), .B(n670), .Z(n668) );
  AND U2192 ( .A(n671), .B(n672), .Z(n670) );
  XNOR U2193 ( .A(n677), .B(n675), .Z(n667) );
  XOR U2194 ( .A(n678), .B(n679), .Z(n677) );
  XOR U2195 ( .A(n680), .B(n681), .Z(n679) );
  XOR U2196 ( .A(n682), .B(n683), .Z(n681) );
  XOR U2197 ( .A(n688), .B(n689), .Z(n680) );
  XOR U2198 ( .A(n694), .B(n695), .Z(n678) );
  XNOR U2199 ( .A(n684), .B(n696), .Z(n695) );
  XOR U2200 ( .A(n692), .B(n690), .Z(n694) );
  XNOR U2201 ( .A(n699), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U2202 ( .A(n697), .B(\_MxM/Y0[30] ), .Z(\_MxM/Y1[29] ) );
  XNOR U2203 ( .A(n700), .B(n701), .Z(n697) );
  XNOR U2204 ( .A(n698), .B(n702), .Z(n700) );
  AND U2205 ( .A(n671), .B(n703), .Z(n702) );
  XOR U2206 ( .A(n674), .B(n701), .Z(n703) );
  XNOR U2207 ( .A(n673), .B(n701), .Z(n674) );
  XOR U2208 ( .A(n687), .B(n696), .Z(n685) );
  IV U2209 ( .A(n686), .Z(n696) );
  XOR U2210 ( .A(n692), .B(n693), .Z(n691) );
  OR U2211 ( .A(n713), .B(n714), .Z(n693) );
  ANDN U2212 ( .A(n722), .B(n723), .Z(n721) );
  XOR U2213 ( .A(\_MxM/Y0[29] ), .B(n724), .Z(n722) );
  XNOR U2214 ( .A(n723), .B(\_MxM/Y0[29] ), .Z(\_MxM/Y1[28] ) );
  XNOR U2215 ( .A(n725), .B(n726), .Z(n723) );
  XNOR U2216 ( .A(n724), .B(n727), .Z(n725) );
  AND U2217 ( .A(n671), .B(n728), .Z(n727) );
  XOR U2218 ( .A(n719), .B(n726), .Z(n728) );
  XNOR U2219 ( .A(n718), .B(n726), .Z(n719) );
  XOR U2220 ( .A(n733), .B(n734), .Z(n708) );
  ANDN U2221 ( .A(n735), .B(n733), .Z(n734) );
  XOR U2222 ( .A(n733), .B(n736), .Z(n735) );
  XOR U2223 ( .A(n737), .B(n738), .Z(n711) );
  IV U2224 ( .A(n710), .Z(n738) );
  XNOR U2225 ( .A(n716), .B(n717), .Z(n712) );
  NANDN U2226 ( .B(n713), .A(n744), .Z(n717) );
  XNOR U2227 ( .A(n715), .B(n745), .Z(n716) );
  ANDN U2228 ( .A(n746), .B(n714), .Z(n745) );
  IV U2229 ( .A(n720), .Z(n724) );
  XNOR U2230 ( .A(n753), .B(\_MxM/Y0[28] ), .Z(\_MxM/Y1[27] ) );
  XNOR U2231 ( .A(n755), .B(n756), .Z(n753) );
  XNOR U2232 ( .A(n754), .B(n757), .Z(n755) );
  AND U2233 ( .A(n671), .B(n758), .Z(n757) );
  XOR U2234 ( .A(n751), .B(n756), .Z(n758) );
  XNOR U2235 ( .A(n750), .B(n756), .Z(n751) );
  XOR U2236 ( .A(n761), .B(n762), .Z(n731) );
  ANDN U2237 ( .A(n763), .B(n761), .Z(n762) );
  XOR U2238 ( .A(n761), .B(n764), .Z(n763) );
  XOR U2239 ( .A(n741), .B(n768), .Z(n736) );
  IV U2240 ( .A(n740), .Z(n768) );
  XOR U2241 ( .A(n773), .B(n743), .Z(n769) );
  NANDN U2242 ( .B(n714), .A(n774), .Z(n743) );
  IV U2243 ( .A(n739), .Z(n773) );
  XNOR U2244 ( .A(n748), .B(n749), .Z(n741) );
  NANDN U2245 ( .B(n713), .A(n778), .Z(n749) );
  XNOR U2246 ( .A(n747), .B(n779), .Z(n748) );
  AND U2247 ( .A(n744), .B(n746), .Z(n779) );
  IV U2248 ( .A(n752), .Z(n754) );
  XNOR U2249 ( .A(n786), .B(\_MxM/Y0[27] ), .Z(\_MxM/Y1[26] ) );
  XNOR U2250 ( .A(n788), .B(n789), .Z(n786) );
  XNOR U2251 ( .A(n787), .B(n790), .Z(n788) );
  AND U2252 ( .A(n671), .B(n791), .Z(n790) );
  XOR U2253 ( .A(n784), .B(n789), .Z(n791) );
  XNOR U2254 ( .A(n783), .B(n789), .Z(n784) );
  XNOR U2255 ( .A(n767), .B(n766), .Z(n764) );
  XOR U2256 ( .A(n796), .B(n797), .Z(n766) );
  XOR U2257 ( .A(n798), .B(n799), .Z(n797) );
  XOR U2258 ( .A(n800), .B(n801), .Z(n799) );
  XNOR U2259 ( .A(n770), .B(n809), .Z(n771) );
  ANDN U2260 ( .A(n810), .B(n714), .Z(n809) );
  XOR U2261 ( .A(n814), .B(n772), .Z(n808) );
  NAND U2262 ( .A(n774), .B(n744), .Z(n772) );
  IV U2263 ( .A(n775), .Z(n814) );
  XNOR U2264 ( .A(n781), .B(n782), .Z(n777) );
  NANDN U2265 ( .B(n713), .A(n818), .Z(n782) );
  XNOR U2266 ( .A(n780), .B(n819), .Z(n781) );
  AND U2267 ( .A(n778), .B(n746), .Z(n819) );
  IV U2268 ( .A(n785), .Z(n787) );
  XNOR U2269 ( .A(n826), .B(\_MxM/Y0[26] ), .Z(\_MxM/Y1[25] ) );
  XNOR U2270 ( .A(n827), .B(n828), .Z(n826) );
  AND U2271 ( .A(n671), .B(n830), .Z(n829) );
  XOR U2272 ( .A(n824), .B(n828), .Z(n830) );
  XNOR U2273 ( .A(n823), .B(n828), .Z(n824) );
  XNOR U2274 ( .A(n835), .B(n802), .Z(n806) );
  XOR U2275 ( .A(n803), .B(n804), .Z(n802) );
  OR U2276 ( .A(n714), .B(n836), .Z(n804) );
  XNOR U2277 ( .A(n798), .B(n805), .Z(n835) );
  XNOR U2278 ( .A(n811), .B(n847), .Z(n812) );
  AND U2279 ( .A(n744), .B(n810), .Z(n847) );
  XOR U2280 ( .A(n851), .B(n813), .Z(n846) );
  NAND U2281 ( .A(n774), .B(n778), .Z(n813) );
  IV U2282 ( .A(n815), .Z(n851) );
  XNOR U2283 ( .A(n821), .B(n822), .Z(n817) );
  NANDN U2284 ( .B(n713), .A(n855), .Z(n822) );
  XNOR U2285 ( .A(n820), .B(n856), .Z(n821) );
  AND U2286 ( .A(n818), .B(n746), .Z(n856) );
  XNOR U2287 ( .A(n863), .B(\_MxM/Y0[25] ), .Z(\_MxM/Y1[24] ) );
  XNOR U2288 ( .A(n864), .B(n865), .Z(n863) );
  AND U2289 ( .A(n671), .B(n867), .Z(n866) );
  XOR U2290 ( .A(n861), .B(n865), .Z(n867) );
  XNOR U2291 ( .A(n860), .B(n865), .Z(n861) );
  XNOR U2292 ( .A(n872), .B(n845), .Z(n841) );
  XNOR U2293 ( .A(n838), .B(n839), .Z(n845) );
  NANDN U2294 ( .B(n836), .A(n744), .Z(n839) );
  XNOR U2295 ( .A(n837), .B(n873), .Z(n838) );
  ANDN U2296 ( .A(n874), .B(n714), .Z(n873) );
  XNOR U2297 ( .A(n844), .B(n840), .Z(n872) );
  XNOR U2298 ( .A(n881), .B(n882), .Z(n844) );
  IV U2299 ( .A(n843), .Z(n882) );
  XNOR U2300 ( .A(n848), .B(n889), .Z(n849) );
  AND U2301 ( .A(n778), .B(n810), .Z(n889) );
  XOR U2302 ( .A(n893), .B(n850), .Z(n888) );
  NAND U2303 ( .A(n774), .B(n818), .Z(n850) );
  IV U2304 ( .A(n852), .Z(n893) );
  XOR U2305 ( .A(n894), .B(n895), .Z(n852) );
  ANDN U2306 ( .A(n896), .B(n897), .Z(n895) );
  XOR U2307 ( .A(n894), .B(n898), .Z(n896) );
  XNOR U2308 ( .A(n858), .B(n859), .Z(n854) );
  NANDN U2309 ( .B(n713), .A(n899), .Z(n859) );
  XNOR U2310 ( .A(n857), .B(n900), .Z(n858) );
  AND U2311 ( .A(n855), .B(n746), .Z(n900) );
  XNOR U2312 ( .A(n907), .B(\_MxM/Y0[24] ), .Z(\_MxM/Y1[23] ) );
  XNOR U2313 ( .A(n908), .B(n909), .Z(n907) );
  AND U2314 ( .A(n671), .B(n911), .Z(n910) );
  XOR U2315 ( .A(n905), .B(n909), .Z(n911) );
  XNOR U2316 ( .A(n904), .B(n909), .Z(n905) );
  XNOR U2317 ( .A(n914), .B(n915), .Z(n870) );
  ANDN U2318 ( .A(n916), .B(n917), .Z(n915) );
  XNOR U2319 ( .A(n914), .B(n918), .Z(n916) );
  XNOR U2320 ( .A(n919), .B(n885), .Z(n879) );
  XNOR U2321 ( .A(n876), .B(n877), .Z(n885) );
  NANDN U2322 ( .B(n836), .A(n778), .Z(n877) );
  XNOR U2323 ( .A(n875), .B(n920), .Z(n876) );
  AND U2324 ( .A(n744), .B(n874), .Z(n920) );
  XNOR U2325 ( .A(n884), .B(n878), .Z(n919) );
  XOR U2326 ( .A(n931), .B(n887), .Z(n927) );
  NANDN U2327 ( .B(n714), .A(n932), .Z(n887) );
  IV U2328 ( .A(n883), .Z(n931) );
  XNOR U2329 ( .A(n890), .B(n937), .Z(n891) );
  AND U2330 ( .A(n818), .B(n810), .Z(n937) );
  XOR U2331 ( .A(n941), .B(n892), .Z(n936) );
  NAND U2332 ( .A(n774), .B(n855), .Z(n892) );
  IV U2333 ( .A(n894), .Z(n941) );
  XNOR U2334 ( .A(n902), .B(n903), .Z(n898) );
  NANDN U2335 ( .B(n713), .A(n945), .Z(n903) );
  XNOR U2336 ( .A(n901), .B(n946), .Z(n902) );
  AND U2337 ( .A(n899), .B(n746), .Z(n946) );
  XNOR U2338 ( .A(n953), .B(\_MxM/Y0[23] ), .Z(\_MxM/Y1[22] ) );
  XNOR U2339 ( .A(n954), .B(n955), .Z(n953) );
  AND U2340 ( .A(n671), .B(n957), .Z(n956) );
  XOR U2341 ( .A(n951), .B(n955), .Z(n957) );
  XNOR U2342 ( .A(n950), .B(n955), .Z(n951) );
  XNOR U2343 ( .A(n918), .B(n917), .Z(n913) );
  XOR U2344 ( .A(n960), .B(n961), .Z(n917) );
  XOR U2345 ( .A(n962), .B(n963), .Z(n961) );
  XOR U2346 ( .A(n966), .B(n967), .Z(n962) );
  XOR U2347 ( .A(n972), .B(n914), .Z(n960) );
  XOR U2348 ( .A(n970), .B(n968), .Z(n972) );
  XNOR U2349 ( .A(n976), .B(n935), .Z(n925) );
  XNOR U2350 ( .A(n922), .B(n923), .Z(n935) );
  NANDN U2351 ( .B(n836), .A(n818), .Z(n923) );
  XNOR U2352 ( .A(n921), .B(n977), .Z(n922) );
  AND U2353 ( .A(n778), .B(n874), .Z(n977) );
  XNOR U2354 ( .A(n934), .B(n924), .Z(n976) );
  XNOR U2355 ( .A(n928), .B(n985), .Z(n929) );
  ANDN U2356 ( .A(n986), .B(n714), .Z(n985) );
  XOR U2357 ( .A(n990), .B(n930), .Z(n984) );
  NAND U2358 ( .A(n932), .B(n744), .Z(n930) );
  IV U2359 ( .A(n933), .Z(n990) );
  XNOR U2360 ( .A(n938), .B(n995), .Z(n939) );
  AND U2361 ( .A(n855), .B(n810), .Z(n995) );
  XOR U2362 ( .A(n999), .B(n940), .Z(n994) );
  NAND U2363 ( .A(n774), .B(n899), .Z(n940) );
  IV U2364 ( .A(n942), .Z(n999) );
  XNOR U2365 ( .A(n948), .B(n949), .Z(n944) );
  NANDN U2366 ( .B(n713), .A(n1003), .Z(n949) );
  XNOR U2367 ( .A(n947), .B(n1004), .Z(n948) );
  AND U2368 ( .A(n945), .B(n746), .Z(n1004) );
  XNOR U2369 ( .A(n1011), .B(\_MxM/Y0[22] ), .Z(\_MxM/Y1[21] ) );
  XNOR U2370 ( .A(n1012), .B(n1013), .Z(n1011) );
  AND U2371 ( .A(n671), .B(n1015), .Z(n1014) );
  XOR U2372 ( .A(n1009), .B(n1013), .Z(n1015) );
  XNOR U2373 ( .A(n1008), .B(n1013), .Z(n1009) );
  XNOR U2374 ( .A(n1018), .B(n965), .Z(n974) );
  XOR U2375 ( .A(n970), .B(n971), .Z(n969) );
  OR U2376 ( .A(n714), .B(n1022), .Z(n971) );
  XNOR U2377 ( .A(n964), .B(n973), .Z(n1018) );
  XNOR U2378 ( .A(n1031), .B(n993), .Z(n982) );
  XNOR U2379 ( .A(n979), .B(n980), .Z(n993) );
  NANDN U2380 ( .B(n836), .A(n855), .Z(n980) );
  XNOR U2381 ( .A(n978), .B(n1032), .Z(n979) );
  AND U2382 ( .A(n818), .B(n874), .Z(n1032) );
  XNOR U2383 ( .A(n992), .B(n981), .Z(n1031) );
  XNOR U2384 ( .A(n987), .B(n1040), .Z(n988) );
  AND U2385 ( .A(n744), .B(n986), .Z(n1040) );
  XOR U2386 ( .A(n1044), .B(n989), .Z(n1039) );
  NAND U2387 ( .A(n932), .B(n778), .Z(n989) );
  IV U2388 ( .A(n991), .Z(n1044) );
  XNOR U2389 ( .A(n996), .B(n1049), .Z(n997) );
  AND U2390 ( .A(n899), .B(n810), .Z(n1049) );
  XOR U2391 ( .A(n1053), .B(n998), .Z(n1048) );
  NAND U2392 ( .A(n774), .B(n945), .Z(n998) );
  IV U2393 ( .A(n1000), .Z(n1053) );
  XNOR U2394 ( .A(n1006), .B(n1007), .Z(n1002) );
  NANDN U2395 ( .B(n713), .A(n1057), .Z(n1007) );
  XNOR U2396 ( .A(n1005), .B(n1058), .Z(n1006) );
  AND U2397 ( .A(n1003), .B(n746), .Z(n1058) );
  XNOR U2398 ( .A(n1065), .B(\_MxM/Y0[21] ), .Z(\_MxM/Y1[20] ) );
  XNOR U2399 ( .A(n1066), .B(n1067), .Z(n1065) );
  AND U2400 ( .A(n671), .B(n1069), .Z(n1068) );
  XOR U2401 ( .A(n1063), .B(n1067), .Z(n1069) );
  XNOR U2402 ( .A(n1062), .B(n1067), .Z(n1063) );
  XNOR U2403 ( .A(n1072), .B(n1030), .Z(n1027) );
  XOR U2404 ( .A(n1073), .B(n1074), .Z(n1020) );
  IV U2405 ( .A(n1019), .Z(n1074) );
  XNOR U2406 ( .A(n1024), .B(n1025), .Z(n1021) );
  NANDN U2407 ( .B(n1022), .A(n744), .Z(n1025) );
  XNOR U2408 ( .A(n1023), .B(n1081), .Z(n1024) );
  ANDN U2409 ( .A(n1082), .B(n714), .Z(n1081) );
  XOR U2410 ( .A(n1089), .B(n1090), .Z(n1029) );
  ANDN U2411 ( .A(n1091), .B(n1089), .Z(n1090) );
  XOR U2412 ( .A(n1089), .B(n1092), .Z(n1091) );
  XNOR U2413 ( .A(n1093), .B(n1047), .Z(n1037) );
  XNOR U2414 ( .A(n1034), .B(n1035), .Z(n1047) );
  NANDN U2415 ( .B(n836), .A(n899), .Z(n1035) );
  XNOR U2416 ( .A(n1033), .B(n1094), .Z(n1034) );
  AND U2417 ( .A(n855), .B(n874), .Z(n1094) );
  XNOR U2418 ( .A(n1046), .B(n1036), .Z(n1093) );
  XNOR U2419 ( .A(n1041), .B(n1102), .Z(n1042) );
  AND U2420 ( .A(n778), .B(n986), .Z(n1102) );
  XOR U2421 ( .A(n1106), .B(n1043), .Z(n1101) );
  NAND U2422 ( .A(n932), .B(n818), .Z(n1043) );
  IV U2423 ( .A(n1045), .Z(n1106) );
  XNOR U2424 ( .A(n1050), .B(n1111), .Z(n1051) );
  AND U2425 ( .A(n945), .B(n810), .Z(n1111) );
  XOR U2426 ( .A(n1115), .B(n1052), .Z(n1110) );
  NAND U2427 ( .A(n774), .B(n1003), .Z(n1052) );
  IV U2428 ( .A(n1054), .Z(n1115) );
  XNOR U2429 ( .A(n1060), .B(n1061), .Z(n1056) );
  NANDN U2430 ( .B(n713), .A(n1119), .Z(n1061) );
  XNOR U2431 ( .A(n1059), .B(n1120), .Z(n1060) );
  AND U2432 ( .A(n1057), .B(n746), .Z(n1120) );
  XNOR U2433 ( .A(n1128), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U2434 ( .A(n1127), .B(\_MxM/Y0[20] ), .Z(\_MxM/Y1[19] ) );
  XNOR U2435 ( .A(n1129), .B(n1130), .Z(n1127) );
  AND U2436 ( .A(n671), .B(n1132), .Z(n1131) );
  XOR U2437 ( .A(n1125), .B(n1130), .Z(n1132) );
  XNOR U2438 ( .A(n1124), .B(n1130), .Z(n1125) );
  XNOR U2439 ( .A(n1135), .B(n1092), .Z(n1087) );
  XOR U2440 ( .A(n1136), .B(n1078), .Z(n1076) );
  IV U2441 ( .A(n1079), .Z(n1078) );
  NANDN U2442 ( .B(n714), .A(n1140), .Z(n1080) );
  XNOR U2443 ( .A(n1084), .B(n1085), .Z(n1077) );
  NANDN U2444 ( .B(n1022), .A(n778), .Z(n1085) );
  XNOR U2445 ( .A(n1083), .B(n1144), .Z(n1084) );
  AND U2446 ( .A(n744), .B(n1082), .Z(n1144) );
  XNOR U2447 ( .A(n1154), .B(n1109), .Z(n1099) );
  XNOR U2448 ( .A(n1096), .B(n1097), .Z(n1109) );
  NANDN U2449 ( .B(n836), .A(n945), .Z(n1097) );
  XNOR U2450 ( .A(n1095), .B(n1155), .Z(n1096) );
  AND U2451 ( .A(n899), .B(n874), .Z(n1155) );
  XNOR U2452 ( .A(n1108), .B(n1098), .Z(n1154) );
  XNOR U2453 ( .A(n1103), .B(n1163), .Z(n1104) );
  AND U2454 ( .A(n818), .B(n986), .Z(n1163) );
  XOR U2455 ( .A(n1167), .B(n1105), .Z(n1162) );
  NAND U2456 ( .A(n932), .B(n855), .Z(n1105) );
  IV U2457 ( .A(n1107), .Z(n1167) );
  XNOR U2458 ( .A(n1112), .B(n1172), .Z(n1113) );
  AND U2459 ( .A(n1003), .B(n810), .Z(n1172) );
  XOR U2460 ( .A(n1176), .B(n1114), .Z(n1171) );
  NAND U2461 ( .A(n774), .B(n1057), .Z(n1114) );
  IV U2462 ( .A(n1116), .Z(n1176) );
  XNOR U2463 ( .A(n1122), .B(n1123), .Z(n1118) );
  NANDN U2464 ( .B(n713), .A(n1180), .Z(n1123) );
  XNOR U2465 ( .A(n1121), .B(n1181), .Z(n1122) );
  AND U2466 ( .A(n1119), .B(n746), .Z(n1181) );
  XNOR U2467 ( .A(n1188), .B(\_MxM/Y0[19] ), .Z(\_MxM/Y1[18] ) );
  XNOR U2468 ( .A(n1189), .B(n1190), .Z(n1188) );
  AND U2469 ( .A(n671), .B(n1192), .Z(n1191) );
  XOR U2470 ( .A(n1186), .B(n1190), .Z(n1192) );
  XNOR U2471 ( .A(n1185), .B(n1190), .Z(n1186) );
  XNOR U2472 ( .A(n1195), .B(n1153), .Z(n1149) );
  XNOR U2473 ( .A(n1137), .B(n1197), .Z(n1138) );
  ANDN U2474 ( .A(n1198), .B(n714), .Z(n1197) );
  XOR U2475 ( .A(n1202), .B(n1139), .Z(n1196) );
  NAND U2476 ( .A(n1140), .B(n744), .Z(n1139) );
  IV U2477 ( .A(n1141), .Z(n1202) );
  XNOR U2478 ( .A(n1146), .B(n1147), .Z(n1143) );
  NANDN U2479 ( .B(n1022), .A(n818), .Z(n1147) );
  XNOR U2480 ( .A(n1145), .B(n1206), .Z(n1146) );
  AND U2481 ( .A(n778), .B(n1082), .Z(n1206) );
  XNOR U2482 ( .A(n1152), .B(n1148), .Z(n1195) );
  XNOR U2483 ( .A(n1213), .B(n1214), .Z(n1152) );
  IV U2484 ( .A(n1151), .Z(n1214) );
  XNOR U2485 ( .A(n1220), .B(n1170), .Z(n1160) );
  XNOR U2486 ( .A(n1157), .B(n1158), .Z(n1170) );
  NANDN U2487 ( .B(n836), .A(n1003), .Z(n1158) );
  XNOR U2488 ( .A(n1156), .B(n1221), .Z(n1157) );
  AND U2489 ( .A(n945), .B(n874), .Z(n1221) );
  XNOR U2490 ( .A(n1169), .B(n1159), .Z(n1220) );
  XNOR U2491 ( .A(n1164), .B(n1229), .Z(n1165) );
  AND U2492 ( .A(n855), .B(n986), .Z(n1229) );
  XOR U2493 ( .A(n1233), .B(n1166), .Z(n1228) );
  NAND U2494 ( .A(n932), .B(n899), .Z(n1166) );
  IV U2495 ( .A(n1168), .Z(n1233) );
  XNOR U2496 ( .A(n1173), .B(n1238), .Z(n1174) );
  AND U2497 ( .A(n1057), .B(n810), .Z(n1238) );
  XOR U2498 ( .A(n1242), .B(n1175), .Z(n1237) );
  NAND U2499 ( .A(n774), .B(n1119), .Z(n1175) );
  IV U2500 ( .A(n1177), .Z(n1242) );
  XNOR U2501 ( .A(n1183), .B(n1184), .Z(n1179) );
  NANDN U2502 ( .B(n713), .A(n1246), .Z(n1184) );
  XNOR U2503 ( .A(n1182), .B(n1247), .Z(n1183) );
  AND U2504 ( .A(n1180), .B(n746), .Z(n1247) );
  ANDN U2505 ( .A(n1248), .B(n1249), .Z(n1182) );
  NANDN U2506 ( .B(n1250), .A(n1251), .Z(n1248) );
  XOR U2507 ( .A(n1255), .B(\_MxM/Y0[18] ), .Z(\_MxM/Y1[17] ) );
  XNOR U2508 ( .A(n1256), .B(n1257), .Z(n1255) );
  AND U2509 ( .A(n671), .B(n1259), .Z(n1258) );
  XOR U2510 ( .A(n1253), .B(n1257), .Z(n1259) );
  XNOR U2511 ( .A(n1252), .B(n1257), .Z(n1253) );
  XNOR U2512 ( .A(n1212), .B(n1211), .Z(n1194) );
  XOR U2513 ( .A(n1262), .B(n1217), .Z(n1211) );
  XNOR U2514 ( .A(n1199), .B(n1264), .Z(n1200) );
  AND U2515 ( .A(n744), .B(n1198), .Z(n1264) );
  XOR U2516 ( .A(n1268), .B(n1201), .Z(n1263) );
  NAND U2517 ( .A(n1140), .B(n778), .Z(n1201) );
  IV U2518 ( .A(n1203), .Z(n1268) );
  XNOR U2519 ( .A(n1208), .B(n1209), .Z(n1205) );
  NANDN U2520 ( .B(n1022), .A(n855), .Z(n1209) );
  XNOR U2521 ( .A(n1207), .B(n1272), .Z(n1208) );
  AND U2522 ( .A(n818), .B(n1082), .Z(n1272) );
  XNOR U2523 ( .A(n1216), .B(n1210), .Z(n1262) );
  XOR U2524 ( .A(n1279), .B(n1218), .Z(n1216) );
  NAND U2525 ( .A(n1282), .B(n1283), .Z(n1219) );
  NANDN U2526 ( .B(n714), .A(n1284), .Z(n1283) );
  OR U2527 ( .A(n1285), .B(n1286), .Z(n1282) );
  XNOR U2528 ( .A(n1290), .B(n1236), .Z(n1226) );
  XNOR U2529 ( .A(n1223), .B(n1224), .Z(n1236) );
  NANDN U2530 ( .B(n836), .A(n1057), .Z(n1224) );
  XNOR U2531 ( .A(n1222), .B(n1291), .Z(n1223) );
  AND U2532 ( .A(n1003), .B(n874), .Z(n1291) );
  XNOR U2533 ( .A(n1235), .B(n1225), .Z(n1290) );
  XNOR U2534 ( .A(n1230), .B(n1299), .Z(n1231) );
  AND U2535 ( .A(n899), .B(n986), .Z(n1299) );
  XOR U2536 ( .A(n1303), .B(n1232), .Z(n1298) );
  NAND U2537 ( .A(n932), .B(n945), .Z(n1232) );
  IV U2538 ( .A(n1234), .Z(n1303) );
  XNOR U2539 ( .A(n1239), .B(n1308), .Z(n1240) );
  AND U2540 ( .A(n1119), .B(n810), .Z(n1308) );
  XOR U2541 ( .A(n1312), .B(n1241), .Z(n1307) );
  NAND U2542 ( .A(n774), .B(n1180), .Z(n1241) );
  IV U2543 ( .A(n1243), .Z(n1312) );
  XNOR U2544 ( .A(n1250), .B(n1251), .Z(n1245) );
  NANDN U2545 ( .B(n713), .A(n1316), .Z(n1251) );
  XOR U2546 ( .A(n1249), .B(n1317), .Z(n1250) );
  AND U2547 ( .A(n1246), .B(n746), .Z(n1317) );
  NAND U2548 ( .A(n1318), .B(n1319), .Z(n1249) );
  NANDN U2549 ( .B(n1320), .A(n1321), .Z(n1318) );
  XOR U2550 ( .A(n1325), .B(\_MxM/Y0[17] ), .Z(\_MxM/Y1[16] ) );
  XNOR U2551 ( .A(n1326), .B(n1327), .Z(n1325) );
  AND U2552 ( .A(n671), .B(n1329), .Z(n1328) );
  XOR U2553 ( .A(n1323), .B(n1327), .Z(n1329) );
  XNOR U2554 ( .A(n1322), .B(n1327), .Z(n1323) );
  XNOR U2555 ( .A(n1278), .B(n1277), .Z(n1261) );
  XOR U2556 ( .A(n1332), .B(n1289), .Z(n1277) );
  XNOR U2557 ( .A(n1265), .B(n1334), .Z(n1266) );
  AND U2558 ( .A(n778), .B(n1198), .Z(n1334) );
  XOR U2559 ( .A(n1338), .B(n1267), .Z(n1333) );
  NAND U2560 ( .A(n1140), .B(n818), .Z(n1267) );
  IV U2561 ( .A(n1269), .Z(n1338) );
  XNOR U2562 ( .A(n1274), .B(n1275), .Z(n1271) );
  NANDN U2563 ( .B(n1022), .A(n899), .Z(n1275) );
  XNOR U2564 ( .A(n1273), .B(n1342), .Z(n1274) );
  AND U2565 ( .A(n855), .B(n1082), .Z(n1342) );
  XNOR U2566 ( .A(n1288), .B(n1276), .Z(n1332) );
  XNOR U2567 ( .A(n1349), .B(n1281), .Z(n1288) );
  XOR U2568 ( .A(n1350), .B(n1285), .Z(n1281) );
  NAND U2569 ( .A(n1284), .B(n744), .Z(n1285) );
  NANDN U2570 ( .B(n714), .A(n1352), .Z(n1351) );
  XNOR U2571 ( .A(n1362), .B(n1306), .Z(n1296) );
  XNOR U2572 ( .A(n1293), .B(n1294), .Z(n1306) );
  NANDN U2573 ( .B(n836), .A(n1119), .Z(n1294) );
  XNOR U2574 ( .A(n1292), .B(n1363), .Z(n1293) );
  AND U2575 ( .A(n1057), .B(n874), .Z(n1363) );
  XNOR U2576 ( .A(n1305), .B(n1295), .Z(n1362) );
  XNOR U2577 ( .A(n1300), .B(n1371), .Z(n1301) );
  AND U2578 ( .A(n945), .B(n986), .Z(n1371) );
  XOR U2579 ( .A(n1375), .B(n1302), .Z(n1370) );
  NAND U2580 ( .A(n932), .B(n1003), .Z(n1302) );
  IV U2581 ( .A(n1304), .Z(n1375) );
  XNOR U2582 ( .A(n1309), .B(n1380), .Z(n1310) );
  AND U2583 ( .A(n1180), .B(n810), .Z(n1380) );
  XOR U2584 ( .A(n1384), .B(n1311), .Z(n1379) );
  NAND U2585 ( .A(n774), .B(n1246), .Z(n1311) );
  IV U2586 ( .A(n1313), .Z(n1384) );
  XNOR U2587 ( .A(n1320), .B(n1321), .Z(n1315) );
  NANDN U2588 ( .B(n713), .A(n1388), .Z(n1321) );
  XNOR U2589 ( .A(n1319), .B(n1389), .Z(n1320) );
  AND U2590 ( .A(n1316), .B(n746), .Z(n1389) );
  AND U2591 ( .A(n1390), .B(n1391), .Z(n1319) );
  NANDN U2592 ( .B(n1392), .A(n1393), .Z(n1390) );
  XOR U2593 ( .A(n1397), .B(\_MxM/Y0[16] ), .Z(\_MxM/Y1[15] ) );
  XNOR U2594 ( .A(n1398), .B(n1399), .Z(n1397) );
  AND U2595 ( .A(n671), .B(n1401), .Z(n1400) );
  XOR U2596 ( .A(n1395), .B(n1399), .Z(n1401) );
  XNOR U2597 ( .A(n1394), .B(n1399), .Z(n1395) );
  XNOR U2598 ( .A(n1348), .B(n1347), .Z(n1331) );
  XOR U2599 ( .A(n1405), .B(n1358), .Z(n1347) );
  XNOR U2600 ( .A(n1335), .B(n1407), .Z(n1336) );
  AND U2601 ( .A(n818), .B(n1198), .Z(n1407) );
  XOR U2602 ( .A(n1411), .B(n1337), .Z(n1406) );
  NAND U2603 ( .A(n1140), .B(n855), .Z(n1337) );
  IV U2604 ( .A(n1339), .Z(n1411) );
  XNOR U2605 ( .A(n1344), .B(n1345), .Z(n1341) );
  NANDN U2606 ( .B(n1022), .A(n945), .Z(n1345) );
  XNOR U2607 ( .A(n1343), .B(n1415), .Z(n1344) );
  AND U2608 ( .A(n899), .B(n1082), .Z(n1415) );
  XNOR U2609 ( .A(n1357), .B(n1346), .Z(n1405) );
  XNOR U2610 ( .A(n1422), .B(n1361), .Z(n1357) );
  NAND U2611 ( .A(n1284), .B(n778), .Z(n1355) );
  XNOR U2612 ( .A(n1353), .B(n1423), .Z(n1354) );
  AND U2613 ( .A(n744), .B(n1352), .Z(n1423) );
  XNOR U2614 ( .A(n1360), .B(n1356), .Z(n1422) );
  AND U2615 ( .A(n1431), .B(n1432), .Z(n1430) );
  NANDN U2616 ( .B(n714), .A(n1433), .Z(n1432) );
  OR U2617 ( .A(n1434), .B(n1435), .Z(n1431) );
  XNOR U2618 ( .A(n1439), .B(n1378), .Z(n1368) );
  XNOR U2619 ( .A(n1365), .B(n1366), .Z(n1378) );
  NANDN U2620 ( .B(n836), .A(n1180), .Z(n1366) );
  XNOR U2621 ( .A(n1364), .B(n1440), .Z(n1365) );
  AND U2622 ( .A(n1119), .B(n874), .Z(n1440) );
  XNOR U2623 ( .A(n1377), .B(n1367), .Z(n1439) );
  XNOR U2624 ( .A(n1372), .B(n1448), .Z(n1373) );
  AND U2625 ( .A(n1003), .B(n986), .Z(n1448) );
  XOR U2626 ( .A(n1452), .B(n1374), .Z(n1447) );
  NAND U2627 ( .A(n932), .B(n1057), .Z(n1374) );
  IV U2628 ( .A(n1376), .Z(n1452) );
  XNOR U2629 ( .A(n1381), .B(n1457), .Z(n1382) );
  AND U2630 ( .A(n1246), .B(n810), .Z(n1457) );
  XOR U2631 ( .A(n1461), .B(n1383), .Z(n1456) );
  NAND U2632 ( .A(n774), .B(n1316), .Z(n1383) );
  IV U2633 ( .A(n1385), .Z(n1461) );
  XNOR U2634 ( .A(n1392), .B(n1393), .Z(n1387) );
  NANDN U2635 ( .B(n713), .A(n1465), .Z(n1393) );
  XNOR U2636 ( .A(n1391), .B(n1466), .Z(n1392) );
  AND U2637 ( .A(n1388), .B(n746), .Z(n1466) );
  ANDN U2638 ( .A(n1467), .B(n1468), .Z(n1391) );
  NANDN U2639 ( .B(n1469), .A(n1470), .Z(n1467) );
  XOR U2640 ( .A(n1474), .B(\_MxM/Y0[15] ), .Z(\_MxM/Y1[14] ) );
  XNOR U2641 ( .A(n1475), .B(n1476), .Z(n1474) );
  AND U2642 ( .A(n671), .B(n1478), .Z(n1477) );
  XOR U2643 ( .A(n1472), .B(n1476), .Z(n1478) );
  XNOR U2644 ( .A(n1471), .B(n1476), .Z(n1472) );
  XOR U2645 ( .A(n1404), .B(n1403), .Z(n1476) );
  XOR U2646 ( .A(n1479), .B(n1480), .Z(n1403) );
  XOR U2647 ( .A(n1481), .B(n1482), .Z(n1480) );
  XOR U2648 ( .A(n1483), .B(n1481), .Z(n1482) );
  XNOR U2649 ( .A(n1421), .B(n1420), .Z(n1404) );
  XOR U2650 ( .A(n1489), .B(n1429), .Z(n1420) );
  XNOR U2651 ( .A(n1408), .B(n1491), .Z(n1409) );
  AND U2652 ( .A(n855), .B(n1198), .Z(n1491) );
  XOR U2653 ( .A(n1495), .B(n1410), .Z(n1490) );
  NAND U2654 ( .A(n1140), .B(n899), .Z(n1410) );
  IV U2655 ( .A(n1412), .Z(n1495) );
  XNOR U2656 ( .A(n1417), .B(n1418), .Z(n1414) );
  NANDN U2657 ( .B(n1022), .A(n1003), .Z(n1418) );
  XNOR U2658 ( .A(n1416), .B(n1499), .Z(n1417) );
  AND U2659 ( .A(n945), .B(n1082), .Z(n1499) );
  XNOR U2660 ( .A(n1428), .B(n1419), .Z(n1489) );
  XNOR U2661 ( .A(n1506), .B(n1438), .Z(n1428) );
  NAND U2662 ( .A(n1284), .B(n818), .Z(n1426) );
  XNOR U2663 ( .A(n1424), .B(n1507), .Z(n1425) );
  AND U2664 ( .A(n778), .B(n1352), .Z(n1507) );
  XNOR U2665 ( .A(n1437), .B(n1427), .Z(n1506) );
  XNOR U2666 ( .A(n1514), .B(n1436), .Z(n1437) );
  XNOR U2667 ( .A(n1518), .B(n1434), .Z(n1514) );
  NAND U2668 ( .A(n1433), .B(n744), .Z(n1434) );
  NANDN U2669 ( .B(n714), .A(n1520), .Z(n1519) );
  XNOR U2670 ( .A(n1524), .B(n1455), .Z(n1445) );
  XNOR U2671 ( .A(n1442), .B(n1443), .Z(n1455) );
  NANDN U2672 ( .B(n836), .A(n1246), .Z(n1443) );
  XNOR U2673 ( .A(n1441), .B(n1525), .Z(n1442) );
  AND U2674 ( .A(n1180), .B(n874), .Z(n1525) );
  XNOR U2675 ( .A(n1454), .B(n1444), .Z(n1524) );
  XNOR U2676 ( .A(n1449), .B(n1533), .Z(n1450) );
  AND U2677 ( .A(n1057), .B(n986), .Z(n1533) );
  XOR U2678 ( .A(n1537), .B(n1451), .Z(n1532) );
  NAND U2679 ( .A(n932), .B(n1119), .Z(n1451) );
  IV U2680 ( .A(n1453), .Z(n1537) );
  XNOR U2681 ( .A(n1458), .B(n1542), .Z(n1459) );
  AND U2682 ( .A(n1316), .B(n810), .Z(n1542) );
  XOR U2683 ( .A(n1546), .B(n1460), .Z(n1541) );
  NAND U2684 ( .A(n774), .B(n1388), .Z(n1460) );
  IV U2685 ( .A(n1462), .Z(n1546) );
  XNOR U2686 ( .A(n1469), .B(n1470), .Z(n1464) );
  NANDN U2687 ( .B(n713), .A(n1550), .Z(n1470) );
  AND U2688 ( .A(n1465), .B(n746), .Z(n1551) );
  NAND U2689 ( .A(n1552), .B(n1553), .Z(n1468) );
  NANDN U2690 ( .B(n1554), .A(n1555), .Z(n1552) );
  XOR U2691 ( .A(n1559), .B(\_MxM/Y0[14] ), .Z(\_MxM/Y1[13] ) );
  XNOR U2692 ( .A(n1560), .B(n1561), .Z(n1559) );
  AND U2693 ( .A(n671), .B(n1563), .Z(n1562) );
  XOR U2694 ( .A(n1557), .B(n1561), .Z(n1563) );
  XNOR U2695 ( .A(n1556), .B(n1561), .Z(n1557) );
  XNOR U2696 ( .A(n1488), .B(n1487), .Z(n1561) );
  XNOR U2697 ( .A(n1564), .B(n1484), .Z(n1487) );
  NAND U2698 ( .A(n1481), .B(n1567), .Z(n1485) );
  AND U2699 ( .A(n1568), .B(n1569), .Z(n1567) );
  NANDN U2700 ( .B(n714), .A(n1570), .Z(n1569) );
  NANDN U2701 ( .B(n1571), .A(n1572), .Z(n1568) );
  AND U2702 ( .A(n1573), .B(n1574), .Z(n1481) );
  NANDN U2703 ( .B(n1575), .A(n1576), .Z(n1574) );
  NANDN U2704 ( .B(n1577), .A(n1578), .Z(n1573) );
  XNOR U2705 ( .A(n1582), .B(n1513), .Z(n1504) );
  XNOR U2706 ( .A(n1492), .B(n1584), .Z(n1493) );
  AND U2707 ( .A(n899), .B(n1198), .Z(n1584) );
  XOR U2708 ( .A(n1588), .B(n1494), .Z(n1583) );
  NAND U2709 ( .A(n1140), .B(n945), .Z(n1494) );
  IV U2710 ( .A(n1496), .Z(n1588) );
  XNOR U2711 ( .A(n1501), .B(n1502), .Z(n1498) );
  NANDN U2712 ( .B(n1022), .A(n1057), .Z(n1502) );
  XNOR U2713 ( .A(n1500), .B(n1592), .Z(n1501) );
  AND U2714 ( .A(n1003), .B(n1082), .Z(n1592) );
  XNOR U2715 ( .A(n1512), .B(n1503), .Z(n1582) );
  XOR U2716 ( .A(n1599), .B(n1517), .Z(n1512) );
  XNOR U2717 ( .A(n1509), .B(n1510), .Z(n1517) );
  NAND U2718 ( .A(n1284), .B(n855), .Z(n1510) );
  XNOR U2719 ( .A(n1508), .B(n1600), .Z(n1509) );
  AND U2720 ( .A(n818), .B(n1352), .Z(n1600) );
  XNOR U2721 ( .A(n1516), .B(n1511), .Z(n1599) );
  XNOR U2722 ( .A(n1521), .B(n1608), .Z(n1522) );
  AND U2723 ( .A(n744), .B(n1520), .Z(n1608) );
  XOR U2724 ( .A(n1612), .B(n1523), .Z(n1607) );
  NAND U2725 ( .A(n1433), .B(n778), .Z(n1523) );
  IV U2726 ( .A(n1515), .Z(n1612) );
  XNOR U2727 ( .A(n1616), .B(n1540), .Z(n1530) );
  XNOR U2728 ( .A(n1527), .B(n1528), .Z(n1540) );
  NANDN U2729 ( .B(n836), .A(n1316), .Z(n1528) );
  XNOR U2730 ( .A(n1526), .B(n1617), .Z(n1527) );
  AND U2731 ( .A(n1246), .B(n874), .Z(n1617) );
  XNOR U2732 ( .A(n1539), .B(n1529), .Z(n1616) );
  XNOR U2733 ( .A(n1534), .B(n1625), .Z(n1535) );
  AND U2734 ( .A(n1119), .B(n986), .Z(n1625) );
  XOR U2735 ( .A(n1629), .B(n1536), .Z(n1624) );
  NAND U2736 ( .A(n932), .B(n1180), .Z(n1536) );
  IV U2737 ( .A(n1538), .Z(n1629) );
  XNOR U2738 ( .A(n1543), .B(n1634), .Z(n1544) );
  AND U2739 ( .A(n1388), .B(n810), .Z(n1634) );
  XOR U2740 ( .A(n1638), .B(n1545), .Z(n1633) );
  NAND U2741 ( .A(n774), .B(n1465), .Z(n1545) );
  IV U2742 ( .A(n1547), .Z(n1638) );
  XNOR U2743 ( .A(n1554), .B(n1555), .Z(n1549) );
  NANDN U2744 ( .B(n713), .A(n1642), .Z(n1555) );
  XNOR U2745 ( .A(n1553), .B(n1643), .Z(n1554) );
  AND U2746 ( .A(n1550), .B(n746), .Z(n1643) );
  ANDN U2747 ( .A(n1644), .B(n1645), .Z(n1553) );
  NANDN U2748 ( .B(n1646), .A(n1647), .Z(n1644) );
  XOR U2749 ( .A(n1651), .B(\_MxM/Y0[13] ), .Z(\_MxM/Y1[12] ) );
  XNOR U2750 ( .A(n1652), .B(n1653), .Z(n1651) );
  AND U2751 ( .A(n671), .B(n1655), .Z(n1654) );
  XOR U2752 ( .A(n1649), .B(n1653), .Z(n1655) );
  XNOR U2753 ( .A(n1648), .B(n1653), .Z(n1649) );
  XNOR U2754 ( .A(n1581), .B(n1580), .Z(n1653) );
  XNOR U2755 ( .A(n1656), .B(n1566), .Z(n1580) );
  XNOR U2756 ( .A(n1572), .B(n1571), .Z(n1566) );
  OR U2757 ( .A(n1657), .B(n1658), .Z(n1571) );
  XNOR U2758 ( .A(n1575), .B(n1576), .Z(n1572) );
  XOR U2759 ( .A(n1662), .B(n1577), .Z(n1575) );
  NAND U2760 ( .A(n744), .B(n1570), .Z(n1577) );
  NANDN U2761 ( .B(n1578), .A(n1663), .Z(n1662) );
  NANDN U2762 ( .B(n714), .A(n1664), .Z(n1663) );
  XNOR U2763 ( .A(n1673), .B(n1606), .Z(n1597) );
  XNOR U2764 ( .A(n1585), .B(n1675), .Z(n1586) );
  AND U2765 ( .A(n945), .B(n1198), .Z(n1675) );
  XOR U2766 ( .A(n1679), .B(n1587), .Z(n1674) );
  NAND U2767 ( .A(n1140), .B(n1003), .Z(n1587) );
  IV U2768 ( .A(n1589), .Z(n1679) );
  XOR U2769 ( .A(n1680), .B(n1681), .Z(n1589) );
  ANDN U2770 ( .A(n1682), .B(n1683), .Z(n1681) );
  XOR U2771 ( .A(n1680), .B(n1684), .Z(n1682) );
  XNOR U2772 ( .A(n1594), .B(n1595), .Z(n1591) );
  NANDN U2773 ( .B(n1022), .A(n1119), .Z(n1595) );
  XNOR U2774 ( .A(n1593), .B(n1685), .Z(n1594) );
  AND U2775 ( .A(n1057), .B(n1082), .Z(n1685) );
  XNOR U2776 ( .A(n1605), .B(n1596), .Z(n1673) );
  XOR U2777 ( .A(n1692), .B(n1615), .Z(n1605) );
  XNOR U2778 ( .A(n1602), .B(n1603), .Z(n1615) );
  NAND U2779 ( .A(n1284), .B(n899), .Z(n1603) );
  XNOR U2780 ( .A(n1601), .B(n1693), .Z(n1602) );
  AND U2781 ( .A(n855), .B(n1352), .Z(n1693) );
  XNOR U2782 ( .A(n1614), .B(n1604), .Z(n1692) );
  XNOR U2783 ( .A(n1609), .B(n1701), .Z(n1610) );
  AND U2784 ( .A(n778), .B(n1520), .Z(n1701) );
  XOR U2785 ( .A(n1705), .B(n1611), .Z(n1700) );
  NAND U2786 ( .A(n1433), .B(n818), .Z(n1611) );
  IV U2787 ( .A(n1613), .Z(n1705) );
  XNOR U2788 ( .A(n1709), .B(n1632), .Z(n1622) );
  XNOR U2789 ( .A(n1619), .B(n1620), .Z(n1632) );
  NANDN U2790 ( .B(n836), .A(n1388), .Z(n1620) );
  XNOR U2791 ( .A(n1618), .B(n1710), .Z(n1619) );
  AND U2792 ( .A(n1316), .B(n874), .Z(n1710) );
  XNOR U2793 ( .A(n1631), .B(n1621), .Z(n1709) );
  XNOR U2794 ( .A(n1626), .B(n1718), .Z(n1627) );
  AND U2795 ( .A(n1180), .B(n986), .Z(n1718) );
  XOR U2796 ( .A(n1722), .B(n1628), .Z(n1717) );
  NAND U2797 ( .A(n932), .B(n1246), .Z(n1628) );
  IV U2798 ( .A(n1630), .Z(n1722) );
  XNOR U2799 ( .A(n1635), .B(n1727), .Z(n1636) );
  AND U2800 ( .A(n1465), .B(n810), .Z(n1727) );
  XOR U2801 ( .A(n1731), .B(n1637), .Z(n1726) );
  NAND U2802 ( .A(n774), .B(n1550), .Z(n1637) );
  IV U2803 ( .A(n1639), .Z(n1731) );
  XOR U2804 ( .A(n1732), .B(n1733), .Z(n1639) );
  ANDN U2805 ( .A(n1734), .B(n1735), .Z(n1733) );
  XOR U2806 ( .A(n1732), .B(n1736), .Z(n1734) );
  XNOR U2807 ( .A(n1646), .B(n1647), .Z(n1641) );
  NANDN U2808 ( .B(n713), .A(n1737), .Z(n1647) );
  AND U2809 ( .A(n1642), .B(n746), .Z(n1738) );
  NAND U2810 ( .A(n1739), .B(n1740), .Z(n1645) );
  NANDN U2811 ( .B(n1741), .A(n1742), .Z(n1739) );
  XOR U2812 ( .A(n1746), .B(\_MxM/Y0[12] ), .Z(\_MxM/Y1[11] ) );
  XNOR U2813 ( .A(n1747), .B(n1748), .Z(n1746) );
  AND U2814 ( .A(n671), .B(n1750), .Z(n1749) );
  XOR U2815 ( .A(n1744), .B(n1748), .Z(n1750) );
  XNOR U2816 ( .A(n1743), .B(n1748), .Z(n1744) );
  XNOR U2817 ( .A(n1670), .B(n1669), .Z(n1748) );
  XNOR U2818 ( .A(n1751), .B(n1672), .Z(n1669) );
  XOR U2819 ( .A(n1658), .B(n1657), .Z(n1672) );
  NANDN U2820 ( .B(n1752), .A(n1753), .Z(n1657) );
  XOR U2821 ( .A(n1661), .B(n1660), .Z(n1658) );
  XOR U2822 ( .A(n1659), .B(n1754), .Z(n1660) );
  AND U2823 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U2824 ( .B(n714), .A(n1757), .Z(n1756) );
  OR U2825 ( .A(n1758), .B(n1759), .Z(n1755) );
  NAND U2826 ( .A(n778), .B(n1570), .Z(n1667) );
  XNOR U2827 ( .A(n1665), .B(n1762), .Z(n1666) );
  AND U2828 ( .A(n1664), .B(n744), .Z(n1762) );
  XNOR U2829 ( .A(n1771), .B(n1699), .Z(n1690) );
  XNOR U2830 ( .A(n1676), .B(n1773), .Z(n1677) );
  AND U2831 ( .A(n1003), .B(n1198), .Z(n1773) );
  XOR U2832 ( .A(n1777), .B(n1678), .Z(n1772) );
  NAND U2833 ( .A(n1140), .B(n1057), .Z(n1678) );
  IV U2834 ( .A(n1680), .Z(n1777) );
  XNOR U2835 ( .A(n1687), .B(n1688), .Z(n1684) );
  NANDN U2836 ( .B(n1022), .A(n1180), .Z(n1688) );
  XNOR U2837 ( .A(n1686), .B(n1781), .Z(n1687) );
  AND U2838 ( .A(n1119), .B(n1082), .Z(n1781) );
  XNOR U2839 ( .A(n1698), .B(n1689), .Z(n1771) );
  XOR U2840 ( .A(n1788), .B(n1708), .Z(n1698) );
  XNOR U2841 ( .A(n1695), .B(n1696), .Z(n1708) );
  NAND U2842 ( .A(n1284), .B(n945), .Z(n1696) );
  XNOR U2843 ( .A(n1694), .B(n1789), .Z(n1695) );
  AND U2844 ( .A(n899), .B(n1352), .Z(n1789) );
  XNOR U2845 ( .A(n1707), .B(n1697), .Z(n1788) );
  XNOR U2846 ( .A(n1702), .B(n1797), .Z(n1703) );
  AND U2847 ( .A(n818), .B(n1520), .Z(n1797) );
  XOR U2848 ( .A(n1801), .B(n1704), .Z(n1796) );
  NAND U2849 ( .A(n1433), .B(n855), .Z(n1704) );
  IV U2850 ( .A(n1706), .Z(n1801) );
  XNOR U2851 ( .A(n1805), .B(n1725), .Z(n1715) );
  XNOR U2852 ( .A(n1712), .B(n1713), .Z(n1725) );
  NANDN U2853 ( .B(n836), .A(n1465), .Z(n1713) );
  XNOR U2854 ( .A(n1711), .B(n1806), .Z(n1712) );
  AND U2855 ( .A(n1388), .B(n874), .Z(n1806) );
  XNOR U2856 ( .A(n1724), .B(n1714), .Z(n1805) );
  XNOR U2857 ( .A(n1719), .B(n1814), .Z(n1720) );
  AND U2858 ( .A(n1246), .B(n986), .Z(n1814) );
  XOR U2859 ( .A(n1818), .B(n1721), .Z(n1813) );
  NAND U2860 ( .A(n932), .B(n1316), .Z(n1721) );
  IV U2861 ( .A(n1723), .Z(n1818) );
  XNOR U2862 ( .A(n1728), .B(n1823), .Z(n1729) );
  AND U2863 ( .A(n1550), .B(n810), .Z(n1823) );
  XOR U2864 ( .A(n1827), .B(n1730), .Z(n1822) );
  NAND U2865 ( .A(n774), .B(n1642), .Z(n1730) );
  IV U2866 ( .A(n1732), .Z(n1827) );
  XNOR U2867 ( .A(n1741), .B(n1742), .Z(n1736) );
  NANDN U2868 ( .B(n713), .A(n1831), .Z(n1742) );
  XNOR U2869 ( .A(n1740), .B(n1832), .Z(n1741) );
  AND U2870 ( .A(n1737), .B(n746), .Z(n1832) );
  ANDN U2871 ( .A(n1833), .B(n1834), .Z(n1740) );
  NANDN U2872 ( .B(n1835), .A(n1836), .Z(n1833) );
  XOR U2873 ( .A(n1840), .B(\_MxM/Y0[11] ), .Z(\_MxM/Y1[10] ) );
  XNOR U2874 ( .A(n1841), .B(n1842), .Z(n1840) );
  AND U2875 ( .A(n671), .B(n1844), .Z(n1843) );
  XOR U2876 ( .A(n1838), .B(n1842), .Z(n1844) );
  XNOR U2877 ( .A(n1837), .B(n1842), .Z(n1838) );
  XNOR U2878 ( .A(n1768), .B(n1767), .Z(n1842) );
  XNOR U2879 ( .A(n1845), .B(n1770), .Z(n1767) );
  XNOR U2880 ( .A(n1752), .B(n1753), .Z(n1770) );
  XOR U2881 ( .A(n1761), .B(n1760), .Z(n1752) );
  XNOR U2882 ( .A(n1849), .B(n1850), .Z(n1760) );
  ANDN U2883 ( .A(n1853), .B(n1854), .Z(n1852) );
  XOR U2884 ( .A(n1851), .B(n1855), .Z(n1853) );
  XNOR U2885 ( .A(n1856), .B(n1758), .Z(n1849) );
  NAND U2886 ( .A(n744), .B(n1757), .Z(n1758) );
  NANDN U2887 ( .B(n714), .A(n1858), .Z(n1857) );
  NAND U2888 ( .A(n818), .B(n1570), .Z(n1765) );
  XNOR U2889 ( .A(n1763), .B(n1862), .Z(n1764) );
  AND U2890 ( .A(n1664), .B(n778), .Z(n1862) );
  XNOR U2891 ( .A(n1871), .B(n1795), .Z(n1786) );
  XNOR U2892 ( .A(n1774), .B(n1873), .Z(n1775) );
  AND U2893 ( .A(n1057), .B(n1198), .Z(n1873) );
  XOR U2894 ( .A(n1877), .B(n1776), .Z(n1872) );
  NAND U2895 ( .A(n1140), .B(n1119), .Z(n1776) );
  IV U2896 ( .A(n1778), .Z(n1877) );
  XNOR U2897 ( .A(n1783), .B(n1784), .Z(n1780) );
  NANDN U2898 ( .B(n1022), .A(n1246), .Z(n1784) );
  XNOR U2899 ( .A(n1782), .B(n1881), .Z(n1783) );
  AND U2900 ( .A(n1180), .B(n1082), .Z(n1881) );
  XNOR U2901 ( .A(n1794), .B(n1785), .Z(n1871) );
  XOR U2902 ( .A(n1888), .B(n1804), .Z(n1794) );
  XNOR U2903 ( .A(n1791), .B(n1792), .Z(n1804) );
  NAND U2904 ( .A(n1284), .B(n1003), .Z(n1792) );
  XNOR U2905 ( .A(n1790), .B(n1889), .Z(n1791) );
  AND U2906 ( .A(n945), .B(n1352), .Z(n1889) );
  XNOR U2907 ( .A(n1803), .B(n1793), .Z(n1888) );
  XNOR U2908 ( .A(n1798), .B(n1897), .Z(n1799) );
  AND U2909 ( .A(n855), .B(n1520), .Z(n1897) );
  XOR U2910 ( .A(n1901), .B(n1800), .Z(n1896) );
  NAND U2911 ( .A(n1433), .B(n899), .Z(n1800) );
  IV U2912 ( .A(n1802), .Z(n1901) );
  XNOR U2913 ( .A(n1905), .B(n1821), .Z(n1811) );
  XNOR U2914 ( .A(n1808), .B(n1809), .Z(n1821) );
  NANDN U2915 ( .B(n836), .A(n1550), .Z(n1809) );
  XNOR U2916 ( .A(n1807), .B(n1906), .Z(n1808) );
  AND U2917 ( .A(n1465), .B(n874), .Z(n1906) );
  XNOR U2918 ( .A(n1820), .B(n1810), .Z(n1905) );
  XNOR U2919 ( .A(n1815), .B(n1914), .Z(n1816) );
  AND U2920 ( .A(n1316), .B(n986), .Z(n1914) );
  XOR U2921 ( .A(n1918), .B(n1817), .Z(n1913) );
  NAND U2922 ( .A(n932), .B(n1388), .Z(n1817) );
  IV U2923 ( .A(n1819), .Z(n1918) );
  XNOR U2924 ( .A(n1824), .B(n1923), .Z(n1825) );
  AND U2925 ( .A(n1642), .B(n810), .Z(n1923) );
  XOR U2926 ( .A(n1927), .B(n1826), .Z(n1922) );
  NAND U2927 ( .A(n774), .B(n1737), .Z(n1826) );
  IV U2928 ( .A(n1828), .Z(n1927) );
  XNOR U2929 ( .A(n1835), .B(n1836), .Z(n1830) );
  NANDN U2930 ( .B(n713), .A(n1931), .Z(n1836) );
  AND U2931 ( .A(n1831), .B(n746), .Z(n1932) );
  NAND U2932 ( .A(n1933), .B(n1934), .Z(n1834) );
  NANDN U2933 ( .B(n1935), .A(n1936), .Z(n1933) );
  XNOR U2934 ( .A(n1940), .B(n1941), .Z(n655) );
  AND U2935 ( .A(n671), .B(n1943), .Z(n1942) );
  XOR U2936 ( .A(n1938), .B(n1941), .Z(n1943) );
  XNOR U2937 ( .A(n1937), .B(n1941), .Z(n1938) );
  XNOR U2938 ( .A(n1868), .B(n1867), .Z(n1941) );
  XNOR U2939 ( .A(n1944), .B(n1870), .Z(n1867) );
  XNOR U2940 ( .A(n1848), .B(n1847), .Z(n1870) );
  XNOR U2941 ( .A(n1846), .B(n1945), .Z(n1847) );
  AND U2942 ( .A(n1946), .B(n1947), .Z(n1945) );
  OR U2943 ( .A(n1948), .B(n1949), .Z(n1947) );
  AND U2944 ( .A(n1950), .B(n1951), .Z(n1946) );
  NANDN U2945 ( .B(n714), .A(n1952), .Z(n1951) );
  NAND U2946 ( .A(n1953), .B(n1954), .Z(n1950) );
  XNOR U2947 ( .A(n1859), .B(n1959), .Z(n1860) );
  AND U2948 ( .A(n1858), .B(n744), .Z(n1959) );
  XOR U2949 ( .A(n1963), .B(n1861), .Z(n1958) );
  NAND U2950 ( .A(n778), .B(n1757), .Z(n1861) );
  IV U2951 ( .A(n1851), .Z(n1963) );
  XNOR U2952 ( .A(n1864), .B(n1865), .Z(n1855) );
  NAND U2953 ( .A(n855), .B(n1570), .Z(n1865) );
  XNOR U2954 ( .A(n1863), .B(n1967), .Z(n1864) );
  AND U2955 ( .A(n1664), .B(n818), .Z(n1967) );
  XNOR U2956 ( .A(n1976), .B(n1895), .Z(n1886) );
  XNOR U2957 ( .A(n1874), .B(n1978), .Z(n1875) );
  AND U2958 ( .A(n1119), .B(n1198), .Z(n1978) );
  XOR U2959 ( .A(n1982), .B(n1876), .Z(n1977) );
  NAND U2960 ( .A(n1140), .B(n1180), .Z(n1876) );
  IV U2961 ( .A(n1878), .Z(n1982) );
  XNOR U2962 ( .A(n1883), .B(n1884), .Z(n1880) );
  NANDN U2963 ( .B(n1022), .A(n1316), .Z(n1884) );
  XNOR U2964 ( .A(n1882), .B(n1986), .Z(n1883) );
  AND U2965 ( .A(n1246), .B(n1082), .Z(n1986) );
  XNOR U2966 ( .A(n1894), .B(n1885), .Z(n1976) );
  XOR U2967 ( .A(n1993), .B(n1904), .Z(n1894) );
  XNOR U2968 ( .A(n1891), .B(n1892), .Z(n1904) );
  NAND U2969 ( .A(n1284), .B(n1057), .Z(n1892) );
  XNOR U2970 ( .A(n1890), .B(n1994), .Z(n1891) );
  AND U2971 ( .A(n1003), .B(n1352), .Z(n1994) );
  XNOR U2972 ( .A(n1903), .B(n1893), .Z(n1993) );
  XNOR U2973 ( .A(n1898), .B(n2002), .Z(n1899) );
  AND U2974 ( .A(n899), .B(n1520), .Z(n2002) );
  XOR U2975 ( .A(n2006), .B(n1900), .Z(n2001) );
  NAND U2976 ( .A(n1433), .B(n945), .Z(n1900) );
  IV U2977 ( .A(n1902), .Z(n2006) );
  XNOR U2978 ( .A(n2010), .B(n1921), .Z(n1911) );
  XNOR U2979 ( .A(n1908), .B(n1909), .Z(n1921) );
  NANDN U2980 ( .B(n836), .A(n1642), .Z(n1909) );
  XNOR U2981 ( .A(n1907), .B(n2011), .Z(n1908) );
  AND U2982 ( .A(n1550), .B(n874), .Z(n2011) );
  XNOR U2983 ( .A(n1920), .B(n1910), .Z(n2010) );
  XNOR U2984 ( .A(n1915), .B(n2019), .Z(n1916) );
  AND U2985 ( .A(n1388), .B(n986), .Z(n2019) );
  XOR U2986 ( .A(n2023), .B(n1917), .Z(n2018) );
  NAND U2987 ( .A(n932), .B(n1465), .Z(n1917) );
  IV U2988 ( .A(n1919), .Z(n2023) );
  XNOR U2989 ( .A(n1924), .B(n2028), .Z(n1925) );
  AND U2990 ( .A(n1737), .B(n810), .Z(n2028) );
  XOR U2991 ( .A(n2032), .B(n1926), .Z(n2027) );
  NAND U2992 ( .A(n774), .B(n1831), .Z(n1926) );
  IV U2993 ( .A(n1928), .Z(n2032) );
  XNOR U2994 ( .A(n1935), .B(n1936), .Z(n1930) );
  NANDN U2995 ( .B(n713), .A(n2036), .Z(n1936) );
  XNOR U2996 ( .A(n1934), .B(n2037), .Z(n1935) );
  AND U2997 ( .A(n1931), .B(n746), .Z(n2037) );
  ANDN U2998 ( .A(n2038), .B(n2039), .Z(n1934) );
  NANDN U2999 ( .B(n2040), .A(n2041), .Z(n2038) );
  XNOR U3000 ( .A(n2045), .B(n2046), .Z(n656) );
  AND U3001 ( .A(n671), .B(n2048), .Z(n2047) );
  XOR U3002 ( .A(n2043), .B(n2046), .Z(n2048) );
  XNOR U3003 ( .A(n2042), .B(n2046), .Z(n2043) );
  XNOR U3004 ( .A(n1973), .B(n1972), .Z(n2046) );
  XNOR U3005 ( .A(n2049), .B(n1975), .Z(n1972) );
  XNOR U3006 ( .A(n1957), .B(n1956), .Z(n1975) );
  XNOR U3007 ( .A(n2050), .B(n1953), .Z(n1956) );
  XNOR U3008 ( .A(n2051), .B(n1948), .Z(n1953) );
  NAND U3009 ( .A(n744), .B(n1952), .Z(n1948) );
  NANDN U3010 ( .B(n714), .A(n2053), .Z(n2052) );
  XNOR U3011 ( .A(n1954), .B(n1955), .Z(n2050) );
  XNOR U3012 ( .A(n1960), .B(n2064), .Z(n1961) );
  AND U3013 ( .A(n1858), .B(n778), .Z(n2064) );
  XOR U3014 ( .A(n2068), .B(n1962), .Z(n2063) );
  NAND U3015 ( .A(n818), .B(n1757), .Z(n1962) );
  IV U3016 ( .A(n1964), .Z(n2068) );
  XNOR U3017 ( .A(n1969), .B(n1970), .Z(n1966) );
  NAND U3018 ( .A(n899), .B(n1570), .Z(n1970) );
  XNOR U3019 ( .A(n1968), .B(n2072), .Z(n1969) );
  AND U3020 ( .A(n1664), .B(n855), .Z(n2072) );
  XNOR U3021 ( .A(n2081), .B(n2000), .Z(n1991) );
  XNOR U3022 ( .A(n1979), .B(n2083), .Z(n1980) );
  AND U3023 ( .A(n1180), .B(n1198), .Z(n2083) );
  XOR U3024 ( .A(n2087), .B(n1981), .Z(n2082) );
  NAND U3025 ( .A(n1140), .B(n1246), .Z(n1981) );
  IV U3026 ( .A(n1983), .Z(n2087) );
  XNOR U3027 ( .A(n1988), .B(n1989), .Z(n1985) );
  NANDN U3028 ( .B(n1022), .A(n1388), .Z(n1989) );
  XNOR U3029 ( .A(n1987), .B(n2091), .Z(n1988) );
  AND U3030 ( .A(n1316), .B(n1082), .Z(n2091) );
  XNOR U3031 ( .A(n1999), .B(n1990), .Z(n2081) );
  XOR U3032 ( .A(n2098), .B(n2009), .Z(n1999) );
  XNOR U3033 ( .A(n1996), .B(n1997), .Z(n2009) );
  NAND U3034 ( .A(n1284), .B(n1119), .Z(n1997) );
  XNOR U3035 ( .A(n1995), .B(n2099), .Z(n1996) );
  AND U3036 ( .A(n1057), .B(n1352), .Z(n2099) );
  XNOR U3037 ( .A(n2008), .B(n1998), .Z(n2098) );
  XNOR U3038 ( .A(n2003), .B(n2107), .Z(n2004) );
  AND U3039 ( .A(n945), .B(n1520), .Z(n2107) );
  XOR U3040 ( .A(n2111), .B(n2005), .Z(n2106) );
  NAND U3041 ( .A(n1433), .B(n1003), .Z(n2005) );
  IV U3042 ( .A(n2007), .Z(n2111) );
  XNOR U3043 ( .A(n2115), .B(n2026), .Z(n2016) );
  XNOR U3044 ( .A(n2013), .B(n2014), .Z(n2026) );
  NANDN U3045 ( .B(n836), .A(n1737), .Z(n2014) );
  XNOR U3046 ( .A(n2012), .B(n2116), .Z(n2013) );
  AND U3047 ( .A(n1642), .B(n874), .Z(n2116) );
  XNOR U3048 ( .A(n2025), .B(n2015), .Z(n2115) );
  XNOR U3049 ( .A(n2020), .B(n2124), .Z(n2021) );
  AND U3050 ( .A(n1465), .B(n986), .Z(n2124) );
  XOR U3051 ( .A(n2128), .B(n2022), .Z(n2123) );
  NAND U3052 ( .A(n932), .B(n1550), .Z(n2022) );
  IV U3053 ( .A(n2024), .Z(n2128) );
  XNOR U3054 ( .A(n2029), .B(n2133), .Z(n2030) );
  AND U3055 ( .A(n1831), .B(n810), .Z(n2133) );
  XOR U3056 ( .A(n2137), .B(n2031), .Z(n2132) );
  NAND U3057 ( .A(n774), .B(n1931), .Z(n2031) );
  IV U3058 ( .A(n2033), .Z(n2137) );
  XNOR U3059 ( .A(n2040), .B(n2041), .Z(n2035) );
  NANDN U3060 ( .B(n713), .A(n2141), .Z(n2041) );
  AND U3061 ( .A(n2036), .B(n746), .Z(n2142) );
  NAND U3062 ( .A(n2143), .B(n2144), .Z(n2039) );
  NANDN U3063 ( .B(n2145), .A(n2146), .Z(n2143) );
  XNOR U3064 ( .A(n2150), .B(n2151), .Z(n657) );
  AND U3065 ( .A(n671), .B(n2153), .Z(n2152) );
  XOR U3066 ( .A(n2148), .B(n2151), .Z(n2153) );
  XNOR U3067 ( .A(n2147), .B(n2151), .Z(n2148) );
  XNOR U3068 ( .A(n2078), .B(n2077), .Z(n2151) );
  XNOR U3069 ( .A(n2154), .B(n2080), .Z(n2077) );
  XNOR U3070 ( .A(n2059), .B(n2058), .Z(n2080) );
  XNOR U3071 ( .A(n2155), .B(n2062), .Z(n2058) );
  XNOR U3072 ( .A(n2055), .B(n2056), .Z(n2062) );
  NAND U3073 ( .A(n778), .B(n1952), .Z(n2056) );
  XNOR U3074 ( .A(n2054), .B(n2156), .Z(n2055) );
  AND U3075 ( .A(n2053), .B(n744), .Z(n2156) );
  XNOR U3076 ( .A(n2061), .B(n2057), .Z(n2155) );
  AND U3077 ( .A(n2164), .B(n2165), .Z(n2163) );
  NANDN U3078 ( .B(n714), .A(n2166), .Z(n2165) );
  OR U3079 ( .A(n2167), .B(n2168), .Z(n2164) );
  XNOR U3080 ( .A(n2065), .B(n2173), .Z(n2066) );
  AND U3081 ( .A(n1858), .B(n818), .Z(n2173) );
  XOR U3082 ( .A(n2177), .B(n2067), .Z(n2172) );
  NAND U3083 ( .A(n855), .B(n1757), .Z(n2067) );
  IV U3084 ( .A(n2069), .Z(n2177) );
  XNOR U3085 ( .A(n2074), .B(n2075), .Z(n2071) );
  NAND U3086 ( .A(n945), .B(n1570), .Z(n2075) );
  XNOR U3087 ( .A(n2073), .B(n2181), .Z(n2074) );
  AND U3088 ( .A(n1664), .B(n899), .Z(n2181) );
  XNOR U3089 ( .A(n2191), .B(n2188), .Z(n2190) );
  XNOR U3090 ( .A(n2192), .B(n2105), .Z(n2096) );
  XNOR U3091 ( .A(n2084), .B(n2194), .Z(n2085) );
  AND U3092 ( .A(n1246), .B(n1198), .Z(n2194) );
  XOR U3093 ( .A(n2198), .B(n2086), .Z(n2193) );
  NAND U3094 ( .A(n1140), .B(n1316), .Z(n2086) );
  IV U3095 ( .A(n2088), .Z(n2198) );
  XNOR U3096 ( .A(n2093), .B(n2094), .Z(n2090) );
  NANDN U3097 ( .B(n1022), .A(n1465), .Z(n2094) );
  XNOR U3098 ( .A(n2092), .B(n2202), .Z(n2093) );
  AND U3099 ( .A(n1388), .B(n1082), .Z(n2202) );
  XNOR U3100 ( .A(n2104), .B(n2095), .Z(n2192) );
  XOR U3101 ( .A(n2209), .B(n2114), .Z(n2104) );
  XNOR U3102 ( .A(n2101), .B(n2102), .Z(n2114) );
  NAND U3103 ( .A(n1284), .B(n1180), .Z(n2102) );
  XNOR U3104 ( .A(n2100), .B(n2210), .Z(n2101) );
  AND U3105 ( .A(n1119), .B(n1352), .Z(n2210) );
  XNOR U3106 ( .A(n2113), .B(n2103), .Z(n2209) );
  XNOR U3107 ( .A(n2108), .B(n2218), .Z(n2109) );
  AND U3108 ( .A(n1003), .B(n1520), .Z(n2218) );
  XOR U3109 ( .A(n2222), .B(n2110), .Z(n2217) );
  NAND U3110 ( .A(n1433), .B(n1057), .Z(n2110) );
  IV U3111 ( .A(n2112), .Z(n2222) );
  XNOR U3112 ( .A(n2226), .B(n2131), .Z(n2121) );
  XNOR U3113 ( .A(n2118), .B(n2119), .Z(n2131) );
  NANDN U3114 ( .B(n836), .A(n1831), .Z(n2119) );
  XNOR U3115 ( .A(n2117), .B(n2227), .Z(n2118) );
  AND U3116 ( .A(n1737), .B(n874), .Z(n2227) );
  XNOR U3117 ( .A(n2130), .B(n2120), .Z(n2226) );
  XNOR U3118 ( .A(n2125), .B(n2235), .Z(n2126) );
  AND U3119 ( .A(n1550), .B(n986), .Z(n2235) );
  XOR U3120 ( .A(n2239), .B(n2127), .Z(n2234) );
  NAND U3121 ( .A(n932), .B(n1642), .Z(n2127) );
  IV U3122 ( .A(n2129), .Z(n2239) );
  XNOR U3123 ( .A(n2134), .B(n2244), .Z(n2135) );
  AND U3124 ( .A(n1931), .B(n810), .Z(n2244) );
  XOR U3125 ( .A(n2245), .B(n2246), .Z(n2134) );
  ANDN U3126 ( .A(n2247), .B(n2248), .Z(n2246) );
  XNOR U3127 ( .A(n2249), .B(n2245), .Z(n2247) );
  XOR U3128 ( .A(n2250), .B(n2136), .Z(n2243) );
  NAND U3129 ( .A(n774), .B(n2036), .Z(n2136) );
  IV U3130 ( .A(n2138), .Z(n2250) );
  XNOR U3131 ( .A(n2145), .B(n2146), .Z(n2140) );
  NANDN U3132 ( .B(n713), .A(n2254), .Z(n2146) );
  XNOR U3133 ( .A(n2144), .B(n2255), .Z(n2145) );
  AND U3134 ( .A(n2141), .B(n746), .Z(n2255) );
  ANDN U3135 ( .A(n2256), .B(n2257), .Z(n2144) );
  NANDN U3136 ( .B(n2258), .A(n2259), .Z(n2256) );
  XNOR U3137 ( .A(n2263), .B(n2264), .Z(n658) );
  AND U3138 ( .A(n671), .B(n2266), .Z(n2265) );
  XOR U3139 ( .A(n2261), .B(n2264), .Z(n2266) );
  XNOR U3140 ( .A(n2260), .B(n2264), .Z(n2261) );
  XNOR U3141 ( .A(n2187), .B(n2186), .Z(n2264) );
  XNOR U3142 ( .A(n2267), .B(n2191), .Z(n2186) );
  XNOR U3143 ( .A(n2162), .B(n2161), .Z(n2191) );
  XNOR U3144 ( .A(n2268), .B(n2171), .Z(n2161) );
  XNOR U3145 ( .A(n2158), .B(n2159), .Z(n2171) );
  NAND U3146 ( .A(n818), .B(n1952), .Z(n2159) );
  XNOR U3147 ( .A(n2157), .B(n2269), .Z(n2158) );
  AND U3148 ( .A(n2053), .B(n778), .Z(n2269) );
  XNOR U3149 ( .A(n2170), .B(n2160), .Z(n2268) );
  XNOR U3150 ( .A(n2276), .B(n2169), .Z(n2170) );
  XNOR U3151 ( .A(n2280), .B(n2167), .Z(n2276) );
  NAND U3152 ( .A(n744), .B(n2166), .Z(n2167) );
  NANDN U3153 ( .B(n714), .A(n2282), .Z(n2281) );
  XNOR U3154 ( .A(n2174), .B(n2287), .Z(n2175) );
  AND U3155 ( .A(n1858), .B(n855), .Z(n2287) );
  XOR U3156 ( .A(n2291), .B(n2176), .Z(n2286) );
  NAND U3157 ( .A(n899), .B(n1757), .Z(n2176) );
  IV U3158 ( .A(n2178), .Z(n2291) );
  XNOR U3159 ( .A(n2183), .B(n2184), .Z(n2180) );
  NAND U3160 ( .A(n1003), .B(n1570), .Z(n2184) );
  XNOR U3161 ( .A(n2182), .B(n2295), .Z(n2183) );
  AND U3162 ( .A(n1664), .B(n945), .Z(n2295) );
  XNOR U3163 ( .A(n2189), .B(n2185), .Z(n2267) );
  XOR U3164 ( .A(n2306), .B(n2307), .Z(n2302) );
  NANDN U3165 ( .B(n2308), .A(n2309), .Z(n2306) );
  XNOR U3166 ( .A(n2310), .B(n2216), .Z(n2207) );
  XNOR U3167 ( .A(n2195), .B(n2312), .Z(n2196) );
  AND U3168 ( .A(n1316), .B(n1198), .Z(n2312) );
  XOR U3169 ( .A(n2316), .B(n2197), .Z(n2311) );
  NAND U3170 ( .A(n1140), .B(n1388), .Z(n2197) );
  IV U3171 ( .A(n2199), .Z(n2316) );
  XNOR U3172 ( .A(n2204), .B(n2205), .Z(n2201) );
  NANDN U3173 ( .B(n1022), .A(n1550), .Z(n2205) );
  XNOR U3174 ( .A(n2203), .B(n2320), .Z(n2204) );
  AND U3175 ( .A(n1465), .B(n1082), .Z(n2320) );
  XNOR U3176 ( .A(n2215), .B(n2206), .Z(n2310) );
  XOR U3177 ( .A(n2327), .B(n2225), .Z(n2215) );
  XNOR U3178 ( .A(n2212), .B(n2213), .Z(n2225) );
  NAND U3179 ( .A(n1284), .B(n1246), .Z(n2213) );
  XNOR U3180 ( .A(n2211), .B(n2328), .Z(n2212) );
  AND U3181 ( .A(n1180), .B(n1352), .Z(n2328) );
  XNOR U3182 ( .A(n2224), .B(n2214), .Z(n2327) );
  XNOR U3183 ( .A(n2219), .B(n2336), .Z(n2220) );
  AND U3184 ( .A(n1057), .B(n1520), .Z(n2336) );
  XOR U3185 ( .A(n2340), .B(n2221), .Z(n2335) );
  NAND U3186 ( .A(n1433), .B(n1119), .Z(n2221) );
  IV U3187 ( .A(n2223), .Z(n2340) );
  XNOR U3188 ( .A(n2344), .B(n2242), .Z(n2232) );
  XNOR U3189 ( .A(n2229), .B(n2230), .Z(n2242) );
  NANDN U3190 ( .B(n836), .A(n1931), .Z(n2230) );
  XNOR U3191 ( .A(n2228), .B(n2345), .Z(n2229) );
  AND U3192 ( .A(n1831), .B(n874), .Z(n2345) );
  XNOR U3193 ( .A(n2241), .B(n2231), .Z(n2344) );
  XNOR U3194 ( .A(n2236), .B(n2353), .Z(n2237) );
  AND U3195 ( .A(n1642), .B(n986), .Z(n2353) );
  XOR U3196 ( .A(n2357), .B(n2238), .Z(n2352) );
  NAND U3197 ( .A(n932), .B(n1737), .Z(n2238) );
  IV U3198 ( .A(n2240), .Z(n2357) );
  XNOR U3199 ( .A(n2245), .B(n2362), .Z(n2248) );
  AND U3200 ( .A(n2036), .B(n810), .Z(n2362) );
  XOR U3201 ( .A(n2366), .B(n2249), .Z(n2361) );
  NAND U3202 ( .A(n774), .B(n2141), .Z(n2249) );
  IV U3203 ( .A(n2251), .Z(n2366) );
  XNOR U3204 ( .A(n2258), .B(n2259), .Z(n2253) );
  NANDN U3205 ( .B(n713), .A(n2370), .Z(n2259) );
  AND U3206 ( .A(n2254), .B(n746), .Z(n2371) );
  NAND U3207 ( .A(n2372), .B(n2373), .Z(n2257) );
  NANDN U3208 ( .B(n2374), .A(n2375), .Z(n2372) );
  XNOR U3209 ( .A(n2379), .B(n2380), .Z(n659) );
  AND U3210 ( .A(n671), .B(n2382), .Z(n2381) );
  XOR U3211 ( .A(n2377), .B(n2380), .Z(n2382) );
  XNOR U3212 ( .A(n2376), .B(n2380), .Z(n2377) );
  XNOR U3213 ( .A(n2301), .B(n2300), .Z(n2380) );
  XNOR U3214 ( .A(n2383), .B(n2305), .Z(n2300) );
  XNOR U3215 ( .A(n2384), .B(n2279), .Z(n2274) );
  XNOR U3216 ( .A(n2271), .B(n2272), .Z(n2279) );
  NAND U3217 ( .A(n855), .B(n1952), .Z(n2272) );
  XNOR U3218 ( .A(n2270), .B(n2385), .Z(n2271) );
  AND U3219 ( .A(n2053), .B(n818), .Z(n2385) );
  XNOR U3220 ( .A(n2278), .B(n2273), .Z(n2384) );
  XNOR U3221 ( .A(n2283), .B(n2393), .Z(n2284) );
  AND U3222 ( .A(n2282), .B(n744), .Z(n2393) );
  XOR U3223 ( .A(n2397), .B(n2285), .Z(n2392) );
  NAND U3224 ( .A(n778), .B(n2166), .Z(n2285) );
  IV U3225 ( .A(n2277), .Z(n2397) );
  XNOR U3226 ( .A(n2288), .B(n2402), .Z(n2289) );
  AND U3227 ( .A(n1858), .B(n899), .Z(n2402) );
  XOR U3228 ( .A(n2406), .B(n2290), .Z(n2401) );
  NAND U3229 ( .A(n945), .B(n1757), .Z(n2290) );
  IV U3230 ( .A(n2292), .Z(n2406) );
  XNOR U3231 ( .A(n2297), .B(n2298), .Z(n2294) );
  NAND U3232 ( .A(n1057), .B(n1570), .Z(n2298) );
  XNOR U3233 ( .A(n2296), .B(n2410), .Z(n2297) );
  AND U3234 ( .A(n1664), .B(n1003), .Z(n2410) );
  XNOR U3235 ( .A(n2304), .B(n2299), .Z(n2383) );
  AND U3236 ( .A(n2307), .B(n2418), .Z(n2417) );
  AND U3237 ( .A(n2419), .B(n2420), .Z(n2418) );
  NANDN U3238 ( .B(n714), .A(n2421), .Z(n2420) );
  NANDN U3239 ( .B(n2422), .A(n2423), .Z(n2419) );
  ANDN U3240 ( .A(n2309), .B(n2308), .Z(n2307) );
  NOR U3241 ( .A(n2424), .B(n2425), .Z(n2308) );
  NANDN U3242 ( .B(n2426), .A(n2427), .Z(n2309) );
  XNOR U3243 ( .A(n2431), .B(n2334), .Z(n2325) );
  XNOR U3244 ( .A(n2313), .B(n2433), .Z(n2314) );
  AND U3245 ( .A(n1388), .B(n1198), .Z(n2433) );
  XOR U3246 ( .A(n2437), .B(n2315), .Z(n2432) );
  NAND U3247 ( .A(n1140), .B(n1465), .Z(n2315) );
  IV U3248 ( .A(n2317), .Z(n2437) );
  XNOR U3249 ( .A(n2322), .B(n2323), .Z(n2319) );
  NANDN U3250 ( .B(n1022), .A(n1642), .Z(n2323) );
  XNOR U3251 ( .A(n2321), .B(n2441), .Z(n2322) );
  AND U3252 ( .A(n1550), .B(n1082), .Z(n2441) );
  XNOR U3253 ( .A(n2333), .B(n2324), .Z(n2431) );
  XOR U3254 ( .A(n2448), .B(n2343), .Z(n2333) );
  XNOR U3255 ( .A(n2330), .B(n2331), .Z(n2343) );
  NAND U3256 ( .A(n1284), .B(n1316), .Z(n2331) );
  XNOR U3257 ( .A(n2329), .B(n2449), .Z(n2330) );
  AND U3258 ( .A(n1246), .B(n1352), .Z(n2449) );
  XNOR U3259 ( .A(n2342), .B(n2332), .Z(n2448) );
  XNOR U3260 ( .A(n2337), .B(n2457), .Z(n2338) );
  AND U3261 ( .A(n1119), .B(n1520), .Z(n2457) );
  XOR U3262 ( .A(n2461), .B(n2339), .Z(n2456) );
  NAND U3263 ( .A(n1433), .B(n1180), .Z(n2339) );
  IV U3264 ( .A(n2341), .Z(n2461) );
  XNOR U3265 ( .A(n2465), .B(n2360), .Z(n2350) );
  XNOR U3266 ( .A(n2347), .B(n2348), .Z(n2360) );
  NANDN U3267 ( .B(n836), .A(n2036), .Z(n2348) );
  XNOR U3268 ( .A(n2346), .B(n2466), .Z(n2347) );
  AND U3269 ( .A(n1931), .B(n874), .Z(n2466) );
  XNOR U3270 ( .A(n2359), .B(n2349), .Z(n2465) );
  XNOR U3271 ( .A(n2354), .B(n2474), .Z(n2355) );
  AND U3272 ( .A(n1737), .B(n986), .Z(n2474) );
  XOR U3273 ( .A(n2478), .B(n2356), .Z(n2473) );
  NAND U3274 ( .A(n932), .B(n1831), .Z(n2356) );
  IV U3275 ( .A(n2358), .Z(n2478) );
  XNOR U3276 ( .A(n2363), .B(n2483), .Z(n2364) );
  AND U3277 ( .A(n2141), .B(n810), .Z(n2483) );
  XOR U3278 ( .A(n2487), .B(n2365), .Z(n2482) );
  NAND U3279 ( .A(n774), .B(n2254), .Z(n2365) );
  IV U3280 ( .A(n2367), .Z(n2487) );
  XNOR U3281 ( .A(n2374), .B(n2375), .Z(n2369) );
  NANDN U3282 ( .B(n713), .A(n2491), .Z(n2375) );
  XNOR U3283 ( .A(n2373), .B(n2492), .Z(n2374) );
  AND U3284 ( .A(n2370), .B(n746), .Z(n2492) );
  ANDN U3285 ( .A(n2493), .B(n2494), .Z(n2373) );
  NANDN U3286 ( .B(n2495), .A(n2496), .Z(n2493) );
  XNOR U3287 ( .A(n2500), .B(n2501), .Z(n660) );
  AND U3288 ( .A(n671), .B(n2503), .Z(n2502) );
  XOR U3289 ( .A(n2498), .B(n2501), .Z(n2503) );
  XNOR U3290 ( .A(n2497), .B(n2501), .Z(n2498) );
  XNOR U3291 ( .A(n2416), .B(n2415), .Z(n2501) );
  XNOR U3292 ( .A(n2504), .B(n2430), .Z(n2415) );
  XNOR U3293 ( .A(n2505), .B(n2400), .Z(n2390) );
  XNOR U3294 ( .A(n2387), .B(n2388), .Z(n2400) );
  NAND U3295 ( .A(n899), .B(n1952), .Z(n2388) );
  XNOR U3296 ( .A(n2386), .B(n2506), .Z(n2387) );
  AND U3297 ( .A(n2053), .B(n855), .Z(n2506) );
  XNOR U3298 ( .A(n2399), .B(n2389), .Z(n2505) );
  XNOR U3299 ( .A(n2394), .B(n2514), .Z(n2395) );
  AND U3300 ( .A(n2282), .B(n778), .Z(n2514) );
  XOR U3301 ( .A(n2518), .B(n2396), .Z(n2513) );
  NAND U3302 ( .A(n818), .B(n2166), .Z(n2396) );
  IV U3303 ( .A(n2398), .Z(n2518) );
  XNOR U3304 ( .A(n2403), .B(n2523), .Z(n2404) );
  AND U3305 ( .A(n1858), .B(n945), .Z(n2523) );
  XOR U3306 ( .A(n2527), .B(n2405), .Z(n2522) );
  NAND U3307 ( .A(n1003), .B(n1757), .Z(n2405) );
  IV U3308 ( .A(n2407), .Z(n2527) );
  XNOR U3309 ( .A(n2412), .B(n2413), .Z(n2409) );
  NAND U3310 ( .A(n1119), .B(n1570), .Z(n2413) );
  XNOR U3311 ( .A(n2411), .B(n2531), .Z(n2412) );
  AND U3312 ( .A(n1664), .B(n1057), .Z(n2531) );
  XNOR U3313 ( .A(n2429), .B(n2414), .Z(n2504) );
  XOR U3314 ( .A(n2538), .B(n2423), .Z(n2429) );
  XNOR U3315 ( .A(n2426), .B(n2427), .Z(n2423) );
  XOR U3316 ( .A(n2542), .B(n2425), .Z(n2426) );
  NAND U3317 ( .A(n744), .B(n2421), .Z(n2425) );
  NANDN U3318 ( .B(n714), .A(n2544), .Z(n2543) );
  OR U3319 ( .A(n2548), .B(n2549), .Z(n2422) );
  XNOR U3320 ( .A(n2553), .B(n2455), .Z(n2446) );
  XNOR U3321 ( .A(n2434), .B(n2555), .Z(n2435) );
  AND U3322 ( .A(n1465), .B(n1198), .Z(n2555) );
  XOR U3323 ( .A(n2559), .B(n2436), .Z(n2554) );
  NAND U3324 ( .A(n1140), .B(n1550), .Z(n2436) );
  IV U3325 ( .A(n2438), .Z(n2559) );
  XNOR U3326 ( .A(n2443), .B(n2444), .Z(n2440) );
  NANDN U3327 ( .B(n1022), .A(n1737), .Z(n2444) );
  XNOR U3328 ( .A(n2442), .B(n2563), .Z(n2443) );
  AND U3329 ( .A(n1642), .B(n1082), .Z(n2563) );
  XNOR U3330 ( .A(n2454), .B(n2445), .Z(n2553) );
  XOR U3331 ( .A(n2570), .B(n2464), .Z(n2454) );
  XNOR U3332 ( .A(n2451), .B(n2452), .Z(n2464) );
  NAND U3333 ( .A(n1284), .B(n1388), .Z(n2452) );
  XNOR U3334 ( .A(n2450), .B(n2571), .Z(n2451) );
  AND U3335 ( .A(n1316), .B(n1352), .Z(n2571) );
  XNOR U3336 ( .A(n2463), .B(n2453), .Z(n2570) );
  XNOR U3337 ( .A(n2458), .B(n2579), .Z(n2459) );
  AND U3338 ( .A(n1180), .B(n1520), .Z(n2579) );
  XOR U3339 ( .A(n2583), .B(n2460), .Z(n2578) );
  NAND U3340 ( .A(n1433), .B(n1246), .Z(n2460) );
  IV U3341 ( .A(n2462), .Z(n2583) );
  XNOR U3342 ( .A(n2587), .B(n2481), .Z(n2471) );
  XNOR U3343 ( .A(n2468), .B(n2469), .Z(n2481) );
  NANDN U3344 ( .B(n836), .A(n2141), .Z(n2469) );
  XNOR U3345 ( .A(n2467), .B(n2588), .Z(n2468) );
  AND U3346 ( .A(n2036), .B(n874), .Z(n2588) );
  XNOR U3347 ( .A(n2480), .B(n2470), .Z(n2587) );
  XNOR U3348 ( .A(n2475), .B(n2596), .Z(n2476) );
  AND U3349 ( .A(n1831), .B(n986), .Z(n2596) );
  XOR U3350 ( .A(n2600), .B(n2477), .Z(n2595) );
  NAND U3351 ( .A(n932), .B(n1931), .Z(n2477) );
  IV U3352 ( .A(n2479), .Z(n2600) );
  XNOR U3353 ( .A(n2484), .B(n2605), .Z(n2485) );
  AND U3354 ( .A(n2254), .B(n810), .Z(n2605) );
  XOR U3355 ( .A(n2609), .B(n2486), .Z(n2604) );
  NAND U3356 ( .A(n774), .B(n2370), .Z(n2486) );
  IV U3357 ( .A(n2488), .Z(n2609) );
  XNOR U3358 ( .A(n2495), .B(n2496), .Z(n2490) );
  NANDN U3359 ( .B(n713), .A(n2613), .Z(n2496) );
  AND U3360 ( .A(n2491), .B(n746), .Z(n2614) );
  NAND U3361 ( .A(n2615), .B(n2616), .Z(n2494) );
  NANDN U3362 ( .B(n2617), .A(n2618), .Z(n2615) );
  XOR U3363 ( .A(n2622), .B(n2623), .Z(n661) );
  AND U3364 ( .A(n671), .B(n2625), .Z(n2624) );
  XNOR U3365 ( .A(n2620), .B(n2623), .Z(n2625) );
  XNOR U3366 ( .A(n2623), .B(n2619), .Z(n2620) );
  OR U3367 ( .A(n2626), .B(n2627), .Z(n2619) );
  XNOR U3368 ( .A(n2537), .B(n2536), .Z(n2623) );
  XNOR U3369 ( .A(n2628), .B(n2552), .Z(n2536) );
  XNOR U3370 ( .A(n2629), .B(n2521), .Z(n2511) );
  XNOR U3371 ( .A(n2508), .B(n2509), .Z(n2521) );
  NAND U3372 ( .A(n945), .B(n1952), .Z(n2509) );
  XNOR U3373 ( .A(n2507), .B(n2630), .Z(n2508) );
  AND U3374 ( .A(n2053), .B(n899), .Z(n2630) );
  XNOR U3375 ( .A(n2520), .B(n2510), .Z(n2629) );
  XNOR U3376 ( .A(n2515), .B(n2638), .Z(n2516) );
  AND U3377 ( .A(n2282), .B(n818), .Z(n2638) );
  XOR U3378 ( .A(n2642), .B(n2517), .Z(n2637) );
  NAND U3379 ( .A(n855), .B(n2166), .Z(n2517) );
  IV U3380 ( .A(n2519), .Z(n2642) );
  XNOR U3381 ( .A(n2524), .B(n2647), .Z(n2525) );
  AND U3382 ( .A(n1858), .B(n1003), .Z(n2647) );
  XOR U3383 ( .A(n2651), .B(n2526), .Z(n2646) );
  NAND U3384 ( .A(n1057), .B(n1757), .Z(n2526) );
  IV U3385 ( .A(n2528), .Z(n2651) );
  XNOR U3386 ( .A(n2533), .B(n2534), .Z(n2530) );
  NAND U3387 ( .A(n1180), .B(n1570), .Z(n2534) );
  XNOR U3388 ( .A(n2532), .B(n2655), .Z(n2533) );
  AND U3389 ( .A(n1664), .B(n1119), .Z(n2655) );
  XNOR U3390 ( .A(n2551), .B(n2535), .Z(n2628) );
  XNOR U3391 ( .A(n2662), .B(n2548), .Z(n2551) );
  XOR U3392 ( .A(n2541), .B(n2540), .Z(n2548) );
  XOR U3393 ( .A(n2539), .B(n2663), .Z(n2540) );
  AND U3394 ( .A(n2664), .B(n2665), .Z(n2663) );
  NANDN U3395 ( .B(n714), .A(n2666), .Z(n2665) );
  OR U3396 ( .A(n2667), .B(n2668), .Z(n2664) );
  NAND U3397 ( .A(n778), .B(n2421), .Z(n2547) );
  XNOR U3398 ( .A(n2545), .B(n2672), .Z(n2546) );
  AND U3399 ( .A(n2544), .B(n744), .Z(n2672) );
  NANDN U3400 ( .B(n2676), .A(n2677), .Z(n2549) );
  XNOR U3401 ( .A(n2681), .B(n2577), .Z(n2568) );
  XNOR U3402 ( .A(n2556), .B(n2683), .Z(n2557) );
  AND U3403 ( .A(n1550), .B(n1198), .Z(n2683) );
  XOR U3404 ( .A(n2687), .B(n2558), .Z(n2682) );
  NAND U3405 ( .A(n1140), .B(n1642), .Z(n2558) );
  IV U3406 ( .A(n2560), .Z(n2687) );
  XNOR U3407 ( .A(n2565), .B(n2566), .Z(n2562) );
  NANDN U3408 ( .B(n1022), .A(n1831), .Z(n2566) );
  XNOR U3409 ( .A(n2564), .B(n2691), .Z(n2565) );
  AND U3410 ( .A(n1737), .B(n1082), .Z(n2691) );
  XNOR U3411 ( .A(n2576), .B(n2567), .Z(n2681) );
  XOR U3412 ( .A(n2698), .B(n2586), .Z(n2576) );
  XNOR U3413 ( .A(n2573), .B(n2574), .Z(n2586) );
  NAND U3414 ( .A(n1284), .B(n1465), .Z(n2574) );
  XNOR U3415 ( .A(n2572), .B(n2699), .Z(n2573) );
  AND U3416 ( .A(n1388), .B(n1352), .Z(n2699) );
  XNOR U3417 ( .A(n2585), .B(n2575), .Z(n2698) );
  XNOR U3418 ( .A(n2580), .B(n2707), .Z(n2581) );
  AND U3419 ( .A(n1246), .B(n1520), .Z(n2707) );
  XOR U3420 ( .A(n2711), .B(n2582), .Z(n2706) );
  NAND U3421 ( .A(n1433), .B(n1316), .Z(n2582) );
  IV U3422 ( .A(n2584), .Z(n2711) );
  XNOR U3423 ( .A(n2715), .B(n2603), .Z(n2593) );
  XNOR U3424 ( .A(n2590), .B(n2591), .Z(n2603) );
  NANDN U3425 ( .B(n836), .A(n2254), .Z(n2591) );
  XNOR U3426 ( .A(n2589), .B(n2716), .Z(n2590) );
  AND U3427 ( .A(n2141), .B(n874), .Z(n2716) );
  XNOR U3428 ( .A(n2602), .B(n2592), .Z(n2715) );
  XNOR U3429 ( .A(n2597), .B(n2724), .Z(n2598) );
  AND U3430 ( .A(n1931), .B(n986), .Z(n2724) );
  XOR U3431 ( .A(n2728), .B(n2599), .Z(n2723) );
  NAND U3432 ( .A(n932), .B(n2036), .Z(n2599) );
  IV U3433 ( .A(n2601), .Z(n2728) );
  XNOR U3434 ( .A(n2606), .B(n2733), .Z(n2607) );
  AND U3435 ( .A(n2370), .B(n810), .Z(n2733) );
  XOR U3436 ( .A(n2737), .B(n2608), .Z(n2732) );
  NAND U3437 ( .A(n774), .B(n2491), .Z(n2608) );
  IV U3438 ( .A(n2610), .Z(n2737) );
  XNOR U3439 ( .A(n2617), .B(n2618), .Z(n2612) );
  NANDN U3440 ( .B(n713), .A(n2741), .Z(n2618) );
  XNOR U3441 ( .A(n2616), .B(n2742), .Z(n2617) );
  AND U3442 ( .A(n2613), .B(n746), .Z(n2742) );
  ANDN U3443 ( .A(n2743), .B(n2744), .Z(n2616) );
  NANDN U3444 ( .B(n2745), .A(n2746), .Z(n2743) );
  XNOR U3445 ( .A(n2748), .B(n2749), .Z(n699) );
  AND U3446 ( .A(n671), .B(n2751), .Z(n2750) );
  XOR U3447 ( .A(n2626), .B(n2752), .Z(n2751) );
  XOR U3448 ( .A(n2752), .B(n2627), .Z(n2626) );
  OR U3449 ( .A(n2753), .B(n2754), .Z(n2627) );
  IV U3450 ( .A(n2749), .Z(n2752) );
  XOR U3451 ( .A(n2661), .B(n2660), .Z(n2749) );
  XNOR U3452 ( .A(n2755), .B(n2680), .Z(n2660) );
  XNOR U3453 ( .A(n2756), .B(n2645), .Z(n2635) );
  XNOR U3454 ( .A(n2632), .B(n2633), .Z(n2645) );
  NAND U3455 ( .A(n1003), .B(n1952), .Z(n2633) );
  XNOR U3456 ( .A(n2631), .B(n2757), .Z(n2632) );
  AND U3457 ( .A(n2053), .B(n945), .Z(n2757) );
  XNOR U3458 ( .A(n2644), .B(n2634), .Z(n2756) );
  XNOR U3459 ( .A(n2639), .B(n2765), .Z(n2640) );
  AND U3460 ( .A(n2282), .B(n855), .Z(n2765) );
  XOR U3461 ( .A(n2769), .B(n2641), .Z(n2764) );
  NAND U3462 ( .A(n899), .B(n2166), .Z(n2641) );
  IV U3463 ( .A(n2643), .Z(n2769) );
  XNOR U3464 ( .A(n2648), .B(n2774), .Z(n2649) );
  AND U3465 ( .A(n1858), .B(n1057), .Z(n2774) );
  XOR U3466 ( .A(n2778), .B(n2650), .Z(n2773) );
  NAND U3467 ( .A(n1119), .B(n1757), .Z(n2650) );
  IV U3468 ( .A(n2652), .Z(n2778) );
  XNOR U3469 ( .A(n2657), .B(n2658), .Z(n2654) );
  NAND U3470 ( .A(n1246), .B(n1570), .Z(n2658) );
  XNOR U3471 ( .A(n2656), .B(n2782), .Z(n2657) );
  AND U3472 ( .A(n1664), .B(n1180), .Z(n2782) );
  XNOR U3473 ( .A(n2679), .B(n2659), .Z(n2755) );
  XNOR U3474 ( .A(n2789), .B(n2676), .Z(n2679) );
  XOR U3475 ( .A(n2671), .B(n2670), .Z(n2676) );
  XNOR U3476 ( .A(n2794), .B(n2667), .Z(n2790) );
  NAND U3477 ( .A(n744), .B(n2666), .Z(n2667) );
  NANDN U3478 ( .B(n714), .A(n2796), .Z(n2795) );
  NAND U3479 ( .A(n818), .B(n2421), .Z(n2675) );
  XNOR U3480 ( .A(n2673), .B(n2800), .Z(n2674) );
  AND U3481 ( .A(n2544), .B(n778), .Z(n2800) );
  XNOR U3482 ( .A(n2677), .B(n2678), .Z(n2789) );
  XNOR U3483 ( .A(n2810), .B(n2705), .Z(n2696) );
  XNOR U3484 ( .A(n2684), .B(n2812), .Z(n2685) );
  AND U3485 ( .A(n1642), .B(n1198), .Z(n2812) );
  XOR U3486 ( .A(n2816), .B(n2686), .Z(n2811) );
  NAND U3487 ( .A(n1140), .B(n1737), .Z(n2686) );
  IV U3488 ( .A(n2688), .Z(n2816) );
  XNOR U3489 ( .A(n2693), .B(n2694), .Z(n2690) );
  NANDN U3490 ( .B(n1022), .A(n1931), .Z(n2694) );
  XNOR U3491 ( .A(n2692), .B(n2820), .Z(n2693) );
  AND U3492 ( .A(n1831), .B(n1082), .Z(n2820) );
  XNOR U3493 ( .A(n2704), .B(n2695), .Z(n2810) );
  XOR U3494 ( .A(n2827), .B(n2714), .Z(n2704) );
  XNOR U3495 ( .A(n2701), .B(n2702), .Z(n2714) );
  NAND U3496 ( .A(n1284), .B(n1550), .Z(n2702) );
  XNOR U3497 ( .A(n2700), .B(n2828), .Z(n2701) );
  AND U3498 ( .A(n1465), .B(n1352), .Z(n2828) );
  XNOR U3499 ( .A(n2713), .B(n2703), .Z(n2827) );
  XNOR U3500 ( .A(n2708), .B(n2836), .Z(n2709) );
  AND U3501 ( .A(n1316), .B(n1520), .Z(n2836) );
  XOR U3502 ( .A(n2840), .B(n2710), .Z(n2835) );
  NAND U3503 ( .A(n1433), .B(n1388), .Z(n2710) );
  IV U3504 ( .A(n2712), .Z(n2840) );
  XNOR U3505 ( .A(n2844), .B(n2731), .Z(n2721) );
  XNOR U3506 ( .A(n2718), .B(n2719), .Z(n2731) );
  NANDN U3507 ( .B(n836), .A(n2370), .Z(n2719) );
  XNOR U3508 ( .A(n2717), .B(n2845), .Z(n2718) );
  AND U3509 ( .A(n2254), .B(n874), .Z(n2845) );
  XNOR U3510 ( .A(n2730), .B(n2720), .Z(n2844) );
  XNOR U3511 ( .A(n2725), .B(n2853), .Z(n2726) );
  AND U3512 ( .A(n2036), .B(n986), .Z(n2853) );
  XOR U3513 ( .A(n2857), .B(n2727), .Z(n2852) );
  NAND U3514 ( .A(n932), .B(n2141), .Z(n2727) );
  IV U3515 ( .A(n2729), .Z(n2857) );
  XNOR U3516 ( .A(n2734), .B(n2862), .Z(n2735) );
  AND U3517 ( .A(n2491), .B(n810), .Z(n2862) );
  XOR U3518 ( .A(n2866), .B(n2736), .Z(n2861) );
  NAND U3519 ( .A(n774), .B(n2613), .Z(n2736) );
  IV U3520 ( .A(n2738), .Z(n2866) );
  XNOR U3521 ( .A(n2745), .B(n2746), .Z(n2740) );
  OR U3522 ( .A(n2870), .B(n713), .Z(n2746) );
  AND U3523 ( .A(n2741), .B(n746), .Z(n2871) );
  NAND U3524 ( .A(n2872), .B(n2873), .Z(n2744) );
  NANDN U3525 ( .B(n2874), .A(n2875), .Z(n2872) );
  XNOR U3526 ( .A(n2877), .B(n2878), .Z(n1128) );
  XOR U3527 ( .A(n2876), .B(n2879), .Z(n2877) );
  AND U3528 ( .A(n671), .B(n2880), .Z(n2879) );
  XOR U3529 ( .A(n2753), .B(n2881), .Z(n2880) );
  XOR U3530 ( .A(n2881), .B(n2754), .Z(n2753) );
  NANDN U3531 ( .B(n2882), .A(n2883), .Z(n2754) );
  IV U3532 ( .A(n2878), .Z(n2881) );
  XOR U3533 ( .A(n2788), .B(n2787), .Z(n2878) );
  XNOR U3534 ( .A(n2884), .B(n2806), .Z(n2787) );
  XNOR U3535 ( .A(n2885), .B(n2772), .Z(n2762) );
  XNOR U3536 ( .A(n2759), .B(n2760), .Z(n2772) );
  NAND U3537 ( .A(n1057), .B(n1952), .Z(n2760) );
  XNOR U3538 ( .A(n2758), .B(n2886), .Z(n2759) );
  AND U3539 ( .A(n2053), .B(n1003), .Z(n2886) );
  XNOR U3540 ( .A(n2771), .B(n2761), .Z(n2885) );
  XNOR U3541 ( .A(n2766), .B(n2894), .Z(n2767) );
  AND U3542 ( .A(n2282), .B(n899), .Z(n2894) );
  XOR U3543 ( .A(n2898), .B(n2768), .Z(n2893) );
  NAND U3544 ( .A(n945), .B(n2166), .Z(n2768) );
  IV U3545 ( .A(n2770), .Z(n2898) );
  XNOR U3546 ( .A(n2775), .B(n2903), .Z(n2776) );
  AND U3547 ( .A(n1858), .B(n1119), .Z(n2903) );
  XOR U3548 ( .A(n2907), .B(n2777), .Z(n2902) );
  NAND U3549 ( .A(n1180), .B(n1757), .Z(n2777) );
  IV U3550 ( .A(n2779), .Z(n2907) );
  XNOR U3551 ( .A(n2784), .B(n2785), .Z(n2781) );
  NAND U3552 ( .A(n1316), .B(n1570), .Z(n2785) );
  XNOR U3553 ( .A(n2783), .B(n2911), .Z(n2784) );
  AND U3554 ( .A(n1664), .B(n1246), .Z(n2911) );
  XNOR U3555 ( .A(n2805), .B(n2786), .Z(n2884) );
  XOR U3556 ( .A(n2918), .B(n2809), .Z(n2805) );
  XNOR U3557 ( .A(n2797), .B(n2920), .Z(n2798) );
  AND U3558 ( .A(n2796), .B(n744), .Z(n2920) );
  XOR U3559 ( .A(n2924), .B(n2799), .Z(n2919) );
  NAND U3560 ( .A(n778), .B(n2666), .Z(n2799) );
  IV U3561 ( .A(n2791), .Z(n2924) );
  XNOR U3562 ( .A(n2802), .B(n2803), .Z(n2793) );
  NAND U3563 ( .A(n855), .B(n2421), .Z(n2803) );
  XNOR U3564 ( .A(n2801), .B(n2928), .Z(n2802) );
  AND U3565 ( .A(n2544), .B(n818), .Z(n2928) );
  XNOR U3566 ( .A(n2808), .B(n2804), .Z(n2918) );
  AND U3567 ( .A(n2936), .B(n2937), .Z(n2935) );
  OR U3568 ( .A(n2938), .B(n2939), .Z(n2937) );
  AND U3569 ( .A(n2940), .B(n2941), .Z(n2936) );
  NANDN U3570 ( .B(n714), .A(n2942), .Z(n2941) );
  NANDN U3571 ( .B(n2943), .A(n2944), .Z(n2940) );
  XNOR U3572 ( .A(n2948), .B(n2834), .Z(n2825) );
  XNOR U3573 ( .A(n2813), .B(n2950), .Z(n2814) );
  AND U3574 ( .A(n1737), .B(n1198), .Z(n2950) );
  XOR U3575 ( .A(n2954), .B(n2815), .Z(n2949) );
  NAND U3576 ( .A(n1140), .B(n1831), .Z(n2815) );
  IV U3577 ( .A(n2817), .Z(n2954) );
  XNOR U3578 ( .A(n2822), .B(n2823), .Z(n2819) );
  NANDN U3579 ( .B(n1022), .A(n2036), .Z(n2823) );
  XNOR U3580 ( .A(n2821), .B(n2958), .Z(n2822) );
  AND U3581 ( .A(n1931), .B(n1082), .Z(n2958) );
  XNOR U3582 ( .A(n2833), .B(n2824), .Z(n2948) );
  XOR U3583 ( .A(n2965), .B(n2843), .Z(n2833) );
  XNOR U3584 ( .A(n2830), .B(n2831), .Z(n2843) );
  NAND U3585 ( .A(n1284), .B(n1642), .Z(n2831) );
  XNOR U3586 ( .A(n2829), .B(n2966), .Z(n2830) );
  AND U3587 ( .A(n1550), .B(n1352), .Z(n2966) );
  XNOR U3588 ( .A(n2842), .B(n2832), .Z(n2965) );
  XNOR U3589 ( .A(n2837), .B(n2974), .Z(n2838) );
  AND U3590 ( .A(n1388), .B(n1520), .Z(n2974) );
  XOR U3591 ( .A(n2978), .B(n2839), .Z(n2973) );
  NAND U3592 ( .A(n1433), .B(n1465), .Z(n2839) );
  IV U3593 ( .A(n2841), .Z(n2978) );
  XNOR U3594 ( .A(n2982), .B(n2860), .Z(n2850) );
  XNOR U3595 ( .A(n2847), .B(n2848), .Z(n2860) );
  NANDN U3596 ( .B(n836), .A(n2491), .Z(n2848) );
  XNOR U3597 ( .A(n2846), .B(n2983), .Z(n2847) );
  AND U3598 ( .A(n2370), .B(n874), .Z(n2983) );
  XNOR U3599 ( .A(n2859), .B(n2849), .Z(n2982) );
  XNOR U3600 ( .A(n2854), .B(n2991), .Z(n2855) );
  AND U3601 ( .A(n2141), .B(n986), .Z(n2991) );
  XOR U3602 ( .A(n2995), .B(n2856), .Z(n2990) );
  NAND U3603 ( .A(n932), .B(n2254), .Z(n2856) );
  IV U3604 ( .A(n2858), .Z(n2995) );
  XNOR U3605 ( .A(n2863), .B(n3000), .Z(n2864) );
  AND U3606 ( .A(n2613), .B(n810), .Z(n3000) );
  XOR U3607 ( .A(n3004), .B(n2865), .Z(n2999) );
  NAND U3608 ( .A(n774), .B(n2741), .Z(n2865) );
  IV U3609 ( .A(n2867), .Z(n3004) );
  XNOR U3610 ( .A(n2874), .B(n2875), .Z(n2869) );
  OR U3611 ( .A(n3008), .B(n713), .Z(n2875) );
  XNOR U3612 ( .A(n2873), .B(n3009), .Z(n2874) );
  ANDN U3613 ( .A(n746), .B(n2870), .Z(n3009) );
  ANDN U3614 ( .A(n3010), .B(n3011), .Z(n2873) );
  NANDN U3615 ( .B(n3012), .A(n3013), .Z(n3010) );
  XOR U3616 ( .A(n3015), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U3617 ( .A(n3016), .B(n3017), .Z(n3015) );
  XNOR U3618 ( .A(n3018), .B(n3014), .Z(n3016) );
  NANDN U3619 ( .B(n2883), .A(\_MxM/Y0[0] ), .Z(n3014) );
  NAND U3620 ( .A(n3019), .B(n671), .Z(n3018) );
  XOR U3621 ( .A(e_input[31]), .B(g_input[31]), .Z(n671) );
  XNOR U3622 ( .A(n2882), .B(n3017), .Z(n3019) );
  XOR U3623 ( .A(n2883), .B(n3017), .Z(n2882) );
  XOR U3624 ( .A(n2917), .B(n2916), .Z(n3017) );
  XNOR U3625 ( .A(n3020), .B(n2934), .Z(n2916) );
  XNOR U3626 ( .A(n3021), .B(n2901), .Z(n2891) );
  XNOR U3627 ( .A(n2888), .B(n2889), .Z(n2901) );
  NAND U3628 ( .A(n1119), .B(n1952), .Z(n2889) );
  XNOR U3629 ( .A(n2887), .B(n3022), .Z(n2888) );
  AND U3630 ( .A(n2053), .B(n1057), .Z(n3022) );
  XNOR U3631 ( .A(n2900), .B(n2890), .Z(n3021) );
  XNOR U3632 ( .A(n2895), .B(n3030), .Z(n2896) );
  AND U3633 ( .A(n2282), .B(n945), .Z(n3030) );
  XOR U3634 ( .A(n3034), .B(n2897), .Z(n3029) );
  NAND U3635 ( .A(n1003), .B(n2166), .Z(n2897) );
  IV U3636 ( .A(n2899), .Z(n3034) );
  XNOR U3637 ( .A(n2904), .B(n3039), .Z(n2905) );
  AND U3638 ( .A(n1858), .B(n1180), .Z(n3039) );
  XOR U3639 ( .A(n3043), .B(n2906), .Z(n3038) );
  NAND U3640 ( .A(n1246), .B(n1757), .Z(n2906) );
  IV U3641 ( .A(n2908), .Z(n3043) );
  XNOR U3642 ( .A(n2913), .B(n2914), .Z(n2910) );
  NAND U3643 ( .A(n1388), .B(n1570), .Z(n2914) );
  XNOR U3644 ( .A(n2912), .B(n3047), .Z(n2913) );
  AND U3645 ( .A(n1664), .B(n1316), .Z(n3047) );
  XNOR U3646 ( .A(n2933), .B(n2915), .Z(n3020) );
  XOR U3647 ( .A(n3054), .B(n2947), .Z(n2933) );
  XNOR U3648 ( .A(n2921), .B(n3056), .Z(n2922) );
  AND U3649 ( .A(n2796), .B(n778), .Z(n3056) );
  XOR U3650 ( .A(n3060), .B(n2923), .Z(n3055) );
  NAND U3651 ( .A(n818), .B(n2666), .Z(n2923) );
  IV U3652 ( .A(n2925), .Z(n3060) );
  XNOR U3653 ( .A(n2930), .B(n2931), .Z(n2927) );
  NAND U3654 ( .A(n899), .B(n2421), .Z(n2931) );
  XNOR U3655 ( .A(n2929), .B(n3064), .Z(n2930) );
  AND U3656 ( .A(n2544), .B(n855), .Z(n3064) );
  XNOR U3657 ( .A(n2946), .B(n2932), .Z(n3054) );
  XNOR U3658 ( .A(n3071), .B(n2943), .Z(n2946) );
  XOR U3659 ( .A(n3072), .B(n2938), .Z(n2943) );
  NAND U3660 ( .A(n744), .B(n2942), .Z(n2938) );
  NANDN U3661 ( .B(n714), .A(n3074), .Z(n3073) );
  XNOR U3662 ( .A(n2944), .B(n2945), .Z(n3071) );
  XNOR U3663 ( .A(n3084), .B(n2972), .Z(n2963) );
  XNOR U3664 ( .A(n2951), .B(n3086), .Z(n2952) );
  AND U3665 ( .A(n1831), .B(n1198), .Z(n3086) );
  XOR U3666 ( .A(n3090), .B(n2953), .Z(n3085) );
  NAND U3667 ( .A(n1140), .B(n1931), .Z(n2953) );
  IV U3668 ( .A(n2955), .Z(n3090) );
  XNOR U3669 ( .A(n2960), .B(n2961), .Z(n2957) );
  NANDN U3670 ( .B(n1022), .A(n2141), .Z(n2961) );
  XNOR U3671 ( .A(n2959), .B(n3094), .Z(n2960) );
  AND U3672 ( .A(n2036), .B(n1082), .Z(n3094) );
  XNOR U3673 ( .A(n2971), .B(n2962), .Z(n3084) );
  XOR U3674 ( .A(n3101), .B(n2981), .Z(n2971) );
  XNOR U3675 ( .A(n2968), .B(n2969), .Z(n2981) );
  NAND U3676 ( .A(n1284), .B(n1737), .Z(n2969) );
  XNOR U3677 ( .A(n2967), .B(n3102), .Z(n2968) );
  AND U3678 ( .A(n1642), .B(n1352), .Z(n3102) );
  XNOR U3679 ( .A(n2980), .B(n2970), .Z(n3101) );
  XNOR U3680 ( .A(n2975), .B(n3110), .Z(n2976) );
  AND U3681 ( .A(n1465), .B(n1520), .Z(n3110) );
  XOR U3682 ( .A(n3114), .B(n2977), .Z(n3109) );
  NAND U3683 ( .A(n1433), .B(n1550), .Z(n2977) );
  IV U3684 ( .A(n2979), .Z(n3114) );
  XNOR U3685 ( .A(n3118), .B(n2998), .Z(n2988) );
  XNOR U3686 ( .A(n2985), .B(n2986), .Z(n2998) );
  NANDN U3687 ( .B(n836), .A(n2613), .Z(n2986) );
  XNOR U3688 ( .A(n2984), .B(n3119), .Z(n2985) );
  AND U3689 ( .A(n2491), .B(n874), .Z(n3119) );
  XNOR U3690 ( .A(n2997), .B(n2987), .Z(n3118) );
  XNOR U3691 ( .A(n2992), .B(n3127), .Z(n2993) );
  AND U3692 ( .A(n2254), .B(n986), .Z(n3127) );
  XOR U3693 ( .A(n3131), .B(n2994), .Z(n3126) );
  NAND U3694 ( .A(n932), .B(n2370), .Z(n2994) );
  IV U3695 ( .A(n2996), .Z(n3131) );
  XNOR U3696 ( .A(n3001), .B(n3136), .Z(n3002) );
  AND U3697 ( .A(n2741), .B(n810), .Z(n3136) );
  XOR U3698 ( .A(n3140), .B(n3003), .Z(n3135) );
  NANDN U3699 ( .B(n2870), .A(n774), .Z(n3003) );
  IV U3700 ( .A(n3005), .Z(n3140) );
  XNOR U3701 ( .A(n3012), .B(n3013), .Z(n3007) );
  NANDN U3702 ( .B(n713), .A(n3144), .Z(n3013) );
  ANDN U3703 ( .A(n746), .B(n3008), .Z(n3145) );
  NAND U3704 ( .A(n3146), .B(n3147), .Z(n3011) );
  NANDN U3705 ( .B(n3148), .A(n3149), .Z(n3146) );
  XOR U3706 ( .A(n3053), .B(n3052), .Z(n2883) );
  XNOR U3707 ( .A(n3150), .B(n3070), .Z(n3052) );
  XNOR U3708 ( .A(n3151), .B(n3037), .Z(n3027) );
  XNOR U3709 ( .A(n3024), .B(n3025), .Z(n3037) );
  NAND U3710 ( .A(n1180), .B(n1952), .Z(n3025) );
  XNOR U3711 ( .A(n3023), .B(n3152), .Z(n3024) );
  AND U3712 ( .A(n2053), .B(n1119), .Z(n3152) );
  XNOR U3713 ( .A(n3036), .B(n3026), .Z(n3151) );
  XNOR U3714 ( .A(n3031), .B(n3160), .Z(n3032) );
  AND U3715 ( .A(n2282), .B(n1003), .Z(n3160) );
  XOR U3716 ( .A(n3164), .B(n3033), .Z(n3159) );
  NAND U3717 ( .A(n1057), .B(n2166), .Z(n3033) );
  IV U3718 ( .A(n3035), .Z(n3164) );
  XNOR U3719 ( .A(n3040), .B(n3169), .Z(n3041) );
  AND U3720 ( .A(n1858), .B(n1246), .Z(n3169) );
  XOR U3721 ( .A(n3173), .B(n3042), .Z(n3168) );
  NAND U3722 ( .A(n1316), .B(n1757), .Z(n3042) );
  IV U3723 ( .A(n3044), .Z(n3173) );
  XNOR U3724 ( .A(n3049), .B(n3050), .Z(n3046) );
  NAND U3725 ( .A(n1465), .B(n1570), .Z(n3050) );
  XNOR U3726 ( .A(n3048), .B(n3177), .Z(n3049) );
  AND U3727 ( .A(n1664), .B(n1388), .Z(n3177) );
  XNOR U3728 ( .A(n3069), .B(n3051), .Z(n3150) );
  XOR U3729 ( .A(n3181), .B(n3182), .Z(n3051) );
  XOR U3730 ( .A(n3183), .B(n3080), .Z(n3069) );
  XNOR U3731 ( .A(n3057), .B(n3185), .Z(n3058) );
  AND U3732 ( .A(n2796), .B(n818), .Z(n3185) );
  XOR U3733 ( .A(n3189), .B(n3059), .Z(n3184) );
  NAND U3734 ( .A(n855), .B(n2666), .Z(n3059) );
  IV U3735 ( .A(n3061), .Z(n3189) );
  XNOR U3736 ( .A(n3066), .B(n3067), .Z(n3063) );
  NAND U3737 ( .A(n945), .B(n2421), .Z(n3067) );
  XNOR U3738 ( .A(n3065), .B(n3193), .Z(n3066) );
  AND U3739 ( .A(n2544), .B(n899), .Z(n3193) );
  XNOR U3740 ( .A(n3079), .B(n3068), .Z(n3183) );
  XOR U3741 ( .A(n3197), .B(n3198), .Z(n3068) );
  AND U3742 ( .A(n3199), .B(n3200), .Z(n3198) );
  XNOR U3743 ( .A(n3201), .B(n3202), .Z(n3200) );
  XOR U3744 ( .A(n3203), .B(n3197), .Z(n3201) );
  XOR U3745 ( .A(n3157), .B(n3204), .Z(n3199) );
  XNOR U3746 ( .A(n3197), .B(n3158), .Z(n3204) );
  XNOR U3747 ( .A(n3170), .B(n3206), .Z(n3171) );
  AND U3748 ( .A(n1858), .B(n1316), .Z(n3206) );
  XOR U3749 ( .A(n3210), .B(n3172), .Z(n3205) );
  NAND U3750 ( .A(n1388), .B(n1757), .Z(n3172) );
  IV U3751 ( .A(n3174), .Z(n3210) );
  XNOR U3752 ( .A(n3179), .B(n3180), .Z(n3176) );
  NAND U3753 ( .A(n1570), .B(n1550), .Z(n3180) );
  XNOR U3754 ( .A(n3178), .B(n3214), .Z(n3179) );
  AND U3755 ( .A(n1664), .B(n1465), .Z(n3214) );
  XOR U3756 ( .A(n3218), .B(n3167), .Z(n3157) );
  XNOR U3757 ( .A(n3154), .B(n3155), .Z(n3167) );
  NAND U3758 ( .A(n1246), .B(n1952), .Z(n3155) );
  XNOR U3759 ( .A(n3153), .B(n3219), .Z(n3154) );
  AND U3760 ( .A(n2053), .B(n1180), .Z(n3219) );
  XNOR U3761 ( .A(n3166), .B(n3156), .Z(n3218) );
  XNOR U3762 ( .A(n3161), .B(n3227), .Z(n3162) );
  AND U3763 ( .A(n2282), .B(n1057), .Z(n3227) );
  XOR U3764 ( .A(n3231), .B(n3163), .Z(n3226) );
  NAND U3765 ( .A(n1119), .B(n2166), .Z(n3163) );
  IV U3766 ( .A(n3165), .Z(n3231) );
  XOR U3767 ( .A(n3235), .B(n3236), .Z(n3197) );
  AND U3768 ( .A(n3237), .B(n3238), .Z(n3236) );
  XNOR U3769 ( .A(n3239), .B(n3240), .Z(n3238) );
  XNOR U3770 ( .A(n3235), .B(n3241), .Z(n3240) );
  XOR U3771 ( .A(n3224), .B(n3242), .Z(n3237) );
  XNOR U3772 ( .A(n3235), .B(n3225), .Z(n3242) );
  XNOR U3773 ( .A(n3207), .B(n3244), .Z(n3208) );
  AND U3774 ( .A(n1858), .B(n1388), .Z(n3244) );
  XOR U3775 ( .A(n3248), .B(n3209), .Z(n3243) );
  NAND U3776 ( .A(n1465), .B(n1757), .Z(n3209) );
  IV U3777 ( .A(n3211), .Z(n3248) );
  XNOR U3778 ( .A(n3216), .B(n3217), .Z(n3213) );
  NAND U3779 ( .A(n1570), .B(n1642), .Z(n3217) );
  XNOR U3780 ( .A(n3215), .B(n3252), .Z(n3216) );
  AND U3781 ( .A(n1550), .B(n1664), .Z(n3252) );
  XOR U3782 ( .A(n3256), .B(n3234), .Z(n3224) );
  XNOR U3783 ( .A(n3221), .B(n3222), .Z(n3234) );
  NAND U3784 ( .A(n1316), .B(n1952), .Z(n3222) );
  XNOR U3785 ( .A(n3220), .B(n3257), .Z(n3221) );
  AND U3786 ( .A(n2053), .B(n1246), .Z(n3257) );
  XNOR U3787 ( .A(n3233), .B(n3223), .Z(n3256) );
  XNOR U3788 ( .A(n3228), .B(n3265), .Z(n3229) );
  AND U3789 ( .A(n2282), .B(n1119), .Z(n3265) );
  XOR U3790 ( .A(n3269), .B(n3230), .Z(n3264) );
  NAND U3791 ( .A(n1180), .B(n2166), .Z(n3230) );
  IV U3792 ( .A(n3232), .Z(n3269) );
  XOR U3793 ( .A(n3273), .B(n3274), .Z(n3235) );
  AND U3794 ( .A(n3275), .B(n3276), .Z(n3274) );
  XNOR U3795 ( .A(n3277), .B(n3278), .Z(n3276) );
  XNOR U3796 ( .A(n3273), .B(n3279), .Z(n3278) );
  XOR U3797 ( .A(n3262), .B(n3280), .Z(n3275) );
  XNOR U3798 ( .A(n3273), .B(n3263), .Z(n3280) );
  XNOR U3799 ( .A(n3245), .B(n3282), .Z(n3246) );
  AND U3800 ( .A(n1858), .B(n1465), .Z(n3282) );
  XOR U3801 ( .A(n3286), .B(n3247), .Z(n3281) );
  NAND U3802 ( .A(n1757), .B(n1550), .Z(n3247) );
  IV U3803 ( .A(n3249), .Z(n3286) );
  XNOR U3804 ( .A(n3254), .B(n3255), .Z(n3251) );
  NAND U3805 ( .A(n1570), .B(n1737), .Z(n3255) );
  XNOR U3806 ( .A(n3253), .B(n3290), .Z(n3254) );
  AND U3807 ( .A(n1642), .B(n1664), .Z(n3290) );
  XOR U3808 ( .A(n3294), .B(n3272), .Z(n3262) );
  XNOR U3809 ( .A(n3259), .B(n3260), .Z(n3272) );
  NAND U3810 ( .A(n1388), .B(n1952), .Z(n3260) );
  XNOR U3811 ( .A(n3258), .B(n3295), .Z(n3259) );
  AND U3812 ( .A(n2053), .B(n1316), .Z(n3295) );
  XNOR U3813 ( .A(n3271), .B(n3261), .Z(n3294) );
  XNOR U3814 ( .A(n3266), .B(n3303), .Z(n3267) );
  AND U3815 ( .A(n2282), .B(n1180), .Z(n3303) );
  XOR U3816 ( .A(n3307), .B(n3268), .Z(n3302) );
  NAND U3817 ( .A(n1246), .B(n2166), .Z(n3268) );
  IV U3818 ( .A(n3270), .Z(n3307) );
  XOR U3819 ( .A(n3311), .B(n3312), .Z(n3273) );
  AND U3820 ( .A(n3313), .B(n3314), .Z(n3312) );
  XNOR U3821 ( .A(n3315), .B(n3316), .Z(n3314) );
  XNOR U3822 ( .A(n3311), .B(n3317), .Z(n3316) );
  XOR U3823 ( .A(n3300), .B(n3318), .Z(n3313) );
  XNOR U3824 ( .A(n3311), .B(n3301), .Z(n3318) );
  XNOR U3825 ( .A(n3283), .B(n3320), .Z(n3284) );
  AND U3826 ( .A(n1550), .B(n1858), .Z(n3320) );
  XOR U3827 ( .A(n3324), .B(n3285), .Z(n3319) );
  NAND U3828 ( .A(n1757), .B(n1642), .Z(n3285) );
  IV U3829 ( .A(n3287), .Z(n3324) );
  XNOR U3830 ( .A(n3292), .B(n3293), .Z(n3289) );
  NAND U3831 ( .A(n1570), .B(n1831), .Z(n3293) );
  XNOR U3832 ( .A(n3291), .B(n3328), .Z(n3292) );
  AND U3833 ( .A(n1737), .B(n1664), .Z(n3328) );
  XOR U3834 ( .A(n3332), .B(n3310), .Z(n3300) );
  XNOR U3835 ( .A(n3297), .B(n3298), .Z(n3310) );
  NAND U3836 ( .A(n1465), .B(n1952), .Z(n3298) );
  XNOR U3837 ( .A(n3296), .B(n3333), .Z(n3297) );
  AND U3838 ( .A(n2053), .B(n1388), .Z(n3333) );
  XNOR U3839 ( .A(n3309), .B(n3299), .Z(n3332) );
  XNOR U3840 ( .A(n3304), .B(n3341), .Z(n3305) );
  AND U3841 ( .A(n2282), .B(n1246), .Z(n3341) );
  XOR U3842 ( .A(n3345), .B(n3306), .Z(n3340) );
  NAND U3843 ( .A(n1316), .B(n2166), .Z(n3306) );
  IV U3844 ( .A(n3308), .Z(n3345) );
  XOR U3845 ( .A(n3349), .B(n3350), .Z(n3311) );
  AND U3846 ( .A(n3351), .B(n3352), .Z(n3350) );
  XNOR U3847 ( .A(n3353), .B(n3354), .Z(n3352) );
  XNOR U3848 ( .A(n3349), .B(n3355), .Z(n3354) );
  XOR U3849 ( .A(n3338), .B(n3356), .Z(n3351) );
  XNOR U3850 ( .A(n3349), .B(n3339), .Z(n3356) );
  XNOR U3851 ( .A(n3321), .B(n3358), .Z(n3322) );
  AND U3852 ( .A(n1642), .B(n1858), .Z(n3358) );
  XOR U3853 ( .A(n3362), .B(n3323), .Z(n3357) );
  NAND U3854 ( .A(n1757), .B(n1737), .Z(n3323) );
  IV U3855 ( .A(n3325), .Z(n3362) );
  XNOR U3856 ( .A(n3330), .B(n3331), .Z(n3327) );
  NAND U3857 ( .A(n1570), .B(n1931), .Z(n3331) );
  XNOR U3858 ( .A(n3329), .B(n3366), .Z(n3330) );
  AND U3859 ( .A(n1831), .B(n1664), .Z(n3366) );
  XOR U3860 ( .A(n3370), .B(n3348), .Z(n3338) );
  XNOR U3861 ( .A(n3335), .B(n3336), .Z(n3348) );
  NAND U3862 ( .A(n1952), .B(n1550), .Z(n3336) );
  XNOR U3863 ( .A(n3334), .B(n3371), .Z(n3335) );
  AND U3864 ( .A(n2053), .B(n1465), .Z(n3371) );
  XNOR U3865 ( .A(n3347), .B(n3337), .Z(n3370) );
  XNOR U3866 ( .A(n3342), .B(n3379), .Z(n3343) );
  AND U3867 ( .A(n2282), .B(n1316), .Z(n3379) );
  XOR U3868 ( .A(n3383), .B(n3344), .Z(n3378) );
  NAND U3869 ( .A(n1388), .B(n2166), .Z(n3344) );
  IV U3870 ( .A(n3346), .Z(n3383) );
  XOR U3871 ( .A(n3387), .B(n3388), .Z(n3349) );
  AND U3872 ( .A(n3389), .B(n3390), .Z(n3388) );
  XNOR U3873 ( .A(n3391), .B(n3392), .Z(n3390) );
  XNOR U3874 ( .A(n3387), .B(n3393), .Z(n3392) );
  XOR U3875 ( .A(n3376), .B(n3394), .Z(n3389) );
  XNOR U3876 ( .A(n3387), .B(n3377), .Z(n3394) );
  XNOR U3877 ( .A(n3359), .B(n3396), .Z(n3360) );
  AND U3878 ( .A(n1737), .B(n1858), .Z(n3396) );
  XOR U3879 ( .A(n3400), .B(n3361), .Z(n3395) );
  NAND U3880 ( .A(n1757), .B(n1831), .Z(n3361) );
  IV U3881 ( .A(n3363), .Z(n3400) );
  XNOR U3882 ( .A(n3368), .B(n3369), .Z(n3365) );
  NAND U3883 ( .A(n1570), .B(n2036), .Z(n3369) );
  XNOR U3884 ( .A(n3367), .B(n3404), .Z(n3368) );
  AND U3885 ( .A(n1931), .B(n1664), .Z(n3404) );
  XOR U3886 ( .A(n3408), .B(n3386), .Z(n3376) );
  XNOR U3887 ( .A(n3373), .B(n3374), .Z(n3386) );
  NAND U3888 ( .A(n1952), .B(n1642), .Z(n3374) );
  XNOR U3889 ( .A(n3372), .B(n3409), .Z(n3373) );
  AND U3890 ( .A(n1550), .B(n2053), .Z(n3409) );
  XNOR U3891 ( .A(n3385), .B(n3375), .Z(n3408) );
  XNOR U3892 ( .A(n3380), .B(n3417), .Z(n3381) );
  AND U3893 ( .A(n2282), .B(n1388), .Z(n3417) );
  XOR U3894 ( .A(n3421), .B(n3382), .Z(n3416) );
  NAND U3895 ( .A(n1465), .B(n2166), .Z(n3382) );
  IV U3896 ( .A(n3384), .Z(n3421) );
  XOR U3897 ( .A(n3425), .B(n3426), .Z(n3387) );
  AND U3898 ( .A(n3427), .B(n3428), .Z(n3426) );
  XNOR U3899 ( .A(n3429), .B(n3430), .Z(n3428) );
  XNOR U3900 ( .A(n3425), .B(n3431), .Z(n3430) );
  XOR U3901 ( .A(n3414), .B(n3432), .Z(n3427) );
  XNOR U3902 ( .A(n3425), .B(n3415), .Z(n3432) );
  XNOR U3903 ( .A(n3397), .B(n3434), .Z(n3398) );
  AND U3904 ( .A(n1831), .B(n1858), .Z(n3434) );
  XOR U3905 ( .A(n3438), .B(n3399), .Z(n3433) );
  NAND U3906 ( .A(n1757), .B(n1931), .Z(n3399) );
  IV U3907 ( .A(n3401), .Z(n3438) );
  XNOR U3908 ( .A(n3406), .B(n3407), .Z(n3403) );
  NAND U3909 ( .A(n1570), .B(n2141), .Z(n3407) );
  XNOR U3910 ( .A(n3405), .B(n3442), .Z(n3406) );
  AND U3911 ( .A(n2036), .B(n1664), .Z(n3442) );
  XOR U3912 ( .A(n3446), .B(n3424), .Z(n3414) );
  XNOR U3913 ( .A(n3411), .B(n3412), .Z(n3424) );
  NAND U3914 ( .A(n1952), .B(n1737), .Z(n3412) );
  XNOR U3915 ( .A(n3410), .B(n3447), .Z(n3411) );
  AND U3916 ( .A(n1642), .B(n2053), .Z(n3447) );
  XNOR U3917 ( .A(n3423), .B(n3413), .Z(n3446) );
  XNOR U3918 ( .A(n3418), .B(n3455), .Z(n3419) );
  AND U3919 ( .A(n2282), .B(n1465), .Z(n3455) );
  XOR U3920 ( .A(n3459), .B(n3420), .Z(n3454) );
  NAND U3921 ( .A(n2166), .B(n1550), .Z(n3420) );
  IV U3922 ( .A(n3422), .Z(n3459) );
  XOR U3923 ( .A(n3463), .B(n3464), .Z(n3425) );
  AND U3924 ( .A(n3465), .B(n3466), .Z(n3464) );
  XNOR U3925 ( .A(n3467), .B(n3468), .Z(n3466) );
  XNOR U3926 ( .A(n3463), .B(n3469), .Z(n3468) );
  XOR U3927 ( .A(n3452), .B(n3470), .Z(n3465) );
  XNOR U3928 ( .A(n3463), .B(n3453), .Z(n3470) );
  XNOR U3929 ( .A(n3435), .B(n3472), .Z(n3436) );
  AND U3930 ( .A(n1931), .B(n1858), .Z(n3472) );
  XOR U3931 ( .A(n3476), .B(n3437), .Z(n3471) );
  NAND U3932 ( .A(n1757), .B(n2036), .Z(n3437) );
  IV U3933 ( .A(n3439), .Z(n3476) );
  XNOR U3934 ( .A(n3444), .B(n3445), .Z(n3441) );
  NAND U3935 ( .A(n1570), .B(n2254), .Z(n3445) );
  XNOR U3936 ( .A(n3443), .B(n3480), .Z(n3444) );
  AND U3937 ( .A(n2141), .B(n1664), .Z(n3480) );
  XOR U3938 ( .A(n3484), .B(n3462), .Z(n3452) );
  XNOR U3939 ( .A(n3449), .B(n3450), .Z(n3462) );
  NAND U3940 ( .A(n1952), .B(n1831), .Z(n3450) );
  XNOR U3941 ( .A(n3448), .B(n3485), .Z(n3449) );
  AND U3942 ( .A(n1737), .B(n2053), .Z(n3485) );
  XNOR U3943 ( .A(n3461), .B(n3451), .Z(n3484) );
  XNOR U3944 ( .A(n3456), .B(n3493), .Z(n3457) );
  AND U3945 ( .A(n1550), .B(n2282), .Z(n3493) );
  XOR U3946 ( .A(n3497), .B(n3458), .Z(n3492) );
  NAND U3947 ( .A(n2166), .B(n1642), .Z(n3458) );
  IV U3948 ( .A(n3460), .Z(n3497) );
  XOR U3949 ( .A(n3501), .B(n3502), .Z(n3463) );
  AND U3950 ( .A(n3503), .B(n3504), .Z(n3502) );
  XNOR U3951 ( .A(n3505), .B(n3506), .Z(n3504) );
  XNOR U3952 ( .A(n3501), .B(n3507), .Z(n3506) );
  XOR U3953 ( .A(n3490), .B(n3508), .Z(n3503) );
  XNOR U3954 ( .A(n3501), .B(n3491), .Z(n3508) );
  XNOR U3955 ( .A(n3473), .B(n3510), .Z(n3474) );
  AND U3956 ( .A(n2036), .B(n1858), .Z(n3510) );
  XOR U3957 ( .A(n3514), .B(n3475), .Z(n3509) );
  NAND U3958 ( .A(n1757), .B(n2141), .Z(n3475) );
  IV U3959 ( .A(n3477), .Z(n3514) );
  XNOR U3960 ( .A(n3482), .B(n3483), .Z(n3479) );
  NAND U3961 ( .A(n1570), .B(n2370), .Z(n3483) );
  XNOR U3962 ( .A(n3481), .B(n3518), .Z(n3482) );
  AND U3963 ( .A(n2254), .B(n1664), .Z(n3518) );
  XOR U3964 ( .A(n3522), .B(n3500), .Z(n3490) );
  XNOR U3965 ( .A(n3487), .B(n3488), .Z(n3500) );
  NAND U3966 ( .A(n1952), .B(n1931), .Z(n3488) );
  XNOR U3967 ( .A(n3486), .B(n3523), .Z(n3487) );
  AND U3968 ( .A(n1831), .B(n2053), .Z(n3523) );
  XNOR U3969 ( .A(n3499), .B(n3489), .Z(n3522) );
  XNOR U3970 ( .A(n3494), .B(n3531), .Z(n3495) );
  AND U3971 ( .A(n1642), .B(n2282), .Z(n3531) );
  XOR U3972 ( .A(n3535), .B(n3496), .Z(n3530) );
  NAND U3973 ( .A(n2166), .B(n1737), .Z(n3496) );
  IV U3974 ( .A(n3498), .Z(n3535) );
  XOR U3975 ( .A(n3539), .B(n3540), .Z(n3501) );
  AND U3976 ( .A(n3541), .B(n3542), .Z(n3540) );
  XNOR U3977 ( .A(n3543), .B(n3544), .Z(n3542) );
  XNOR U3978 ( .A(n3539), .B(n3545), .Z(n3544) );
  XOR U3979 ( .A(n3528), .B(n3546), .Z(n3541) );
  XNOR U3980 ( .A(n3539), .B(n3529), .Z(n3546) );
  XNOR U3981 ( .A(n3511), .B(n3548), .Z(n3512) );
  AND U3982 ( .A(n2141), .B(n1858), .Z(n3548) );
  XOR U3983 ( .A(n3552), .B(n3513), .Z(n3547) );
  NAND U3984 ( .A(n1757), .B(n2254), .Z(n3513) );
  IV U3985 ( .A(n3515), .Z(n3552) );
  XNOR U3986 ( .A(n3520), .B(n3521), .Z(n3517) );
  NAND U3987 ( .A(n1570), .B(n2491), .Z(n3521) );
  XNOR U3988 ( .A(n3519), .B(n3556), .Z(n3520) );
  AND U3989 ( .A(n2370), .B(n1664), .Z(n3556) );
  XOR U3990 ( .A(n3560), .B(n3538), .Z(n3528) );
  XNOR U3991 ( .A(n3525), .B(n3526), .Z(n3538) );
  NAND U3992 ( .A(n1952), .B(n2036), .Z(n3526) );
  XNOR U3993 ( .A(n3524), .B(n3561), .Z(n3525) );
  AND U3994 ( .A(n1931), .B(n2053), .Z(n3561) );
  XNOR U3995 ( .A(n3537), .B(n3527), .Z(n3560) );
  XNOR U3996 ( .A(n3532), .B(n3569), .Z(n3533) );
  AND U3997 ( .A(n1737), .B(n2282), .Z(n3569) );
  XOR U3998 ( .A(n3573), .B(n3534), .Z(n3568) );
  NAND U3999 ( .A(n2166), .B(n1831), .Z(n3534) );
  IV U4000 ( .A(n3536), .Z(n3573) );
  XOR U4001 ( .A(n3577), .B(n3578), .Z(n3539) );
  AND U4002 ( .A(n3579), .B(n3580), .Z(n3578) );
  XNOR U4003 ( .A(n3581), .B(n3582), .Z(n3580) );
  XNOR U4004 ( .A(n3577), .B(n3583), .Z(n3582) );
  XOR U4005 ( .A(n3566), .B(n3584), .Z(n3579) );
  XNOR U4006 ( .A(n3577), .B(n3567), .Z(n3584) );
  XNOR U4007 ( .A(n3549), .B(n3586), .Z(n3550) );
  AND U4008 ( .A(n2254), .B(n1858), .Z(n3586) );
  XOR U4009 ( .A(n3590), .B(n3551), .Z(n3585) );
  NAND U4010 ( .A(n1757), .B(n2370), .Z(n3551) );
  IV U4011 ( .A(n3553), .Z(n3590) );
  XNOR U4012 ( .A(n3558), .B(n3559), .Z(n3555) );
  NAND U4013 ( .A(n1570), .B(n2613), .Z(n3559) );
  XNOR U4014 ( .A(n3557), .B(n3594), .Z(n3558) );
  AND U4015 ( .A(n2491), .B(n1664), .Z(n3594) );
  XOR U4016 ( .A(n3598), .B(n3576), .Z(n3566) );
  XNOR U4017 ( .A(n3563), .B(n3564), .Z(n3576) );
  NAND U4018 ( .A(n1952), .B(n2141), .Z(n3564) );
  XNOR U4019 ( .A(n3562), .B(n3599), .Z(n3563) );
  AND U4020 ( .A(n2036), .B(n2053), .Z(n3599) );
  XNOR U4021 ( .A(n3575), .B(n3565), .Z(n3598) );
  XNOR U4022 ( .A(n3570), .B(n3607), .Z(n3571) );
  AND U4023 ( .A(n1831), .B(n2282), .Z(n3607) );
  XOR U4024 ( .A(n3611), .B(n3572), .Z(n3606) );
  NAND U4025 ( .A(n2166), .B(n1931), .Z(n3572) );
  IV U4026 ( .A(n3574), .Z(n3611) );
  XOR U4027 ( .A(n3615), .B(n3616), .Z(n3577) );
  AND U4028 ( .A(n3617), .B(n3618), .Z(n3616) );
  XNOR U4029 ( .A(n3619), .B(n3620), .Z(n3618) );
  XNOR U4030 ( .A(n3615), .B(n3621), .Z(n3620) );
  XOR U4031 ( .A(n3604), .B(n3622), .Z(n3617) );
  XNOR U4032 ( .A(n3615), .B(n3605), .Z(n3622) );
  XNOR U4033 ( .A(n3587), .B(n3624), .Z(n3588) );
  AND U4034 ( .A(n2370), .B(n1858), .Z(n3624) );
  XOR U4035 ( .A(n3628), .B(n3589), .Z(n3623) );
  NAND U4036 ( .A(n1757), .B(n2491), .Z(n3589) );
  IV U4037 ( .A(n3591), .Z(n3628) );
  XNOR U4038 ( .A(n3596), .B(n3597), .Z(n3593) );
  NAND U4039 ( .A(n1570), .B(n2741), .Z(n3597) );
  XNOR U4040 ( .A(n3595), .B(n3632), .Z(n3596) );
  AND U4041 ( .A(n2613), .B(n1664), .Z(n3632) );
  XOR U4042 ( .A(n3636), .B(n3614), .Z(n3604) );
  XNOR U4043 ( .A(n3601), .B(n3602), .Z(n3614) );
  NAND U4044 ( .A(n1952), .B(n2254), .Z(n3602) );
  XNOR U4045 ( .A(n3600), .B(n3637), .Z(n3601) );
  AND U4046 ( .A(n2141), .B(n2053), .Z(n3637) );
  XNOR U4047 ( .A(n3613), .B(n3603), .Z(n3636) );
  XNOR U4048 ( .A(n3608), .B(n3645), .Z(n3609) );
  AND U4049 ( .A(n1931), .B(n2282), .Z(n3645) );
  XOR U4050 ( .A(n3649), .B(n3610), .Z(n3644) );
  NAND U4051 ( .A(n2166), .B(n2036), .Z(n3610) );
  IV U4052 ( .A(n3612), .Z(n3649) );
  XOR U4053 ( .A(n3653), .B(n3654), .Z(n3615) );
  AND U4054 ( .A(n3655), .B(n3656), .Z(n3654) );
  XNOR U4055 ( .A(n3657), .B(n3658), .Z(n3656) );
  XNOR U4056 ( .A(n3653), .B(n3659), .Z(n3658) );
  XOR U4057 ( .A(n3642), .B(n3660), .Z(n3655) );
  XNOR U4058 ( .A(n3653), .B(n3643), .Z(n3660) );
  XNOR U4059 ( .A(n3625), .B(n3662), .Z(n3626) );
  AND U4060 ( .A(n2491), .B(n1858), .Z(n3662) );
  XOR U4061 ( .A(n3666), .B(n3627), .Z(n3661) );
  NAND U4062 ( .A(n1757), .B(n2613), .Z(n3627) );
  IV U4063 ( .A(n3629), .Z(n3666) );
  XNOR U4064 ( .A(n3634), .B(n3635), .Z(n3631) );
  NANDN U4065 ( .B(n2870), .A(n1570), .Z(n3635) );
  XNOR U4066 ( .A(n3633), .B(n3670), .Z(n3634) );
  AND U4067 ( .A(n2741), .B(n1664), .Z(n3670) );
  XOR U4068 ( .A(n3674), .B(n3652), .Z(n3642) );
  XNOR U4069 ( .A(n3639), .B(n3640), .Z(n3652) );
  NAND U4070 ( .A(n1952), .B(n2370), .Z(n3640) );
  XNOR U4071 ( .A(n3638), .B(n3675), .Z(n3639) );
  AND U4072 ( .A(n2254), .B(n2053), .Z(n3675) );
  XNOR U4073 ( .A(n3651), .B(n3641), .Z(n3674) );
  XNOR U4074 ( .A(n3646), .B(n3683), .Z(n3647) );
  AND U4075 ( .A(n2036), .B(n2282), .Z(n3683) );
  XOR U4076 ( .A(n3687), .B(n3648), .Z(n3682) );
  NAND U4077 ( .A(n2166), .B(n2141), .Z(n3648) );
  IV U4078 ( .A(n3650), .Z(n3687) );
  XOR U4079 ( .A(n3691), .B(n3692), .Z(n3653) );
  AND U4080 ( .A(n3693), .B(n3694), .Z(n3692) );
  XNOR U4081 ( .A(n3695), .B(n3696), .Z(n3694) );
  XNOR U4082 ( .A(n3691), .B(n3697), .Z(n3696) );
  XOR U4083 ( .A(n3680), .B(n3698), .Z(n3693) );
  XNOR U4084 ( .A(n3691), .B(n3681), .Z(n3698) );
  XNOR U4085 ( .A(n3663), .B(n3700), .Z(n3664) );
  AND U4086 ( .A(n2613), .B(n1858), .Z(n3700) );
  XOR U4087 ( .A(n3704), .B(n3665), .Z(n3699) );
  NAND U4088 ( .A(n1757), .B(n2741), .Z(n3665) );
  IV U4089 ( .A(n3667), .Z(n3704) );
  XNOR U4090 ( .A(n3672), .B(n3673), .Z(n3669) );
  NANDN U4091 ( .B(n3008), .A(n1570), .Z(n3673) );
  XNOR U4092 ( .A(n3671), .B(n3708), .Z(n3672) );
  ANDN U4093 ( .A(n1664), .B(n2870), .Z(n3708) );
  XOR U4094 ( .A(n3712), .B(n3690), .Z(n3680) );
  XNOR U4095 ( .A(n3677), .B(n3678), .Z(n3690) );
  NAND U4096 ( .A(n1952), .B(n2491), .Z(n3678) );
  XNOR U4097 ( .A(n3676), .B(n3713), .Z(n3677) );
  AND U4098 ( .A(n2370), .B(n2053), .Z(n3713) );
  XNOR U4099 ( .A(n3689), .B(n3679), .Z(n3712) );
  XNOR U4100 ( .A(n3684), .B(n3721), .Z(n3685) );
  AND U4101 ( .A(n2141), .B(n2282), .Z(n3721) );
  XOR U4102 ( .A(n3725), .B(n3686), .Z(n3720) );
  NAND U4103 ( .A(n2166), .B(n2254), .Z(n3686) );
  IV U4104 ( .A(n3688), .Z(n3725) );
  XOR U4105 ( .A(n3729), .B(n3730), .Z(n3691) );
  AND U4106 ( .A(n3731), .B(n3732), .Z(n3730) );
  XNOR U4107 ( .A(n3733), .B(n3734), .Z(n3732) );
  XNOR U4108 ( .A(n3729), .B(n3735), .Z(n3734) );
  XOR U4109 ( .A(n3718), .B(n3736), .Z(n3731) );
  XNOR U4110 ( .A(n3729), .B(n3719), .Z(n3736) );
  XNOR U4111 ( .A(n3701), .B(n3738), .Z(n3702) );
  AND U4112 ( .A(n2741), .B(n1858), .Z(n3738) );
  XOR U4113 ( .A(n3742), .B(n3703), .Z(n3737) );
  NANDN U4114 ( .B(n2870), .A(n1757), .Z(n3703) );
  IV U4115 ( .A(n3705), .Z(n3742) );
  XNOR U4116 ( .A(n3710), .B(n3711), .Z(n3707) );
  NAND U4117 ( .A(n1570), .B(n3144), .Z(n3711) );
  XNOR U4118 ( .A(n3709), .B(n3746), .Z(n3710) );
  ANDN U4119 ( .A(n1664), .B(n3008), .Z(n3746) );
  XOR U4120 ( .A(n3750), .B(n3728), .Z(n3718) );
  XNOR U4121 ( .A(n3715), .B(n3716), .Z(n3728) );
  NAND U4122 ( .A(n1952), .B(n2613), .Z(n3716) );
  XNOR U4123 ( .A(n3714), .B(n3751), .Z(n3715) );
  AND U4124 ( .A(n2491), .B(n2053), .Z(n3751) );
  XNOR U4125 ( .A(n3727), .B(n3717), .Z(n3750) );
  XNOR U4126 ( .A(n3722), .B(n3759), .Z(n3723) );
  AND U4127 ( .A(n2254), .B(n2282), .Z(n3759) );
  XOR U4128 ( .A(n3763), .B(n3724), .Z(n3758) );
  NAND U4129 ( .A(n2166), .B(n2370), .Z(n3724) );
  IV U4130 ( .A(n3726), .Z(n3763) );
  XNOR U4131 ( .A(n3768), .B(n3769), .Z(n3182) );
  XOR U4132 ( .A(n3770), .B(n3767), .Z(n3768) );
  XNOR U4133 ( .A(n3771), .B(n3766), .Z(n3756) );
  XNOR U4134 ( .A(n3753), .B(n3754), .Z(n3766) );
  NAND U4135 ( .A(n1952), .B(n2741), .Z(n3754) );
  XNOR U4136 ( .A(n3752), .B(n3772), .Z(n3753) );
  AND U4137 ( .A(n2613), .B(n2053), .Z(n3772) );
  XNOR U4138 ( .A(n3776), .B(n3773), .Z(n3775) );
  XNOR U4139 ( .A(n3765), .B(n3755), .Z(n3771) );
  XOR U4140 ( .A(n3777), .B(n3778), .Z(n3755) );
  XNOR U4141 ( .A(n3760), .B(n3780), .Z(n3761) );
  AND U4142 ( .A(n2370), .B(n2282), .Z(n3780) );
  XNOR U4143 ( .A(n3784), .B(n3781), .Z(n3783) );
  XOR U4144 ( .A(n3785), .B(n3762), .Z(n3779) );
  NAND U4145 ( .A(n2166), .B(n2491), .Z(n3762) );
  IV U4146 ( .A(n3764), .Z(n3785) );
  XNOR U4147 ( .A(n3786), .B(n3787), .Z(n3764) );
  AND U4148 ( .A(n3788), .B(n3789), .Z(n3787) );
  XOR U4149 ( .A(n3782), .B(n3790), .Z(n3789) );
  XNOR U4150 ( .A(n3784), .B(n3786), .Z(n3790) );
  NAND U4151 ( .A(n2166), .B(n2613), .Z(n3784) );
  XOR U4152 ( .A(n3781), .B(n3791), .Z(n3782) );
  AND U4153 ( .A(n2491), .B(n2282), .Z(n3791) );
  XNOR U4154 ( .A(n3795), .B(n3792), .Z(n3794) );
  XOR U4155 ( .A(n3774), .B(n3796), .Z(n3788) );
  XNOR U4156 ( .A(n3776), .B(n3786), .Z(n3796) );
  NANDN U4157 ( .B(n2870), .A(n1952), .Z(n3776) );
  XOR U4158 ( .A(n3773), .B(n3797), .Z(n3774) );
  AND U4159 ( .A(n2741), .B(n2053), .Z(n3797) );
  XNOR U4160 ( .A(n3801), .B(n3798), .Z(n3800) );
  XOR U4161 ( .A(n3802), .B(n3803), .Z(n3786) );
  AND U4162 ( .A(n3804), .B(n3805), .Z(n3803) );
  XOR U4163 ( .A(n3793), .B(n3806), .Z(n3805) );
  XNOR U4164 ( .A(n3795), .B(n3802), .Z(n3806) );
  NAND U4165 ( .A(n2166), .B(n2741), .Z(n3795) );
  XOR U4166 ( .A(n3792), .B(n3807), .Z(n3793) );
  AND U4167 ( .A(n2613), .B(n2282), .Z(n3807) );
  XNOR U4168 ( .A(n3811), .B(n3808), .Z(n3810) );
  XOR U4169 ( .A(n3799), .B(n3812), .Z(n3804) );
  XNOR U4170 ( .A(n3801), .B(n3802), .Z(n3812) );
  NANDN U4171 ( .B(n3008), .A(n1952), .Z(n3801) );
  XOR U4172 ( .A(n3798), .B(n3813), .Z(n3799) );
  ANDN U4173 ( .A(n2053), .B(n2870), .Z(n3813) );
  XNOR U4174 ( .A(n3817), .B(n3814), .Z(n3816) );
  XOR U4175 ( .A(n3818), .B(n3819), .Z(n3802) );
  AND U4176 ( .A(n3820), .B(n3821), .Z(n3819) );
  XOR U4177 ( .A(n3809), .B(n3822), .Z(n3821) );
  XNOR U4178 ( .A(n3811), .B(n3818), .Z(n3822) );
  NANDN U4179 ( .B(n2870), .A(n2166), .Z(n3811) );
  XOR U4180 ( .A(n3808), .B(n3823), .Z(n3809) );
  AND U4181 ( .A(n2741), .B(n2282), .Z(n3823) );
  XOR U4182 ( .A(n3815), .B(n3827), .Z(n3820) );
  XNOR U4183 ( .A(n3817), .B(n3818), .Z(n3827) );
  NAND U4184 ( .A(n1952), .B(n3144), .Z(n3817) );
  XOR U4185 ( .A(n3814), .B(n3828), .Z(n3815) );
  ANDN U4186 ( .A(n2053), .B(n3008), .Z(n3828) );
  NAND U4187 ( .A(n1952), .B(n3833), .Z(n3831) );
  XNOR U4188 ( .A(n3829), .B(n3834), .Z(n3830) );
  AND U4189 ( .A(n3144), .B(n2053), .Z(n3834) );
  AND U4190 ( .A(n3835), .B(g_input[0]), .Z(n3829) );
  NANDN U4191 ( .B(n1952), .A(n3836), .Z(n3835) );
  NAND U4192 ( .A(n3833), .B(n2053), .Z(n3836) );
  XNOR U4193 ( .A(n3824), .B(n3840), .Z(n3825) );
  ANDN U4194 ( .A(n2282), .B(n2870), .Z(n3840) );
  XOR U4195 ( .A(n3843), .B(n3841), .Z(n3842) );
  ANDN U4196 ( .A(n2282), .B(n3008), .Z(n3843) );
  AND U4197 ( .A(n3144), .B(n2166), .Z(n3844) );
  XOR U4198 ( .A(n3848), .B(n3826), .Z(n3839) );
  NANDN U4199 ( .B(n3008), .A(n2166), .Z(n3826) );
  IV U4200 ( .A(n3832), .Z(n3848) );
  NAND U4201 ( .A(n2166), .B(n3833), .Z(n3847) );
  XNOR U4202 ( .A(n3845), .B(n3849), .Z(n3846) );
  AND U4203 ( .A(n3144), .B(n2282), .Z(n3849) );
  AND U4204 ( .A(n3850), .B(g_input[0]), .Z(n3845) );
  NANDN U4205 ( .B(n2166), .A(n3851), .Z(n3850) );
  NAND U4206 ( .A(n3833), .B(n2282), .Z(n3851) );
  XNOR U4207 ( .A(n3739), .B(n3855), .Z(n3740) );
  ANDN U4208 ( .A(n1858), .B(n2870), .Z(n3855) );
  XOR U4209 ( .A(n3858), .B(n3856), .Z(n3857) );
  ANDN U4210 ( .A(n1858), .B(n3008), .Z(n3858) );
  AND U4211 ( .A(n3144), .B(n1757), .Z(n3859) );
  XOR U4212 ( .A(n3863), .B(n3741), .Z(n3854) );
  NANDN U4213 ( .B(n3008), .A(n1757), .Z(n3741) );
  IV U4214 ( .A(n3743), .Z(n3863) );
  NAND U4215 ( .A(n1757), .B(n3833), .Z(n3862) );
  XNOR U4216 ( .A(n3860), .B(n3864), .Z(n3861) );
  AND U4217 ( .A(n3144), .B(n1858), .Z(n3864) );
  AND U4218 ( .A(n3865), .B(g_input[0]), .Z(n3860) );
  NANDN U4219 ( .B(n1757), .A(n3866), .Z(n3865) );
  NAND U4220 ( .A(n3833), .B(n1858), .Z(n3866) );
  XNOR U4221 ( .A(n3748), .B(n3749), .Z(n3745) );
  NAND U4222 ( .A(n1570), .B(n3833), .Z(n3749) );
  XNOR U4223 ( .A(n3747), .B(n3869), .Z(n3748) );
  AND U4224 ( .A(n3144), .B(n1664), .Z(n3869) );
  AND U4225 ( .A(n3870), .B(g_input[0]), .Z(n3747) );
  NANDN U4226 ( .B(n1570), .A(n3871), .Z(n3870) );
  NAND U4227 ( .A(n3833), .B(n1664), .Z(n3871) );
  XOR U4228 ( .A(n3874), .B(n3875), .Z(n3767) );
  XNOR U4229 ( .A(n3876), .B(n3083), .Z(n3079) );
  NAND U4230 ( .A(n778), .B(n2942), .Z(n3077) );
  XNOR U4231 ( .A(n3075), .B(n3877), .Z(n3076) );
  AND U4232 ( .A(n3074), .B(n744), .Z(n3877) );
  XNOR U4233 ( .A(n3082), .B(n3078), .Z(n3876) );
  XNOR U4234 ( .A(n3186), .B(n3883), .Z(n3187) );
  AND U4235 ( .A(n2796), .B(n855), .Z(n3883) );
  XOR U4236 ( .A(n3887), .B(n3188), .Z(n3882) );
  NAND U4237 ( .A(n899), .B(n2666), .Z(n3188) );
  IV U4238 ( .A(n3190), .Z(n3887) );
  XNOR U4239 ( .A(n3195), .B(n3196), .Z(n3192) );
  NAND U4240 ( .A(n1003), .B(n2421), .Z(n3196) );
  XNOR U4241 ( .A(n3194), .B(n3891), .Z(n3195) );
  AND U4242 ( .A(n2544), .B(n945), .Z(n3891) );
  XOR U4243 ( .A(n3895), .B(n3896), .Z(n3203) );
  XNOR U4244 ( .A(n3897), .B(n3881), .Z(n3895) );
  XOR U4245 ( .A(n3899), .B(n3900), .Z(n3241) );
  XNOR U4246 ( .A(n3901), .B(n3898), .Z(n3899) );
  XNOR U4247 ( .A(n3884), .B(n3903), .Z(n3885) );
  AND U4248 ( .A(n2796), .B(n899), .Z(n3903) );
  XOR U4249 ( .A(n3907), .B(n3886), .Z(n3902) );
  NAND U4250 ( .A(n945), .B(n2666), .Z(n3886) );
  IV U4251 ( .A(n3888), .Z(n3907) );
  XNOR U4252 ( .A(n3893), .B(n3894), .Z(n3890) );
  NAND U4253 ( .A(n1057), .B(n2421), .Z(n3894) );
  XNOR U4254 ( .A(n3892), .B(n3911), .Z(n3893) );
  AND U4255 ( .A(n2544), .B(n1003), .Z(n3911) );
  XOR U4256 ( .A(n3916), .B(n3917), .Z(n3279) );
  XNOR U4257 ( .A(n3918), .B(n3915), .Z(n3916) );
  XNOR U4258 ( .A(n3904), .B(n3920), .Z(n3905) );
  AND U4259 ( .A(n2796), .B(n945), .Z(n3920) );
  XOR U4260 ( .A(n3924), .B(n3906), .Z(n3919) );
  NAND U4261 ( .A(n1003), .B(n2666), .Z(n3906) );
  IV U4262 ( .A(n3908), .Z(n3924) );
  XNOR U4263 ( .A(n3913), .B(n3914), .Z(n3910) );
  NAND U4264 ( .A(n1119), .B(n2421), .Z(n3914) );
  XNOR U4265 ( .A(n3912), .B(n3928), .Z(n3913) );
  AND U4266 ( .A(n2544), .B(n1057), .Z(n3928) );
  XOR U4267 ( .A(n3933), .B(n3934), .Z(n3317) );
  XNOR U4268 ( .A(n3935), .B(n3932), .Z(n3933) );
  XNOR U4269 ( .A(n3921), .B(n3937), .Z(n3922) );
  AND U4270 ( .A(n2796), .B(n1003), .Z(n3937) );
  XOR U4271 ( .A(n3941), .B(n3923), .Z(n3936) );
  NAND U4272 ( .A(n1057), .B(n2666), .Z(n3923) );
  IV U4273 ( .A(n3925), .Z(n3941) );
  XNOR U4274 ( .A(n3930), .B(n3931), .Z(n3927) );
  NAND U4275 ( .A(n1180), .B(n2421), .Z(n3931) );
  XNOR U4276 ( .A(n3929), .B(n3945), .Z(n3930) );
  AND U4277 ( .A(n2544), .B(n1119), .Z(n3945) );
  XOR U4278 ( .A(n3950), .B(n3951), .Z(n3355) );
  XNOR U4279 ( .A(n3952), .B(n3949), .Z(n3950) );
  XNOR U4280 ( .A(n3938), .B(n3954), .Z(n3939) );
  AND U4281 ( .A(n2796), .B(n1057), .Z(n3954) );
  XOR U4282 ( .A(n3958), .B(n3940), .Z(n3953) );
  NAND U4283 ( .A(n1119), .B(n2666), .Z(n3940) );
  IV U4284 ( .A(n3942), .Z(n3958) );
  XNOR U4285 ( .A(n3947), .B(n3948), .Z(n3944) );
  NAND U4286 ( .A(n1246), .B(n2421), .Z(n3948) );
  XNOR U4287 ( .A(n3946), .B(n3962), .Z(n3947) );
  AND U4288 ( .A(n2544), .B(n1180), .Z(n3962) );
  XOR U4289 ( .A(n3967), .B(n3968), .Z(n3393) );
  XNOR U4290 ( .A(n3969), .B(n3966), .Z(n3967) );
  XNOR U4291 ( .A(n3955), .B(n3971), .Z(n3956) );
  AND U4292 ( .A(n2796), .B(n1119), .Z(n3971) );
  XOR U4293 ( .A(n3975), .B(n3957), .Z(n3970) );
  NAND U4294 ( .A(n1180), .B(n2666), .Z(n3957) );
  IV U4295 ( .A(n3959), .Z(n3975) );
  XNOR U4296 ( .A(n3964), .B(n3965), .Z(n3961) );
  NAND U4297 ( .A(n1316), .B(n2421), .Z(n3965) );
  XNOR U4298 ( .A(n3963), .B(n3979), .Z(n3964) );
  AND U4299 ( .A(n2544), .B(n1246), .Z(n3979) );
  XOR U4300 ( .A(n3984), .B(n3985), .Z(n3431) );
  XNOR U4301 ( .A(n3986), .B(n3983), .Z(n3984) );
  XNOR U4302 ( .A(n3972), .B(n3988), .Z(n3973) );
  AND U4303 ( .A(n2796), .B(n1180), .Z(n3988) );
  XOR U4304 ( .A(n3992), .B(n3974), .Z(n3987) );
  NAND U4305 ( .A(n1246), .B(n2666), .Z(n3974) );
  IV U4306 ( .A(n3976), .Z(n3992) );
  XNOR U4307 ( .A(n3981), .B(n3982), .Z(n3978) );
  NAND U4308 ( .A(n1388), .B(n2421), .Z(n3982) );
  XNOR U4309 ( .A(n3980), .B(n3996), .Z(n3981) );
  AND U4310 ( .A(n2544), .B(n1316), .Z(n3996) );
  XOR U4311 ( .A(n4001), .B(n4002), .Z(n3469) );
  XNOR U4312 ( .A(n4003), .B(n4000), .Z(n4001) );
  XNOR U4313 ( .A(n3989), .B(n4005), .Z(n3990) );
  AND U4314 ( .A(n2796), .B(n1246), .Z(n4005) );
  XOR U4315 ( .A(n4009), .B(n3991), .Z(n4004) );
  NAND U4316 ( .A(n1316), .B(n2666), .Z(n3991) );
  IV U4317 ( .A(n3993), .Z(n4009) );
  XNOR U4318 ( .A(n3998), .B(n3999), .Z(n3995) );
  NAND U4319 ( .A(n1465), .B(n2421), .Z(n3999) );
  XNOR U4320 ( .A(n3997), .B(n4013), .Z(n3998) );
  AND U4321 ( .A(n2544), .B(n1388), .Z(n4013) );
  XOR U4322 ( .A(n4018), .B(n4019), .Z(n3507) );
  XNOR U4323 ( .A(n4020), .B(n4017), .Z(n4018) );
  XNOR U4324 ( .A(n4006), .B(n4022), .Z(n4007) );
  AND U4325 ( .A(n2796), .B(n1316), .Z(n4022) );
  XOR U4326 ( .A(n4026), .B(n4008), .Z(n4021) );
  NAND U4327 ( .A(n1388), .B(n2666), .Z(n4008) );
  IV U4328 ( .A(n4010), .Z(n4026) );
  XNOR U4329 ( .A(n4015), .B(n4016), .Z(n4012) );
  NAND U4330 ( .A(n1550), .B(n2421), .Z(n4016) );
  XNOR U4331 ( .A(n4014), .B(n4030), .Z(n4015) );
  AND U4332 ( .A(n2544), .B(n1465), .Z(n4030) );
  XOR U4333 ( .A(n4035), .B(n4036), .Z(n3545) );
  XNOR U4334 ( .A(n4037), .B(n4034), .Z(n4035) );
  XNOR U4335 ( .A(n4023), .B(n4039), .Z(n4024) );
  AND U4336 ( .A(n2796), .B(n1388), .Z(n4039) );
  XOR U4337 ( .A(n4043), .B(n4025), .Z(n4038) );
  NAND U4338 ( .A(n1465), .B(n2666), .Z(n4025) );
  IV U4339 ( .A(n4027), .Z(n4043) );
  XNOR U4340 ( .A(n4032), .B(n4033), .Z(n4029) );
  NAND U4341 ( .A(n1642), .B(n2421), .Z(n4033) );
  XNOR U4342 ( .A(n4031), .B(n4047), .Z(n4032) );
  AND U4343 ( .A(n2544), .B(n1550), .Z(n4047) );
  XOR U4344 ( .A(n4052), .B(n4053), .Z(n3583) );
  XNOR U4345 ( .A(n4054), .B(n4051), .Z(n4052) );
  XNOR U4346 ( .A(n4040), .B(n4056), .Z(n4041) );
  AND U4347 ( .A(n2796), .B(n1465), .Z(n4056) );
  XOR U4348 ( .A(n4060), .B(n4042), .Z(n4055) );
  NAND U4349 ( .A(n1550), .B(n2666), .Z(n4042) );
  IV U4350 ( .A(n4044), .Z(n4060) );
  XNOR U4351 ( .A(n4049), .B(n4050), .Z(n4046) );
  NAND U4352 ( .A(n1737), .B(n2421), .Z(n4050) );
  XNOR U4353 ( .A(n4048), .B(n4064), .Z(n4049) );
  AND U4354 ( .A(n2544), .B(n1642), .Z(n4064) );
  XOR U4355 ( .A(n4069), .B(n4070), .Z(n3621) );
  XNOR U4356 ( .A(n4071), .B(n4068), .Z(n4069) );
  XNOR U4357 ( .A(n4057), .B(n4073), .Z(n4058) );
  AND U4358 ( .A(n2796), .B(n1550), .Z(n4073) );
  XOR U4359 ( .A(n4077), .B(n4059), .Z(n4072) );
  NAND U4360 ( .A(n1642), .B(n2666), .Z(n4059) );
  IV U4361 ( .A(n4061), .Z(n4077) );
  XNOR U4362 ( .A(n4066), .B(n4067), .Z(n4063) );
  NAND U4363 ( .A(n1831), .B(n2421), .Z(n4067) );
  XNOR U4364 ( .A(n4065), .B(n4081), .Z(n4066) );
  AND U4365 ( .A(n2544), .B(n1737), .Z(n4081) );
  XOR U4366 ( .A(n4086), .B(n4087), .Z(n3659) );
  XNOR U4367 ( .A(n4088), .B(n4085), .Z(n4086) );
  XNOR U4368 ( .A(n4074), .B(n4090), .Z(n4075) );
  AND U4369 ( .A(n2796), .B(n1642), .Z(n4090) );
  XOR U4370 ( .A(n4094), .B(n4076), .Z(n4089) );
  NAND U4371 ( .A(n1737), .B(n2666), .Z(n4076) );
  IV U4372 ( .A(n4078), .Z(n4094) );
  XNOR U4373 ( .A(n4083), .B(n4084), .Z(n4080) );
  NAND U4374 ( .A(n1931), .B(n2421), .Z(n4084) );
  XNOR U4375 ( .A(n4082), .B(n4098), .Z(n4083) );
  AND U4376 ( .A(n2544), .B(n1831), .Z(n4098) );
  XOR U4377 ( .A(n4103), .B(n4104), .Z(n3697) );
  XNOR U4378 ( .A(n4105), .B(n4102), .Z(n4103) );
  XNOR U4379 ( .A(n4091), .B(n4107), .Z(n4092) );
  AND U4380 ( .A(n2796), .B(n1737), .Z(n4107) );
  XOR U4381 ( .A(n4111), .B(n4093), .Z(n4106) );
  NAND U4382 ( .A(n1831), .B(n2666), .Z(n4093) );
  IV U4383 ( .A(n4095), .Z(n4111) );
  XNOR U4384 ( .A(n4100), .B(n4101), .Z(n4097) );
  NAND U4385 ( .A(n2036), .B(n2421), .Z(n4101) );
  XNOR U4386 ( .A(n4099), .B(n4115), .Z(n4100) );
  AND U4387 ( .A(n2544), .B(n1931), .Z(n4115) );
  XOR U4388 ( .A(n4120), .B(n4121), .Z(n3735) );
  XNOR U4389 ( .A(n4122), .B(n4119), .Z(n4120) );
  XNOR U4390 ( .A(n4108), .B(n4124), .Z(n4109) );
  AND U4391 ( .A(n2796), .B(n1831), .Z(n4124) );
  XOR U4392 ( .A(n4128), .B(n4110), .Z(n4123) );
  NAND U4393 ( .A(n1931), .B(n2666), .Z(n4110) );
  IV U4394 ( .A(n4112), .Z(n4128) );
  XNOR U4395 ( .A(n4117), .B(n4118), .Z(n4114) );
  NAND U4396 ( .A(n2141), .B(n2421), .Z(n4118) );
  XNOR U4397 ( .A(n4116), .B(n4132), .Z(n4117) );
  AND U4398 ( .A(n2544), .B(n2036), .Z(n4132) );
  XOR U4399 ( .A(n4137), .B(n4138), .Z(n3770) );
  XNOR U4400 ( .A(n4139), .B(n4136), .Z(n4137) );
  XNOR U4401 ( .A(n4125), .B(n4141), .Z(n4126) );
  AND U4402 ( .A(n2796), .B(n1931), .Z(n4141) );
  XOR U4403 ( .A(n4145), .B(n4127), .Z(n4140) );
  NAND U4404 ( .A(n2036), .B(n2666), .Z(n4127) );
  IV U4405 ( .A(n4129), .Z(n4145) );
  XNOR U4406 ( .A(n4134), .B(n4135), .Z(n4131) );
  NAND U4407 ( .A(n2254), .B(n2421), .Z(n4135) );
  XNOR U4408 ( .A(n4133), .B(n4149), .Z(n4134) );
  AND U4409 ( .A(n2544), .B(n2141), .Z(n4149) );
  XOR U4410 ( .A(n4153), .B(n4154), .Z(n4136) );
  AND U4411 ( .A(n4155), .B(n4156), .Z(n4154) );
  XOR U4412 ( .A(n4157), .B(n4158), .Z(n4156) );
  XOR U4413 ( .A(n4153), .B(n4159), .Z(n4158) );
  XOR U4414 ( .A(n4147), .B(n4160), .Z(n4155) );
  XOR U4415 ( .A(n4153), .B(n4148), .Z(n4160) );
  NAND U4416 ( .A(n2421), .B(n2370), .Z(n4152) );
  XNOR U4417 ( .A(n4150), .B(n4161), .Z(n4151) );
  AND U4418 ( .A(n2544), .B(n2254), .Z(n4161) );
  XNOR U4419 ( .A(n4142), .B(n4166), .Z(n4143) );
  AND U4420 ( .A(n2796), .B(n2036), .Z(n4166) );
  XOR U4421 ( .A(n4170), .B(n4144), .Z(n4165) );
  NAND U4422 ( .A(n2141), .B(n2666), .Z(n4144) );
  IV U4423 ( .A(n4146), .Z(n4170) );
  XOR U4424 ( .A(n4174), .B(n4175), .Z(n4153) );
  AND U4425 ( .A(n4176), .B(n4177), .Z(n4175) );
  XOR U4426 ( .A(n4178), .B(n4179), .Z(n4177) );
  XOR U4427 ( .A(n4174), .B(n4180), .Z(n4179) );
  XOR U4428 ( .A(n4172), .B(n4181), .Z(n4176) );
  XOR U4429 ( .A(n4174), .B(n4173), .Z(n4181) );
  NAND U4430 ( .A(n2421), .B(n2491), .Z(n4164) );
  XNOR U4431 ( .A(n4162), .B(n4182), .Z(n4163) );
  AND U4432 ( .A(n2370), .B(n2544), .Z(n4182) );
  XNOR U4433 ( .A(n4167), .B(n4187), .Z(n4168) );
  AND U4434 ( .A(n2796), .B(n2141), .Z(n4187) );
  XOR U4435 ( .A(n4191), .B(n4169), .Z(n4186) );
  NAND U4436 ( .A(n2254), .B(n2666), .Z(n4169) );
  IV U4437 ( .A(n4171), .Z(n4191) );
  XOR U4438 ( .A(n4195), .B(n4196), .Z(n4174) );
  AND U4439 ( .A(n4197), .B(n4198), .Z(n4196) );
  XOR U4440 ( .A(n4199), .B(n4200), .Z(n4198) );
  XOR U4441 ( .A(n4195), .B(n4201), .Z(n4200) );
  XOR U4442 ( .A(n4193), .B(n4202), .Z(n4197) );
  XOR U4443 ( .A(n4195), .B(n4194), .Z(n4202) );
  NAND U4444 ( .A(n2421), .B(n2613), .Z(n4185) );
  XNOR U4445 ( .A(n4183), .B(n4203), .Z(n4184) );
  AND U4446 ( .A(n2491), .B(n2544), .Z(n4203) );
  XNOR U4447 ( .A(n4188), .B(n4208), .Z(n4189) );
  AND U4448 ( .A(n2796), .B(n2254), .Z(n4208) );
  XOR U4449 ( .A(n4212), .B(n4190), .Z(n4207) );
  NAND U4450 ( .A(n2666), .B(n2370), .Z(n4190) );
  IV U4451 ( .A(n4192), .Z(n4212) );
  XOR U4452 ( .A(n4216), .B(n4217), .Z(n4195) );
  AND U4453 ( .A(n4218), .B(n4219), .Z(n4217) );
  XOR U4454 ( .A(n4220), .B(n4221), .Z(n4219) );
  XOR U4455 ( .A(n4216), .B(n4222), .Z(n4221) );
  XOR U4456 ( .A(n4214), .B(n4223), .Z(n4218) );
  XOR U4457 ( .A(n4216), .B(n4215), .Z(n4223) );
  NAND U4458 ( .A(n2421), .B(n2741), .Z(n4206) );
  XNOR U4459 ( .A(n4204), .B(n4224), .Z(n4205) );
  AND U4460 ( .A(n2613), .B(n2544), .Z(n4224) );
  XNOR U4461 ( .A(n4209), .B(n4229), .Z(n4210) );
  AND U4462 ( .A(n2370), .B(n2796), .Z(n4229) );
  XOR U4463 ( .A(n4233), .B(n4211), .Z(n4228) );
  NAND U4464 ( .A(n2666), .B(n2491), .Z(n4211) );
  IV U4465 ( .A(n4213), .Z(n4233) );
  XOR U4466 ( .A(n4237), .B(n4238), .Z(n4216) );
  AND U4467 ( .A(n4239), .B(n4240), .Z(n4238) );
  XOR U4468 ( .A(n4241), .B(n4242), .Z(n4240) );
  XOR U4469 ( .A(n4237), .B(n4243), .Z(n4242) );
  XOR U4470 ( .A(n4235), .B(n4244), .Z(n4239) );
  XOR U4471 ( .A(n4237), .B(n4236), .Z(n4244) );
  NANDN U4472 ( .B(n2870), .A(n2421), .Z(n4227) );
  XNOR U4473 ( .A(n4225), .B(n4245), .Z(n4226) );
  AND U4474 ( .A(n2741), .B(n2544), .Z(n4245) );
  XNOR U4475 ( .A(n4230), .B(n4250), .Z(n4231) );
  AND U4476 ( .A(n2491), .B(n2796), .Z(n4250) );
  XOR U4477 ( .A(n4254), .B(n4232), .Z(n4249) );
  NAND U4478 ( .A(n2666), .B(n2613), .Z(n4232) );
  IV U4479 ( .A(n4234), .Z(n4254) );
  XOR U4480 ( .A(n4258), .B(n4259), .Z(n4237) );
  AND U4481 ( .A(n4260), .B(n4261), .Z(n4259) );
  XOR U4482 ( .A(n4262), .B(n4263), .Z(n4261) );
  XOR U4483 ( .A(n4258), .B(n4264), .Z(n4263) );
  XOR U4484 ( .A(n4256), .B(n4265), .Z(n4260) );
  XOR U4485 ( .A(n4258), .B(n4257), .Z(n4265) );
  NANDN U4486 ( .B(n3008), .A(n2421), .Z(n4248) );
  XNOR U4487 ( .A(n4246), .B(n4266), .Z(n4247) );
  ANDN U4488 ( .A(n2544), .B(n2870), .Z(n4266) );
  XNOR U4489 ( .A(n4251), .B(n4271), .Z(n4252) );
  AND U4490 ( .A(n2613), .B(n2796), .Z(n4271) );
  XOR U4491 ( .A(n4275), .B(n4253), .Z(n4270) );
  NAND U4492 ( .A(n2666), .B(n2741), .Z(n4253) );
  IV U4493 ( .A(n4255), .Z(n4275) );
  XOR U4494 ( .A(n4279), .B(n4280), .Z(n4258) );
  AND U4495 ( .A(n4281), .B(n4282), .Z(n4280) );
  XOR U4496 ( .A(n4283), .B(n4284), .Z(n4282) );
  XOR U4497 ( .A(n4279), .B(n4285), .Z(n4284) );
  XOR U4498 ( .A(n4277), .B(n4286), .Z(n4281) );
  XOR U4499 ( .A(n4279), .B(n4278), .Z(n4286) );
  NAND U4500 ( .A(n2421), .B(n3144), .Z(n4269) );
  XNOR U4501 ( .A(n4267), .B(n4287), .Z(n4268) );
  ANDN U4502 ( .A(n2544), .B(n3008), .Z(n4287) );
  XNOR U4503 ( .A(n4272), .B(n4292), .Z(n4273) );
  AND U4504 ( .A(n2741), .B(n2796), .Z(n4292) );
  XOR U4505 ( .A(n4296), .B(n4274), .Z(n4291) );
  NANDN U4506 ( .B(n2870), .A(n2666), .Z(n4274) );
  IV U4507 ( .A(n4276), .Z(n4296) );
  XOR U4508 ( .A(n4301), .B(n4302), .Z(n3875) );
  XNOR U4509 ( .A(n4303), .B(n4300), .Z(n4301) );
  XNOR U4510 ( .A(n4293), .B(n4305), .Z(n4294) );
  ANDN U4511 ( .A(n2796), .B(n2870), .Z(n4305) );
  XOR U4512 ( .A(n4308), .B(n4306), .Z(n4307) );
  ANDN U4513 ( .A(n2796), .B(n3008), .Z(n4308) );
  AND U4514 ( .A(n3144), .B(n2666), .Z(n4309) );
  XOR U4515 ( .A(n4313), .B(n4295), .Z(n4304) );
  NANDN U4516 ( .B(n3008), .A(n2666), .Z(n4295) );
  IV U4517 ( .A(n4297), .Z(n4313) );
  NAND U4518 ( .A(n2666), .B(n3833), .Z(n4312) );
  XNOR U4519 ( .A(n4310), .B(n4314), .Z(n4311) );
  AND U4520 ( .A(n3144), .B(n2796), .Z(n4314) );
  AND U4521 ( .A(n4315), .B(g_input[0]), .Z(n4310) );
  NANDN U4522 ( .B(n2666), .A(n4316), .Z(n4315) );
  NAND U4523 ( .A(n3833), .B(n2796), .Z(n4316) );
  XNOR U4524 ( .A(n4289), .B(n4290), .Z(n4299) );
  NAND U4525 ( .A(n2421), .B(n3833), .Z(n4290) );
  XNOR U4526 ( .A(n4288), .B(n4319), .Z(n4289) );
  AND U4527 ( .A(n3144), .B(n2544), .Z(n4319) );
  AND U4528 ( .A(n4320), .B(g_input[0]), .Z(n4288) );
  NANDN U4529 ( .B(n2421), .A(n4321), .Z(n4320) );
  NAND U4530 ( .A(n3833), .B(n2544), .Z(n4321) );
  XOR U4531 ( .A(n4324), .B(n4325), .Z(n4300) );
  AND U4532 ( .A(n4327), .B(n4328), .Z(n4326) );
  NANDN U4533 ( .B(n714), .A(n4329), .Z(n4328) );
  OR U4534 ( .A(n4330), .B(n4331), .Z(n4327) );
  XNOR U4535 ( .A(n4333), .B(n4332), .Z(n3897) );
  XNOR U4536 ( .A(n4334), .B(n4330), .Z(n4333) );
  NAND U4537 ( .A(n744), .B(n4329), .Z(n4330) );
  NANDN U4538 ( .B(n714), .A(e_input[0]), .Z(n4335) );
  NANDN U4539 ( .B(n4336), .A(n4337), .Z(n714) );
  AND U4540 ( .A(n4338), .B(g_input[31]), .Z(n4337) );
  NAND U4541 ( .A(n818), .B(n2942), .Z(n3880) );
  XNOR U4542 ( .A(n3878), .B(n4342), .Z(n3879) );
  AND U4543 ( .A(n3074), .B(n778), .Z(n4342) );
  NAND U4544 ( .A(n855), .B(n2942), .Z(n4345) );
  XNOR U4545 ( .A(n4343), .B(n4347), .Z(n4344) );
  AND U4546 ( .A(n3074), .B(n818), .Z(n4347) );
  XNOR U4547 ( .A(n4339), .B(n4352), .Z(n4340) );
  AND U4548 ( .A(n744), .B(e_input[0]), .Z(n4352) );
  XNOR U4549 ( .A(n4338), .B(g_input[30]), .Z(n4336) );
  NOR U4550 ( .A(n4353), .B(n4354), .Z(n4338) );
  XOR U4551 ( .A(n4358), .B(n4341), .Z(n4351) );
  NAND U4552 ( .A(n778), .B(n4329), .Z(n4341) );
  IV U4553 ( .A(n4346), .Z(n4358) );
  NAND U4554 ( .A(n899), .B(n2942), .Z(n4350) );
  XNOR U4555 ( .A(n4348), .B(n4360), .Z(n4349) );
  AND U4556 ( .A(n3074), .B(n855), .Z(n4360) );
  XNOR U4557 ( .A(n4355), .B(n4365), .Z(n4356) );
  AND U4558 ( .A(n778), .B(e_input[0]), .Z(n4365) );
  XOR U4559 ( .A(n4353), .B(g_input[29]), .Z(n4354) );
  NANDN U4560 ( .B(n4366), .A(n4367), .Z(n4353) );
  XOR U4561 ( .A(n4371), .B(n4357), .Z(n4364) );
  NAND U4562 ( .A(n818), .B(n4329), .Z(n4357) );
  IV U4563 ( .A(n4359), .Z(n4371) );
  NAND U4564 ( .A(n945), .B(n2942), .Z(n4363) );
  XNOR U4565 ( .A(n4361), .B(n4373), .Z(n4362) );
  AND U4566 ( .A(n3074), .B(n899), .Z(n4373) );
  XNOR U4567 ( .A(n4368), .B(n4378), .Z(n4369) );
  AND U4568 ( .A(n818), .B(e_input[0]), .Z(n4378) );
  XNOR U4569 ( .A(n4367), .B(g_input[28]), .Z(n4366) );
  NOR U4570 ( .A(n4379), .B(n4380), .Z(n4367) );
  XOR U4571 ( .A(n4384), .B(n4370), .Z(n4377) );
  NAND U4572 ( .A(n855), .B(n4329), .Z(n4370) );
  IV U4573 ( .A(n4372), .Z(n4384) );
  NAND U4574 ( .A(n1003), .B(n2942), .Z(n4376) );
  XNOR U4575 ( .A(n4374), .B(n4386), .Z(n4375) );
  AND U4576 ( .A(n3074), .B(n945), .Z(n4386) );
  XNOR U4577 ( .A(n4381), .B(n4391), .Z(n4382) );
  AND U4578 ( .A(n855), .B(e_input[0]), .Z(n4391) );
  XOR U4579 ( .A(n4379), .B(g_input[27]), .Z(n4380) );
  NANDN U4580 ( .B(n4392), .A(n4393), .Z(n4379) );
  XOR U4581 ( .A(n4397), .B(n4383), .Z(n4390) );
  NAND U4582 ( .A(n899), .B(n4329), .Z(n4383) );
  IV U4583 ( .A(n4385), .Z(n4397) );
  NAND U4584 ( .A(n1057), .B(n2942), .Z(n4389) );
  XNOR U4585 ( .A(n4387), .B(n4399), .Z(n4388) );
  AND U4586 ( .A(n3074), .B(n1003), .Z(n4399) );
  XNOR U4587 ( .A(n4394), .B(n4404), .Z(n4395) );
  AND U4588 ( .A(n899), .B(e_input[0]), .Z(n4404) );
  XNOR U4589 ( .A(n4393), .B(g_input[26]), .Z(n4392) );
  NOR U4590 ( .A(n4405), .B(n4406), .Z(n4393) );
  XOR U4591 ( .A(n4410), .B(n4396), .Z(n4403) );
  NAND U4592 ( .A(n945), .B(n4329), .Z(n4396) );
  IV U4593 ( .A(n4398), .Z(n4410) );
  NAND U4594 ( .A(n1119), .B(n2942), .Z(n4402) );
  XNOR U4595 ( .A(n4400), .B(n4412), .Z(n4401) );
  AND U4596 ( .A(n3074), .B(n1057), .Z(n4412) );
  XNOR U4597 ( .A(n4407), .B(n4417), .Z(n4408) );
  AND U4598 ( .A(n945), .B(e_input[0]), .Z(n4417) );
  XOR U4599 ( .A(n4405), .B(g_input[25]), .Z(n4406) );
  NANDN U4600 ( .B(n4418), .A(n4419), .Z(n4405) );
  XOR U4601 ( .A(n4423), .B(n4409), .Z(n4416) );
  NAND U4602 ( .A(n1003), .B(n4329), .Z(n4409) );
  IV U4603 ( .A(n4411), .Z(n4423) );
  NAND U4604 ( .A(n1180), .B(n2942), .Z(n4415) );
  XNOR U4605 ( .A(n4413), .B(n4425), .Z(n4414) );
  AND U4606 ( .A(n3074), .B(n1119), .Z(n4425) );
  XNOR U4607 ( .A(n4420), .B(n4430), .Z(n4421) );
  AND U4608 ( .A(n1003), .B(e_input[0]), .Z(n4430) );
  XNOR U4609 ( .A(n4419), .B(g_input[24]), .Z(n4418) );
  NOR U4610 ( .A(n4431), .B(n4432), .Z(n4419) );
  XOR U4611 ( .A(n4436), .B(n4422), .Z(n4429) );
  NAND U4612 ( .A(n1057), .B(n4329), .Z(n4422) );
  IV U4613 ( .A(n4424), .Z(n4436) );
  NAND U4614 ( .A(n1246), .B(n2942), .Z(n4428) );
  XNOR U4615 ( .A(n4426), .B(n4438), .Z(n4427) );
  AND U4616 ( .A(n3074), .B(n1180), .Z(n4438) );
  XNOR U4617 ( .A(n4433), .B(n4443), .Z(n4434) );
  AND U4618 ( .A(n1057), .B(e_input[0]), .Z(n4443) );
  XOR U4619 ( .A(n4431), .B(g_input[23]), .Z(n4432) );
  NANDN U4620 ( .B(n4444), .A(n4445), .Z(n4431) );
  XOR U4621 ( .A(n4449), .B(n4435), .Z(n4442) );
  NAND U4622 ( .A(n1119), .B(n4329), .Z(n4435) );
  IV U4623 ( .A(n4437), .Z(n4449) );
  NAND U4624 ( .A(n1316), .B(n2942), .Z(n4441) );
  XNOR U4625 ( .A(n4439), .B(n4451), .Z(n4440) );
  AND U4626 ( .A(n3074), .B(n1246), .Z(n4451) );
  XNOR U4627 ( .A(n4446), .B(n4456), .Z(n4447) );
  AND U4628 ( .A(n1119), .B(e_input[0]), .Z(n4456) );
  XNOR U4629 ( .A(n4445), .B(g_input[22]), .Z(n4444) );
  NOR U4630 ( .A(n4457), .B(n4458), .Z(n4445) );
  XOR U4631 ( .A(n4462), .B(n4448), .Z(n4455) );
  NAND U4632 ( .A(n1180), .B(n4329), .Z(n4448) );
  IV U4633 ( .A(n4450), .Z(n4462) );
  NAND U4634 ( .A(n1388), .B(n2942), .Z(n4454) );
  XNOR U4635 ( .A(n4452), .B(n4464), .Z(n4453) );
  AND U4636 ( .A(n3074), .B(n1316), .Z(n4464) );
  XNOR U4637 ( .A(n4459), .B(n4469), .Z(n4460) );
  AND U4638 ( .A(n1180), .B(e_input[0]), .Z(n4469) );
  XOR U4639 ( .A(n4457), .B(g_input[21]), .Z(n4458) );
  NANDN U4640 ( .B(n4470), .A(n4471), .Z(n4457) );
  XOR U4641 ( .A(n4475), .B(n4461), .Z(n4468) );
  NAND U4642 ( .A(n1246), .B(n4329), .Z(n4461) );
  IV U4643 ( .A(n4463), .Z(n4475) );
  NAND U4644 ( .A(n1465), .B(n2942), .Z(n4467) );
  XNOR U4645 ( .A(n4465), .B(n4477), .Z(n4466) );
  AND U4646 ( .A(n3074), .B(n1388), .Z(n4477) );
  XNOR U4647 ( .A(n4472), .B(n4482), .Z(n4473) );
  AND U4648 ( .A(n1246), .B(e_input[0]), .Z(n4482) );
  XNOR U4649 ( .A(n4471), .B(g_input[20]), .Z(n4470) );
  NOR U4650 ( .A(n4483), .B(n4484), .Z(n4471) );
  XOR U4651 ( .A(n4488), .B(n4474), .Z(n4481) );
  NAND U4652 ( .A(n1316), .B(n4329), .Z(n4474) );
  IV U4653 ( .A(n4476), .Z(n4488) );
  NAND U4654 ( .A(n1550), .B(n2942), .Z(n4480) );
  XNOR U4655 ( .A(n4478), .B(n4490), .Z(n4479) );
  AND U4656 ( .A(n3074), .B(n1465), .Z(n4490) );
  XNOR U4657 ( .A(n4485), .B(n4495), .Z(n4486) );
  AND U4658 ( .A(n1316), .B(e_input[0]), .Z(n4495) );
  XOR U4659 ( .A(n4483), .B(g_input[19]), .Z(n4484) );
  NANDN U4660 ( .B(n4496), .A(n4497), .Z(n4483) );
  XOR U4661 ( .A(n4501), .B(n4487), .Z(n4494) );
  NAND U4662 ( .A(n1388), .B(n4329), .Z(n4487) );
  IV U4663 ( .A(n4489), .Z(n4501) );
  NAND U4664 ( .A(n1642), .B(n2942), .Z(n4493) );
  XNOR U4665 ( .A(n4491), .B(n4503), .Z(n4492) );
  AND U4666 ( .A(n3074), .B(n1550), .Z(n4503) );
  XNOR U4667 ( .A(n4498), .B(n4508), .Z(n4499) );
  AND U4668 ( .A(n1388), .B(e_input[0]), .Z(n4508) );
  XNOR U4669 ( .A(n4497), .B(g_input[18]), .Z(n4496) );
  NOR U4670 ( .A(n4509), .B(n4510), .Z(n4497) );
  XOR U4671 ( .A(n4514), .B(n4500), .Z(n4507) );
  NAND U4672 ( .A(n1465), .B(n4329), .Z(n4500) );
  IV U4673 ( .A(n4502), .Z(n4514) );
  NAND U4674 ( .A(n1737), .B(n2942), .Z(n4506) );
  XNOR U4675 ( .A(n4504), .B(n4516), .Z(n4505) );
  AND U4676 ( .A(n3074), .B(n1642), .Z(n4516) );
  XNOR U4677 ( .A(n4511), .B(n4521), .Z(n4512) );
  AND U4678 ( .A(n1465), .B(e_input[0]), .Z(n4521) );
  XOR U4679 ( .A(n4509), .B(g_input[17]), .Z(n4510) );
  NANDN U4680 ( .B(n4522), .A(n4523), .Z(n4509) );
  XOR U4681 ( .A(n4527), .B(n4513), .Z(n4520) );
  NAND U4682 ( .A(n1550), .B(n4329), .Z(n4513) );
  IV U4683 ( .A(n4515), .Z(n4527) );
  XOR U4684 ( .A(n4528), .B(n4529), .Z(n4515) );
  AND U4685 ( .A(n4139), .B(n4530), .Z(n4529) );
  XNOR U4686 ( .A(n4528), .B(n4138), .Z(n4530) );
  NAND U4687 ( .A(n1831), .B(n2942), .Z(n4519) );
  XNOR U4688 ( .A(n4517), .B(n4531), .Z(n4518) );
  AND U4689 ( .A(n3074), .B(n1737), .Z(n4531) );
  XNOR U4690 ( .A(n4524), .B(n4536), .Z(n4525) );
  AND U4691 ( .A(n1550), .B(e_input[0]), .Z(n4536) );
  XOR U4692 ( .A(n4540), .B(n4526), .Z(n4535) );
  NAND U4693 ( .A(n1642), .B(n4329), .Z(n4526) );
  IV U4694 ( .A(n4528), .Z(n4540) );
  NAND U4695 ( .A(n1931), .B(n2942), .Z(n4534) );
  XNOR U4696 ( .A(n4532), .B(n4542), .Z(n4533) );
  AND U4697 ( .A(n3074), .B(n1831), .Z(n4542) );
  XNOR U4698 ( .A(n4537), .B(n4547), .Z(n4538) );
  AND U4699 ( .A(n1642), .B(e_input[0]), .Z(n4547) );
  XOR U4700 ( .A(n4551), .B(n4539), .Z(n4546) );
  NAND U4701 ( .A(n1737), .B(n4329), .Z(n4539) );
  IV U4702 ( .A(n4541), .Z(n4551) );
  NAND U4703 ( .A(n2036), .B(n2942), .Z(n4545) );
  XNOR U4704 ( .A(n4543), .B(n4553), .Z(n4544) );
  AND U4705 ( .A(n3074), .B(n1931), .Z(n4553) );
  XNOR U4706 ( .A(n4548), .B(n4558), .Z(n4549) );
  AND U4707 ( .A(n1737), .B(e_input[0]), .Z(n4558) );
  XOR U4708 ( .A(n4562), .B(n4550), .Z(n4557) );
  NAND U4709 ( .A(n1831), .B(n4329), .Z(n4550) );
  IV U4710 ( .A(n4552), .Z(n4562) );
  NAND U4711 ( .A(n2141), .B(n2942), .Z(n4556) );
  XNOR U4712 ( .A(n4554), .B(n4564), .Z(n4555) );
  AND U4713 ( .A(n3074), .B(n2036), .Z(n4564) );
  XNOR U4714 ( .A(n4559), .B(n4569), .Z(n4560) );
  AND U4715 ( .A(n1831), .B(e_input[0]), .Z(n4569) );
  XOR U4716 ( .A(n4573), .B(n4561), .Z(n4568) );
  NAND U4717 ( .A(n1931), .B(n4329), .Z(n4561) );
  IV U4718 ( .A(n4563), .Z(n4573) );
  NAND U4719 ( .A(n2254), .B(n2942), .Z(n4567) );
  XNOR U4720 ( .A(n4565), .B(n4575), .Z(n4566) );
  AND U4721 ( .A(n3074), .B(n2141), .Z(n4575) );
  XNOR U4722 ( .A(n4570), .B(n4580), .Z(n4571) );
  AND U4723 ( .A(n1931), .B(e_input[0]), .Z(n4580) );
  XOR U4724 ( .A(n4584), .B(n4572), .Z(n4579) );
  NAND U4725 ( .A(n2036), .B(n4329), .Z(n4572) );
  IV U4726 ( .A(n4574), .Z(n4584) );
  NAND U4727 ( .A(n2370), .B(n2942), .Z(n4578) );
  XNOR U4728 ( .A(n4576), .B(n4586), .Z(n4577) );
  AND U4729 ( .A(n3074), .B(n2254), .Z(n4586) );
  XNOR U4730 ( .A(n4581), .B(n4591), .Z(n4582) );
  AND U4731 ( .A(n2036), .B(e_input[0]), .Z(n4591) );
  XOR U4732 ( .A(n4595), .B(n4583), .Z(n4590) );
  NAND U4733 ( .A(n2141), .B(n4329), .Z(n4583) );
  IV U4734 ( .A(n4585), .Z(n4595) );
  NAND U4735 ( .A(n2491), .B(n2942), .Z(n4589) );
  XNOR U4736 ( .A(n4587), .B(n4597), .Z(n4588) );
  AND U4737 ( .A(n3074), .B(n2370), .Z(n4597) );
  XNOR U4738 ( .A(n4592), .B(n4602), .Z(n4593) );
  AND U4739 ( .A(n2141), .B(e_input[0]), .Z(n4602) );
  XOR U4740 ( .A(n4606), .B(n4594), .Z(n4601) );
  NAND U4741 ( .A(n2254), .B(n4329), .Z(n4594) );
  IV U4742 ( .A(n4596), .Z(n4606) );
  NAND U4743 ( .A(n2613), .B(n2942), .Z(n4600) );
  XNOR U4744 ( .A(n4598), .B(n4608), .Z(n4599) );
  AND U4745 ( .A(n3074), .B(n2491), .Z(n4608) );
  XNOR U4746 ( .A(n4603), .B(n4613), .Z(n4604) );
  AND U4747 ( .A(n2254), .B(e_input[0]), .Z(n4613) );
  XOR U4748 ( .A(n4617), .B(n4605), .Z(n4612) );
  NAND U4749 ( .A(n2370), .B(n4329), .Z(n4605) );
  IV U4750 ( .A(n4607), .Z(n4617) );
  NAND U4751 ( .A(n2741), .B(n2942), .Z(n4611) );
  XNOR U4752 ( .A(n4609), .B(n4619), .Z(n4610) );
  AND U4753 ( .A(n3074), .B(n2613), .Z(n4619) );
  XNOR U4754 ( .A(n4623), .B(n4620), .Z(n4622) );
  XNOR U4755 ( .A(n4614), .B(n4625), .Z(n4615) );
  AND U4756 ( .A(n2370), .B(e_input[0]), .Z(n4625) );
  XNOR U4757 ( .A(n4629), .B(n4626), .Z(n4628) );
  XOR U4758 ( .A(n4630), .B(n4616), .Z(n4624) );
  NAND U4759 ( .A(n2491), .B(n4329), .Z(n4616) );
  IV U4760 ( .A(n4618), .Z(n4630) );
  XNOR U4761 ( .A(n4631), .B(n4632), .Z(n4618) );
  AND U4762 ( .A(n4633), .B(n4634), .Z(n4632) );
  XOR U4763 ( .A(n4627), .B(n4635), .Z(n4634) );
  XNOR U4764 ( .A(n4629), .B(n4631), .Z(n4635) );
  NAND U4765 ( .A(n2613), .B(n4329), .Z(n4629) );
  XOR U4766 ( .A(n4626), .B(n4636), .Z(n4627) );
  AND U4767 ( .A(n2491), .B(e_input[0]), .Z(n4636) );
  XNOR U4768 ( .A(n4640), .B(n4637), .Z(n4639) );
  XOR U4769 ( .A(n4621), .B(n4641), .Z(n4633) );
  XNOR U4770 ( .A(n4623), .B(n4631), .Z(n4641) );
  NANDN U4771 ( .B(n2870), .A(n2942), .Z(n4623) );
  XOR U4772 ( .A(n4620), .B(n4642), .Z(n4621) );
  AND U4773 ( .A(n3074), .B(n2741), .Z(n4642) );
  XNOR U4774 ( .A(n4646), .B(n4643), .Z(n4645) );
  XOR U4775 ( .A(n4647), .B(n4648), .Z(n4631) );
  AND U4776 ( .A(n4649), .B(n4650), .Z(n4648) );
  XOR U4777 ( .A(n4638), .B(n4651), .Z(n4650) );
  XNOR U4778 ( .A(n4640), .B(n4647), .Z(n4651) );
  NAND U4779 ( .A(n2741), .B(n4329), .Z(n4640) );
  XOR U4780 ( .A(n4637), .B(n4652), .Z(n4638) );
  AND U4781 ( .A(n2613), .B(e_input[0]), .Z(n4652) );
  XNOR U4782 ( .A(n4656), .B(n4653), .Z(n4655) );
  XOR U4783 ( .A(n4644), .B(n4657), .Z(n4649) );
  XNOR U4784 ( .A(n4646), .B(n4647), .Z(n4657) );
  NANDN U4785 ( .B(n3008), .A(n2942), .Z(n4646) );
  XOR U4786 ( .A(n4643), .B(n4658), .Z(n4644) );
  ANDN U4787 ( .A(n3074), .B(n2870), .Z(n4658) );
  XNOR U4788 ( .A(n4662), .B(n4659), .Z(n4661) );
  XOR U4789 ( .A(n4663), .B(n4664), .Z(n4647) );
  AND U4790 ( .A(n4665), .B(n4666), .Z(n4664) );
  XOR U4791 ( .A(n4654), .B(n4667), .Z(n4666) );
  XNOR U4792 ( .A(n4656), .B(n4663), .Z(n4667) );
  NANDN U4793 ( .B(n2870), .A(n4329), .Z(n4656) );
  XOR U4794 ( .A(n4653), .B(n4668), .Z(n4654) );
  AND U4795 ( .A(n2741), .B(e_input[0]), .Z(n4668) );
  XOR U4796 ( .A(n4660), .B(n4672), .Z(n4665) );
  XNOR U4797 ( .A(n4662), .B(n4663), .Z(n4672) );
  NAND U4798 ( .A(n2942), .B(n3144), .Z(n4662) );
  XOR U4799 ( .A(n4659), .B(n4673), .Z(n4660) );
  ANDN U4800 ( .A(n3074), .B(n3008), .Z(n4673) );
  NAND U4801 ( .A(n2942), .B(n3833), .Z(n4676) );
  XNOR U4802 ( .A(n4674), .B(n4678), .Z(n4675) );
  AND U4803 ( .A(n3144), .B(n3074), .Z(n4678) );
  AND U4804 ( .A(n4679), .B(g_input[0]), .Z(n4674) );
  NANDN U4805 ( .B(n2942), .A(n4680), .Z(n4679) );
  NAND U4806 ( .A(n3833), .B(n3074), .Z(n4680) );
  XNOR U4807 ( .A(n4669), .B(n4684), .Z(n4670) );
  ANDN U4808 ( .A(e_input[0]), .B(n2870), .Z(n4684) );
  XOR U4809 ( .A(n4687), .B(n4685), .Z(n4686) );
  ANDN U4810 ( .A(e_input[0]), .B(n3008), .Z(n4687) );
  AND U4811 ( .A(n4329), .B(n3144), .Z(n4688) );
  XOR U4812 ( .A(n4692), .B(n4671), .Z(n4683) );
  NANDN U4813 ( .B(n3008), .A(n4329), .Z(n4671) );
  IV U4814 ( .A(n4677), .Z(n4692) );
  NAND U4815 ( .A(n4329), .B(n3833), .Z(n4691) );
  XNOR U4816 ( .A(n4689), .B(n4693), .Z(n4690) );
  AND U4817 ( .A(n3144), .B(e_input[0]), .Z(n4693) );
  AND U4818 ( .A(n4694), .B(g_input[0]), .Z(n4689) );
  NANDN U4819 ( .B(n4329), .A(n4695), .Z(n4694) );
  NAND U4820 ( .A(n3833), .B(e_input[0]), .Z(n4695) );
  XNOR U4821 ( .A(n4697), .B(n3108), .Z(n3099) );
  XNOR U4822 ( .A(n3087), .B(n4699), .Z(n3088) );
  AND U4823 ( .A(n1931), .B(n1198), .Z(n4699) );
  XOR U4824 ( .A(n4703), .B(n3089), .Z(n4698) );
  NAND U4825 ( .A(n1140), .B(n2036), .Z(n3089) );
  IV U4826 ( .A(n3091), .Z(n4703) );
  XNOR U4827 ( .A(n3096), .B(n3097), .Z(n3093) );
  NANDN U4828 ( .B(n1022), .A(n2254), .Z(n3097) );
  XNOR U4829 ( .A(n3095), .B(n4707), .Z(n3096) );
  AND U4830 ( .A(n2141), .B(n1082), .Z(n4707) );
  XNOR U4831 ( .A(n3107), .B(n3098), .Z(n4697) );
  XOR U4832 ( .A(n4711), .B(n4712), .Z(n3098) );
  XOR U4833 ( .A(n4713), .B(n3117), .Z(n3107) );
  XNOR U4834 ( .A(n3104), .B(n3105), .Z(n3117) );
  NAND U4835 ( .A(n1284), .B(n1831), .Z(n3105) );
  XNOR U4836 ( .A(n3103), .B(n4714), .Z(n3104) );
  AND U4837 ( .A(n1737), .B(n1352), .Z(n4714) );
  XNOR U4838 ( .A(n3116), .B(n3106), .Z(n4713) );
  XOR U4839 ( .A(n4718), .B(n4719), .Z(n3106) );
  AND U4840 ( .A(n4720), .B(n4721), .Z(n4719) );
  XOR U4841 ( .A(n4722), .B(n4723), .Z(n4721) );
  XOR U4842 ( .A(n4718), .B(n4724), .Z(n4723) );
  XOR U4843 ( .A(n4705), .B(n4725), .Z(n4720) );
  XOR U4844 ( .A(n4718), .B(n4706), .Z(n4725) );
  NANDN U4845 ( .B(n1022), .A(n2370), .Z(n4710) );
  XNOR U4846 ( .A(n4708), .B(n4726), .Z(n4709) );
  AND U4847 ( .A(n2254), .B(n1082), .Z(n4726) );
  XNOR U4848 ( .A(n4700), .B(n4731), .Z(n4701) );
  AND U4849 ( .A(n2036), .B(n1198), .Z(n4731) );
  XOR U4850 ( .A(n4735), .B(n4702), .Z(n4730) );
  NAND U4851 ( .A(n1140), .B(n2141), .Z(n4702) );
  IV U4852 ( .A(n4704), .Z(n4735) );
  XOR U4853 ( .A(n4739), .B(n4740), .Z(n4718) );
  AND U4854 ( .A(n4741), .B(n4742), .Z(n4740) );
  XOR U4855 ( .A(n4743), .B(n4744), .Z(n4742) );
  XOR U4856 ( .A(n4739), .B(n4745), .Z(n4744) );
  XOR U4857 ( .A(n4737), .B(n4746), .Z(n4741) );
  XOR U4858 ( .A(n4739), .B(n4738), .Z(n4746) );
  NANDN U4859 ( .B(n1022), .A(n2491), .Z(n4729) );
  XNOR U4860 ( .A(n4727), .B(n4747), .Z(n4728) );
  AND U4861 ( .A(n2370), .B(n1082), .Z(n4747) );
  XNOR U4862 ( .A(n4732), .B(n4752), .Z(n4733) );
  AND U4863 ( .A(n2141), .B(n1198), .Z(n4752) );
  XOR U4864 ( .A(n4756), .B(n4734), .Z(n4751) );
  NAND U4865 ( .A(n1140), .B(n2254), .Z(n4734) );
  IV U4866 ( .A(n4736), .Z(n4756) );
  XOR U4867 ( .A(n4760), .B(n4761), .Z(n4739) );
  AND U4868 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR U4869 ( .A(n4764), .B(n4765), .Z(n4763) );
  XOR U4870 ( .A(n4760), .B(n4766), .Z(n4765) );
  XOR U4871 ( .A(n4758), .B(n4767), .Z(n4762) );
  XOR U4872 ( .A(n4760), .B(n4759), .Z(n4767) );
  NANDN U4873 ( .B(n1022), .A(n2613), .Z(n4750) );
  XNOR U4874 ( .A(n4748), .B(n4768), .Z(n4749) );
  AND U4875 ( .A(n2491), .B(n1082), .Z(n4768) );
  XNOR U4876 ( .A(n4753), .B(n4773), .Z(n4754) );
  AND U4877 ( .A(n2254), .B(n1198), .Z(n4773) );
  XOR U4878 ( .A(n4777), .B(n4755), .Z(n4772) );
  NAND U4879 ( .A(n1140), .B(n2370), .Z(n4755) );
  IV U4880 ( .A(n4757), .Z(n4777) );
  XOR U4881 ( .A(n4781), .B(n4782), .Z(n4760) );
  AND U4882 ( .A(n4783), .B(n4784), .Z(n4782) );
  XOR U4883 ( .A(n4785), .B(n4786), .Z(n4784) );
  XOR U4884 ( .A(n4781), .B(n4787), .Z(n4786) );
  XOR U4885 ( .A(n4779), .B(n4788), .Z(n4783) );
  XOR U4886 ( .A(n4781), .B(n4780), .Z(n4788) );
  NANDN U4887 ( .B(n1022), .A(n2741), .Z(n4771) );
  XNOR U4888 ( .A(n4769), .B(n4789), .Z(n4770) );
  AND U4889 ( .A(n2613), .B(n1082), .Z(n4789) );
  XNOR U4890 ( .A(n4774), .B(n4794), .Z(n4775) );
  AND U4891 ( .A(n2370), .B(n1198), .Z(n4794) );
  XOR U4892 ( .A(n4798), .B(n4776), .Z(n4793) );
  NAND U4893 ( .A(n1140), .B(n2491), .Z(n4776) );
  IV U4894 ( .A(n4778), .Z(n4798) );
  XOR U4895 ( .A(n4802), .B(n4803), .Z(n4781) );
  AND U4896 ( .A(n4804), .B(n4805), .Z(n4803) );
  XOR U4897 ( .A(n4806), .B(n4807), .Z(n4805) );
  XOR U4898 ( .A(n4802), .B(n4808), .Z(n4807) );
  XOR U4899 ( .A(n4800), .B(n4809), .Z(n4804) );
  XOR U4900 ( .A(n4802), .B(n4801), .Z(n4809) );
  OR U4901 ( .A(n1022), .B(n2870), .Z(n4792) );
  XNOR U4902 ( .A(n4790), .B(n4810), .Z(n4791) );
  AND U4903 ( .A(n2741), .B(n1082), .Z(n4810) );
  XNOR U4904 ( .A(n4795), .B(n4815), .Z(n4796) );
  AND U4905 ( .A(n2491), .B(n1198), .Z(n4815) );
  XOR U4906 ( .A(n4819), .B(n4797), .Z(n4814) );
  NAND U4907 ( .A(n1140), .B(n2613), .Z(n4797) );
  IV U4908 ( .A(n4799), .Z(n4819) );
  XOR U4909 ( .A(n4823), .B(n4824), .Z(n4802) );
  AND U4910 ( .A(n4825), .B(n4826), .Z(n4824) );
  XOR U4911 ( .A(n4827), .B(n4828), .Z(n4826) );
  XOR U4912 ( .A(n4823), .B(n4829), .Z(n4828) );
  XOR U4913 ( .A(n4821), .B(n4830), .Z(n4825) );
  XOR U4914 ( .A(n4823), .B(n4822), .Z(n4830) );
  OR U4915 ( .A(n1022), .B(n3008), .Z(n4813) );
  XNOR U4916 ( .A(n4811), .B(n4831), .Z(n4812) );
  ANDN U4917 ( .A(n1082), .B(n2870), .Z(n4831) );
  XNOR U4918 ( .A(n4816), .B(n4836), .Z(n4817) );
  AND U4919 ( .A(n2613), .B(n1198), .Z(n4836) );
  XOR U4920 ( .A(n4840), .B(n4818), .Z(n4835) );
  NAND U4921 ( .A(n1140), .B(n2741), .Z(n4818) );
  IV U4922 ( .A(n4820), .Z(n4840) );
  XOR U4923 ( .A(n4844), .B(n4845), .Z(n4823) );
  AND U4924 ( .A(n4846), .B(n4847), .Z(n4845) );
  XOR U4925 ( .A(n4848), .B(n4849), .Z(n4847) );
  XOR U4926 ( .A(n4844), .B(n4850), .Z(n4849) );
  XOR U4927 ( .A(n4842), .B(n4851), .Z(n4846) );
  XOR U4928 ( .A(n4844), .B(n4843), .Z(n4851) );
  NANDN U4929 ( .B(n1022), .A(n3144), .Z(n4834) );
  XNOR U4930 ( .A(n4832), .B(n4852), .Z(n4833) );
  ANDN U4931 ( .A(n1082), .B(n3008), .Z(n4852) );
  XNOR U4932 ( .A(n4837), .B(n4857), .Z(n4838) );
  AND U4933 ( .A(n2741), .B(n1198), .Z(n4857) );
  XOR U4934 ( .A(n4861), .B(n4839), .Z(n4856) );
  NANDN U4935 ( .B(n2870), .A(n1140), .Z(n4839) );
  IV U4936 ( .A(n4841), .Z(n4861) );
  XOR U4937 ( .A(n4866), .B(n4867), .Z(n4712) );
  XNOR U4938 ( .A(n4868), .B(n4865), .Z(n4866) );
  XNOR U4939 ( .A(n4858), .B(n4870), .Z(n4859) );
  ANDN U4940 ( .A(n1198), .B(n2870), .Z(n4870) );
  XOR U4941 ( .A(n4873), .B(n4871), .Z(n4872) );
  ANDN U4942 ( .A(n1198), .B(n3008), .Z(n4873) );
  AND U4943 ( .A(n3144), .B(n1140), .Z(n4874) );
  XOR U4944 ( .A(n4878), .B(n4860), .Z(n4869) );
  NANDN U4945 ( .B(n3008), .A(n1140), .Z(n4860) );
  IV U4946 ( .A(n4862), .Z(n4878) );
  NAND U4947 ( .A(n1140), .B(n3833), .Z(n4877) );
  XNOR U4948 ( .A(n4875), .B(n4879), .Z(n4876) );
  AND U4949 ( .A(n3144), .B(n1198), .Z(n4879) );
  AND U4950 ( .A(n4880), .B(g_input[0]), .Z(n4875) );
  NANDN U4951 ( .B(n1140), .A(n4881), .Z(n4880) );
  NAND U4952 ( .A(n3833), .B(n1198), .Z(n4881) );
  XNOR U4953 ( .A(n4854), .B(n4855), .Z(n4864) );
  NANDN U4954 ( .B(n1022), .A(n3833), .Z(n4855) );
  XNOR U4955 ( .A(n4853), .B(n4884), .Z(n4854) );
  AND U4956 ( .A(n3144), .B(n1082), .Z(n4884) );
  AND U4957 ( .A(n4885), .B(g_input[0]), .Z(n4853) );
  NAND U4958 ( .A(n4886), .B(n1022), .Z(n4885) );
  NAND U4959 ( .A(n3833), .B(n1082), .Z(n4886) );
  XOR U4960 ( .A(n4889), .B(n4890), .Z(n4865) );
  XNOR U4961 ( .A(n3111), .B(n4892), .Z(n3112) );
  AND U4962 ( .A(n1550), .B(n1520), .Z(n4892) );
  XNOR U4963 ( .A(n4523), .B(g_input[16]), .Z(n4522) );
  NOR U4964 ( .A(n4893), .B(n4894), .Z(n4523) );
  XOR U4965 ( .A(n4898), .B(n3113), .Z(n4891) );
  NAND U4966 ( .A(n1433), .B(n1642), .Z(n3113) );
  IV U4967 ( .A(n3115), .Z(n4898) );
  NAND U4968 ( .A(n1284), .B(n1931), .Z(n4717) );
  XNOR U4969 ( .A(n4715), .B(n4900), .Z(n4716) );
  AND U4970 ( .A(n1831), .B(n1352), .Z(n4900) );
  XNOR U4971 ( .A(n4895), .B(n4905), .Z(n4896) );
  AND U4972 ( .A(n1642), .B(n1520), .Z(n4905) );
  XOR U4973 ( .A(n4893), .B(g_input[15]), .Z(n4894) );
  NANDN U4974 ( .B(n4906), .A(n4907), .Z(n4893) );
  XOR U4975 ( .A(n4911), .B(n4897), .Z(n4904) );
  NAND U4976 ( .A(n1433), .B(n1737), .Z(n4897) );
  IV U4977 ( .A(n4899), .Z(n4911) );
  NAND U4978 ( .A(n1284), .B(n2036), .Z(n4903) );
  XNOR U4979 ( .A(n4901), .B(n4913), .Z(n4902) );
  AND U4980 ( .A(n1931), .B(n1352), .Z(n4913) );
  XNOR U4981 ( .A(n4908), .B(n4918), .Z(n4909) );
  AND U4982 ( .A(n1737), .B(n1520), .Z(n4918) );
  XNOR U4983 ( .A(n4907), .B(g_input[14]), .Z(n4906) );
  NOR U4984 ( .A(n4919), .B(n4920), .Z(n4907) );
  XOR U4985 ( .A(n4924), .B(n4910), .Z(n4917) );
  NAND U4986 ( .A(n1433), .B(n1831), .Z(n4910) );
  IV U4987 ( .A(n4912), .Z(n4924) );
  NAND U4988 ( .A(n1284), .B(n2141), .Z(n4916) );
  XNOR U4989 ( .A(n4914), .B(n4926), .Z(n4915) );
  AND U4990 ( .A(n2036), .B(n1352), .Z(n4926) );
  XNOR U4991 ( .A(n4921), .B(n4931), .Z(n4922) );
  AND U4992 ( .A(n1831), .B(n1520), .Z(n4931) );
  XOR U4993 ( .A(n4919), .B(g_input[13]), .Z(n4920) );
  NANDN U4994 ( .B(n4932), .A(n4933), .Z(n4919) );
  XOR U4995 ( .A(n4937), .B(n4923), .Z(n4930) );
  NAND U4996 ( .A(n1433), .B(n1931), .Z(n4923) );
  IV U4997 ( .A(n4925), .Z(n4937) );
  NAND U4998 ( .A(n1284), .B(n2254), .Z(n4929) );
  XNOR U4999 ( .A(n4927), .B(n4939), .Z(n4928) );
  AND U5000 ( .A(n2141), .B(n1352), .Z(n4939) );
  XNOR U5001 ( .A(n4934), .B(n4944), .Z(n4935) );
  AND U5002 ( .A(n1931), .B(n1520), .Z(n4944) );
  XNOR U5003 ( .A(n4933), .B(g_input[12]), .Z(n4932) );
  NOR U5004 ( .A(n4945), .B(n4946), .Z(n4933) );
  XOR U5005 ( .A(n4950), .B(n4936), .Z(n4943) );
  NAND U5006 ( .A(n1433), .B(n2036), .Z(n4936) );
  IV U5007 ( .A(n4938), .Z(n4950) );
  NAND U5008 ( .A(n1284), .B(n2370), .Z(n4942) );
  XNOR U5009 ( .A(n4940), .B(n4952), .Z(n4941) );
  AND U5010 ( .A(n2254), .B(n1352), .Z(n4952) );
  XNOR U5011 ( .A(n4947), .B(n4957), .Z(n4948) );
  AND U5012 ( .A(n2036), .B(n1520), .Z(n4957) );
  XOR U5013 ( .A(n4945), .B(g_input[11]), .Z(n4946) );
  NANDN U5014 ( .B(n4958), .A(n4959), .Z(n4945) );
  XOR U5015 ( .A(n4963), .B(n4949), .Z(n4956) );
  NAND U5016 ( .A(n1433), .B(n2141), .Z(n4949) );
  IV U5017 ( .A(n4951), .Z(n4963) );
  NAND U5018 ( .A(n1284), .B(n2491), .Z(n4955) );
  XNOR U5019 ( .A(n4953), .B(n4965), .Z(n4954) );
  AND U5020 ( .A(n2370), .B(n1352), .Z(n4965) );
  XNOR U5021 ( .A(n4960), .B(n4970), .Z(n4961) );
  AND U5022 ( .A(n2141), .B(n1520), .Z(n4970) );
  XNOR U5023 ( .A(n4959), .B(g_input[10]), .Z(n4958) );
  NOR U5024 ( .A(n4971), .B(n4972), .Z(n4959) );
  XOR U5025 ( .A(n4976), .B(n4962), .Z(n4969) );
  NAND U5026 ( .A(n1433), .B(n2254), .Z(n4962) );
  IV U5027 ( .A(n4964), .Z(n4976) );
  NAND U5028 ( .A(n1284), .B(n2613), .Z(n4968) );
  XNOR U5029 ( .A(n4966), .B(n4978), .Z(n4967) );
  AND U5030 ( .A(n2491), .B(n1352), .Z(n4978) );
  XNOR U5031 ( .A(n4973), .B(n4983), .Z(n4974) );
  AND U5032 ( .A(n2254), .B(n1520), .Z(n4983) );
  XOR U5033 ( .A(n4971), .B(g_input[9]), .Z(n4972) );
  NANDN U5034 ( .B(n4984), .A(n4985), .Z(n4971) );
  XOR U5035 ( .A(n4989), .B(n4975), .Z(n4982) );
  NAND U5036 ( .A(n1433), .B(n2370), .Z(n4975) );
  IV U5037 ( .A(n4977), .Z(n4989) );
  NAND U5038 ( .A(n1284), .B(n2741), .Z(n4981) );
  XNOR U5039 ( .A(n4979), .B(n4991), .Z(n4980) );
  AND U5040 ( .A(n2613), .B(n1352), .Z(n4991) );
  XNOR U5041 ( .A(n4995), .B(n4992), .Z(n4994) );
  XNOR U5042 ( .A(n4986), .B(n4997), .Z(n4987) );
  AND U5043 ( .A(n2370), .B(n1520), .Z(n4997) );
  XNOR U5044 ( .A(n5001), .B(n4998), .Z(n5000) );
  XOR U5045 ( .A(n5002), .B(n4988), .Z(n4996) );
  NAND U5046 ( .A(n1433), .B(n2491), .Z(n4988) );
  IV U5047 ( .A(n4990), .Z(n5002) );
  XNOR U5048 ( .A(n5003), .B(n5004), .Z(n4990) );
  AND U5049 ( .A(n5005), .B(n5006), .Z(n5004) );
  XOR U5050 ( .A(n4999), .B(n5007), .Z(n5006) );
  XNOR U5051 ( .A(n5001), .B(n5003), .Z(n5007) );
  NAND U5052 ( .A(n1433), .B(n2613), .Z(n5001) );
  XOR U5053 ( .A(n4998), .B(n5008), .Z(n4999) );
  AND U5054 ( .A(n2491), .B(n1520), .Z(n5008) );
  XNOR U5055 ( .A(n5012), .B(n5009), .Z(n5011) );
  XOR U5056 ( .A(n4993), .B(n5013), .Z(n5005) );
  XNOR U5057 ( .A(n4995), .B(n5003), .Z(n5013) );
  NANDN U5058 ( .B(n2870), .A(n1284), .Z(n4995) );
  XOR U5059 ( .A(n4992), .B(n5014), .Z(n4993) );
  AND U5060 ( .A(n2741), .B(n1352), .Z(n5014) );
  XNOR U5061 ( .A(n5018), .B(n5015), .Z(n5017) );
  XOR U5062 ( .A(n5019), .B(n5020), .Z(n5003) );
  AND U5063 ( .A(n5021), .B(n5022), .Z(n5020) );
  XOR U5064 ( .A(n5010), .B(n5023), .Z(n5022) );
  XNOR U5065 ( .A(n5012), .B(n5019), .Z(n5023) );
  NAND U5066 ( .A(n1433), .B(n2741), .Z(n5012) );
  XOR U5067 ( .A(n5009), .B(n5024), .Z(n5010) );
  AND U5068 ( .A(n2613), .B(n1520), .Z(n5024) );
  XNOR U5069 ( .A(n5028), .B(n5025), .Z(n5027) );
  XOR U5070 ( .A(n5016), .B(n5029), .Z(n5021) );
  XNOR U5071 ( .A(n5018), .B(n5019), .Z(n5029) );
  NANDN U5072 ( .B(n3008), .A(n1284), .Z(n5018) );
  XOR U5073 ( .A(n5015), .B(n5030), .Z(n5016) );
  ANDN U5074 ( .A(n1352), .B(n2870), .Z(n5030) );
  XNOR U5075 ( .A(n5034), .B(n5031), .Z(n5033) );
  XOR U5076 ( .A(n5035), .B(n5036), .Z(n5019) );
  AND U5077 ( .A(n5037), .B(n5038), .Z(n5036) );
  XOR U5078 ( .A(n5026), .B(n5039), .Z(n5038) );
  XNOR U5079 ( .A(n5028), .B(n5035), .Z(n5039) );
  NANDN U5080 ( .B(n2870), .A(n1433), .Z(n5028) );
  XOR U5081 ( .A(n5025), .B(n5040), .Z(n5026) );
  AND U5082 ( .A(n2741), .B(n1520), .Z(n5040) );
  XOR U5083 ( .A(n5032), .B(n5044), .Z(n5037) );
  XNOR U5084 ( .A(n5034), .B(n5035), .Z(n5044) );
  NAND U5085 ( .A(n1284), .B(n3144), .Z(n5034) );
  XOR U5086 ( .A(n5031), .B(n5045), .Z(n5032) );
  ANDN U5087 ( .A(n1352), .B(n3008), .Z(n5045) );
  NAND U5088 ( .A(n1284), .B(n3833), .Z(n5048) );
  XNOR U5089 ( .A(n5046), .B(n5050), .Z(n5047) );
  AND U5090 ( .A(n3144), .B(n1352), .Z(n5050) );
  AND U5091 ( .A(n5051), .B(g_input[0]), .Z(n5046) );
  NANDN U5092 ( .B(n1284), .A(n5052), .Z(n5051) );
  NAND U5093 ( .A(n3833), .B(n1352), .Z(n5052) );
  XNOR U5094 ( .A(n5041), .B(n5056), .Z(n5042) );
  ANDN U5095 ( .A(n1520), .B(n2870), .Z(n5056) );
  XOR U5096 ( .A(n5059), .B(n5057), .Z(n5058) );
  ANDN U5097 ( .A(n1520), .B(n3008), .Z(n5059) );
  AND U5098 ( .A(n3144), .B(n1433), .Z(n5060) );
  XOR U5099 ( .A(n5064), .B(n5043), .Z(n5055) );
  NANDN U5100 ( .B(n3008), .A(n1433), .Z(n5043) );
  IV U5101 ( .A(n5049), .Z(n5064) );
  NAND U5102 ( .A(n1433), .B(n3833), .Z(n5063) );
  XNOR U5103 ( .A(n5061), .B(n5065), .Z(n5062) );
  AND U5104 ( .A(n3144), .B(n1520), .Z(n5065) );
  AND U5105 ( .A(n5066), .B(g_input[0]), .Z(n5061) );
  NANDN U5106 ( .B(n1433), .A(n5067), .Z(n5066) );
  NAND U5107 ( .A(n3833), .B(n1520), .Z(n5067) );
  XNOR U5108 ( .A(n5070), .B(n3134), .Z(n3124) );
  XNOR U5109 ( .A(n3121), .B(n3122), .Z(n3134) );
  NANDN U5110 ( .B(n836), .A(n2741), .Z(n3122) );
  XNOR U5111 ( .A(n3120), .B(n5071), .Z(n3121) );
  AND U5112 ( .A(n2613), .B(n874), .Z(n5071) );
  XNOR U5113 ( .A(n5075), .B(n5072), .Z(n5074) );
  XNOR U5114 ( .A(n3133), .B(n3123), .Z(n5070) );
  XOR U5115 ( .A(n5076), .B(n5077), .Z(n3123) );
  XNOR U5116 ( .A(n3128), .B(n5079), .Z(n3129) );
  AND U5117 ( .A(n2370), .B(n986), .Z(n5079) );
  XNOR U5118 ( .A(n4985), .B(g_input[8]), .Z(n4984) );
  NOR U5119 ( .A(n5080), .B(n5081), .Z(n4985) );
  XNOR U5120 ( .A(n5085), .B(n5082), .Z(n5084) );
  XOR U5121 ( .A(n5086), .B(n3130), .Z(n5078) );
  NAND U5122 ( .A(n932), .B(n2491), .Z(n3130) );
  IV U5123 ( .A(n3132), .Z(n5086) );
  XNOR U5124 ( .A(n5087), .B(n5088), .Z(n3132) );
  AND U5125 ( .A(n5089), .B(n5090), .Z(n5088) );
  XOR U5126 ( .A(n5083), .B(n5091), .Z(n5090) );
  XNOR U5127 ( .A(n5085), .B(n5087), .Z(n5091) );
  NAND U5128 ( .A(n932), .B(n2613), .Z(n5085) );
  XOR U5129 ( .A(n5082), .B(n5092), .Z(n5083) );
  AND U5130 ( .A(n2491), .B(n986), .Z(n5092) );
  XOR U5131 ( .A(n5080), .B(g_input[7]), .Z(n5081) );
  NANDN U5132 ( .B(n5093), .A(n5094), .Z(n5080) );
  XNOR U5133 ( .A(n5098), .B(n5095), .Z(n5097) );
  XOR U5134 ( .A(n5073), .B(n5099), .Z(n5089) );
  XNOR U5135 ( .A(n5075), .B(n5087), .Z(n5099) );
  OR U5136 ( .A(n836), .B(n2870), .Z(n5075) );
  XOR U5137 ( .A(n5072), .B(n5100), .Z(n5073) );
  AND U5138 ( .A(n2741), .B(n874), .Z(n5100) );
  XNOR U5139 ( .A(n5104), .B(n5101), .Z(n5103) );
  XOR U5140 ( .A(n5105), .B(n5106), .Z(n5087) );
  AND U5141 ( .A(n5107), .B(n5108), .Z(n5106) );
  XOR U5142 ( .A(n5096), .B(n5109), .Z(n5108) );
  XNOR U5143 ( .A(n5098), .B(n5105), .Z(n5109) );
  NAND U5144 ( .A(n932), .B(n2741), .Z(n5098) );
  XOR U5145 ( .A(n5095), .B(n5110), .Z(n5096) );
  AND U5146 ( .A(n2613), .B(n986), .Z(n5110) );
  XNOR U5147 ( .A(n5094), .B(g_input[6]), .Z(n5093) );
  NOR U5148 ( .A(n5111), .B(n5112), .Z(n5094) );
  XNOR U5149 ( .A(n5116), .B(n5113), .Z(n5115) );
  XOR U5150 ( .A(n5102), .B(n5117), .Z(n5107) );
  XNOR U5151 ( .A(n5104), .B(n5105), .Z(n5117) );
  OR U5152 ( .A(n836), .B(n3008), .Z(n5104) );
  XOR U5153 ( .A(n5101), .B(n5118), .Z(n5102) );
  ANDN U5154 ( .A(n874), .B(n2870), .Z(n5118) );
  XNOR U5155 ( .A(n5122), .B(n5119), .Z(n5121) );
  XOR U5156 ( .A(n5123), .B(n5124), .Z(n5105) );
  AND U5157 ( .A(n5125), .B(n5126), .Z(n5124) );
  XOR U5158 ( .A(n5114), .B(n5127), .Z(n5126) );
  XNOR U5159 ( .A(n5116), .B(n5123), .Z(n5127) );
  NANDN U5160 ( .B(n2870), .A(n932), .Z(n5116) );
  XOR U5161 ( .A(n5113), .B(n5128), .Z(n5114) );
  AND U5162 ( .A(n2741), .B(n986), .Z(n5128) );
  XOR U5163 ( .A(n5111), .B(g_input[5]), .Z(n5112) );
  NANDN U5164 ( .B(n5129), .A(n5130), .Z(n5111) );
  XOR U5165 ( .A(n5120), .B(n5134), .Z(n5125) );
  XNOR U5166 ( .A(n5122), .B(n5123), .Z(n5134) );
  NANDN U5167 ( .B(n836), .A(n3144), .Z(n5122) );
  XOR U5168 ( .A(n5119), .B(n5135), .Z(n5120) );
  ANDN U5169 ( .A(n874), .B(n3008), .Z(n5135) );
  NANDN U5170 ( .B(n836), .A(n3833), .Z(n5138) );
  XNOR U5171 ( .A(n5136), .B(n5140), .Z(n5137) );
  AND U5172 ( .A(n3144), .B(n874), .Z(n5140) );
  AND U5173 ( .A(n5141), .B(g_input[0]), .Z(n5136) );
  NAND U5174 ( .A(n5142), .B(n836), .Z(n5141) );
  NAND U5175 ( .A(n3833), .B(n874), .Z(n5142) );
  XNOR U5176 ( .A(n5131), .B(n5146), .Z(n5132) );
  ANDN U5177 ( .A(n986), .B(n2870), .Z(n5146) );
  XOR U5178 ( .A(n5149), .B(n5147), .Z(n5148) );
  ANDN U5179 ( .A(n986), .B(n3008), .Z(n5149) );
  AND U5180 ( .A(n3144), .B(n932), .Z(n5150) );
  XOR U5181 ( .A(n5154), .B(n5133), .Z(n5145) );
  NANDN U5182 ( .B(n3008), .A(n932), .Z(n5133) );
  IV U5183 ( .A(n5139), .Z(n5154) );
  NAND U5184 ( .A(n932), .B(n3833), .Z(n5153) );
  XNOR U5185 ( .A(n5151), .B(n5155), .Z(n5152) );
  AND U5186 ( .A(n3144), .B(n986), .Z(n5155) );
  AND U5187 ( .A(n5156), .B(g_input[0]), .Z(n5151) );
  NANDN U5188 ( .B(n932), .A(n5157), .Z(n5156) );
  NAND U5189 ( .A(n3833), .B(n986), .Z(n5157) );
  XNOR U5190 ( .A(n3137), .B(n5161), .Z(n3138) );
  ANDN U5191 ( .A(n810), .B(n2870), .Z(n5161) );
  XNOR U5192 ( .A(n5130), .B(g_input[4]), .Z(n5129) );
  NOR U5193 ( .A(n5162), .B(n5163), .Z(n5130) );
  XOR U5194 ( .A(n5166), .B(n5164), .Z(n5165) );
  ANDN U5195 ( .A(n810), .B(n3008), .Z(n5166) );
  AND U5196 ( .A(n3144), .B(n774), .Z(n5167) );
  XOR U5197 ( .A(n5171), .B(n3139), .Z(n5160) );
  NANDN U5198 ( .B(n3008), .A(n774), .Z(n3139) );
  NANDN U5199 ( .B(n5172), .A(n5173), .Z(n5162) );
  IV U5200 ( .A(n3141), .Z(n5171) );
  NAND U5201 ( .A(n774), .B(n3833), .Z(n5170) );
  XNOR U5202 ( .A(n5168), .B(n5174), .Z(n5169) );
  AND U5203 ( .A(n3144), .B(n810), .Z(n5174) );
  AND U5204 ( .A(n5175), .B(g_input[0]), .Z(n5168) );
  NANDN U5205 ( .B(n774), .A(n5176), .Z(n5175) );
  NAND U5206 ( .A(n3833), .B(n810), .Z(n5176) );
  XNOR U5207 ( .A(n3148), .B(n3149), .Z(n3143) );
  NANDN U5208 ( .B(n713), .A(n3833), .Z(n3149) );
  XNOR U5209 ( .A(n3147), .B(n5179), .Z(n3148) );
  AND U5210 ( .A(n3144), .B(n746), .Z(n5179) );
  XNOR U5211 ( .A(n5173), .B(g_input[2]), .Z(n5172) );
  AND U5212 ( .A(n5181), .B(g_input[0]), .Z(n3147) );
  NAND U5213 ( .A(n5182), .B(n713), .Z(n5181) );
  NANDN U5214 ( .B(n5183), .A(n5184), .Z(n713) );
  ANDN U5215 ( .A(e_input[31]), .B(n5185), .Z(n5184) );
  NAND U5216 ( .A(n3833), .B(n746), .Z(n5182) );
  XOR U5217 ( .A(n5185), .B(e_input[30]), .Z(n5183) );
  OR U5218 ( .A(n5178), .B(n5186), .Z(n5185) );
  XOR U5219 ( .A(n5186), .B(e_input[29]), .Z(n5178) );
  OR U5220 ( .A(n5177), .B(n5187), .Z(n5186) );
  XOR U5221 ( .A(n5187), .B(e_input[28]), .Z(n5177) );
  OR U5222 ( .A(n5143), .B(n5188), .Z(n5187) );
  XOR U5223 ( .A(n5188), .B(e_input[27]), .Z(n5143) );
  OR U5224 ( .A(n5144), .B(n5189), .Z(n5188) );
  XOR U5225 ( .A(n5189), .B(e_input[26]), .Z(n5144) );
  OR U5226 ( .A(n5159), .B(n5190), .Z(n5189) );
  XOR U5227 ( .A(n5190), .B(e_input[25]), .Z(n5159) );
  OR U5228 ( .A(n5158), .B(n5191), .Z(n5190) );
  XOR U5229 ( .A(n5191), .B(e_input[24]), .Z(n5158) );
  OR U5230 ( .A(n4887), .B(n5192), .Z(n5191) );
  XOR U5231 ( .A(n5192), .B(e_input[23]), .Z(n4887) );
  OR U5232 ( .A(n4888), .B(n5193), .Z(n5192) );
  XOR U5233 ( .A(n5193), .B(e_input[22]), .Z(n4888) );
  OR U5234 ( .A(n4883), .B(n5194), .Z(n5193) );
  XOR U5235 ( .A(n5194), .B(e_input[21]), .Z(n4883) );
  OR U5236 ( .A(n4882), .B(n5195), .Z(n5194) );
  XOR U5237 ( .A(n5195), .B(e_input[20]), .Z(n4882) );
  OR U5238 ( .A(n5054), .B(n5196), .Z(n5195) );
  XOR U5239 ( .A(n5196), .B(e_input[19]), .Z(n5054) );
  OR U5240 ( .A(n5053), .B(n5197), .Z(n5196) );
  XOR U5241 ( .A(n5197), .B(e_input[18]), .Z(n5053) );
  OR U5242 ( .A(n5069), .B(n5198), .Z(n5197) );
  XOR U5243 ( .A(n5198), .B(e_input[17]), .Z(n5069) );
  OR U5244 ( .A(n5068), .B(n5199), .Z(n5198) );
  XOR U5245 ( .A(n5199), .B(e_input[16]), .Z(n5068) );
  OR U5246 ( .A(n3873), .B(n5200), .Z(n5199) );
  XOR U5247 ( .A(n5200), .B(e_input[15]), .Z(n3873) );
  OR U5248 ( .A(n3872), .B(n5201), .Z(n5200) );
  XOR U5249 ( .A(n5201), .B(e_input[14]), .Z(n3872) );
  OR U5250 ( .A(n3868), .B(n5202), .Z(n5201) );
  XOR U5251 ( .A(n5202), .B(e_input[13]), .Z(n3868) );
  OR U5252 ( .A(n3867), .B(n5203), .Z(n5202) );
  XOR U5253 ( .A(n5203), .B(e_input[12]), .Z(n3867) );
  OR U5254 ( .A(n3838), .B(n5204), .Z(n5203) );
  XOR U5255 ( .A(n5204), .B(e_input[11]), .Z(n3838) );
  OR U5256 ( .A(n3837), .B(n5205), .Z(n5204) );
  XOR U5257 ( .A(n5205), .B(e_input[10]), .Z(n3837) );
  OR U5258 ( .A(n3853), .B(n5206), .Z(n5205) );
  XOR U5259 ( .A(n5206), .B(e_input[9]), .Z(n3853) );
  OR U5260 ( .A(n3852), .B(n5207), .Z(n5206) );
  XOR U5261 ( .A(n5207), .B(e_input[8]), .Z(n3852) );
  OR U5262 ( .A(n4323), .B(n5208), .Z(n5207) );
  XOR U5263 ( .A(n5208), .B(e_input[7]), .Z(n4323) );
  OR U5264 ( .A(n4322), .B(n5209), .Z(n5208) );
  XOR U5265 ( .A(n5209), .B(e_input[6]), .Z(n4322) );
  OR U5266 ( .A(n4318), .B(n5210), .Z(n5209) );
  XOR U5267 ( .A(n5210), .B(e_input[5]), .Z(n4318) );
  OR U5268 ( .A(n4317), .B(n5211), .Z(n5210) );
  XOR U5269 ( .A(n5211), .B(e_input[4]), .Z(n4317) );
  OR U5270 ( .A(n4682), .B(n5212), .Z(n5211) );
  XOR U5271 ( .A(n5212), .B(e_input[3]), .Z(n4682) );
  OR U5272 ( .A(n4681), .B(n5213), .Z(n5212) );
  XOR U5273 ( .A(n5213), .B(e_input[2]), .Z(n4681) );
  NANDN U5274 ( .B(e_input[0]), .A(n4696), .Z(n5213) );
  XNOR U5275 ( .A(e_input[0]), .B(e_input[1]), .Z(n4696) );
  XOR U5276 ( .A(g_input[0]), .B(g_input[1]), .Z(n5180) );
  AND U5277 ( .A(n5214), .B(n5215), .Z(\_MxM/N23 ) );
  XOR U5278 ( .A(\_MxM/n[9] ), .B(\_MxM/add_43/carry[9] ), .Z(n5215) );
  AND U5279 ( .A(\_MxM/N12 ), .B(n5214), .Z(\_MxM/N22 ) );
  AND U5280 ( .A(\_MxM/N11 ), .B(n5214), .Z(\_MxM/N21 ) );
  AND U5281 ( .A(\_MxM/N10 ), .B(n5214), .Z(\_MxM/N20 ) );
  AND U5282 ( .A(\_MxM/N9 ), .B(n5214), .Z(\_MxM/N19 ) );
  AND U5283 ( .A(\_MxM/N8 ), .B(n5214), .Z(\_MxM/N18 ) );
  AND U5284 ( .A(\_MxM/N7 ), .B(n5214), .Z(\_MxM/N17 ) );
  AND U5285 ( .A(\_MxM/N6 ), .B(n5214), .Z(\_MxM/N16 ) );
  AND U5286 ( .A(\_MxM/N5 ), .B(n5214), .Z(\_MxM/N15 ) );
  NAND U5287 ( .A(n5216), .B(n5217), .Z(n5214) );
  AND U5288 ( .A(n5218), .B(n5219), .Z(n5217) );
  AND U5289 ( .A(\_MxM/n[1] ), .B(n5220), .Z(n5219) );
  NOR U5290 ( .A(\_MxM/N14 ), .B(n654), .Z(n5220) );
  OR U5291 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n654) );
  AND U5292 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n5218) );
  AND U5293 ( .A(n5221), .B(n5222), .Z(n5216) );
  AND U5294 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n5222) );
  AND U5295 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n5221) );
  IV U5296 ( .A(\_MxM/n[0] ), .Z(\_MxM/N14 ) );
endmodule

