
module MxM_TG_W16_N10000 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MxM/n104 , \_MxM/n101 , \_MxM/n98 , \_MxM/n95 , \_MxM/n92 ,
         \_MxM/n89 , \_MxM/n86 , \_MxM/n83 , \_MxM/n80 , \_MxM/n77 ,
         \_MxM/n74 , \_MxM/n71 , \_MxM/n68 , \_MxM/n65 , \_MxM/n62 ,
         \_MxM/n59 , \_MxM/N31 , \_MxM/N30 , \_MxM/N29 , \_MxM/N28 ,
         \_MxM/N27 , \_MxM/N26 , \_MxM/N25 , \_MxM/N24 , \_MxM/N23 ,
         \_MxM/N22 , \_MxM/N21 , \_MxM/N20 , \_MxM/N19 , \_MxM/N18 ,
         \_MxM/N16 , \_MxM/N15 , \_MxM/N14 , \_MxM/N13 , \_MxM/N12 ,
         \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/N7 , \_MxM/N6 ,
         \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] ,
         \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] ,
         \_MxM/n[9] , \_MxM/n[10] , \_MxM/n[11] , \_MxM/n[12] , \_MxM/n[13] ,
         \_MxM/Y1[0] , \_MxM/Y1[1] , \_MxM/Y1[2] , \_MxM/Y1[3] , \_MxM/Y1[4] ,
         \_MxM/Y1[5] , \_MxM/Y1[6] , \_MxM/Y1[7] , \_MxM/Y1[8] , \_MxM/Y1[9] ,
         \_MxM/Y1[10] , \_MxM/Y1[11] , \_MxM/Y1[12] , \_MxM/Y1[13] ,
         \_MxM/Y1[14] , \_MxM/Y1[15] , \_MxM/Y0[15] , \_MxM/Y0[14] ,
         \_MxM/Y0[13] , \_MxM/Y0[12] , \_MxM/Y0[11] , \_MxM/Y0[10] ,
         \_MxM/Y0[9] , \_MxM/Y0[8] , \_MxM/Y0[7] , \_MxM/Y0[6] , \_MxM/Y0[5] ,
         \_MxM/Y0[4] , \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] , \_MxM/Y0[0] ,
         \_MxM/add_43/carry[13] , \_MxM/add_43/carry[12] ,
         \_MxM/add_43/carry[11] , \_MxM/add_43/carry[10] ,
         \_MxM/add_43/carry[9] , \_MxM/add_43/carry[8] ,
         \_MxM/add_43/carry[7] , \_MxM/add_43/carry[6] ,
         \_MxM/add_43/carry[5] , \_MxM/add_43/carry[4] ,
         \_MxM/add_43/carry[3] , \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386;

  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n59 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/Y1[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n62 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/Y1[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n65 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/Y1[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n68 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/Y1[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n71 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/Y1[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n74 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/Y1[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n77 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/Y1[9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n80 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/Y1[8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n83 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n86 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n89 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n92 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n95 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n98 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n101 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n104 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[13]  ( .D(\_MxM/N31 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[13] ) );
  DFF \_MxM/n_reg[12]  ( .D(\_MxM/N30 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[12] ) );
  DFF \_MxM/n_reg[11]  ( .D(\_MxM/N29 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[11] ) );
  DFF \_MxM/n_reg[10]  ( .D(\_MxM/N28 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[10] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N27 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N26 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N25 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N24 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_43/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_43/carry[6] ), .COUT(\_MxM/add_43/carry[7] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_43/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_43/carry[7] ), .COUT(\_MxM/add_43/carry[8] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_43/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_43/carry[8] ), .COUT(\_MxM/add_43/carry[9] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_43/U1_1_9  ( .IN0(\_MxM/n[9] ), .IN1(\_MxM/add_43/carry[9] ), .COUT(\_MxM/add_43/carry[10] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_43/U1_1_10  ( .IN0(\_MxM/n[10] ), .IN1(
        \_MxM/add_43/carry[10] ), .COUT(\_MxM/add_43/carry[11] ), .SUM(
        \_MxM/N14 ) );
  HADDER \_MxM/add_43/U1_1_11  ( .IN0(\_MxM/n[11] ), .IN1(
        \_MxM/add_43/carry[11] ), .COUT(\_MxM/add_43/carry[12] ), .SUM(
        \_MxM/N15 ) );
  HADDER \_MxM/add_43/U1_1_12  ( .IN0(\_MxM/n[12] ), .IN1(
        \_MxM/add_43/carry[12] ), .COUT(\_MxM/add_43/carry[13] ), .SUM(
        \_MxM/N16 ) );
  MUX U1 ( .IN0(n1), .IN1(n1303), .SEL(n1304), .F(n1284) );
  IV U2 ( .A(n1305), .Z(n1) );
  MUX U3 ( .IN0(n2), .IN1(n848), .SEL(n849), .F(n827) );
  IV U4 ( .A(n850), .Z(n2) );
  XOR U5 ( .A(n1068), .B(n1058), .Z(n868) );
  MUX U6 ( .IN0(n1002), .IN1(n1005), .SEL(n1003), .F(n987) );
  XOR U7 ( .A(n1040), .B(n1041), .Z(n843) );
  MUX U8 ( .IN0(n3), .IN1(n563), .SEL(n564), .F(n502) );
  IV U9 ( .A(n565), .Z(n3) );
  MUX U10 ( .IN0(e_input[12]), .IN1(n1355), .SEL(e_input[15]), .F(n230) );
  MUX U11 ( .IN0(n1284), .IN1(n1302), .SEL(n1286), .F(n1264) );
  XOR U12 ( .A(n1050), .B(n1051), .Z(n866) );
  MUX U13 ( .IN0(n4), .IN1(n808), .SEL(n809), .F(n741) );
  IV U14 ( .A(n810), .Z(n4) );
  XOR U15 ( .A(n851), .B(n833), .Z(n837) );
  MUX U16 ( .IN0(n1045), .IN1(n5), .SEL(n1044), .F(n1034) );
  IV U17 ( .A(n1043), .Z(n5) );
  MUX U18 ( .IN0(e_input[8]), .IN1(n1331), .SEL(e_input[15]), .F(n389) );
  XNOR U19 ( .A(n1333), .B(n783), .Z(n787) );
  MUX U20 ( .IN0(n6), .IN1(n1089), .SEL(n1090), .F(n1072) );
  IV U21 ( .A(n1091), .Z(n6) );
  MUX U22 ( .IN0(n1233), .IN1(n1263), .SEL(n1235), .F(n761) );
  XOR U23 ( .A(n809), .B(n810), .Z(n806) );
  MUX U24 ( .IN0(n7), .IN1(n1039), .SEL(n1040), .F(n815) );
  IV U25 ( .A(n1041), .Z(n7) );
  MUX U26 ( .IN0(n8), .IN1(n444), .SEL(n445), .F(n390) );
  IV U27 ( .A(n446), .Z(n8) );
  MUX U28 ( .IN0(n605), .IN1(n9), .SEL(n604), .F(n540) );
  IV U29 ( .A(n603), .Z(n9) );
  MUX U30 ( .IN0(e_input[13]), .IN1(n1356), .SEL(e_input[15]), .F(n195) );
  MUX U31 ( .IN0(n10), .IN1(n1049), .SEL(n1050), .F(n1039) );
  IV U32 ( .A(n1051), .Z(n10) );
  MUX U33 ( .IN0(n11), .IN1(n1057), .SEL(n1058), .F(n1043) );
  IV U34 ( .A(n1059), .Z(n11) );
  MUX U35 ( .IN0(n12), .IN1(n741), .SEL(n742), .F(n671) );
  IV U36 ( .A(n743), .Z(n12) );
  MUX U37 ( .IN0(n13), .IN1(n733), .SEL(n734), .F(n663) );
  IV U38 ( .A(n735), .Z(n13) );
  MUX U39 ( .IN0(n14), .IN1(n555), .SEL(n556), .F(n494) );
  IV U40 ( .A(n557), .Z(n14) );
  MUX U41 ( .IN0(e_input[9]), .IN1(n1332), .SEL(e_input[15]), .F(n342) );
  MUX U42 ( .IN0(n580), .IN1(n578), .SEL(n579), .F(n517) );
  MUX U43 ( .IN0(n233), .IN1(n15), .SEL(n232), .F(n197) );
  IV U44 ( .A(n231), .Z(n15) );
  MUX U45 ( .IN0(n16), .IN1(n1201), .SEL(n1202), .F(n1184) );
  IV U46 ( .A(n1203), .Z(n16) );
  XOR U47 ( .A(n828), .B(n829), .Z(n838) );
  MUX U48 ( .IN0(n17), .IN1(n761), .SEL(n762), .F(n692) );
  IV U49 ( .A(n763), .Z(n17) );
  MUX U50 ( .IN0(n18), .IN1(n700), .SEL(n701), .F(n626) );
  IV U51 ( .A(n702), .Z(n18) );
  MUX U52 ( .IN0(n19), .IN1(n663), .SEL(n664), .F(n603) );
  IV U53 ( .A(n665), .Z(n19) );
  MUX U54 ( .IN0(g_input[11]), .IN1(n1088), .SEL(g_input[15]), .F(n274) );
  XOR U55 ( .A(n752), .B(n753), .Z(n758) );
  MUX U56 ( .IN0(n506), .IN1(n508), .SEL(n507), .F(n448) );
  MUX U57 ( .IN0(n543), .IN1(n20), .SEL(n542), .F(n477) );
  IV U58 ( .A(n541), .Z(n20) );
  XNOR U59 ( .A(n778), .B(n712), .Z(n716) );
  XOR U60 ( .A(n849), .B(n850), .Z(n861) );
  MUX U61 ( .IN0(g_input[1]), .IN1(n1358), .SEL(g_input[15]), .F(n1012) );
  XOR U62 ( .A(n1042), .B(n1034), .Z(n824) );
  MUX U63 ( .IN0(g_input[2]), .IN1(n1349), .SEL(g_input[15]), .F(n789) );
  MUX U64 ( .IN0(n21), .IN1(n618), .SEL(n619), .F(n555) );
  IV U65 ( .A(n620), .Z(n21) );
  MUX U66 ( .IN0(n22), .IN1(n502), .SEL(n503), .F(n444) );
  IV U67 ( .A(n504), .Z(n22) );
  MUX U68 ( .IN0(g_input[10]), .IN1(n1104), .SEL(g_input[15]), .F(n314) );
  MUX U69 ( .IN0(n753), .IN1(n23), .SEL(n752), .F(n681) );
  IV U70 ( .A(n751), .Z(n23) );
  MUX U71 ( .IN0(n461), .IN1(n459), .SEL(n460), .F(n401) );
  MUX U72 ( .IN0(n384), .IN1(n386), .SEL(n385), .F(n24) );
  IV U73 ( .A(n24), .Z(n345) );
  XNOR U74 ( .A(n731), .B(n664), .Z(n668) );
  XNOR U75 ( .A(n707), .B(n640), .Z(n644) );
  MUX U76 ( .IN0(n1219), .IN1(n1222), .SEL(n1220), .F(n1201) );
  XOR U77 ( .A(n1304), .B(n1305), .Z(n1237) );
  XOR U78 ( .A(n816), .B(n817), .Z(n822) );
  MUX U79 ( .IN0(n25), .IN1(n671), .SEL(n672), .F(n607) );
  IV U80 ( .A(n673), .Z(n25) );
  MUX U81 ( .IN0(g_input[9]), .IN1(n1124), .SEL(g_input[15]), .F(n357) );
  XNOR U82 ( .A(n796), .B(n734), .Z(n738) );
  MUX U83 ( .IN0(n448), .IN1(n450), .SEL(n449), .F(n384) );
  MUX U84 ( .IN0(n403), .IN1(n401), .SEL(n402), .F(n354) );
  MUX U85 ( .IN0(n392), .IN1(n26), .SEL(n391), .F(n344) );
  IV U86 ( .A(n390), .Z(n26) );
  XNOR U87 ( .A(n635), .B(n575), .Z(n579) );
  NAND U88 ( .A(n540), .B(n601), .Z(n600) );
  MUX U89 ( .IN0(n27), .IN1(n996), .SEL(n812), .F(n969) );
  IV U90 ( .A(n811), .Z(n27) );
  MUX U91 ( .IN0(n1167), .IN1(n1183), .SEL(n1169), .F(n1156) );
  MUX U92 ( .IN0(n28), .IN1(n815), .SEL(n816), .F(n751) );
  IV U93 ( .A(n817), .Z(n28) );
  MUX U94 ( .IN0(n29), .IN1(n607), .SEL(n608), .F(n545) );
  IV U95 ( .A(n609), .Z(n29) );
  XOR U96 ( .A(n721), .B(n790), .Z(n722) );
  MUX U97 ( .IN0(n356), .IN1(n354), .SEL(n355), .F(n311) );
  MUX U98 ( .IN0(e_input[10]), .IN1(n1310), .SEL(e_input[15]), .F(n293) );
  XOR U99 ( .A(n596), .B(n541), .Z(n542) );
  XNOR U100 ( .A(n570), .B(n514), .Z(n518) );
  XOR U101 ( .A(n442), .B(n391), .Z(n385) );
  MUX U102 ( .IN0(n431), .IN1(n433), .SEL(n432), .F(n30) );
  IV U103 ( .A(n30), .Z(n372) );
  XOR U104 ( .A(n587), .B(n590), .Z(n588) );
  MUX U105 ( .IN0(n939), .IN1(n31), .SEL(n940), .F(n912) );
  IV U106 ( .A(n941), .Z(n31) );
  MUX U107 ( .IN0(n32), .IN1(n1072), .SEL(n1073), .F(n1057) );
  IV U108 ( .A(n1074), .Z(n32) );
  XOR U109 ( .A(n1135), .B(n1136), .Z(n998) );
  MUX U110 ( .IN0(n632), .IN1(n634), .SEL(n633), .F(n567) );
  XOR U111 ( .A(n465), .B(n521), .Z(n466) );
  MUX U112 ( .IN0(e_input[6]), .IN1(n1021), .SEL(e_input[15]), .F(n482) );
  MUX U113 ( .IN0(n33), .IN1(n333), .SEL(n334), .F(n294) );
  IV U114 ( .A(n335), .Z(n33) );
  XNOR U115 ( .A(n661), .B(n604), .Z(n598) );
  MUX U116 ( .IN0(n34), .IN1(n558), .SEL(n559), .F(n497) );
  IV U117 ( .A(n560), .Z(n34) );
  XNOR U118 ( .A(n509), .B(n456), .Z(n460) );
  NAND U119 ( .A(n344), .B(n388), .Z(n387) );
  XOR U120 ( .A(n526), .B(n529), .Z(n527) );
  MUX U121 ( .IN0(n35), .IN1(n1125), .SEL(n1126), .F(n1106) );
  IV U122 ( .A(n1127), .Z(n35) );
  MUX U123 ( .IN0(n36), .IN1(n1023), .SEL(n1024), .F(n1195) );
  IV U124 ( .A(n1211), .Z(n36) );
  MUX U125 ( .IN0(n1150), .IN1(n1172), .SEL(n1152), .F(n1132) );
  XOR U126 ( .A(n830), .B(n801), .Z(n805) );
  MUX U127 ( .IN0(g_input[3]), .IN1(n1336), .SEL(g_input[15]), .F(n37) );
  IV U128 ( .A(n37), .Z(n718) );
  MUX U129 ( .IN0(n38), .IN1(n692), .SEL(n693), .F(n618) );
  IV U130 ( .A(n694), .Z(n38) );
  MUX U131 ( .IN0(n788), .IN1(n786), .SEL(n787), .F(n715) );
  XOR U132 ( .A(n584), .B(n647), .Z(n585) );
  MUX U133 ( .IN0(n567), .IN1(n569), .SEL(n568), .F(n506) );
  MUX U134 ( .IN0(n273), .IN1(n271), .SEL(n272), .F(n223) );
  MUX U135 ( .IN0(g_input[12]), .IN1(n1070), .SEL(g_input[15]), .F(n234) );
  XOR U136 ( .A(n484), .B(n485), .Z(n479) );
  MUX U137 ( .IN0(n39), .IN1(n439), .SEL(n440), .F(n380) );
  IV U138 ( .A(n441), .Z(n39) );
  XNOR U139 ( .A(n451), .B(n398), .Z(n402) );
  XNOR U140 ( .A(n300), .B(n339), .Z(n301) );
  MUX U141 ( .IN0(n674), .IN1(n40), .SEL(n675), .F(n610) );
  IV U142 ( .A(n676), .Z(n40) );
  MUX U143 ( .IN0(n41), .IN1(n320), .SEL(n114), .F(n280) );
  IV U144 ( .A(\_MxM/Y0[8] ), .Z(n41) );
  XOR U145 ( .A(n468), .B(n471), .Z(n469) );
  MUX U146 ( .IN0(n1093), .IN1(n42), .SEL(n921), .F(n1076) );
  IV U147 ( .A(n919), .Z(n42) );
  MUX U148 ( .IN0(e_input[1]), .IN1(n43), .SEL(e_input[15]), .F(n1029) );
  IV U149 ( .A(n1230), .Z(n43) );
  MUX U150 ( .IN0(n836), .IN1(n44), .SEL(n837), .F(n804) );
  IV U151 ( .A(n838), .Z(n44) );
  XNOR U152 ( .A(n1009), .B(n1010), .Z(n993) );
  MUX U153 ( .IN0(n775), .IN1(n777), .SEL(n776), .F(n704) );
  MUX U154 ( .IN0(e_input[2]), .IN1(n1215), .SEL(e_input[15]), .F(n750) );
  MUX U155 ( .IN0(n519), .IN1(n517), .SEL(n518), .F(n459) );
  XOR U156 ( .A(n360), .B(n405), .Z(n361) );
  MUX U157 ( .IN0(n45), .IN1(n754), .SEL(n755), .F(n687) );
  IV U158 ( .A(n756), .Z(n45) );
  MUX U159 ( .IN0(n46), .IN1(n695), .SEL(n696), .F(n621) );
  IV U160 ( .A(n697), .Z(n46) );
  XOR U161 ( .A(n561), .B(n503), .Z(n507) );
  MUX U162 ( .IN0(n47), .IN1(n483), .SEL(n484), .F(n430) );
  IV U163 ( .A(n485), .Z(n47) );
  MUX U164 ( .IN0(n48), .IN1(n380), .SEL(n381), .F(n336) );
  IV U165 ( .A(n382), .Z(n48) );
  NAND U166 ( .A(n254), .B(n292), .Z(n291) );
  XNOR U167 ( .A(n303), .B(n268), .Z(n272) );
  MUX U168 ( .IN0(n49), .IN1(n552), .SEL(n551), .F(n489) );
  IV U169 ( .A(n550), .Z(n49) );
  MUX U170 ( .IN0(n50), .IN1(n206), .SEL(n207), .F(n176) );
  IV U171 ( .A(\_MxM/Y0[11] ), .Z(n50) );
  XOR U172 ( .A(n410), .B(n413), .Z(n411) );
  MUX U173 ( .IN0(n966), .IN1(n51), .SEL(n967), .F(n939) );
  IV U174 ( .A(n968), .Z(n51) );
  MUX U175 ( .IN0(n1129), .IN1(n52), .SEL(n975), .F(n1112) );
  IV U176 ( .A(n973), .Z(n52) );
  MUX U177 ( .IN0(n859), .IN1(n53), .SEL(n860), .F(n836) );
  IV U178 ( .A(n861), .Z(n53) );
  MUX U179 ( .IN0(n1061), .IN1(n54), .SEL(n868), .F(n1047) );
  IV U180 ( .A(n866), .Z(n54) );
  XOR U181 ( .A(n1217), .B(n1202), .Z(n1024) );
  MUX U182 ( .IN0(e_input[4]), .IN1(n1016), .SEL(e_input[15]), .F(n602) );
  XOR U183 ( .A(n1239), .B(n772), .Z(n776) );
  MUX U184 ( .IN0(n669), .IN1(n667), .SEL(n668), .F(n597) );
  MUX U185 ( .IN0(n55), .IN1(n545), .SEL(n546), .F(n483) );
  IV U186 ( .A(n547), .Z(n55) );
  MUX U187 ( .IN0(e_input[11]), .IN1(n1311), .SEL(e_input[15]), .F(n257) );
  MUX U188 ( .IN0(n56), .IN1(n621), .SEL(n622), .F(n558) );
  IV U189 ( .A(n623), .Z(n56) );
  XNOR U190 ( .A(n263), .B(n232), .Z(n226) );
  MUX U191 ( .IN0(n57), .IN1(n260), .SEL(n261), .F(n218) );
  IV U192 ( .A(n262), .Z(n57) );
  MUX U193 ( .IN0(e_input[14]), .IN1(n1361), .SEL(e_input[15]), .F(n165) );
  XNOR U194 ( .A(n613), .B(n677), .Z(n614) );
  MUX U195 ( .IN0(n489), .IN1(n491), .SEL(n490), .F(n431) );
  MUX U196 ( .IN0(n58), .IN1(n652), .SEL(n120), .F(n587) );
  IV U197 ( .A(\_MxM/Y0[2] ), .Z(n58) );
  XNOR U198 ( .A(n176), .B(n177), .Z(n134) );
  XOR U199 ( .A(n364), .B(n370), .Z(n115) );
  MUX U200 ( .IN0(n1112), .IN1(n59), .SEL(n948), .F(n1093) );
  IV U201 ( .A(n946), .Z(n59) );
  MUX U202 ( .IN0(n60), .IN1(n1223), .SEL(n1224), .F(n1219) );
  IV U203 ( .A(n1225), .Z(n60) );
  MUX U204 ( .IN0(n1047), .IN1(n61), .SEL(n845), .F(n1035) );
  IV U205 ( .A(n843), .Z(n61) );
  MUX U206 ( .IN0(n804), .IN1(n62), .SEL(n805), .F(n737) );
  IV U207 ( .A(n806), .Z(n62) );
  XNOR U208 ( .A(n1000), .B(n990), .Z(n994) );
  MUX U209 ( .IN0(g_input[5]), .IN1(n1276), .SEL(g_input[15]), .F(n581) );
  MUX U210 ( .IN0(n717), .IN1(n715), .SEL(n716), .F(n643) );
  MUX U211 ( .IN0(n347), .IN1(n63), .SEL(n346), .F(n300) );
  IV U212 ( .A(n345), .Z(n63) );
  XOR U213 ( .A(n277), .B(n315), .Z(n278) );
  MUX U214 ( .IN0(n64), .IN1(n764), .SEL(n765), .F(n695) );
  IV U215 ( .A(n766), .Z(n64) );
  NAND U216 ( .A(n681), .B(n749), .Z(n748) );
  XOR U217 ( .A(n698), .B(n629), .Z(n633) );
  XOR U218 ( .A(n546), .B(n547), .Z(n543) );
  MUX U219 ( .IN0(n65), .IN1(n497), .SEL(n498), .F(n439) );
  IV U220 ( .A(n499), .Z(n65) );
  XNOR U221 ( .A(n393), .B(n351), .Z(n355) );
  MUX U222 ( .IN0(n66), .IN1(n297), .SEL(n298), .F(n260) );
  IV U223 ( .A(n299), .Z(n66) );
  MUX U224 ( .IN0(n296), .IN1(n67), .SEL(n295), .F(n254) );
  IV U225 ( .A(n294), .Z(n67) );
  XNOR U226 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U227 ( .A(n599), .B(n598), .Z(n615) );
  XNOR U228 ( .A(n227), .B(n226), .Z(n220) );
  XOR U229 ( .A(n476), .B(n424), .Z(n432) );
  MUX U230 ( .IN0(n68), .IN1(n526), .SEL(n118), .F(n468) );
  IV U231 ( .A(\_MxM/Y0[4] ), .Z(n68) );
  MUX U232 ( .IN0(\_MxM/Y0[13] ), .IN1(n134), .SEL(n133), .F(n130) );
  XOR U233 ( .A(n280), .B(n283), .Z(n281) );
  XOR U234 ( .A(n1154), .B(n1145), .Z(n999) );
  MUX U235 ( .IN0(n69), .IN1(n436), .SEL(n437), .F(n377) );
  IV U236 ( .A(n438), .Z(n69) );
  MUX U237 ( .IN0(e_input[3]), .IN1(n1216), .SEL(e_input[15]), .F(n684) );
  MUX U238 ( .IN0(n645), .IN1(n643), .SEL(n644), .F(n578) );
  MUX U239 ( .IN0(e_input[5]), .IN1(n1017), .SEL(e_input[15]), .F(n538) );
  MUX U240 ( .IN0(n313), .IN1(n311), .SEL(n312), .F(n271) );
  XOR U241 ( .A(n767), .B(n701), .Z(n705) );
  XNOR U242 ( .A(n788), .B(n787), .Z(n766) );
  MUX U243 ( .IN0(n689), .IN1(n70), .SEL(n688), .F(n613) );
  IV U244 ( .A(n687), .Z(n70) );
  MUX U245 ( .IN0(e_input[7]), .IN1(n1022), .SEL(e_input[15]), .F(n422) );
  MUX U246 ( .IN0(n302), .IN1(n300), .SEL(n301), .F(n71) );
  IV U247 ( .A(n71), .Z(n259) );
  NAND U248 ( .A(n197), .B(n229), .Z(n228) );
  XOR U249 ( .A(n203), .B(n235), .Z(n204) );
  MUX U250 ( .IN0(n610), .IN1(n72), .SEL(n611), .F(n550) );
  IV U251 ( .A(n612), .Z(n72) );
  XNOR U252 ( .A(n403), .B(n402), .Z(n382) );
  MUX U253 ( .IN0(n220), .IN1(n73), .SEL(n219), .F(n191) );
  IV U254 ( .A(n218), .Z(n73) );
  XNOR U255 ( .A(n499), .B(n498), .Z(n491) );
  MUX U256 ( .IN0(n74), .IN1(n468), .SEL(n117), .F(n410) );
  IV U257 ( .A(\_MxM/Y0[5] ), .Z(n74) );
  MUX U258 ( .IN0(n75), .IN1(n280), .SEL(n113), .F(n240) );
  IV U259 ( .A(\_MxM/Y0[9] ), .Z(n75) );
  MUX U260 ( .IN0(n76), .IN1(n128), .SEL(n127), .F(n132) );
  IV U261 ( .A(n135), .Z(n76) );
  MUX U262 ( .IN0(n912), .IN1(n77), .SEL(n913), .F(n885) );
  IV U263 ( .A(n914), .Z(n77) );
  MUX U264 ( .IN0(n1191), .IN1(n1205), .SEL(n1193), .F(n1173) );
  XNOR U265 ( .A(n1224), .B(n1225), .Z(n1211) );
  XOR U266 ( .A(n1335), .B(g_input[3]), .Z(n1336) );
  MUX U267 ( .IN0(g_input[6]), .IN1(n1255), .SEL(g_input[15]), .F(n520) );
  MUX U268 ( .IN0(n78), .IN1(n494), .SEL(n495), .F(n436) );
  IV U269 ( .A(n496), .Z(n78) );
  MUX U270 ( .IN0(g_input[7]), .IN1(n1242), .SEL(g_input[15]), .F(n462) );
  MUX U271 ( .IN0(g_input[8]), .IN1(n1140), .SEL(g_input[15]), .F(n404) );
  XNOR U272 ( .A(n1035), .B(n1036), .Z(n1025) );
  XNOR U273 ( .A(n995), .B(n994), .Z(n811) );
  MUX U274 ( .IN0(n599), .IN1(n597), .SEL(n598), .F(n541) );
  XNOR U275 ( .A(n739), .B(n738), .Z(n756) );
  XOR U276 ( .A(n624), .B(n564), .Z(n568) );
  MUX U277 ( .IN0(n79), .IN1(n336), .SEL(n337), .F(n297) );
  IV U278 ( .A(n338), .Z(n79) );
  XNOR U279 ( .A(n348), .B(n308), .Z(n312) );
  MUX U280 ( .IN0(g_input[13]), .IN1(n1056), .SEL(g_input[15]), .F(n200) );
  XNOR U281 ( .A(n669), .B(n668), .Z(n689) );
  XNOR U282 ( .A(n766), .B(n765), .Z(n746) );
  XNOR U283 ( .A(n645), .B(n644), .Z(n623) );
  XNOR U284 ( .A(n580), .B(n579), .Z(n560) );
  AND U285 ( .A(n160), .B(n141), .Z(n159) );
  XNOR U286 ( .A(n697), .B(n696), .Z(n676) );
  XNOR U287 ( .A(n489), .B(n488), .Z(n534) );
  MUX U288 ( .IN0(n80), .IN1(n587), .SEL(n119), .F(n526) );
  IV U289 ( .A(\_MxM/Y0[3] ), .Z(n80) );
  XNOR U290 ( .A(n441), .B(n440), .Z(n433) );
  XNOR U291 ( .A(n382), .B(n381), .Z(n374) );
  MUX U292 ( .IN0(n81), .IN1(n363), .SEL(n115), .F(n320) );
  IV U293 ( .A(\_MxM/Y0[7] ), .Z(n81) );
  XNOR U294 ( .A(n190), .B(n191), .Z(n189) );
  XOR U295 ( .A(n240), .B(n243), .Z(n241) );
  MUX U296 ( .IN0(\_MxM/Y0[14] ), .IN1(n130), .SEL(n131), .F(n124) );
  MUX U297 ( .IN0(n995), .IN1(n993), .SEL(n994), .F(n966) );
  MUX U298 ( .IN0(n1148), .IN1(n82), .SEL(n999), .F(n1129) );
  IV U299 ( .A(n998), .Z(n82) );
  MUX U300 ( .IN0(n83), .IN1(n1237), .SEL(n1238), .F(n1288) );
  IV U301 ( .A(n1306), .Z(n83) );
  MUX U302 ( .IN0(n885), .IN1(n84), .SEL(n886), .F(n859) );
  IV U303 ( .A(n887), .Z(n84) );
  NOR U304 ( .A(g_input[0]), .B(n1358), .Z(n1350) );
  MUX U305 ( .IN0(n1076), .IN1(n85), .SEL(n894), .F(n1061) );
  IV U306 ( .A(n892), .Z(n85) );
  MUX U307 ( .IN0(n86), .IN1(n827), .SEL(n828), .F(n808) );
  IV U308 ( .A(n829), .Z(n86) );
  MUX U309 ( .IN0(n87), .IN1(n832), .SEL(n833), .F(n798) );
  IV U310 ( .A(n834), .Z(n87) );
  MUX U311 ( .IN0(n1156), .IN1(n1166), .SEL(n1158), .F(n1142) );
  XOR U312 ( .A(n1209), .B(n1210), .Z(n1023) );
  MUX U313 ( .IN0(g_input[4]), .IN1(n1294), .SEL(g_input[15]), .F(n88) );
  IV U314 ( .A(n88), .Z(n646) );
  MUX U315 ( .IN0(n89), .IN1(n350), .SEL(n351), .F(n305) );
  IV U316 ( .A(n352), .Z(n89) );
  MUX U317 ( .IN0(n90), .IN1(n377), .SEL(n378), .F(n333) );
  IV U318 ( .A(n379), .Z(n90) );
  MUX U319 ( .IN0(n739), .IN1(n737), .SEL(n738), .F(n667) );
  MUX U320 ( .IN0(n704), .IN1(n706), .SEL(n705), .F(n632) );
  MUX U321 ( .IN0(n758), .IN1(n1025), .SEL(n757), .F(n686) );
  XOR U322 ( .A(n500), .B(n445), .Z(n449) );
  MUX U323 ( .IN0(n479), .IN1(n477), .SEL(n478), .F(n428) );
  XNOR U324 ( .A(n717), .B(n716), .Z(n697) );
  MUX U325 ( .IN0(n744), .IN1(n91), .SEL(n745), .F(n674) );
  IV U326 ( .A(n746), .Z(n91) );
  MUX U327 ( .IN0(n615), .IN1(n613), .SEL(n614), .F(n92) );
  IV U328 ( .A(n92), .Z(n549) );
  XNOR U329 ( .A(n519), .B(n518), .Z(n499) );
  XNOR U330 ( .A(n461), .B(n460), .Z(n441) );
  XNOR U331 ( .A(n356), .B(n355), .Z(n338) );
  XNOR U332 ( .A(n313), .B(n312), .Z(n299) );
  XNOR U333 ( .A(n273), .B(n272), .Z(n262) );
  MUX U334 ( .IN0(n199), .IN1(n222), .SEL(n198), .F(n171) );
  MUX U335 ( .IN0(g_input[14]), .IN1(n1030), .SEL(g_input[15]), .F(n166) );
  XNOR U336 ( .A(n623), .B(n622), .Z(n612) );
  XNOR U337 ( .A(n560), .B(n559), .Z(n552) );
  MUX U338 ( .IN0(n372), .IN1(n93), .SEL(n373), .F(n330) );
  IV U339 ( .A(n374), .Z(n93) );
  MUX U340 ( .IN0(n94), .IN1(n410), .SEL(n116), .F(n363) );
  IV U341 ( .A(\_MxM/Y0[6] ), .Z(n94) );
  MUX U342 ( .IN0(n95), .IN1(n240), .SEL(n112), .F(n206) );
  IV U343 ( .A(\_MxM/Y0[10] ), .Z(n95) );
  MUX U344 ( .IN0(n724), .IN1(n96), .SEL(n725), .F(n652) );
  IV U345 ( .A(\_MxM/Y0[1] ), .Z(n96) );
  XNOR U346 ( .A(n189), .B(n188), .Z(n210) );
  MUX U347 ( .IN0(\_MxM/Y0[15] ), .IN1(n124), .SEL(n125), .F(n97) );
  IV U348 ( .A(n97), .Z(n121) );
  MUX U349 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n98), .F(\_MxM/n98 ) );
  MUX U350 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n98), .F(\_MxM/n95 ) );
  MUX U351 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n98), .F(\_MxM/n92 ) );
  MUX U352 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n98), .F(\_MxM/n89 ) );
  MUX U353 ( .IN0(\_MxM/Y1[6] ), .IN1(o[6]), .SEL(n98), .F(\_MxM/n86 ) );
  MUX U354 ( .IN0(\_MxM/Y1[7] ), .IN1(o[7]), .SEL(n98), .F(\_MxM/n83 ) );
  MUX U355 ( .IN0(\_MxM/Y1[8] ), .IN1(o[8]), .SEL(n98), .F(\_MxM/n80 ) );
  MUX U356 ( .IN0(\_MxM/Y1[9] ), .IN1(o[9]), .SEL(n98), .F(\_MxM/n77 ) );
  MUX U357 ( .IN0(\_MxM/Y1[10] ), .IN1(o[10]), .SEL(n98), .F(\_MxM/n74 ) );
  MUX U358 ( .IN0(\_MxM/Y1[11] ), .IN1(o[11]), .SEL(n98), .F(\_MxM/n71 ) );
  MUX U359 ( .IN0(\_MxM/Y1[12] ), .IN1(o[12]), .SEL(n98), .F(\_MxM/n68 ) );
  MUX U360 ( .IN0(\_MxM/Y1[13] ), .IN1(o[13]), .SEL(n98), .F(\_MxM/n65 ) );
  MUX U361 ( .IN0(\_MxM/Y1[14] ), .IN1(o[14]), .SEL(n98), .F(\_MxM/n62 ) );
  MUX U362 ( .IN0(\_MxM/Y1[15] ), .IN1(o[15]), .SEL(n98), .F(\_MxM/n59 ) );
  IV U363 ( .A(n99), .Z(n98) );
  MUX U364 ( .IN0(o[0]), .IN1(\_MxM/Y1[0] ), .SEL(n99), .F(\_MxM/n104 ) );
  MUX U365 ( .IN0(o[1]), .IN1(\_MxM/Y1[1] ), .SEL(n99), .F(\_MxM/n101 ) );
  AND U366 ( .A(n100), .B(n101), .Z(n99) );
  AND U367 ( .A(n102), .B(n103), .Z(n101) );
  ANDN U368 ( .A(n104), .B(\_MxM/n[3] ), .Z(n103) );
  NOR U369 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n104) );
  ANDN U370 ( .A(n105), .B(\_MxM/n[13] ), .Z(n102) );
  NOR U371 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n105) );
  AND U372 ( .A(n106), .B(n107), .Z(n100) );
  ANDN U373 ( .A(n108), .B(\_MxM/n[10] ), .Z(n107) );
  ANDN U374 ( .A(n109), .B(n110), .Z(n106) );
  NOR U375 ( .A(\_MxM/n[0] ), .B(n111), .Z(n109) );
  XNOR U376 ( .A(n112), .B(\_MxM/Y0[10] ), .Z(\_MxM/Y1[9] ) );
  XNOR U377 ( .A(n113), .B(\_MxM/Y0[9] ), .Z(\_MxM/Y1[8] ) );
  XNOR U378 ( .A(n114), .B(\_MxM/Y0[8] ), .Z(\_MxM/Y1[7] ) );
  XNOR U379 ( .A(n115), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XNOR U380 ( .A(n116), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XNOR U381 ( .A(n117), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U382 ( .A(n118), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U383 ( .A(n119), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U384 ( .A(n120), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U385 ( .A(n121), .B(n122), .Z(\_MxM/Y1[15] ) );
  XNOR U386 ( .A(\_MxM/Y0[15] ), .B(n123), .Z(n122) );
  XNOR U387 ( .A(n125), .B(\_MxM/Y0[15] ), .Z(\_MxM/Y1[14] ) );
  XOR U388 ( .A(n124), .B(n123), .Z(n125) );
  NAND U389 ( .A(n126), .B(n127), .Z(n123) );
  OR U390 ( .A(n128), .B(n129), .Z(n126) );
  XNOR U391 ( .A(n131), .B(\_MxM/Y0[14] ), .Z(\_MxM/Y1[13] ) );
  XNOR U392 ( .A(n132), .B(n130), .Z(n131) );
  XNOR U393 ( .A(n129), .B(n135), .Z(n128) );
  OR U394 ( .A(n136), .B(n137), .Z(n129) );
  AND U395 ( .A(n138), .B(n139), .Z(n135) );
  OR U396 ( .A(n140), .B(n141), .Z(n139) );
  AND U397 ( .A(n142), .B(n143), .Z(n138) );
  OR U398 ( .A(n144), .B(n145), .Z(n143) );
  OR U399 ( .A(n146), .B(n147), .Z(n142) );
  XNOR U400 ( .A(n133), .B(\_MxM/Y0[13] ), .Z(\_MxM/Y1[12] ) );
  XNOR U401 ( .A(n148), .B(n149), .Z(n133) );
  XNOR U402 ( .A(n134), .B(n150), .Z(n148) );
  AND U403 ( .A(n127), .B(n151), .Z(n150) );
  XOR U404 ( .A(n136), .B(n152), .Z(n151) );
  XOR U405 ( .A(n152), .B(n137), .Z(n136) );
  OR U406 ( .A(n153), .B(n154), .Z(n137) );
  IV U407 ( .A(n149), .Z(n152) );
  XNOR U408 ( .A(n147), .B(n146), .Z(n149) );
  OR U409 ( .A(n155), .B(n156), .Z(n146) );
  AND U410 ( .A(n157), .B(n158), .Z(n147) );
  XNOR U411 ( .A(n140), .B(n159), .Z(n158) );
  NAND U412 ( .A(n161), .B(n162), .Z(n141) );
  NANDN U413 ( .B(n163), .A(n164), .Z(n161) );
  NANDN U414 ( .B(n144), .A(n165), .Z(n160) );
  NANDN U415 ( .B(n145), .A(n166), .Z(n140) );
  AND U416 ( .A(n167), .B(n168), .Z(n157) );
  OR U417 ( .A(n169), .B(n170), .Z(n168) );
  XNOR U418 ( .A(n171), .B(n172), .Z(n167) );
  ANDN U419 ( .A(n173), .B(n174), .Z(n172) );
  XOR U420 ( .A(n171), .B(n175), .Z(n173) );
  ANDN U421 ( .A(n178), .B(n179), .Z(n177) );
  XOR U422 ( .A(\_MxM/Y0[12] ), .B(n180), .Z(n178) );
  XNOR U423 ( .A(n179), .B(\_MxM/Y0[12] ), .Z(\_MxM/Y1[11] ) );
  XNOR U424 ( .A(n181), .B(n182), .Z(n179) );
  XNOR U425 ( .A(n180), .B(n183), .Z(n181) );
  AND U426 ( .A(n127), .B(n184), .Z(n183) );
  XOR U427 ( .A(n153), .B(n185), .Z(n184) );
  XOR U428 ( .A(n185), .B(n154), .Z(n153) );
  OR U429 ( .A(n186), .B(n187), .Z(n154) );
  IV U430 ( .A(n182), .Z(n185) );
  XNOR U431 ( .A(n156), .B(n155), .Z(n182) );
  OR U432 ( .A(n188), .B(n189), .Z(n155) );
  XNOR U433 ( .A(n170), .B(n169), .Z(n156) );
  OR U434 ( .A(n190), .B(n191), .Z(n169) );
  XOR U435 ( .A(n175), .B(n174), .Z(n170) );
  XOR U436 ( .A(n171), .B(n192), .Z(n174) );
  AND U437 ( .A(n193), .B(n194), .Z(n192) );
  NANDN U438 ( .B(n144), .A(n195), .Z(n194) );
  OR U439 ( .A(n196), .B(n197), .Z(n193) );
  XOR U440 ( .A(n163), .B(n164), .Z(n175) );
  NANDN U441 ( .B(n145), .A(n200), .Z(n164) );
  XNOR U442 ( .A(n162), .B(n201), .Z(n163) );
  AND U443 ( .A(n166), .B(n165), .Z(n201) );
  ANDN U444 ( .A(n202), .B(n203), .Z(n162) );
  NANDN U445 ( .B(n204), .A(n205), .Z(n202) );
  IV U446 ( .A(n176), .Z(n180) );
  XNOR U447 ( .A(n207), .B(\_MxM/Y0[11] ), .Z(\_MxM/Y1[10] ) );
  XNOR U448 ( .A(n209), .B(n210), .Z(n207) );
  XNOR U449 ( .A(n208), .B(n211), .Z(n209) );
  AND U450 ( .A(n127), .B(n212), .Z(n211) );
  XOR U451 ( .A(n186), .B(n213), .Z(n212) );
  XOR U452 ( .A(n213), .B(n187), .Z(n186) );
  OR U453 ( .A(n214), .B(n215), .Z(n187) );
  IV U454 ( .A(n210), .Z(n213) );
  OR U455 ( .A(n216), .B(n217), .Z(n188) );
  XOR U456 ( .A(n199), .B(n198), .Z(n190) );
  XNOR U457 ( .A(n221), .B(n222), .Z(n198) );
  ANDN U458 ( .A(n225), .B(n226), .Z(n224) );
  XOR U459 ( .A(n223), .B(n227), .Z(n225) );
  XNOR U460 ( .A(n228), .B(n196), .Z(n221) );
  NAND U461 ( .A(n195), .B(n166), .Z(n196) );
  NANDN U462 ( .B(n144), .A(n230), .Z(n229) );
  XOR U463 ( .A(n204), .B(n205), .Z(n199) );
  NANDN U464 ( .B(n145), .A(n234), .Z(n205) );
  AND U465 ( .A(n200), .B(n165), .Z(n235) );
  NAND U466 ( .A(n236), .B(n237), .Z(n203) );
  NANDN U467 ( .B(n238), .A(n239), .Z(n236) );
  IV U468 ( .A(n206), .Z(n208) );
  XNOR U469 ( .A(n241), .B(n242), .Z(n112) );
  AND U470 ( .A(n127), .B(n244), .Z(n243) );
  XOR U471 ( .A(n214), .B(n245), .Z(n244) );
  XOR U472 ( .A(n245), .B(n215), .Z(n214) );
  OR U473 ( .A(n246), .B(n247), .Z(n215) );
  IV U474 ( .A(n242), .Z(n245) );
  XNOR U475 ( .A(n217), .B(n216), .Z(n242) );
  OR U476 ( .A(n248), .B(n249), .Z(n216) );
  XNOR U477 ( .A(n220), .B(n219), .Z(n217) );
  XOR U478 ( .A(n218), .B(n250), .Z(n219) );
  AND U479 ( .A(n251), .B(n252), .Z(n250) );
  OR U480 ( .A(n253), .B(n254), .Z(n252) );
  AND U481 ( .A(n255), .B(n256), .Z(n251) );
  NANDN U482 ( .B(n144), .A(n257), .Z(n256) );
  NAND U483 ( .A(n258), .B(n259), .Z(n255) );
  XNOR U484 ( .A(n231), .B(n264), .Z(n232) );
  AND U485 ( .A(n166), .B(n230), .Z(n264) );
  XOR U486 ( .A(n265), .B(n266), .Z(n231) );
  ANDN U487 ( .A(n267), .B(n268), .Z(n266) );
  XNOR U488 ( .A(n269), .B(n265), .Z(n267) );
  XOR U489 ( .A(n270), .B(n233), .Z(n263) );
  NAND U490 ( .A(n195), .B(n200), .Z(n233) );
  IV U491 ( .A(n223), .Z(n270) );
  XNOR U492 ( .A(n238), .B(n239), .Z(n227) );
  NANDN U493 ( .B(n145), .A(n274), .Z(n239) );
  XNOR U494 ( .A(n237), .B(n275), .Z(n238) );
  AND U495 ( .A(n234), .B(n165), .Z(n275) );
  ANDN U496 ( .A(n276), .B(n277), .Z(n237) );
  NANDN U497 ( .B(n278), .A(n279), .Z(n276) );
  XNOR U498 ( .A(n281), .B(n282), .Z(n113) );
  AND U499 ( .A(n127), .B(n284), .Z(n283) );
  XOR U500 ( .A(n246), .B(n285), .Z(n284) );
  XOR U501 ( .A(n285), .B(n247), .Z(n246) );
  OR U502 ( .A(n286), .B(n287), .Z(n247) );
  IV U503 ( .A(n282), .Z(n285) );
  XNOR U504 ( .A(n249), .B(n248), .Z(n282) );
  OR U505 ( .A(n288), .B(n289), .Z(n248) );
  XNOR U506 ( .A(n262), .B(n261), .Z(n249) );
  XOR U507 ( .A(n290), .B(n258), .Z(n261) );
  XNOR U508 ( .A(n291), .B(n253), .Z(n258) );
  NAND U509 ( .A(n257), .B(n166), .Z(n253) );
  NANDN U510 ( .B(n144), .A(n293), .Z(n292) );
  XNOR U511 ( .A(n259), .B(n260), .Z(n290) );
  XNOR U512 ( .A(n265), .B(n304), .Z(n268) );
  AND U513 ( .A(n200), .B(n230), .Z(n304) );
  XOR U514 ( .A(n305), .B(n306), .Z(n265) );
  ANDN U515 ( .A(n307), .B(n308), .Z(n306) );
  XNOR U516 ( .A(n309), .B(n305), .Z(n307) );
  XOR U517 ( .A(n310), .B(n269), .Z(n303) );
  NAND U518 ( .A(n195), .B(n234), .Z(n269) );
  IV U519 ( .A(n271), .Z(n310) );
  XNOR U520 ( .A(n278), .B(n279), .Z(n273) );
  NANDN U521 ( .B(n145), .A(n314), .Z(n279) );
  AND U522 ( .A(n274), .B(n165), .Z(n315) );
  NAND U523 ( .A(n316), .B(n317), .Z(n277) );
  NANDN U524 ( .B(n318), .A(n319), .Z(n316) );
  XNOR U525 ( .A(n321), .B(n322), .Z(n114) );
  XNOR U526 ( .A(n323), .B(n324), .Z(n321) );
  AND U527 ( .A(n127), .B(n325), .Z(n324) );
  XOR U528 ( .A(n286), .B(n326), .Z(n325) );
  XOR U529 ( .A(n326), .B(n287), .Z(n286) );
  OR U530 ( .A(n327), .B(n328), .Z(n287) );
  IV U531 ( .A(n322), .Z(n326) );
  XNOR U532 ( .A(n289), .B(n288), .Z(n322) );
  NANDN U533 ( .B(n329), .A(n330), .Z(n288) );
  XNOR U534 ( .A(n299), .B(n298), .Z(n289) );
  XOR U535 ( .A(n331), .B(n302), .Z(n298) );
  XNOR U536 ( .A(n295), .B(n296), .Z(n302) );
  NAND U537 ( .A(n257), .B(n200), .Z(n296) );
  XNOR U538 ( .A(n294), .B(n332), .Z(n295) );
  AND U539 ( .A(n166), .B(n293), .Z(n332) );
  XNOR U540 ( .A(n301), .B(n297), .Z(n331) );
  AND U541 ( .A(n340), .B(n341), .Z(n339) );
  NANDN U542 ( .B(n144), .A(n342), .Z(n341) );
  OR U543 ( .A(n343), .B(n344), .Z(n340) );
  XNOR U544 ( .A(n305), .B(n349), .Z(n308) );
  AND U545 ( .A(n234), .B(n230), .Z(n349) );
  XOR U546 ( .A(n353), .B(n309), .Z(n348) );
  NAND U547 ( .A(n195), .B(n274), .Z(n309) );
  IV U548 ( .A(n311), .Z(n353) );
  XNOR U549 ( .A(n318), .B(n319), .Z(n313) );
  NANDN U550 ( .B(n145), .A(n357), .Z(n319) );
  XNOR U551 ( .A(n317), .B(n358), .Z(n318) );
  AND U552 ( .A(n314), .B(n165), .Z(n358) );
  ANDN U553 ( .A(n359), .B(n360), .Z(n317) );
  NANDN U554 ( .B(n361), .A(n362), .Z(n359) );
  IV U555 ( .A(n320), .Z(n323) );
  XNOR U556 ( .A(n365), .B(n366), .Z(n364) );
  AND U557 ( .A(n127), .B(n367), .Z(n366) );
  XOR U558 ( .A(n327), .B(n370), .Z(n367) );
  XOR U559 ( .A(n370), .B(n328), .Z(n327) );
  OR U560 ( .A(n368), .B(n369), .Z(n328) );
  XNOR U561 ( .A(n329), .B(n330), .Z(n370) );
  XNOR U562 ( .A(n338), .B(n337), .Z(n329) );
  XOR U563 ( .A(n375), .B(n347), .Z(n337) );
  XNOR U564 ( .A(n334), .B(n335), .Z(n347) );
  NAND U565 ( .A(n257), .B(n234), .Z(n335) );
  XNOR U566 ( .A(n333), .B(n376), .Z(n334) );
  AND U567 ( .A(n200), .B(n293), .Z(n376) );
  XNOR U568 ( .A(n346), .B(n336), .Z(n375) );
  XNOR U569 ( .A(n383), .B(n345), .Z(n346) );
  XNOR U570 ( .A(n387), .B(n343), .Z(n383) );
  NAND U571 ( .A(n342), .B(n166), .Z(n343) );
  NANDN U572 ( .B(n144), .A(n389), .Z(n388) );
  XNOR U573 ( .A(n350), .B(n394), .Z(n351) );
  AND U574 ( .A(n274), .B(n230), .Z(n394) );
  XOR U575 ( .A(n395), .B(n396), .Z(n350) );
  ANDN U576 ( .A(n397), .B(n398), .Z(n396) );
  XNOR U577 ( .A(n399), .B(n395), .Z(n397) );
  XOR U578 ( .A(n400), .B(n352), .Z(n393) );
  NAND U579 ( .A(n195), .B(n314), .Z(n352) );
  IV U580 ( .A(n354), .Z(n400) );
  XNOR U581 ( .A(n361), .B(n362), .Z(n356) );
  NANDN U582 ( .B(n145), .A(n404), .Z(n362) );
  AND U583 ( .A(n357), .B(n165), .Z(n405) );
  NAND U584 ( .A(n406), .B(n407), .Z(n360) );
  NANDN U585 ( .B(n408), .A(n409), .Z(n406) );
  IV U586 ( .A(n363), .Z(n365) );
  XNOR U587 ( .A(n411), .B(n412), .Z(n116) );
  AND U588 ( .A(n127), .B(n414), .Z(n413) );
  XOR U589 ( .A(n368), .B(n415), .Z(n414) );
  XOR U590 ( .A(n415), .B(n369), .Z(n368) );
  OR U591 ( .A(n416), .B(n417), .Z(n369) );
  IV U592 ( .A(n412), .Z(n415) );
  XOR U593 ( .A(n374), .B(n373), .Z(n412) );
  XNOR U594 ( .A(n372), .B(n418), .Z(n373) );
  AND U595 ( .A(n371), .B(n419), .Z(n418) );
  AND U596 ( .A(n420), .B(n421), .Z(n419) );
  NANDN U597 ( .B(n144), .A(n422), .Z(n421) );
  OR U598 ( .A(n423), .B(n424), .Z(n420) );
  AND U599 ( .A(n425), .B(n426), .Z(n371) );
  NANDN U600 ( .B(n427), .A(n428), .Z(n426) );
  NANDN U601 ( .B(n429), .A(n430), .Z(n425) );
  XNOR U602 ( .A(n434), .B(n386), .Z(n381) );
  XNOR U603 ( .A(n378), .B(n379), .Z(n386) );
  NAND U604 ( .A(n257), .B(n274), .Z(n379) );
  XNOR U605 ( .A(n377), .B(n435), .Z(n378) );
  AND U606 ( .A(n234), .B(n293), .Z(n435) );
  XNOR U607 ( .A(n385), .B(n380), .Z(n434) );
  XNOR U608 ( .A(n390), .B(n443), .Z(n391) );
  AND U609 ( .A(n166), .B(n389), .Z(n443) );
  XOR U610 ( .A(n447), .B(n392), .Z(n442) );
  NAND U611 ( .A(n342), .B(n200), .Z(n392) );
  IV U612 ( .A(n384), .Z(n447) );
  XNOR U613 ( .A(n395), .B(n452), .Z(n398) );
  AND U614 ( .A(n314), .B(n230), .Z(n452) );
  XOR U615 ( .A(n453), .B(n454), .Z(n395) );
  ANDN U616 ( .A(n455), .B(n456), .Z(n454) );
  XNOR U617 ( .A(n457), .B(n453), .Z(n455) );
  XOR U618 ( .A(n458), .B(n399), .Z(n451) );
  NAND U619 ( .A(n195), .B(n357), .Z(n399) );
  IV U620 ( .A(n401), .Z(n458) );
  XNOR U621 ( .A(n408), .B(n409), .Z(n403) );
  NANDN U622 ( .B(n145), .A(n462), .Z(n409) );
  XNOR U623 ( .A(n407), .B(n463), .Z(n408) );
  AND U624 ( .A(n404), .B(n165), .Z(n463) );
  ANDN U625 ( .A(n464), .B(n465), .Z(n407) );
  NANDN U626 ( .B(n466), .A(n467), .Z(n464) );
  XNOR U627 ( .A(n469), .B(n470), .Z(n117) );
  AND U628 ( .A(n127), .B(n472), .Z(n471) );
  XOR U629 ( .A(n416), .B(n473), .Z(n472) );
  XOR U630 ( .A(n473), .B(n417), .Z(n416) );
  OR U631 ( .A(n474), .B(n475), .Z(n417) );
  IV U632 ( .A(n470), .Z(n473) );
  XOR U633 ( .A(n433), .B(n432), .Z(n470) );
  XOR U634 ( .A(n427), .B(n428), .Z(n424) );
  XOR U635 ( .A(n480), .B(n429), .Z(n427) );
  NAND U636 ( .A(n166), .B(n422), .Z(n429) );
  NANDN U637 ( .B(n430), .A(n481), .Z(n480) );
  NANDN U638 ( .B(n144), .A(n482), .Z(n481) );
  XOR U639 ( .A(n486), .B(n423), .Z(n476) );
  OR U640 ( .A(n487), .B(n488), .Z(n423) );
  IV U641 ( .A(n431), .Z(n486) );
  XNOR U642 ( .A(n492), .B(n450), .Z(n440) );
  XNOR U643 ( .A(n437), .B(n438), .Z(n450) );
  NAND U644 ( .A(n257), .B(n314), .Z(n438) );
  XNOR U645 ( .A(n436), .B(n493), .Z(n437) );
  AND U646 ( .A(n274), .B(n293), .Z(n493) );
  XNOR U647 ( .A(n449), .B(n439), .Z(n492) );
  XNOR U648 ( .A(n444), .B(n501), .Z(n445) );
  AND U649 ( .A(n200), .B(n389), .Z(n501) );
  XOR U650 ( .A(n505), .B(n446), .Z(n500) );
  NAND U651 ( .A(n342), .B(n234), .Z(n446) );
  IV U652 ( .A(n448), .Z(n505) );
  XNOR U653 ( .A(n453), .B(n510), .Z(n456) );
  AND U654 ( .A(n357), .B(n230), .Z(n510) );
  XOR U655 ( .A(n511), .B(n512), .Z(n453) );
  ANDN U656 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U657 ( .A(n515), .B(n511), .Z(n513) );
  XOR U658 ( .A(n516), .B(n457), .Z(n509) );
  NAND U659 ( .A(n195), .B(n404), .Z(n457) );
  IV U660 ( .A(n459), .Z(n516) );
  XNOR U661 ( .A(n466), .B(n467), .Z(n461) );
  NANDN U662 ( .B(n145), .A(n520), .Z(n467) );
  AND U663 ( .A(n462), .B(n165), .Z(n521) );
  NAND U664 ( .A(n522), .B(n523), .Z(n465) );
  NANDN U665 ( .B(n524), .A(n525), .Z(n522) );
  XNOR U666 ( .A(n527), .B(n528), .Z(n118) );
  AND U667 ( .A(n127), .B(n530), .Z(n529) );
  XOR U668 ( .A(n474), .B(n531), .Z(n530) );
  XOR U669 ( .A(n531), .B(n475), .Z(n474) );
  OR U670 ( .A(n532), .B(n533), .Z(n475) );
  IV U671 ( .A(n528), .Z(n531) );
  XOR U672 ( .A(n491), .B(n490), .Z(n528) );
  XOR U673 ( .A(n534), .B(n487), .Z(n490) );
  XOR U674 ( .A(n479), .B(n478), .Z(n487) );
  XOR U675 ( .A(n477), .B(n535), .Z(n478) );
  AND U676 ( .A(n536), .B(n537), .Z(n535) );
  NANDN U677 ( .B(n144), .A(n538), .Z(n537) );
  OR U678 ( .A(n539), .B(n540), .Z(n536) );
  NAND U679 ( .A(n200), .B(n422), .Z(n485) );
  XNOR U680 ( .A(n483), .B(n544), .Z(n484) );
  AND U681 ( .A(n482), .B(n166), .Z(n544) );
  NANDN U682 ( .B(n548), .A(n549), .Z(n488) );
  XNOR U683 ( .A(n553), .B(n508), .Z(n498) );
  XNOR U684 ( .A(n495), .B(n496), .Z(n508) );
  NAND U685 ( .A(n257), .B(n357), .Z(n496) );
  XNOR U686 ( .A(n494), .B(n554), .Z(n495) );
  AND U687 ( .A(n314), .B(n293), .Z(n554) );
  XNOR U688 ( .A(n507), .B(n497), .Z(n553) );
  XNOR U689 ( .A(n502), .B(n562), .Z(n503) );
  AND U690 ( .A(n234), .B(n389), .Z(n562) );
  XOR U691 ( .A(n566), .B(n504), .Z(n561) );
  NAND U692 ( .A(n342), .B(n274), .Z(n504) );
  IV U693 ( .A(n506), .Z(n566) );
  XNOR U694 ( .A(n511), .B(n571), .Z(n514) );
  AND U695 ( .A(n404), .B(n230), .Z(n571) );
  XOR U696 ( .A(n572), .B(n573), .Z(n511) );
  ANDN U697 ( .A(n574), .B(n575), .Z(n573) );
  XNOR U698 ( .A(n576), .B(n572), .Z(n574) );
  XOR U699 ( .A(n577), .B(n515), .Z(n570) );
  NAND U700 ( .A(n195), .B(n462), .Z(n515) );
  IV U701 ( .A(n517), .Z(n577) );
  XNOR U702 ( .A(n524), .B(n525), .Z(n519) );
  NANDN U703 ( .B(n145), .A(n581), .Z(n525) );
  XNOR U704 ( .A(n523), .B(n582), .Z(n524) );
  AND U705 ( .A(n520), .B(n165), .Z(n582) );
  ANDN U706 ( .A(n583), .B(n584), .Z(n523) );
  NANDN U707 ( .B(n585), .A(n586), .Z(n583) );
  XNOR U708 ( .A(n588), .B(n589), .Z(n119) );
  AND U709 ( .A(n127), .B(n591), .Z(n590) );
  XOR U710 ( .A(n532), .B(n592), .Z(n591) );
  XOR U711 ( .A(n592), .B(n533), .Z(n532) );
  OR U712 ( .A(n593), .B(n594), .Z(n533) );
  IV U713 ( .A(n589), .Z(n592) );
  XOR U714 ( .A(n552), .B(n551), .Z(n589) );
  XOR U715 ( .A(n595), .B(n548), .Z(n551) );
  XOR U716 ( .A(n543), .B(n542), .Z(n548) );
  XNOR U717 ( .A(n600), .B(n539), .Z(n596) );
  NAND U718 ( .A(n166), .B(n538), .Z(n539) );
  NANDN U719 ( .B(n144), .A(n602), .Z(n601) );
  NAND U720 ( .A(n234), .B(n422), .Z(n547) );
  XNOR U721 ( .A(n545), .B(n606), .Z(n546) );
  AND U722 ( .A(n482), .B(n200), .Z(n606) );
  XNOR U723 ( .A(n549), .B(n550), .Z(n595) );
  XNOR U724 ( .A(n616), .B(n569), .Z(n559) );
  XNOR U725 ( .A(n556), .B(n557), .Z(n569) );
  NAND U726 ( .A(n257), .B(n404), .Z(n557) );
  XNOR U727 ( .A(n555), .B(n617), .Z(n556) );
  AND U728 ( .A(n357), .B(n293), .Z(n617) );
  XNOR U729 ( .A(n568), .B(n558), .Z(n616) );
  XNOR U730 ( .A(n563), .B(n625), .Z(n564) );
  AND U731 ( .A(n274), .B(n389), .Z(n625) );
  XOR U732 ( .A(n626), .B(n627), .Z(n563) );
  ANDN U733 ( .A(n628), .B(n629), .Z(n627) );
  XNOR U734 ( .A(n630), .B(n626), .Z(n628) );
  XOR U735 ( .A(n631), .B(n565), .Z(n624) );
  NAND U736 ( .A(n342), .B(n314), .Z(n565) );
  IV U737 ( .A(n567), .Z(n631) );
  XNOR U738 ( .A(n572), .B(n636), .Z(n575) );
  AND U739 ( .A(n462), .B(n230), .Z(n636) );
  XOR U740 ( .A(n637), .B(n638), .Z(n572) );
  ANDN U741 ( .A(n639), .B(n640), .Z(n638) );
  XNOR U742 ( .A(n641), .B(n637), .Z(n639) );
  XOR U743 ( .A(n642), .B(n576), .Z(n635) );
  NAND U744 ( .A(n195), .B(n520), .Z(n576) );
  IV U745 ( .A(n578), .Z(n642) );
  XNOR U746 ( .A(n585), .B(n586), .Z(n580) );
  OR U747 ( .A(n646), .B(n145), .Z(n586) );
  AND U748 ( .A(n581), .B(n165), .Z(n647) );
  NAND U749 ( .A(n648), .B(n649), .Z(n584) );
  NANDN U750 ( .B(n650), .A(n651), .Z(n648) );
  XNOR U751 ( .A(n653), .B(n654), .Z(n120) );
  XOR U752 ( .A(n652), .B(n655), .Z(n653) );
  AND U753 ( .A(n127), .B(n656), .Z(n655) );
  XOR U754 ( .A(n593), .B(n657), .Z(n656) );
  XOR U755 ( .A(n657), .B(n594), .Z(n593) );
  NANDN U756 ( .B(n658), .A(n659), .Z(n594) );
  IV U757 ( .A(n654), .Z(n657) );
  XOR U758 ( .A(n612), .B(n611), .Z(n654) );
  XNOR U759 ( .A(n660), .B(n615), .Z(n611) );
  XNOR U760 ( .A(n603), .B(n662), .Z(n604) );
  AND U761 ( .A(n602), .B(n166), .Z(n662) );
  XOR U762 ( .A(n666), .B(n605), .Z(n661) );
  NAND U763 ( .A(n200), .B(n538), .Z(n605) );
  IV U764 ( .A(n597), .Z(n666) );
  XNOR U765 ( .A(n608), .B(n609), .Z(n599) );
  NAND U766 ( .A(n274), .B(n422), .Z(n609) );
  XNOR U767 ( .A(n607), .B(n670), .Z(n608) );
  AND U768 ( .A(n482), .B(n234), .Z(n670) );
  XNOR U769 ( .A(n614), .B(n610), .Z(n660) );
  AND U770 ( .A(n678), .B(n679), .Z(n677) );
  OR U771 ( .A(n680), .B(n681), .Z(n679) );
  AND U772 ( .A(n682), .B(n683), .Z(n678) );
  NANDN U773 ( .B(n144), .A(n684), .Z(n683) );
  NANDN U774 ( .B(n685), .A(n686), .Z(n682) );
  XNOR U775 ( .A(n690), .B(n634), .Z(n622) );
  XNOR U776 ( .A(n619), .B(n620), .Z(n634) );
  NAND U777 ( .A(n257), .B(n462), .Z(n620) );
  XNOR U778 ( .A(n618), .B(n691), .Z(n619) );
  AND U779 ( .A(n404), .B(n293), .Z(n691) );
  XNOR U780 ( .A(n633), .B(n621), .Z(n690) );
  XNOR U781 ( .A(n626), .B(n699), .Z(n629) );
  AND U782 ( .A(n314), .B(n389), .Z(n699) );
  XOR U783 ( .A(n703), .B(n630), .Z(n698) );
  NAND U784 ( .A(n342), .B(n357), .Z(n630) );
  IV U785 ( .A(n632), .Z(n703) );
  XNOR U786 ( .A(n637), .B(n708), .Z(n640) );
  AND U787 ( .A(n520), .B(n230), .Z(n708) );
  XOR U788 ( .A(n709), .B(n710), .Z(n637) );
  ANDN U789 ( .A(n711), .B(n712), .Z(n710) );
  XNOR U790 ( .A(n713), .B(n709), .Z(n711) );
  XOR U791 ( .A(n714), .B(n641), .Z(n707) );
  NAND U792 ( .A(n195), .B(n581), .Z(n641) );
  IV U793 ( .A(n643), .Z(n714) );
  XNOR U794 ( .A(n650), .B(n651), .Z(n645) );
  OR U795 ( .A(n718), .B(n145), .Z(n651) );
  XNOR U796 ( .A(n649), .B(n719), .Z(n650) );
  ANDN U797 ( .A(n165), .B(n646), .Z(n719) );
  ANDN U798 ( .A(n720), .B(n721), .Z(n649) );
  NANDN U799 ( .B(n722), .A(n723), .Z(n720) );
  XOR U800 ( .A(n725), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U801 ( .A(n726), .B(n727), .Z(n725) );
  XNOR U802 ( .A(n728), .B(n724), .Z(n726) );
  NANDN U803 ( .B(n659), .A(\_MxM/Y0[0] ), .Z(n724) );
  NAND U804 ( .A(n729), .B(n127), .Z(n728) );
  XOR U805 ( .A(e_input[15]), .B(g_input[15]), .Z(n127) );
  XNOR U806 ( .A(n658), .B(n727), .Z(n729) );
  XOR U807 ( .A(n659), .B(n727), .Z(n658) );
  XOR U808 ( .A(n676), .B(n675), .Z(n727) );
  XNOR U809 ( .A(n730), .B(n689), .Z(n675) );
  XNOR U810 ( .A(n663), .B(n732), .Z(n664) );
  AND U811 ( .A(n602), .B(n200), .Z(n732) );
  XOR U812 ( .A(n736), .B(n665), .Z(n731) );
  NAND U813 ( .A(n234), .B(n538), .Z(n665) );
  IV U814 ( .A(n667), .Z(n736) );
  XNOR U815 ( .A(n672), .B(n673), .Z(n669) );
  NAND U816 ( .A(n314), .B(n422), .Z(n673) );
  XNOR U817 ( .A(n671), .B(n740), .Z(n672) );
  AND U818 ( .A(n482), .B(n274), .Z(n740) );
  XNOR U819 ( .A(n688), .B(n674), .Z(n730) );
  XNOR U820 ( .A(n747), .B(n685), .Z(n688) );
  XOR U821 ( .A(n748), .B(n680), .Z(n685) );
  NAND U822 ( .A(n166), .B(n684), .Z(n680) );
  NANDN U823 ( .B(n144), .A(n750), .Z(n749) );
  XNOR U824 ( .A(n686), .B(n687), .Z(n747) );
  XNOR U825 ( .A(n759), .B(n706), .Z(n696) );
  XNOR U826 ( .A(n693), .B(n694), .Z(n706) );
  NAND U827 ( .A(n257), .B(n520), .Z(n694) );
  XNOR U828 ( .A(n692), .B(n760), .Z(n693) );
  AND U829 ( .A(n462), .B(n293), .Z(n760) );
  XNOR U830 ( .A(n705), .B(n695), .Z(n759) );
  XNOR U831 ( .A(n700), .B(n768), .Z(n701) );
  AND U832 ( .A(n357), .B(n389), .Z(n768) );
  XOR U833 ( .A(n769), .B(n770), .Z(n700) );
  ANDN U834 ( .A(n771), .B(n772), .Z(n770) );
  XNOR U835 ( .A(n773), .B(n769), .Z(n771) );
  XOR U836 ( .A(n774), .B(n702), .Z(n767) );
  NAND U837 ( .A(n342), .B(n404), .Z(n702) );
  IV U838 ( .A(n704), .Z(n774) );
  XNOR U839 ( .A(n709), .B(n779), .Z(n712) );
  AND U840 ( .A(n581), .B(n230), .Z(n779) );
  XOR U841 ( .A(n780), .B(n781), .Z(n709) );
  ANDN U842 ( .A(n782), .B(n783), .Z(n781) );
  XNOR U843 ( .A(n784), .B(n780), .Z(n782) );
  XOR U844 ( .A(n785), .B(n713), .Z(n778) );
  NANDN U845 ( .B(n646), .A(n195), .Z(n713) );
  IV U846 ( .A(n715), .Z(n785) );
  XNOR U847 ( .A(n722), .B(n723), .Z(n717) );
  NANDN U848 ( .B(n145), .A(n789), .Z(n723) );
  ANDN U849 ( .A(n165), .B(n718), .Z(n790) );
  NAND U850 ( .A(n791), .B(n792), .Z(n721) );
  NANDN U851 ( .B(n793), .A(n794), .Z(n791) );
  XOR U852 ( .A(n746), .B(n745), .Z(n659) );
  XNOR U853 ( .A(n795), .B(n756), .Z(n745) );
  XNOR U854 ( .A(n733), .B(n797), .Z(n734) );
  AND U855 ( .A(n602), .B(n234), .Z(n797) );
  XOR U856 ( .A(n798), .B(n799), .Z(n733) );
  ANDN U857 ( .A(n800), .B(n801), .Z(n799) );
  XNOR U858 ( .A(n802), .B(n798), .Z(n800) );
  XOR U859 ( .A(n803), .B(n735), .Z(n796) );
  NAND U860 ( .A(n274), .B(n538), .Z(n735) );
  IV U861 ( .A(n737), .Z(n803) );
  XNOR U862 ( .A(n742), .B(n743), .Z(n739) );
  NAND U863 ( .A(n357), .B(n422), .Z(n743) );
  XNOR U864 ( .A(n741), .B(n807), .Z(n742) );
  AND U865 ( .A(n482), .B(n314), .Z(n807) );
  XNOR U866 ( .A(n755), .B(n744), .Z(n795) );
  XOR U867 ( .A(n811), .B(n812), .Z(n744) );
  XNOR U868 ( .A(n813), .B(n758), .Z(n755) );
  NAND U869 ( .A(n200), .B(n684), .Z(n753) );
  XNOR U870 ( .A(n751), .B(n814), .Z(n752) );
  AND U871 ( .A(n750), .B(n166), .Z(n814) );
  XNOR U872 ( .A(n757), .B(n754), .Z(n813) );
  XOR U873 ( .A(n818), .B(n819), .Z(n754) );
  AND U874 ( .A(n820), .B(n821), .Z(n819) );
  XOR U875 ( .A(n822), .B(n823), .Z(n821) );
  XOR U876 ( .A(n818), .B(n824), .Z(n823) );
  XOR U877 ( .A(n805), .B(n825), .Z(n820) );
  XOR U878 ( .A(n818), .B(n806), .Z(n825) );
  NAND U879 ( .A(n422), .B(n404), .Z(n810) );
  XNOR U880 ( .A(n808), .B(n826), .Z(n809) );
  AND U881 ( .A(n482), .B(n357), .Z(n826) );
  XNOR U882 ( .A(n798), .B(n831), .Z(n801) );
  AND U883 ( .A(n602), .B(n274), .Z(n831) );
  XOR U884 ( .A(n835), .B(n802), .Z(n830) );
  NAND U885 ( .A(n314), .B(n538), .Z(n802) );
  IV U886 ( .A(n804), .Z(n835) );
  XOR U887 ( .A(n839), .B(n840), .Z(n818) );
  AND U888 ( .A(n841), .B(n842), .Z(n840) );
  XOR U889 ( .A(n843), .B(n844), .Z(n842) );
  XOR U890 ( .A(n839), .B(n845), .Z(n844) );
  XOR U891 ( .A(n837), .B(n846), .Z(n841) );
  XOR U892 ( .A(n839), .B(n838), .Z(n846) );
  NAND U893 ( .A(n422), .B(n462), .Z(n829) );
  XNOR U894 ( .A(n827), .B(n847), .Z(n828) );
  AND U895 ( .A(n404), .B(n482), .Z(n847) );
  XNOR U896 ( .A(n832), .B(n852), .Z(n833) );
  AND U897 ( .A(n602), .B(n314), .Z(n852) );
  XOR U898 ( .A(n853), .B(n854), .Z(n832) );
  ANDN U899 ( .A(n855), .B(n856), .Z(n854) );
  XNOR U900 ( .A(n857), .B(n853), .Z(n855) );
  XOR U901 ( .A(n858), .B(n834), .Z(n851) );
  NAND U902 ( .A(n357), .B(n538), .Z(n834) );
  IV U903 ( .A(n836), .Z(n858) );
  XOR U904 ( .A(n862), .B(n863), .Z(n839) );
  AND U905 ( .A(n864), .B(n865), .Z(n863) );
  XOR U906 ( .A(n866), .B(n867), .Z(n865) );
  XOR U907 ( .A(n862), .B(n868), .Z(n867) );
  XOR U908 ( .A(n860), .B(n869), .Z(n864) );
  XOR U909 ( .A(n862), .B(n861), .Z(n869) );
  NAND U910 ( .A(n422), .B(n520), .Z(n850) );
  XNOR U911 ( .A(n848), .B(n870), .Z(n849) );
  AND U912 ( .A(n462), .B(n482), .Z(n870) );
  XOR U913 ( .A(n871), .B(n872), .Z(n848) );
  ANDN U914 ( .A(n873), .B(n874), .Z(n872) );
  XNOR U915 ( .A(n875), .B(n871), .Z(n873) );
  XNOR U916 ( .A(n876), .B(n877), .Z(n860) );
  IV U917 ( .A(n856), .Z(n877) );
  XNOR U918 ( .A(n853), .B(n878), .Z(n856) );
  AND U919 ( .A(n602), .B(n357), .Z(n878) );
  XOR U920 ( .A(n879), .B(n880), .Z(n853) );
  ANDN U921 ( .A(n881), .B(n882), .Z(n880) );
  XNOR U922 ( .A(n883), .B(n879), .Z(n881) );
  XOR U923 ( .A(n884), .B(n857), .Z(n876) );
  NAND U924 ( .A(n538), .B(n404), .Z(n857) );
  IV U925 ( .A(n859), .Z(n884) );
  XOR U926 ( .A(n888), .B(n889), .Z(n862) );
  AND U927 ( .A(n890), .B(n891), .Z(n889) );
  XOR U928 ( .A(n892), .B(n893), .Z(n891) );
  XOR U929 ( .A(n888), .B(n894), .Z(n893) );
  XOR U930 ( .A(n886), .B(n895), .Z(n890) );
  XOR U931 ( .A(n888), .B(n887), .Z(n895) );
  XNOR U932 ( .A(n896), .B(n875), .Z(n887) );
  NAND U933 ( .A(n422), .B(n581), .Z(n875) );
  IV U934 ( .A(n874), .Z(n896) );
  XNOR U935 ( .A(n871), .B(n897), .Z(n874) );
  AND U936 ( .A(n520), .B(n482), .Z(n897) );
  XOR U937 ( .A(n898), .B(n899), .Z(n871) );
  ANDN U938 ( .A(n900), .B(n901), .Z(n899) );
  XNOR U939 ( .A(n902), .B(n898), .Z(n900) );
  XNOR U940 ( .A(n903), .B(n904), .Z(n886) );
  IV U941 ( .A(n882), .Z(n904) );
  XNOR U942 ( .A(n879), .B(n905), .Z(n882) );
  AND U943 ( .A(n404), .B(n602), .Z(n905) );
  XOR U944 ( .A(n906), .B(n907), .Z(n879) );
  ANDN U945 ( .A(n908), .B(n909), .Z(n907) );
  XNOR U946 ( .A(n910), .B(n906), .Z(n908) );
  XOR U947 ( .A(n911), .B(n883), .Z(n903) );
  NAND U948 ( .A(n538), .B(n462), .Z(n883) );
  IV U949 ( .A(n885), .Z(n911) );
  XOR U950 ( .A(n915), .B(n916), .Z(n888) );
  AND U951 ( .A(n917), .B(n918), .Z(n916) );
  XOR U952 ( .A(n919), .B(n920), .Z(n918) );
  XOR U953 ( .A(n915), .B(n921), .Z(n920) );
  XOR U954 ( .A(n913), .B(n922), .Z(n917) );
  XOR U955 ( .A(n915), .B(n914), .Z(n922) );
  XNOR U956 ( .A(n923), .B(n902), .Z(n914) );
  NANDN U957 ( .B(n646), .A(n422), .Z(n902) );
  IV U958 ( .A(n901), .Z(n923) );
  XNOR U959 ( .A(n898), .B(n924), .Z(n901) );
  AND U960 ( .A(n581), .B(n482), .Z(n924) );
  XOR U961 ( .A(n925), .B(n926), .Z(n898) );
  ANDN U962 ( .A(n927), .B(n928), .Z(n926) );
  XNOR U963 ( .A(n929), .B(n925), .Z(n927) );
  XNOR U964 ( .A(n930), .B(n931), .Z(n913) );
  IV U965 ( .A(n909), .Z(n931) );
  XNOR U966 ( .A(n906), .B(n932), .Z(n909) );
  AND U967 ( .A(n462), .B(n602), .Z(n932) );
  XOR U968 ( .A(n933), .B(n934), .Z(n906) );
  ANDN U969 ( .A(n935), .B(n936), .Z(n934) );
  XNOR U970 ( .A(n937), .B(n933), .Z(n935) );
  XOR U971 ( .A(n938), .B(n910), .Z(n930) );
  NAND U972 ( .A(n538), .B(n520), .Z(n910) );
  IV U973 ( .A(n912), .Z(n938) );
  XOR U974 ( .A(n942), .B(n943), .Z(n915) );
  AND U975 ( .A(n944), .B(n945), .Z(n943) );
  XOR U976 ( .A(n946), .B(n947), .Z(n945) );
  XOR U977 ( .A(n942), .B(n948), .Z(n947) );
  XOR U978 ( .A(n940), .B(n949), .Z(n944) );
  XOR U979 ( .A(n942), .B(n941), .Z(n949) );
  XNOR U980 ( .A(n950), .B(n929), .Z(n941) );
  NANDN U981 ( .B(n718), .A(n422), .Z(n929) );
  IV U982 ( .A(n928), .Z(n950) );
  XNOR U983 ( .A(n925), .B(n951), .Z(n928) );
  ANDN U984 ( .A(n482), .B(n646), .Z(n951) );
  XOR U985 ( .A(n952), .B(n953), .Z(n925) );
  ANDN U986 ( .A(n954), .B(n955), .Z(n953) );
  XNOR U987 ( .A(n956), .B(n952), .Z(n954) );
  XNOR U988 ( .A(n957), .B(n958), .Z(n940) );
  IV U989 ( .A(n936), .Z(n958) );
  XNOR U990 ( .A(n933), .B(n959), .Z(n936) );
  AND U991 ( .A(n520), .B(n602), .Z(n959) );
  XOR U992 ( .A(n960), .B(n961), .Z(n933) );
  ANDN U993 ( .A(n962), .B(n963), .Z(n961) );
  XNOR U994 ( .A(n964), .B(n960), .Z(n962) );
  XOR U995 ( .A(n965), .B(n937), .Z(n957) );
  NAND U996 ( .A(n538), .B(n581), .Z(n937) );
  IV U997 ( .A(n939), .Z(n965) );
  XOR U998 ( .A(n969), .B(n970), .Z(n942) );
  AND U999 ( .A(n971), .B(n972), .Z(n970) );
  XOR U1000 ( .A(n973), .B(n974), .Z(n972) );
  XOR U1001 ( .A(n969), .B(n975), .Z(n974) );
  XOR U1002 ( .A(n967), .B(n976), .Z(n971) );
  XOR U1003 ( .A(n969), .B(n968), .Z(n976) );
  XNOR U1004 ( .A(n977), .B(n956), .Z(n968) );
  NAND U1005 ( .A(n422), .B(n789), .Z(n956) );
  IV U1006 ( .A(n955), .Z(n977) );
  XNOR U1007 ( .A(n952), .B(n978), .Z(n955) );
  ANDN U1008 ( .A(n482), .B(n718), .Z(n978) );
  XOR U1009 ( .A(n979), .B(n980), .Z(n952) );
  ANDN U1010 ( .A(n981), .B(n982), .Z(n980) );
  XNOR U1011 ( .A(n983), .B(n979), .Z(n981) );
  XNOR U1012 ( .A(n984), .B(n985), .Z(n967) );
  IV U1013 ( .A(n963), .Z(n985) );
  XNOR U1014 ( .A(n960), .B(n986), .Z(n963) );
  AND U1015 ( .A(n581), .B(n602), .Z(n986) );
  XOR U1016 ( .A(n987), .B(n988), .Z(n960) );
  ANDN U1017 ( .A(n989), .B(n990), .Z(n988) );
  XNOR U1018 ( .A(n991), .B(n987), .Z(n989) );
  XOR U1019 ( .A(n992), .B(n964), .Z(n984) );
  NANDN U1020 ( .B(n646), .A(n538), .Z(n964) );
  IV U1021 ( .A(n966), .Z(n992) );
  XOR U1022 ( .A(n997), .B(n998), .Z(n812) );
  XNOR U1023 ( .A(n999), .B(n996), .Z(n997) );
  XNOR U1024 ( .A(n987), .B(n1001), .Z(n990) );
  ANDN U1025 ( .A(n602), .B(n646), .Z(n1001) );
  XOR U1026 ( .A(n1004), .B(n1002), .Z(n1003) );
  ANDN U1027 ( .A(n602), .B(n718), .Z(n1004) );
  AND U1028 ( .A(n789), .B(n538), .Z(n1005) );
  XOR U1029 ( .A(n1006), .B(n1007), .Z(n1002) );
  ANDN U1030 ( .A(n1008), .B(n1009), .Z(n1007) );
  XNOR U1031 ( .A(n1010), .B(n1006), .Z(n1008) );
  XOR U1032 ( .A(n1011), .B(n991), .Z(n1000) );
  NANDN U1033 ( .B(n718), .A(n538), .Z(n991) );
  IV U1034 ( .A(n993), .Z(n1011) );
  NAND U1035 ( .A(n538), .B(n1012), .Z(n1010) );
  XNOR U1036 ( .A(n1006), .B(n1013), .Z(n1009) );
  AND U1037 ( .A(n789), .B(n602), .Z(n1013) );
  AND U1038 ( .A(n1014), .B(g_input[0]), .Z(n1006) );
  NANDN U1039 ( .B(n538), .A(n1015), .Z(n1014) );
  NAND U1040 ( .A(n1012), .B(n602), .Z(n1015) );
  XNOR U1041 ( .A(n982), .B(n983), .Z(n995) );
  NAND U1042 ( .A(n422), .B(n1012), .Z(n983) );
  XNOR U1043 ( .A(n979), .B(n1018), .Z(n982) );
  AND U1044 ( .A(n789), .B(n482), .Z(n1018) );
  AND U1045 ( .A(n1019), .B(g_input[0]), .Z(n979) );
  NANDN U1046 ( .B(n422), .A(n1020), .Z(n1019) );
  NAND U1047 ( .A(n1012), .B(n482), .Z(n1020) );
  XOR U1048 ( .A(n1023), .B(n1024), .Z(n996) );
  XOR U1049 ( .A(n1025), .B(n1026), .Z(n757) );
  AND U1050 ( .A(n1027), .B(n1028), .Z(n1026) );
  NANDN U1051 ( .B(n144), .A(n1029), .Z(n1028) );
  NANDN U1052 ( .B(n1030), .A(n1031), .Z(n144) );
  AND U1053 ( .A(n1032), .B(g_input[15]), .Z(n1031) );
  OR U1054 ( .A(n1033), .B(n1034), .Z(n1027) );
  AND U1055 ( .A(n824), .B(n1037), .Z(n1036) );
  XNOR U1056 ( .A(n1035), .B(n822), .Z(n1037) );
  NAND U1057 ( .A(n234), .B(n684), .Z(n817) );
  XNOR U1058 ( .A(n815), .B(n1038), .Z(n816) );
  AND U1059 ( .A(n750), .B(n200), .Z(n1038) );
  XOR U1060 ( .A(n1046), .B(n1033), .Z(n1042) );
  NAND U1061 ( .A(n166), .B(n1029), .Z(n1033) );
  IV U1062 ( .A(n1035), .Z(n1046) );
  NAND U1063 ( .A(n274), .B(n684), .Z(n1041) );
  XNOR U1064 ( .A(n1039), .B(n1048), .Z(n1040) );
  AND U1065 ( .A(n750), .B(n234), .Z(n1048) );
  XNOR U1066 ( .A(n1052), .B(n1053), .Z(n845) );
  IV U1067 ( .A(n1044), .Z(n1053) );
  XNOR U1068 ( .A(n1043), .B(n1054), .Z(n1044) );
  AND U1069 ( .A(n166), .B(e_input[0]), .Z(n1054) );
  XNOR U1070 ( .A(n1032), .B(g_input[14]), .Z(n1030) );
  NOR U1071 ( .A(n1055), .B(n1056), .Z(n1032) );
  XOR U1072 ( .A(n1060), .B(n1045), .Z(n1052) );
  NAND U1073 ( .A(n200), .B(n1029), .Z(n1045) );
  IV U1074 ( .A(n1047), .Z(n1060) );
  NAND U1075 ( .A(n314), .B(n684), .Z(n1051) );
  XNOR U1076 ( .A(n1049), .B(n1062), .Z(n1050) );
  AND U1077 ( .A(n750), .B(n274), .Z(n1062) );
  XOR U1078 ( .A(n1063), .B(n1064), .Z(n1049) );
  ANDN U1079 ( .A(n1065), .B(n1066), .Z(n1064) );
  XNOR U1080 ( .A(n1067), .B(n1063), .Z(n1065) );
  XNOR U1081 ( .A(n1057), .B(n1069), .Z(n1058) );
  AND U1082 ( .A(n200), .B(e_input[0]), .Z(n1069) );
  XOR U1083 ( .A(n1055), .B(g_input[13]), .Z(n1056) );
  NANDN U1084 ( .B(n1070), .A(n1071), .Z(n1055) );
  XOR U1085 ( .A(n1075), .B(n1059), .Z(n1068) );
  NAND U1086 ( .A(n234), .B(n1029), .Z(n1059) );
  IV U1087 ( .A(n1061), .Z(n1075) );
  XNOR U1088 ( .A(n1077), .B(n1067), .Z(n892) );
  NAND U1089 ( .A(n357), .B(n684), .Z(n1067) );
  IV U1090 ( .A(n1066), .Z(n1077) );
  XNOR U1091 ( .A(n1063), .B(n1078), .Z(n1066) );
  AND U1092 ( .A(n750), .B(n314), .Z(n1078) );
  XOR U1093 ( .A(n1079), .B(n1080), .Z(n1063) );
  ANDN U1094 ( .A(n1081), .B(n1082), .Z(n1080) );
  XNOR U1095 ( .A(n1083), .B(n1079), .Z(n1081) );
  XNOR U1096 ( .A(n1084), .B(n1085), .Z(n894) );
  IV U1097 ( .A(n1073), .Z(n1085) );
  XNOR U1098 ( .A(n1072), .B(n1086), .Z(n1073) );
  AND U1099 ( .A(n234), .B(e_input[0]), .Z(n1086) );
  XNOR U1100 ( .A(n1071), .B(g_input[12]), .Z(n1070) );
  NOR U1101 ( .A(n1087), .B(n1088), .Z(n1071) );
  XOR U1102 ( .A(n1092), .B(n1074), .Z(n1084) );
  NAND U1103 ( .A(n274), .B(n1029), .Z(n1074) );
  IV U1104 ( .A(n1076), .Z(n1092) );
  XNOR U1105 ( .A(n1094), .B(n1083), .Z(n919) );
  NAND U1106 ( .A(n404), .B(n684), .Z(n1083) );
  IV U1107 ( .A(n1082), .Z(n1094) );
  XNOR U1108 ( .A(n1079), .B(n1095), .Z(n1082) );
  AND U1109 ( .A(n750), .B(n357), .Z(n1095) );
  XOR U1110 ( .A(n1096), .B(n1097), .Z(n1079) );
  ANDN U1111 ( .A(n1098), .B(n1099), .Z(n1097) );
  XNOR U1112 ( .A(n1100), .B(n1096), .Z(n1098) );
  XNOR U1113 ( .A(n1101), .B(n1102), .Z(n921) );
  IV U1114 ( .A(n1090), .Z(n1102) );
  XNOR U1115 ( .A(n1089), .B(n1103), .Z(n1090) );
  AND U1116 ( .A(n274), .B(e_input[0]), .Z(n1103) );
  XOR U1117 ( .A(n1087), .B(g_input[11]), .Z(n1088) );
  NANDN U1118 ( .B(n1104), .A(n1105), .Z(n1087) );
  XOR U1119 ( .A(n1106), .B(n1107), .Z(n1089) );
  ANDN U1120 ( .A(n1108), .B(n1109), .Z(n1107) );
  XNOR U1121 ( .A(n1110), .B(n1106), .Z(n1108) );
  XOR U1122 ( .A(n1111), .B(n1091), .Z(n1101) );
  NAND U1123 ( .A(n314), .B(n1029), .Z(n1091) );
  IV U1124 ( .A(n1093), .Z(n1111) );
  XNOR U1125 ( .A(n1113), .B(n1100), .Z(n946) );
  NAND U1126 ( .A(n462), .B(n684), .Z(n1100) );
  IV U1127 ( .A(n1099), .Z(n1113) );
  XNOR U1128 ( .A(n1096), .B(n1114), .Z(n1099) );
  AND U1129 ( .A(n750), .B(n404), .Z(n1114) );
  XOR U1130 ( .A(n1115), .B(n1116), .Z(n1096) );
  ANDN U1131 ( .A(n1117), .B(n1118), .Z(n1116) );
  XNOR U1132 ( .A(n1119), .B(n1115), .Z(n1117) );
  XNOR U1133 ( .A(n1120), .B(n1121), .Z(n948) );
  IV U1134 ( .A(n1109), .Z(n1121) );
  XNOR U1135 ( .A(n1106), .B(n1122), .Z(n1109) );
  AND U1136 ( .A(n314), .B(e_input[0]), .Z(n1122) );
  XNOR U1137 ( .A(n1105), .B(g_input[10]), .Z(n1104) );
  NOR U1138 ( .A(n1123), .B(n1124), .Z(n1105) );
  XOR U1139 ( .A(n1128), .B(n1110), .Z(n1120) );
  NAND U1140 ( .A(n357), .B(n1029), .Z(n1110) );
  IV U1141 ( .A(n1112), .Z(n1128) );
  XNOR U1142 ( .A(n1130), .B(n1119), .Z(n973) );
  NAND U1143 ( .A(n520), .B(n684), .Z(n1119) );
  IV U1144 ( .A(n1118), .Z(n1130) );
  XNOR U1145 ( .A(n1115), .B(n1131), .Z(n1118) );
  AND U1146 ( .A(n750), .B(n462), .Z(n1131) );
  XOR U1147 ( .A(n1132), .B(n1133), .Z(n1115) );
  ANDN U1148 ( .A(n1134), .B(n1135), .Z(n1133) );
  XNOR U1149 ( .A(n1136), .B(n1132), .Z(n1134) );
  XNOR U1150 ( .A(n1137), .B(n1138), .Z(n975) );
  IV U1151 ( .A(n1126), .Z(n1138) );
  XNOR U1152 ( .A(n1125), .B(n1139), .Z(n1126) );
  AND U1153 ( .A(n357), .B(e_input[0]), .Z(n1139) );
  XOR U1154 ( .A(n1123), .B(g_input[9]), .Z(n1124) );
  NANDN U1155 ( .B(n1140), .A(n1141), .Z(n1123) );
  XOR U1156 ( .A(n1142), .B(n1143), .Z(n1125) );
  ANDN U1157 ( .A(n1144), .B(n1145), .Z(n1143) );
  XNOR U1158 ( .A(n1146), .B(n1142), .Z(n1144) );
  XOR U1159 ( .A(n1147), .B(n1127), .Z(n1137) );
  NAND U1160 ( .A(n404), .B(n1029), .Z(n1127) );
  IV U1161 ( .A(n1129), .Z(n1147) );
  NAND U1162 ( .A(n581), .B(n684), .Z(n1136) );
  XNOR U1163 ( .A(n1132), .B(n1149), .Z(n1135) );
  AND U1164 ( .A(n750), .B(n520), .Z(n1149) );
  XNOR U1165 ( .A(n1153), .B(n1150), .Z(n1152) );
  XNOR U1166 ( .A(n1142), .B(n1155), .Z(n1145) );
  AND U1167 ( .A(n404), .B(e_input[0]), .Z(n1155) );
  XNOR U1168 ( .A(n1159), .B(n1156), .Z(n1158) );
  XOR U1169 ( .A(n1160), .B(n1146), .Z(n1154) );
  NAND U1170 ( .A(n462), .B(n1029), .Z(n1146) );
  IV U1171 ( .A(n1148), .Z(n1160) );
  XNOR U1172 ( .A(n1161), .B(n1162), .Z(n1148) );
  AND U1173 ( .A(n1163), .B(n1164), .Z(n1162) );
  XOR U1174 ( .A(n1157), .B(n1165), .Z(n1164) );
  XNOR U1175 ( .A(n1159), .B(n1161), .Z(n1165) );
  NAND U1176 ( .A(n520), .B(n1029), .Z(n1159) );
  XOR U1177 ( .A(n1156), .B(n1166), .Z(n1157) );
  AND U1178 ( .A(n462), .B(e_input[0]), .Z(n1166) );
  XNOR U1179 ( .A(n1170), .B(n1167), .Z(n1169) );
  XOR U1180 ( .A(n1151), .B(n1171), .Z(n1163) );
  XNOR U1181 ( .A(n1153), .B(n1161), .Z(n1171) );
  NANDN U1182 ( .B(n646), .A(n684), .Z(n1153) );
  XOR U1183 ( .A(n1150), .B(n1172), .Z(n1151) );
  AND U1184 ( .A(n750), .B(n581), .Z(n1172) );
  XOR U1185 ( .A(n1173), .B(n1174), .Z(n1150) );
  AND U1186 ( .A(n1175), .B(n1176), .Z(n1174) );
  XNOR U1187 ( .A(n1177), .B(n1173), .Z(n1176) );
  XOR U1188 ( .A(n1178), .B(n1179), .Z(n1161) );
  AND U1189 ( .A(n1180), .B(n1181), .Z(n1179) );
  XOR U1190 ( .A(n1168), .B(n1182), .Z(n1181) );
  XNOR U1191 ( .A(n1170), .B(n1178), .Z(n1182) );
  NAND U1192 ( .A(n581), .B(n1029), .Z(n1170) );
  XOR U1193 ( .A(n1167), .B(n1183), .Z(n1168) );
  AND U1194 ( .A(n520), .B(e_input[0]), .Z(n1183) );
  XOR U1195 ( .A(n1184), .B(n1185), .Z(n1167) );
  AND U1196 ( .A(n1186), .B(n1187), .Z(n1185) );
  XNOR U1197 ( .A(n1188), .B(n1184), .Z(n1187) );
  XOR U1198 ( .A(n1175), .B(n1189), .Z(n1180) );
  XNOR U1199 ( .A(n1177), .B(n1178), .Z(n1189) );
  NANDN U1200 ( .B(n718), .A(n684), .Z(n1177) );
  XOR U1201 ( .A(n1173), .B(n1190), .Z(n1175) );
  ANDN U1202 ( .A(n750), .B(n646), .Z(n1190) );
  XNOR U1203 ( .A(n1194), .B(n1191), .Z(n1193) );
  XOR U1204 ( .A(n1195), .B(n1196), .Z(n1178) );
  AND U1205 ( .A(n1197), .B(n1198), .Z(n1196) );
  XOR U1206 ( .A(n1186), .B(n1199), .Z(n1198) );
  XNOR U1207 ( .A(n1188), .B(n1195), .Z(n1199) );
  NANDN U1208 ( .B(n646), .A(n1029), .Z(n1188) );
  XOR U1209 ( .A(n1184), .B(n1200), .Z(n1186) );
  AND U1210 ( .A(n581), .B(e_input[0]), .Z(n1200) );
  XOR U1211 ( .A(n1192), .B(n1204), .Z(n1197) );
  XNOR U1212 ( .A(n1194), .B(n1195), .Z(n1204) );
  NAND U1213 ( .A(n684), .B(n789), .Z(n1194) );
  XOR U1214 ( .A(n1191), .B(n1205), .Z(n1192) );
  ANDN U1215 ( .A(n750), .B(n718), .Z(n1205) );
  XOR U1216 ( .A(n1206), .B(n1207), .Z(n1191) );
  ANDN U1217 ( .A(n1208), .B(n1209), .Z(n1207) );
  XNOR U1218 ( .A(n1210), .B(n1206), .Z(n1208) );
  NAND U1219 ( .A(n684), .B(n1012), .Z(n1210) );
  XNOR U1220 ( .A(n1206), .B(n1212), .Z(n1209) );
  AND U1221 ( .A(n789), .B(n750), .Z(n1212) );
  AND U1222 ( .A(n1213), .B(g_input[0]), .Z(n1206) );
  NANDN U1223 ( .B(n684), .A(n1214), .Z(n1213) );
  NAND U1224 ( .A(n1012), .B(n750), .Z(n1214) );
  XNOR U1225 ( .A(n1201), .B(n1218), .Z(n1202) );
  ANDN U1226 ( .A(e_input[0]), .B(n646), .Z(n1218) );
  XOR U1227 ( .A(n1221), .B(n1219), .Z(n1220) );
  ANDN U1228 ( .A(e_input[0]), .B(n718), .Z(n1221) );
  AND U1229 ( .A(n1029), .B(n789), .Z(n1222) );
  XOR U1230 ( .A(n1226), .B(n1203), .Z(n1217) );
  NANDN U1231 ( .B(n718), .A(n1029), .Z(n1203) );
  IV U1232 ( .A(n1211), .Z(n1226) );
  NAND U1233 ( .A(n1029), .B(n1012), .Z(n1225) );
  XNOR U1234 ( .A(n1223), .B(n1227), .Z(n1224) );
  AND U1235 ( .A(n789), .B(e_input[0]), .Z(n1227) );
  AND U1236 ( .A(n1228), .B(g_input[0]), .Z(n1223) );
  NANDN U1237 ( .B(n1029), .A(n1229), .Z(n1228) );
  NAND U1238 ( .A(n1012), .B(e_input[0]), .Z(n1229) );
  XNOR U1239 ( .A(n1231), .B(n777), .Z(n765) );
  XNOR U1240 ( .A(n762), .B(n763), .Z(n777) );
  NAND U1241 ( .A(n257), .B(n581), .Z(n763) );
  XNOR U1242 ( .A(n761), .B(n1232), .Z(n762) );
  AND U1243 ( .A(n520), .B(n293), .Z(n1232) );
  XNOR U1244 ( .A(n1236), .B(n1233), .Z(n1235) );
  XNOR U1245 ( .A(n776), .B(n764), .Z(n1231) );
  XOR U1246 ( .A(n1237), .B(n1238), .Z(n764) );
  XNOR U1247 ( .A(n769), .B(n1240), .Z(n772) );
  AND U1248 ( .A(n404), .B(n389), .Z(n1240) );
  XNOR U1249 ( .A(n1141), .B(g_input[8]), .Z(n1140) );
  NOR U1250 ( .A(n1241), .B(n1242), .Z(n1141) );
  XOR U1251 ( .A(n1243), .B(n1244), .Z(n769) );
  AND U1252 ( .A(n1245), .B(n1246), .Z(n1244) );
  XNOR U1253 ( .A(n1247), .B(n1243), .Z(n1246) );
  XOR U1254 ( .A(n1248), .B(n773), .Z(n1239) );
  NAND U1255 ( .A(n342), .B(n462), .Z(n773) );
  IV U1256 ( .A(n775), .Z(n1248) );
  XNOR U1257 ( .A(n1249), .B(n1250), .Z(n775) );
  AND U1258 ( .A(n1251), .B(n1252), .Z(n1250) );
  XOR U1259 ( .A(n1245), .B(n1253), .Z(n1252) );
  XNOR U1260 ( .A(n1247), .B(n1249), .Z(n1253) );
  NAND U1261 ( .A(n342), .B(n520), .Z(n1247) );
  XOR U1262 ( .A(n1243), .B(n1254), .Z(n1245) );
  AND U1263 ( .A(n462), .B(n389), .Z(n1254) );
  XOR U1264 ( .A(n1241), .B(g_input[7]), .Z(n1242) );
  NANDN U1265 ( .B(n1255), .A(n1256), .Z(n1241) );
  XOR U1266 ( .A(n1257), .B(n1258), .Z(n1243) );
  AND U1267 ( .A(n1259), .B(n1260), .Z(n1258) );
  XNOR U1268 ( .A(n1261), .B(n1257), .Z(n1260) );
  XOR U1269 ( .A(n1234), .B(n1262), .Z(n1251) );
  XNOR U1270 ( .A(n1236), .B(n1249), .Z(n1262) );
  NANDN U1271 ( .B(n646), .A(n257), .Z(n1236) );
  XOR U1272 ( .A(n1233), .B(n1263), .Z(n1234) );
  AND U1273 ( .A(n581), .B(n293), .Z(n1263) );
  XOR U1274 ( .A(n1264), .B(n1265), .Z(n1233) );
  AND U1275 ( .A(n1266), .B(n1267), .Z(n1265) );
  XNOR U1276 ( .A(n1268), .B(n1264), .Z(n1267) );
  XOR U1277 ( .A(n1269), .B(n1270), .Z(n1249) );
  AND U1278 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U1279 ( .A(n1259), .B(n1273), .Z(n1272) );
  XNOR U1280 ( .A(n1261), .B(n1269), .Z(n1273) );
  NAND U1281 ( .A(n342), .B(n581), .Z(n1261) );
  XOR U1282 ( .A(n1257), .B(n1274), .Z(n1259) );
  AND U1283 ( .A(n520), .B(n389), .Z(n1274) );
  XNOR U1284 ( .A(n1256), .B(g_input[6]), .Z(n1255) );
  NOR U1285 ( .A(n1275), .B(n1276), .Z(n1256) );
  XOR U1286 ( .A(n1277), .B(n1278), .Z(n1257) );
  AND U1287 ( .A(n1279), .B(n1280), .Z(n1278) );
  XNOR U1288 ( .A(n1281), .B(n1277), .Z(n1280) );
  XOR U1289 ( .A(n1266), .B(n1282), .Z(n1271) );
  XNOR U1290 ( .A(n1268), .B(n1269), .Z(n1282) );
  NANDN U1291 ( .B(n718), .A(n257), .Z(n1268) );
  XOR U1292 ( .A(n1264), .B(n1283), .Z(n1266) );
  ANDN U1293 ( .A(n293), .B(n646), .Z(n1283) );
  XNOR U1294 ( .A(n1287), .B(n1284), .Z(n1286) );
  XOR U1295 ( .A(n1288), .B(n1289), .Z(n1269) );
  AND U1296 ( .A(n1290), .B(n1291), .Z(n1289) );
  XOR U1297 ( .A(n1279), .B(n1292), .Z(n1291) );
  XNOR U1298 ( .A(n1281), .B(n1288), .Z(n1292) );
  NANDN U1299 ( .B(n646), .A(n342), .Z(n1281) );
  XOR U1300 ( .A(n1277), .B(n1293), .Z(n1279) );
  AND U1301 ( .A(n581), .B(n389), .Z(n1293) );
  XOR U1302 ( .A(n1275), .B(g_input[5]), .Z(n1276) );
  NANDN U1303 ( .B(n1294), .A(n1295), .Z(n1275) );
  XOR U1304 ( .A(n1296), .B(n1297), .Z(n1277) );
  ANDN U1305 ( .A(n1298), .B(n1299), .Z(n1297) );
  XNOR U1306 ( .A(n1300), .B(n1296), .Z(n1298) );
  XOR U1307 ( .A(n1285), .B(n1301), .Z(n1290) );
  XNOR U1308 ( .A(n1287), .B(n1288), .Z(n1301) );
  NAND U1309 ( .A(n257), .B(n789), .Z(n1287) );
  XOR U1310 ( .A(n1284), .B(n1302), .Z(n1285) );
  ANDN U1311 ( .A(n293), .B(n718), .Z(n1302) );
  NAND U1312 ( .A(n257), .B(n1012), .Z(n1305) );
  XNOR U1313 ( .A(n1303), .B(n1307), .Z(n1304) );
  AND U1314 ( .A(n789), .B(n293), .Z(n1307) );
  AND U1315 ( .A(n1308), .B(g_input[0]), .Z(n1303) );
  NANDN U1316 ( .B(n257), .A(n1309), .Z(n1308) );
  NAND U1317 ( .A(n1012), .B(n293), .Z(n1309) );
  XNOR U1318 ( .A(n1312), .B(n1313), .Z(n1238) );
  IV U1319 ( .A(n1299), .Z(n1313) );
  XNOR U1320 ( .A(n1296), .B(n1314), .Z(n1299) );
  ANDN U1321 ( .A(n389), .B(n646), .Z(n1314) );
  XOR U1322 ( .A(n1315), .B(n1316), .Z(n1296) );
  AND U1323 ( .A(n1317), .B(n1318), .Z(n1316) );
  XOR U1324 ( .A(n1319), .B(n1315), .Z(n1318) );
  ANDN U1325 ( .A(n389), .B(n718), .Z(n1319) );
  XOR U1326 ( .A(n1320), .B(n1315), .Z(n1317) );
  AND U1327 ( .A(n789), .B(n342), .Z(n1320) );
  XOR U1328 ( .A(n1321), .B(n1322), .Z(n1315) );
  ANDN U1329 ( .A(n1323), .B(n1324), .Z(n1322) );
  XNOR U1330 ( .A(n1325), .B(n1321), .Z(n1323) );
  XOR U1331 ( .A(n1326), .B(n1300), .Z(n1312) );
  NANDN U1332 ( .B(n718), .A(n342), .Z(n1300) );
  IV U1333 ( .A(n1306), .Z(n1326) );
  XOR U1334 ( .A(n1327), .B(n1325), .Z(n1306) );
  NAND U1335 ( .A(n342), .B(n1012), .Z(n1325) );
  IV U1336 ( .A(n1324), .Z(n1327) );
  XNOR U1337 ( .A(n1321), .B(n1328), .Z(n1324) );
  AND U1338 ( .A(n789), .B(n389), .Z(n1328) );
  AND U1339 ( .A(n1329), .B(g_input[0]), .Z(n1321) );
  NANDN U1340 ( .B(n342), .A(n1330), .Z(n1329) );
  NAND U1341 ( .A(n1012), .B(n389), .Z(n1330) );
  XNOR U1342 ( .A(n780), .B(n1334), .Z(n783) );
  ANDN U1343 ( .A(n230), .B(n646), .Z(n1334) );
  XNOR U1344 ( .A(n1295), .B(g_input[4]), .Z(n1294) );
  NOR U1345 ( .A(n1335), .B(n1336), .Z(n1295) );
  XOR U1346 ( .A(n1337), .B(n1338), .Z(n780) );
  AND U1347 ( .A(n1339), .B(n1340), .Z(n1338) );
  XOR U1348 ( .A(n1341), .B(n1337), .Z(n1340) );
  ANDN U1349 ( .A(n230), .B(n718), .Z(n1341) );
  XOR U1350 ( .A(n1342), .B(n1337), .Z(n1339) );
  AND U1351 ( .A(n789), .B(n195), .Z(n1342) );
  XOR U1352 ( .A(n1343), .B(n1344), .Z(n1337) );
  ANDN U1353 ( .A(n1345), .B(n1346), .Z(n1344) );
  XNOR U1354 ( .A(n1347), .B(n1343), .Z(n1345) );
  XOR U1355 ( .A(n1348), .B(n784), .Z(n1333) );
  NANDN U1356 ( .B(n718), .A(n195), .Z(n784) );
  NANDN U1357 ( .B(n1349), .A(n1350), .Z(n1335) );
  IV U1358 ( .A(n786), .Z(n1348) );
  XOR U1359 ( .A(n1351), .B(n1347), .Z(n786) );
  NAND U1360 ( .A(n195), .B(n1012), .Z(n1347) );
  IV U1361 ( .A(n1346), .Z(n1351) );
  XNOR U1362 ( .A(n1343), .B(n1352), .Z(n1346) );
  AND U1363 ( .A(n789), .B(n230), .Z(n1352) );
  AND U1364 ( .A(n1353), .B(g_input[0]), .Z(n1343) );
  NANDN U1365 ( .B(n195), .A(n1354), .Z(n1353) );
  NAND U1366 ( .A(n1012), .B(n230), .Z(n1354) );
  XNOR U1367 ( .A(n793), .B(n794), .Z(n788) );
  NANDN U1368 ( .B(n145), .A(n1012), .Z(n794) );
  XNOR U1369 ( .A(n792), .B(n1357), .Z(n793) );
  AND U1370 ( .A(n789), .B(n165), .Z(n1357) );
  XNOR U1371 ( .A(n1350), .B(g_input[2]), .Z(n1349) );
  AND U1372 ( .A(n1359), .B(g_input[0]), .Z(n792) );
  NAND U1373 ( .A(n1360), .B(n145), .Z(n1359) );
  NANDN U1374 ( .B(n1361), .A(n1362), .Z(n145) );
  ANDN U1375 ( .A(e_input[15]), .B(n1363), .Z(n1362) );
  NAND U1376 ( .A(n1012), .B(n165), .Z(n1360) );
  XOR U1377 ( .A(n1363), .B(e_input[14]), .Z(n1361) );
  OR U1378 ( .A(n1356), .B(n1364), .Z(n1363) );
  XOR U1379 ( .A(n1364), .B(e_input[13]), .Z(n1356) );
  OR U1380 ( .A(n1355), .B(n1365), .Z(n1364) );
  XOR U1381 ( .A(n1365), .B(e_input[12]), .Z(n1355) );
  OR U1382 ( .A(n1311), .B(n1366), .Z(n1365) );
  XOR U1383 ( .A(n1366), .B(e_input[11]), .Z(n1311) );
  OR U1384 ( .A(n1310), .B(n1367), .Z(n1366) );
  XOR U1385 ( .A(n1367), .B(e_input[10]), .Z(n1310) );
  OR U1386 ( .A(n1332), .B(n1368), .Z(n1367) );
  XOR U1387 ( .A(n1368), .B(e_input[9]), .Z(n1332) );
  OR U1388 ( .A(n1331), .B(n1369), .Z(n1368) );
  XOR U1389 ( .A(n1369), .B(e_input[8]), .Z(n1331) );
  OR U1390 ( .A(n1022), .B(n1370), .Z(n1369) );
  XOR U1391 ( .A(n1370), .B(e_input[7]), .Z(n1022) );
  OR U1392 ( .A(n1021), .B(n1371), .Z(n1370) );
  XOR U1393 ( .A(n1371), .B(e_input[6]), .Z(n1021) );
  OR U1394 ( .A(n1017), .B(n1372), .Z(n1371) );
  XOR U1395 ( .A(n1372), .B(e_input[5]), .Z(n1017) );
  OR U1396 ( .A(n1016), .B(n1373), .Z(n1372) );
  XOR U1397 ( .A(n1373), .B(e_input[4]), .Z(n1016) );
  OR U1398 ( .A(n1216), .B(n1374), .Z(n1373) );
  XOR U1399 ( .A(n1374), .B(e_input[3]), .Z(n1216) );
  OR U1400 ( .A(n1215), .B(n1375), .Z(n1374) );
  XOR U1401 ( .A(n1375), .B(e_input[2]), .Z(n1215) );
  NANDN U1402 ( .B(e_input[0]), .A(n1230), .Z(n1375) );
  XNOR U1403 ( .A(e_input[0]), .B(e_input[1]), .Z(n1230) );
  XOR U1404 ( .A(g_input[0]), .B(g_input[1]), .Z(n1358) );
  AND U1405 ( .A(n1376), .B(n1377), .Z(\_MxM/N31 ) );
  XOR U1406 ( .A(\_MxM/n[13] ), .B(\_MxM/add_43/carry[13] ), .Z(n1377) );
  AND U1407 ( .A(\_MxM/N16 ), .B(n1376), .Z(\_MxM/N30 ) );
  AND U1408 ( .A(\_MxM/N15 ), .B(n1376), .Z(\_MxM/N29 ) );
  AND U1409 ( .A(\_MxM/N14 ), .B(n1376), .Z(\_MxM/N28 ) );
  AND U1410 ( .A(\_MxM/N13 ), .B(n1376), .Z(\_MxM/N27 ) );
  AND U1411 ( .A(\_MxM/N12 ), .B(n1376), .Z(\_MxM/N26 ) );
  AND U1412 ( .A(\_MxM/N11 ), .B(n1376), .Z(\_MxM/N25 ) );
  AND U1413 ( .A(\_MxM/N10 ), .B(n1376), .Z(\_MxM/N24 ) );
  AND U1414 ( .A(\_MxM/N9 ), .B(n1376), .Z(\_MxM/N23 ) );
  AND U1415 ( .A(\_MxM/N8 ), .B(n1376), .Z(\_MxM/N22 ) );
  AND U1416 ( .A(\_MxM/N7 ), .B(n1376), .Z(\_MxM/N21 ) );
  AND U1417 ( .A(\_MxM/N6 ), .B(n1376), .Z(\_MxM/N20 ) );
  AND U1418 ( .A(\_MxM/N5 ), .B(n1376), .Z(\_MxM/N19 ) );
  NAND U1419 ( .A(n1378), .B(n1379), .Z(n1376) );
  AND U1420 ( .A(n1380), .B(n1381), .Z(n1379) );
  ANDN U1421 ( .A(n108), .B(\_MxM/N18 ), .Z(n1381) );
  NOR U1422 ( .A(\_MxM/n[12] ), .B(\_MxM/n[11] ), .Z(n108) );
  AND U1423 ( .A(\_MxM/n[10] ), .B(n1382), .Z(n1380) );
  NOR U1424 ( .A(n110), .B(n111), .Z(n1382) );
  OR U1425 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n111) );
  OR U1426 ( .A(\_MxM/n[5] ), .B(\_MxM/n[4] ), .Z(n110) );
  AND U1427 ( .A(n1383), .B(n1384), .Z(n1378) );
  AND U1428 ( .A(\_MxM/n[2] ), .B(n1385), .Z(n1384) );
  AND U1429 ( .A(\_MxM/n[1] ), .B(\_MxM/n[13] ), .Z(n1385) );
  AND U1430 ( .A(\_MxM/n[9] ), .B(n1386), .Z(n1383) );
  AND U1431 ( .A(\_MxM/n[8] ), .B(\_MxM/n[3] ), .Z(n1386) );
  IV U1432 ( .A(\_MxM/n[0] ), .Z(\_MxM/N18 ) );
endmodule

