
module MxM_TG_W32_N1000 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MxM/n341 , \_MxM/n340 , \_MxM/n339 , \_MxM/n338 , \_MxM/n337 ,
         \_MxM/n336 , \_MxM/n335 , \_MxM/n334 , \_MxM/n333 , \_MxM/n332 ,
         \_MxM/n331 , \_MxM/n330 , \_MxM/n329 , \_MxM/n328 , \_MxM/n327 ,
         \_MxM/n326 , \_MxM/n325 , \_MxM/n324 , \_MxM/n323 , \_MxM/n322 ,
         \_MxM/n321 , \_MxM/n320 , \_MxM/n319 , \_MxM/n318 , \_MxM/n317 ,
         \_MxM/n316 , \_MxM/n315 , \_MxM/n314 , \_MxM/n313 , \_MxM/n312 ,
         \_MxM/n311 , \_MxM/n310 , \_MxM/n309 , \_MxM/n308 , \_MxM/n307 ,
         \_MxM/n306 , \_MxM/n305 , \_MxM/n304 , \_MxM/n303 , \_MxM/n302 ,
         \_MxM/n301 , \_MxM/n300 , \_MxM/n299 , \_MxM/n298 , \_MxM/n297 ,
         \_MxM/n296 , \_MxM/n295 , \_MxM/n294 , \_MxM/n293 , \_MxM/n292 ,
         \_MxM/n291 , \_MxM/n290 , \_MxM/n289 , \_MxM/n288 , \_MxM/n287 ,
         \_MxM/n286 , \_MxM/n285 , \_MxM/n284 , \_MxM/n283 , \_MxM/n282 ,
         \_MxM/n281 , \_MxM/n280 , \_MxM/n279 , \_MxM/n278 , \_MxM/N24 ,
         \_MxM/N23 , \_MxM/N22 , \_MxM/N21 , \_MxM/N20 , \_MxM/N19 ,
         \_MxM/N18 , \_MxM/N17 , \_MxM/N16 , \_MxM/N15 , \_MxM/N13 ,
         \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/N7 ,
         \_MxM/N6 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] ,
         \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] ,
         \_MxM/n[9] , \_MxM/Y0[0] , \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] ,
         \_MxM/Y0[4] , \_MxM/Y0[5] , \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/Y0[8] ,
         \_MxM/Y0[9] , \_MxM/Y0[10] , \_MxM/Y0[11] , \_MxM/Y0[12] ,
         \_MxM/Y0[13] , \_MxM/Y0[14] , \_MxM/Y0[15] , \_MxM/Y0[16] ,
         \_MxM/Y0[17] , \_MxM/Y0[18] , \_MxM/Y0[19] , \_MxM/Y0[20] ,
         \_MxM/Y0[21] , \_MxM/Y0[22] , \_MxM/Y0[23] , \_MxM/Y0[24] ,
         \_MxM/Y0[25] , \_MxM/Y0[26] , \_MxM/Y0[27] , \_MxM/Y0[28] ,
         \_MxM/Y0[29] , \_MxM/Y0[30] , \_MxM/Y0[31] , \_MxM/add_39/carry[9] ,
         \_MxM/add_39/carry[8] , \_MxM/add_39/carry[7] ,
         \_MxM/add_39/carry[6] , \_MxM/add_39/carry[5] ,
         \_MxM/add_39/carry[4] , \_MxM/add_39/carry[3] ,
         \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n278 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n279 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n280 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n281 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n282 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n283 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n284 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n285 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n286 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n287 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n288 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n289 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n290 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n291 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n292 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n293 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y_reg[16]  ( .D(\_MxM/n294 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[16]) );
  DFF \_MxM/Y_reg[17]  ( .D(\_MxM/n295 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[17]) );
  DFF \_MxM/Y_reg[18]  ( .D(\_MxM/n296 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[18]) );
  DFF \_MxM/Y_reg[19]  ( .D(\_MxM/n297 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[19]) );
  DFF \_MxM/Y_reg[20]  ( .D(\_MxM/n298 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[20]) );
  DFF \_MxM/Y_reg[21]  ( .D(\_MxM/n299 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[21]) );
  DFF \_MxM/Y_reg[22]  ( .D(\_MxM/n300 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[22]) );
  DFF \_MxM/Y_reg[23]  ( .D(\_MxM/n301 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[23]) );
  DFF \_MxM/Y_reg[24]  ( .D(\_MxM/n302 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[24]) );
  DFF \_MxM/Y_reg[25]  ( .D(\_MxM/n303 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[25]) );
  DFF \_MxM/Y_reg[26]  ( .D(\_MxM/n304 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[26]) );
  DFF \_MxM/Y_reg[27]  ( .D(\_MxM/n305 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[27]) );
  DFF \_MxM/Y_reg[28]  ( .D(\_MxM/n306 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[28]) );
  DFF \_MxM/Y_reg[29]  ( .D(\_MxM/n307 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[29]) );
  DFF \_MxM/Y_reg[30]  ( .D(\_MxM/n308 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[30]) );
  DFF \_MxM/Y_reg[31]  ( .D(\_MxM/n309 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[31]) );
  DFF \_MxM/Y0_reg[31]  ( .D(\_MxM/n310 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[31] ) );
  DFF \_MxM/Y0_reg[30]  ( .D(\_MxM/n311 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[30] ) );
  DFF \_MxM/Y0_reg[29]  ( .D(\_MxM/n312 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[29] ) );
  DFF \_MxM/Y0_reg[28]  ( .D(\_MxM/n313 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[28] ) );
  DFF \_MxM/Y0_reg[27]  ( .D(\_MxM/n314 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[27] ) );
  DFF \_MxM/Y0_reg[26]  ( .D(\_MxM/n315 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[26] ) );
  DFF \_MxM/Y0_reg[25]  ( .D(\_MxM/n316 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[25] ) );
  DFF \_MxM/Y0_reg[24]  ( .D(\_MxM/n317 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[24] ) );
  DFF \_MxM/Y0_reg[23]  ( .D(\_MxM/n318 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[23] ) );
  DFF \_MxM/Y0_reg[22]  ( .D(\_MxM/n319 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[22] ) );
  DFF \_MxM/Y0_reg[21]  ( .D(\_MxM/n320 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[21] ) );
  DFF \_MxM/Y0_reg[20]  ( .D(\_MxM/n321 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[20] ) );
  DFF \_MxM/Y0_reg[19]  ( .D(\_MxM/n322 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[19] ) );
  DFF \_MxM/Y0_reg[18]  ( .D(\_MxM/n323 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[18] ) );
  DFF \_MxM/Y0_reg[17]  ( .D(\_MxM/n324 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[17] ) );
  DFF \_MxM/Y0_reg[16]  ( .D(\_MxM/n325 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[16] ) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/n326 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/n327 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/n328 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/n329 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/n330 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/n331 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/n332 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/n333 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n334 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n335 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n336 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n337 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n338 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n339 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n340 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n341 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N24 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N13 ) );
  MUX U1 ( .IN0(n3698), .IN1(n1), .SEL(n3699), .F(n3652) );
  IV U2 ( .A(n3700), .Z(n1) );
  MUX U3 ( .IN0(n3526), .IN1(n3528), .SEL(n3527), .F(n3480) );
  MUX U4 ( .IN0(n4299), .IN1(n4301), .SEL(n4300), .F(n4275) );
  MUX U5 ( .IN0(n3351), .IN1(n3353), .SEL(n3352), .F(n3305) );
  XNOR U6 ( .A(n4287), .B(n4286), .Z(n4302) );
  XNOR U7 ( .A(n4670), .B(n4668), .Z(n4675) );
  MUX U8 ( .IN0(n3255), .IN1(n3257), .SEL(n3256), .F(n3212) );
  MUX U9 ( .IN0(n5003), .IN1(n5005), .SEL(n5004), .F(n4991) );
  MUX U10 ( .IN0(n4861), .IN1(n2), .SEL(n4862), .F(n4841) );
  IV U11 ( .A(n4863), .Z(n2) );
  MUX U12 ( .IN0(n5010), .IN1(n3), .SEL(n5011), .F(n4998) );
  IV U13 ( .A(n5012), .Z(n3) );
  MUX U14 ( .IN0(n4220), .IN1(n4), .SEL(n4221), .F(n4200) );
  IV U15 ( .A(n4222), .Z(n4) );
  XNOR U16 ( .A(n3208), .B(n3207), .Z(n3244) );
  MUX U17 ( .IN0(n4625), .IN1(n5), .SEL(n4626), .F(n4615) );
  IV U18 ( .A(n4627), .Z(n5) );
  XNOR U19 ( .A(n3233), .B(n3231), .Z(n3268) );
  XNOR U20 ( .A(n4396), .B(n4394), .Z(n4403) );
  NANDN U21 ( .B(n1283), .A(n3009), .Z(n18) );
  MUX U22 ( .IN0(n3085), .IN1(n3087), .SEL(n3086), .F(n3046) );
  MUX U23 ( .IN0(n3078), .IN1(n6), .SEL(n3079), .F(n3039) );
  IV U24 ( .A(n3080), .Z(n6) );
  MUX U25 ( .IN0(n3090), .IN1(n3092), .SEL(n3091), .F(n3019) );
  MUX U26 ( .IN0(n994), .IN1(n7), .SEL(n995), .F(n925) );
  IV U27 ( .A(n996), .Z(n7) );
  MUX U28 ( .IN0(n1291), .IN1(n1293), .SEL(n1292), .F(n1207) );
  MUX U29 ( .IN0(n1346), .IN1(n8), .SEL(n1347), .F(n1255) );
  IV U30 ( .A(n1348), .Z(n8) );
  MUX U31 ( .IN0(n1394), .IN1(n9), .SEL(n1395), .F(n1299) );
  IV U32 ( .A(n1396), .Z(n9) );
  MUX U33 ( .IN0(n1499), .IN1(n10), .SEL(n1500), .F(n1402) );
  IV U34 ( .A(n1501), .Z(n10) );
  MUX U35 ( .IN0(n1758), .IN1(n1760), .SEL(n1759), .F(n1657) );
  MUX U36 ( .IN0(n1874), .IN1(n11), .SEL(n1875), .F(n1766) );
  IV U37 ( .A(n1876), .Z(n11) );
  MUX U38 ( .IN0(n2047), .IN1(n12), .SEL(n2048), .F(n1938) );
  IV U39 ( .A(n2049), .Z(n12) );
  MUX U40 ( .IN0(g_input[29]), .IN1(n4371), .SEL(g_input[31]), .F(n13) );
  IV U41 ( .A(n13), .Z(n618) );
  MUX U42 ( .IN0(n14), .IN1(n4360), .SEL(g_input[31]), .F(n574) );
  IV U43 ( .A(g_input[30]), .Z(n14) );
  MUX U44 ( .IN0(n4922), .IN1(n4924), .SEL(n4923), .F(n4898) );
  MUX U45 ( .IN0(n4672), .IN1(n4674), .SEL(n4673), .F(n4657) );
  XNOR U46 ( .A(n5044), .B(n5042), .Z(n5049) );
  MUX U47 ( .IN0(n4255), .IN1(n4257), .SEL(n4256), .F(n4235) );
  MUX U48 ( .IN0(n4260), .IN1(n15), .SEL(n4261), .F(n4240) );
  IV U49 ( .A(n4262), .Z(n15) );
  XNOR U50 ( .A(n4910), .B(n4909), .Z(n4925) );
  MUX U51 ( .IN0(n4991), .IN1(n4993), .SEL(n4992), .F(n4979) );
  MUX U52 ( .IN0(n4841), .IN1(n16), .SEL(n4842), .F(n4821) );
  IV U53 ( .A(n4843), .Z(n16) );
  MUX U54 ( .IN0(n4998), .IN1(n17), .SEL(n4999), .F(n4986) );
  IV U55 ( .A(n5000), .Z(n17) );
  MUX U56 ( .IN0(n3170), .IN1(n3172), .SEL(n3171), .F(n3125) );
  XNOR U57 ( .A(n4628), .B(n4627), .Z(n4633) );
  MUX U58 ( .IN0(n4620), .IN1(n4622), .SEL(n4621), .F(n4610) );
  MUX U59 ( .IN0(n5115), .IN1(n18), .SEL(n5116), .F(n5104) );
  XNOR U60 ( .A(n3121), .B(n3120), .Z(n3159) );
  MUX U61 ( .IN0(n4605), .IN1(n19), .SEL(n4606), .F(n4592) );
  IV U62 ( .A(n4607), .Z(n19) );
  MUX U63 ( .IN0(n3039), .IN1(n20), .SEL(n3040), .F(n2909) );
  IV U64 ( .A(n3041), .Z(n20) );
  MUX U65 ( .IN0(n1146), .IN1(n21), .SEL(n1147), .F(n1066) );
  IV U66 ( .A(n1148), .Z(n21) );
  MUX U67 ( .IN0(n1207), .IN1(n1209), .SEL(n1208), .F(n1126) );
  MUX U68 ( .IN0(n1264), .IN1(n1266), .SEL(n1265), .F(n1182) );
  MUX U69 ( .IN0(n1579), .IN1(n1581), .SEL(n1580), .F(n1483) );
  MUX U70 ( .IN0(n1587), .IN1(n22), .SEL(n1588), .F(n1491) );
  IV U71 ( .A(n1589), .Z(n22) );
  MUX U72 ( .IN0(n1595), .IN1(n23), .SEL(n1596), .F(n1499) );
  IV U73 ( .A(n1597), .Z(n23) );
  MUX U74 ( .IN0(n1642), .IN1(n24), .SEL(n1643), .F(n1542) );
  IV U75 ( .A(n1644), .Z(n24) );
  MUX U76 ( .IN0(n1839), .IN1(n1841), .SEL(n1840), .F(n1731) );
  MUX U77 ( .IN0(n1981), .IN1(n25), .SEL(n1982), .F(n1874) );
  IV U78 ( .A(n1983), .Z(n25) );
  MUX U79 ( .IN0(n2161), .IN1(n26), .SEL(n2162), .F(n2047) );
  IV U80 ( .A(n2163), .Z(n26) );
  MUX U81 ( .IN0(n2787), .IN1(n27), .SEL(n2788), .F(n2662) );
  IV U82 ( .A(n2789), .Z(n27) );
  MUX U83 ( .IN0(n694), .IN1(n28), .SEL(n695), .F(n648) );
  IV U84 ( .A(n696), .Z(n28) );
  MUX U85 ( .IN0(n2942), .IN1(n2944), .SEL(n2943), .F(n2803) );
  MUX U86 ( .IN0(n29), .IN1(n729), .SEL(n728), .F(n691) );
  IV U87 ( .A(n727), .Z(n29) );
  MUX U88 ( .IN0(n3706), .IN1(n3708), .SEL(n3707), .F(n3662) );
  MUX U89 ( .IN0(n4684), .IN1(n4686), .SEL(n4685), .F(n4672) );
  XNOR U90 ( .A(n4682), .B(n4681), .Z(n4687) );
  MUX U91 ( .IN0(n4876), .IN1(n4878), .SEL(n4877), .F(n4856) );
  MUX U92 ( .IN0(n5024), .IN1(n30), .SEL(n5025), .F(n5010) );
  IV U93 ( .A(n5026), .Z(n30) );
  MUX U94 ( .IN0(n4235), .IN1(n4237), .SEL(n4236), .F(n4215) );
  MUX U95 ( .IN0(n4240), .IN1(n31), .SEL(n4241), .F(n4220) );
  IV U96 ( .A(n4242), .Z(n31) );
  MUX U97 ( .IN0(n3219), .IN1(n3221), .SEL(n3220), .F(n3175) );
  XNOR U98 ( .A(n4844), .B(n4843), .Z(n4859) );
  MUX U99 ( .IN0(n4979), .IN1(n4981), .SEL(n4980), .F(n4967) );
  XNOR U100 ( .A(n4989), .B(n4988), .Z(n4994) );
  NANDN U101 ( .B(n2039), .A(n3009), .Z(n44) );
  MUX U102 ( .IN0(n4615), .IN1(n32), .SEL(n4616), .F(n4605) );
  IV U103 ( .A(n4617), .Z(n32) );
  MUX U104 ( .IN0(n4610), .IN1(n4612), .SEL(n4611), .F(n4600) );
  XNOR U105 ( .A(n3081), .B(n3080), .Z(n3114) );
  MUX U106 ( .IN0(n1386), .IN1(n1388), .SEL(n1387), .F(n1291) );
  MUX U107 ( .IN0(n1683), .IN1(n33), .SEL(n1684), .F(n1587) );
  IV U108 ( .A(n1685), .Z(n33) );
  MUX U109 ( .IN0(n1691), .IN1(n34), .SEL(n1692), .F(n1595) );
  IV U110 ( .A(n1693), .Z(n34) );
  MUX U111 ( .IN0(n1649), .IN1(n1651), .SEL(n1650), .F(n1551) );
  MUX U112 ( .IN0(n1657), .IN1(n1659), .SEL(n1658), .F(n1559) );
  MUX U113 ( .IN0(n1743), .IN1(n35), .SEL(n1744), .F(n1642) );
  IV U114 ( .A(n1745), .Z(n35) );
  MUX U115 ( .IN0(n1776), .IN1(n1778), .SEL(n1777), .F(n1675) );
  MUX U116 ( .IN0(n1947), .IN1(n1949), .SEL(n1948), .F(n1839) );
  MUX U117 ( .IN0(n2089), .IN1(n36), .SEL(n2090), .F(n1981) );
  IV U118 ( .A(n2091), .Z(n36) );
  MUX U119 ( .IN0(n2257), .IN1(n2259), .SEL(n2258), .F(n2138) );
  MUX U120 ( .IN0(n2395), .IN1(n37), .SEL(n2396), .F(n2275) );
  IV U121 ( .A(n2397), .Z(n37) );
  MUX U122 ( .IN0(n2925), .IN1(n38), .SEL(n2926), .F(n2787) );
  IV U123 ( .A(n2927), .Z(n38) );
  MUX U124 ( .IN0(n720), .IN1(n722), .SEL(n721), .F(n678) );
  MUX U125 ( .IN0(n610), .IN1(n39), .SEL(n611), .F(n564) );
  IV U126 ( .A(n612), .Z(n39) );
  MUX U127 ( .IN0(n40), .IN1(n956), .SEL(n955), .F(n891) );
  IV U128 ( .A(n954), .Z(n40) );
  MUX U129 ( .IN0(n5046), .IN1(n5048), .SEL(n5047), .F(n5029) );
  MUX U130 ( .IN0(n4927), .IN1(n41), .SEL(n4928), .F(n4905) );
  IV U131 ( .A(n4929), .Z(n41) );
  MUX U132 ( .IN0(n4745), .IN1(n4747), .SEL(n4746), .F(n4729) );
  MUX U133 ( .IN0(n4856), .IN1(n4858), .SEL(n4857), .F(n4836) );
  MUX U134 ( .IN0(n4630), .IN1(n4632), .SEL(n4631), .F(n4620) );
  XNOR U135 ( .A(n4412), .B(n4411), .Z(n4419) );
  MUX U136 ( .IN0(n4195), .IN1(n4197), .SEL(n4196), .F(n4175) );
  XNOR U137 ( .A(n4223), .B(n4222), .Z(n4238) );
  MUX U138 ( .IN0(n4821), .IN1(n42), .SEL(n4822), .F(n4801) );
  IV U139 ( .A(n4823), .Z(n42) );
  MUX U140 ( .IN0(n4986), .IN1(n43), .SEL(n4987), .F(n4974) );
  IV U141 ( .A(n4988), .Z(n43) );
  MUX U142 ( .IN0(n3791), .IN1(n44), .SEL(n3792), .F(n3780) );
  MUX U143 ( .IN0(n4967), .IN1(n4969), .SEL(n4968), .F(n4784) );
  MUX U144 ( .IN0(n4156), .IN1(n45), .SEL(n4157), .F(n4135) );
  IV U145 ( .A(n4158), .Z(n45) );
  XNOR U146 ( .A(n4608), .B(n4607), .Z(n4613) );
  MUX U147 ( .IN0(n3046), .IN1(n3048), .SEL(n3047), .F(n2916) );
  MUX U148 ( .IN0(n1455), .IN1(n1457), .SEL(n1456), .F(n1353) );
  MUX U149 ( .IN0(n1491), .IN1(n46), .SEL(n1492), .F(n1394) );
  IV U150 ( .A(n1493), .Z(n46) );
  MUX U151 ( .IN0(n1483), .IN1(n1485), .SEL(n1484), .F(n1386) );
  MUX U152 ( .IN0(n1792), .IN1(n47), .SEL(n1793), .F(n1691) );
  IV U153 ( .A(n1794), .Z(n47) );
  MUX U154 ( .IN0(n1965), .IN1(n1967), .SEL(n1966), .F(n1858) );
  MUX U155 ( .IN0(n1958), .IN1(n48), .SEL(n1959), .F(n1851) );
  IV U156 ( .A(n1960), .Z(n48) );
  MUX U157 ( .IN0(n1997), .IN1(n49), .SEL(n1998), .F(n1890) );
  IV U158 ( .A(n1999), .Z(n49) );
  MUX U159 ( .IN0(n2054), .IN1(n2056), .SEL(n2055), .F(n1947) );
  MUX U160 ( .IN0(n2208), .IN1(n50), .SEL(n2209), .F(n2089) );
  IV U161 ( .A(n2210), .Z(n50) );
  MUX U162 ( .IN0(n2625), .IN1(n2627), .SEL(n2626), .F(n2501) );
  MUX U163 ( .IN0(n2633), .IN1(n51), .SEL(n2634), .F(n2509) );
  IV U164 ( .A(n2635), .Z(n51) );
  MUX U165 ( .IN0(g_input[28]), .IN1(n4389), .SEL(g_input[31]), .F(n52) );
  IV U166 ( .A(n52), .Z(n658) );
  MUX U167 ( .IN0(n678), .IN1(n680), .SEL(n679), .F(n637) );
  XNOR U168 ( .A(n959), .B(n956), .Z(n1019) );
  MUX U169 ( .IN0(n5109), .IN1(n5111), .SEL(n5110), .F(n5093) );
  MUX U170 ( .IN0(n53), .IN1(n4724), .SEL(n4725), .F(n4710) );
  IV U171 ( .A(n4726), .Z(n53) );
  XNOR U172 ( .A(n4243), .B(n4242), .Z(n4258) );
  MUX U173 ( .IN0(n5187), .IN1(n54), .SEL(n5188), .F(n5169) );
  IV U174 ( .A(n5189), .Z(n54) );
  MUX U175 ( .IN0(n4836), .IN1(n4838), .SEL(n4837), .F(n4816) );
  MUX U176 ( .IN0(n4175), .IN1(n4177), .SEL(n4176), .F(n4163) );
  NANDN U177 ( .B(n2534), .A(n3009), .Z(n67) );
  MUX U178 ( .IN0(n4180), .IN1(n55), .SEL(n4181), .F(n4156) );
  IV U179 ( .A(n4182), .Z(n55) );
  XNOR U180 ( .A(n3890), .B(n3888), .Z(n3903) );
  XNOR U181 ( .A(n4824), .B(n4823), .Z(n4839) );
  MUX U182 ( .IN0(n4974), .IN1(n56), .SEL(n4975), .F(n4962) );
  IV U183 ( .A(n4976), .Z(n56) );
  MUX U184 ( .IN0(n4600), .IN1(n4602), .SEL(n4601), .F(n4583) );
  MUX U185 ( .IN0(n4770), .IN1(n57), .SEL(n4771), .F(n2956) );
  IV U186 ( .A(n4772), .Z(n57) );
  MUX U187 ( .IN0(n1402), .IN1(n58), .SEL(n1403), .F(n1309) );
  IV U188 ( .A(n1404), .Z(n58) );
  MUX U189 ( .IN0(n1551), .IN1(n1553), .SEL(n1552), .F(n1455) );
  MUX U190 ( .IN0(n1675), .IN1(n1677), .SEL(n1676), .F(n1579) );
  MUX U191 ( .IN0(n1851), .IN1(n59), .SEL(n1852), .F(n1743) );
  IV U192 ( .A(n1853), .Z(n59) );
  MUX U193 ( .IN0(n2005), .IN1(n60), .SEL(n2006), .F(n1898) );
  IV U194 ( .A(n2007), .Z(n60) );
  MUX U195 ( .IN0(n2105), .IN1(n61), .SEL(n2106), .F(n1997) );
  IV U196 ( .A(n2107), .Z(n61) );
  MUX U197 ( .IN0(n2200), .IN1(n2202), .SEL(n2201), .F(n2081) );
  MUX U198 ( .IN0(n2192), .IN1(n2194), .SEL(n2193), .F(n2073) );
  MUX U199 ( .IN0(n2282), .IN1(n2284), .SEL(n2283), .F(n2168) );
  MUX U200 ( .IN0(n2575), .IN1(n62), .SEL(n2576), .F(n2450) );
  IV U201 ( .A(n2577), .Z(n62) );
  MUX U202 ( .IN0(n659), .IN1(n661), .SEL(n660), .F(n619) );
  MUX U203 ( .IN0(n1031), .IN1(n1033), .SEL(n1032), .F(n963) );
  MUX U204 ( .IN0(g_input[25]), .IN1(n4438), .SEL(g_input[31]), .F(n63) );
  IV U205 ( .A(n63), .Z(n803) );
  MUX U206 ( .IN0(n2030), .IN1(n2032), .SEL(n2031), .F(n1925) );
  XNOR U207 ( .A(n790), .B(n789), .Z(n845) );
  XNOR U208 ( .A(n290), .B(n1280), .Z(n1203) );
  AND U209 ( .A(n559), .B(n561), .Z(n530) );
  MUX U210 ( .IN0(n4740), .IN1(n64), .SEL(n4741), .F(n4724) );
  IV U211 ( .A(n4742), .Z(n64) );
  XNOR U212 ( .A(n4886), .B(n4885), .Z(n4903) );
  MUX U213 ( .IN0(n3785), .IN1(n3787), .SEL(n3786), .F(n3771) );
  MUX U214 ( .IN0(n4200), .IN1(n65), .SEL(n4201), .F(n4180) );
  IV U215 ( .A(n4202), .Z(n65) );
  XNOR U216 ( .A(n3166), .B(n3165), .Z(n3201) );
  MUX U217 ( .IN0(n66), .IN1(n5169), .SEL(n5170), .F(n5153) );
  IV U218 ( .A(n5171), .Z(n66) );
  MUX U219 ( .IN0(n4816), .IN1(n4818), .SEL(n4817), .F(n4796) );
  MUX U220 ( .IN0(n4318), .IN1(n67), .SEL(n4319), .F(n4304) );
  XNOR U221 ( .A(n4618), .B(n4617), .Z(n4623) );
  MUX U222 ( .IN0(n4801), .IN1(n68), .SEL(n4802), .F(n4770) );
  IV U223 ( .A(n4803), .Z(n68) );
  XNOR U224 ( .A(n3148), .B(n3146), .Z(n3183) );
  MUX U225 ( .IN0(n4962), .IN1(n69), .SEL(n4963), .F(n2979) );
  IV U226 ( .A(n4964), .Z(n69) );
  MUX U227 ( .IN0(n1898), .IN1(n70), .SEL(n1899), .F(n1792) );
  IV U228 ( .A(n1900), .Z(n70) );
  MUX U229 ( .IN0(n2336), .IN1(n2338), .SEL(n2337), .F(n2216) );
  MUX U230 ( .IN0(n2466), .IN1(n71), .SEL(n2467), .F(n2344) );
  IV U231 ( .A(n2468), .Z(n71) );
  MUX U232 ( .IN0(n2474), .IN1(n72), .SEL(n2475), .F(n2352) );
  IV U233 ( .A(n2476), .Z(n72) );
  MUX U234 ( .IN0(g_input[22]), .IN1(n4489), .SEL(g_input[31]), .F(n73) );
  IV U235 ( .A(n73), .Z(n1002) );
  MUX U236 ( .IN0(g_input[24]), .IN1(n4455), .SEL(g_input[31]), .F(n74) );
  IV U237 ( .A(n74), .Z(n867) );
  MUX U238 ( .IN0(g_input[17]), .IN1(n4574), .SEL(g_input[31]), .F(n75) );
  IV U239 ( .A(n75), .Z(n1410) );
  MUX U240 ( .IN0(g_input[19]), .IN1(n4540), .SEL(g_input[31]), .F(n76) );
  IV U241 ( .A(n76), .Z(n1235) );
  MUX U242 ( .IN0(g_input[26]), .IN1(n4422), .SEL(g_input[31]), .F(n77) );
  IV U243 ( .A(n77), .Z(n744) );
  MUX U244 ( .IN0(g_input[27]), .IN1(n4406), .SEL(g_input[31]), .F(n78) );
  IV U245 ( .A(n78), .Z(n702) );
  MUX U246 ( .IN0(n864), .IN1(n862), .SEL(n863), .F(n798) );
  MUX U247 ( .IN0(n2541), .IN1(n2543), .SEL(n2542), .F(n2415) );
  XNOR U248 ( .A(n1027), .B(n1026), .Z(n1093) );
  XOR U249 ( .A(n1371), .B(n1286), .Z(n1287) );
  ANDN U250 ( .A(n581), .B(n561), .Z(n550) );
  XNOR U251 ( .A(n5013), .B(n5012), .Z(n5020) );
  MUX U252 ( .IN0(n3780), .IN1(n79), .SEL(n3781), .F(n3766) );
  IV U253 ( .A(n3782), .Z(n79) );
  MUX U254 ( .IN0(n4755), .IN1(n4757), .SEL(n4756), .F(n4751) );
  MUX U255 ( .IN0(n80), .IN1(n5088), .SEL(n5089), .F(n5074) );
  IV U256 ( .A(n5090), .Z(n80) );
  MUX U257 ( .IN0(n81), .IN1(n4710), .SEL(n4711), .F(n4701) );
  IV U258 ( .A(n4712), .Z(n81) );
  XNOR U259 ( .A(n4203), .B(n4202), .Z(n4218) );
  NANDN U260 ( .B(n5201), .A(n3009), .Z(n97) );
  MUX U261 ( .IN0(n4796), .IN1(n4798), .SEL(n4797), .F(n4777) );
  XNOR U262 ( .A(n4977), .B(n4976), .Z(n4982) );
  XNOR U263 ( .A(n4804), .B(n4803), .Z(n4819) );
  XNOR U264 ( .A(n3042), .B(n3041), .Z(n3076) );
  MUX U265 ( .IN0(n1890), .IN1(n82), .SEL(n1891), .F(n1784) );
  IV U266 ( .A(n1892), .Z(n82) );
  MUX U267 ( .IN0(n2185), .IN1(n83), .SEL(n2186), .F(n2066) );
  IV U268 ( .A(n2187), .Z(n83) );
  MUX U269 ( .IN0(n2377), .IN1(n2379), .SEL(n2378), .F(n2257) );
  MUX U270 ( .IN0(n2599), .IN1(n84), .SEL(n2600), .F(n2474) );
  IV U271 ( .A(n2601), .Z(n84) );
  MUX U272 ( .IN0(g_input[12]), .IN1(n4997), .SEL(g_input[31]), .F(n85) );
  IV U273 ( .A(n85), .Z(n1906) );
  MUX U274 ( .IN0(n2794), .IN1(n2796), .SEL(n2795), .F(n2669) );
  MUX U275 ( .IN0(g_input[20]), .IN1(n4523), .SEL(g_input[31]), .F(n86) );
  IV U276 ( .A(n86), .Z(n1154) );
  MUX U277 ( .IN0(n2763), .IN1(n87), .SEL(n2764), .F(n2633) );
  IV U278 ( .A(n2765), .Z(n87) );
  MUX U279 ( .IN0(g_input[15]), .IN1(n4961), .SEL(g_input[31]), .F(n88) );
  IV U280 ( .A(n88), .Z(n1603) );
  MUX U281 ( .IN0(g_input[23]), .IN1(n4472), .SEL(g_input[31]), .F(n89) );
  IV U282 ( .A(n89), .Z(n935) );
  MUX U283 ( .IN0(g_input[21]), .IN1(n4506), .SEL(g_input[31]), .F(n90) );
  IV U284 ( .A(n90), .Z(n1076) );
  MUX U285 ( .IN0(n776), .IN1(n778), .SEL(n777), .F(n720) );
  MUX U286 ( .IN0(n932), .IN1(n930), .SEL(n931), .F(n862) );
  MUX U287 ( .IN0(n991), .IN1(n989), .SEL(n990), .F(n920) );
  MUX U288 ( .IN0(n1180), .IN1(n1178), .SEL(n1179), .F(n1100) );
  MUX U289 ( .IN0(n91), .IN1(n1314), .SEL(n1315), .F(n1230) );
  IV U290 ( .A(n1316), .Z(n91) );
  MUX U291 ( .IN0(n1945), .IN1(n1943), .SEL(n1944), .F(n1835) );
  MUX U292 ( .IN0(n92), .IN1(n2235), .SEL(n2236), .F(n2116) );
  IV U293 ( .A(n2237), .Z(n92) );
  MUX U294 ( .IN0(n655), .IN1(n653), .SEL(n654), .F(n613) );
  MUX U295 ( .IN0(n963), .IN1(n965), .SEL(n964), .F(n894) );
  MUX U296 ( .IN0(n93), .IN1(n1131), .SEL(n1132), .F(n1051) );
  IV U297 ( .A(n1133), .Z(n93) );
  XOR U298 ( .A(n348), .B(n1620), .Z(n1524) );
  MUX U299 ( .IN0(n1925), .IN1(n1927), .SEL(n1926), .F(n1818) );
  ANDN U300 ( .A(n550), .B(n532), .Z(n521) );
  AND U301 ( .A(n590), .B(n592), .Z(n559) );
  MUX U302 ( .IN0(n1342), .IN1(n1340), .SEL(n1341), .F(n1249) );
  MUX U303 ( .IN0(n5104), .IN1(n94), .SEL(n5105), .F(n5088) );
  IV U304 ( .A(n5106), .Z(n94) );
  MUX U305 ( .IN0(n4215), .IN1(n4217), .SEL(n4216), .F(n4195) );
  MUX U306 ( .IN0(n5192), .IN1(n5194), .SEL(n5193), .F(n5174) );
  XNOR U307 ( .A(n5001), .B(n5000), .Z(n5006) );
  MUX U308 ( .IN0(n95), .IN1(n3766), .SEL(n3767), .F(n3752) );
  IV U309 ( .A(n3768), .Z(n95) );
  MUX U310 ( .IN0(n96), .IN1(n4701), .SEL(n4702), .F(n4689) );
  IV U311 ( .A(n4703), .Z(n96) );
  MUX U312 ( .IN0(n5198), .IN1(n97), .SEL(n5199), .F(n5187) );
  MUX U313 ( .IN0(n4777), .IN1(n4779), .SEL(n4778), .F(n2963) );
  MUX U314 ( .IN0(n2113), .IN1(n98), .SEL(n2114), .F(n2005) );
  IV U315 ( .A(n2115), .Z(n98) );
  MUX U316 ( .IN0(n2081), .IN1(n2083), .SEL(n2082), .F(n1973) );
  MUX U317 ( .IN0(n2275), .IN1(n99), .SEL(n2276), .F(n2161) );
  IV U318 ( .A(n2277), .Z(n99) );
  MUX U319 ( .IN0(n2450), .IN1(n100), .SEL(n2451), .F(n2328) );
  IV U320 ( .A(n2452), .Z(n100) );
  MUX U321 ( .IN0(n2402), .IN1(n2404), .SEL(n2403), .F(n2282) );
  MUX U322 ( .IN0(n2715), .IN1(n2717), .SEL(n2716), .F(n2583) );
  MUX U323 ( .IN0(n2723), .IN1(n101), .SEL(n2724), .F(n2591) );
  IV U324 ( .A(n2725), .Z(n101) );
  MUX U325 ( .IN0(g_input[16]), .IN1(n4591), .SEL(g_input[31]), .F(n102) );
  IV U326 ( .A(n102), .Z(n1507) );
  MUX U327 ( .IN0(g_input[18]), .IN1(n4557), .SEL(g_input[31]), .F(n103) );
  IV U328 ( .A(n103), .Z(n1319) );
  MUX U329 ( .IN0(g_input[14]), .IN1(n4973), .SEL(g_input[31]), .F(n104) );
  IV U330 ( .A(n104), .Z(n1699) );
  MUX U331 ( .IN0(n2755), .IN1(n2757), .SEL(n2756), .F(n2625) );
  MUX U332 ( .IN0(g_input[13]), .IN1(n4985), .SEL(g_input[31]), .F(n105) );
  IV U333 ( .A(n105), .Z(n1800) );
  MUX U334 ( .IN0(n2901), .IN1(n106), .SEL(n2902), .F(n2763) );
  IV U335 ( .A(n2903), .Z(n106) );
  XNOR U336 ( .A(n3059), .B(n3058), .Z(n3838) );
  MUX U337 ( .IN0(n795), .IN1(n107), .SEL(n796), .F(n736) );
  IV U338 ( .A(n797), .Z(n107) );
  MUX U339 ( .IN0(n1029), .IN1(n1027), .SEL(n1028), .F(n959) );
  MUX U340 ( .IN0(n108), .IN1(n1071), .SEL(n1072), .F(n997) );
  IV U341 ( .A(n1073), .Z(n108) );
  MUX U342 ( .IN0(n1731), .IN1(n1733), .SEL(n1732), .F(n1630) );
  MUX U343 ( .IN0(n1351), .IN1(n1349), .SEL(n1350), .F(n1260) );
  MUX U344 ( .IN0(n1399), .IN1(n1397), .SEL(n1398), .F(n1304) );
  MUX U345 ( .IN0(n1895), .IN1(n1893), .SEL(n1894), .F(n1787) );
  MUX U346 ( .IN0(n1856), .IN1(n1854), .SEL(n1855), .F(n1746) );
  MUX U347 ( .IN0(n1879), .IN1(n1877), .SEL(n1878), .F(n1771) );
  MUX U348 ( .IN0(n2310), .IN1(n2308), .SEL(n2309), .F(n2188) );
  MUX U349 ( .IN0(n2471), .IN1(n2469), .SEL(n2470), .F(n2347) );
  MUX U350 ( .IN0(n109), .IN1(n2477), .SEL(n2478), .F(n2355) );
  IV U351 ( .A(n2479), .Z(n109) );
  MUX U352 ( .IN0(n688), .IN1(n686), .SEL(n687), .F(n643) );
  MUX U353 ( .IN0(n699), .IN1(n697), .SEL(n698), .F(n653) );
  XNOR U354 ( .A(n852), .B(n851), .Z(n913) );
  MUX U355 ( .IN0(n110), .IN1(n1294), .SEL(n1295), .F(n1210) );
  IV U356 ( .A(n1296), .Z(n110) );
  XNOR U357 ( .A(n1372), .B(n1382), .Z(n1471) );
  MUX U358 ( .IN0(n1825), .IN1(n111), .SEL(n1826), .F(n1714) );
  IV U359 ( .A(n1827), .Z(n111) );
  XOR U360 ( .A(n563), .B(n540), .Z(n537) );
  MUX U361 ( .IN0(n637), .IN1(n639), .SEL(n638), .F(n112) );
  IV U362 ( .A(n112), .Z(n603) );
  AND U363 ( .A(n671), .B(n673), .Z(n631) );
  NOR U364 ( .A(n1338), .B(n1339), .Z(n1337) );
  NANDN U365 ( .B(n509), .A(n521), .Z(n489) );
  MUX U366 ( .IN0(n524), .IN1(\_MxM/Y0[29] ), .SEL(n525), .F(n501) );
  MUX U367 ( .IN0(n4122), .IN1(n4120), .SEL(n4121), .F(n4099) );
  MUX U368 ( .IN0(n5058), .IN1(n4935), .SEL(n4936), .F(n5044) );
  MUX U369 ( .IN0(n5118), .IN1(n5120), .SEL(n5119), .F(n5115) );
  MUX U370 ( .IN0(n113), .IN1(n4715), .SEL(n4716), .F(n4696) );
  IV U371 ( .A(n4717), .Z(n113) );
  MUX U372 ( .IN0(n114), .IN1(n5074), .SEL(n5075), .F(n5065) );
  IV U373 ( .A(n5076), .Z(n114) );
  NANDN U374 ( .B(n4942), .A(n3009), .Z(n135) );
  MUX U375 ( .IN0(n4163), .IN1(n4165), .SEL(n4164), .F(n4145) );
  XNOR U376 ( .A(n4183), .B(n4182), .Z(n4198) );
  MUX U377 ( .IN0(n115), .IN1(n5142), .SEL(n5143), .F(n2995) );
  IV U378 ( .A(n5144), .Z(n115) );
  XNOR U379 ( .A(n4965), .B(n4964), .Z(n4970) );
  XNOR U380 ( .A(n4694), .B(n4693), .Z(n4699) );
  MUX U381 ( .IN0(n1858), .IN1(n1860), .SEL(n1859), .F(n1750) );
  MUX U382 ( .IN0(n1973), .IN1(n1975), .SEL(n1974), .F(n1866) );
  MUX U383 ( .IN0(n2216), .IN1(n2218), .SEL(n2217), .F(n2097) );
  MUX U384 ( .IN0(n2224), .IN1(n116), .SEL(n2225), .F(n2105) );
  IV U385 ( .A(n2226), .Z(n116) );
  MUX U386 ( .IN0(n2168), .IN1(n2170), .SEL(n2169), .F(n2054) );
  MUX U387 ( .IN0(n2305), .IN1(n117), .SEL(n2306), .F(n2185) );
  IV U388 ( .A(n2307), .Z(n117) );
  MUX U389 ( .IN0(n2501), .IN1(n2503), .SEL(n2502), .F(n2377) );
  MUX U390 ( .IN0(n2509), .IN1(n118), .SEL(n2510), .F(n2385) );
  IV U391 ( .A(n2511), .Z(n118) );
  MUX U392 ( .IN0(n2648), .IN1(n2650), .SEL(n2649), .F(n2524) );
  MUX U393 ( .IN0(n2699), .IN1(n2701), .SEL(n2700), .F(n2567) );
  MUX U394 ( .IN0(n2707), .IN1(n119), .SEL(n2708), .F(n2575) );
  IV U395 ( .A(n2709), .Z(n119) );
  MUX U396 ( .IN0(n2823), .IN1(n2825), .SEL(n2824), .F(n2691) );
  MUX U397 ( .IN0(n2816), .IN1(n120), .SEL(n2817), .F(n2684) );
  IV U398 ( .A(n2818), .Z(n120) );
  MUX U399 ( .IN0(n2863), .IN1(n121), .SEL(n2864), .F(n2731) );
  IV U400 ( .A(n2865), .Z(n121) );
  MUX U401 ( .IN0(n2771), .IN1(n122), .SEL(n2772), .F(n2641) );
  IV U402 ( .A(n2773), .Z(n122) );
  MUX U403 ( .IN0(n4775), .IN1(n4773), .SEL(n4774), .F(n2959) );
  MUX U404 ( .IN0(n3044), .IN1(n3042), .SEL(n3043), .F(n2912) );
  XNOR U405 ( .A(n3034), .B(n3033), .Z(n3096) );
  MUX U406 ( .IN0(n703), .IN1(n705), .SEL(n704), .F(n659) );
  MUX U407 ( .IN0(n1306), .IN1(n1304), .SEL(n1305), .F(n1220) );
  MUX U408 ( .IN0(n123), .IN1(n1694), .SEL(n1695), .F(n1598) );
  IV U409 ( .A(n1696), .Z(n123) );
  MUX U410 ( .IN0(n1672), .IN1(n1670), .SEL(n1671), .F(n1574) );
  MUX U411 ( .IN0(n1963), .IN1(n1961), .SEL(n1962), .F(n1854) );
  MUX U412 ( .IN0(n2002), .IN1(n2000), .SEL(n2001), .F(n1893) );
  MUX U413 ( .IN0(n2042), .IN1(n2044), .SEL(n2043), .F(n124) );
  IV U414 ( .A(n124), .Z(n1932) );
  MUX U415 ( .IN0(n2213), .IN1(n2211), .SEL(n2212), .F(n2092) );
  MUX U416 ( .IN0(n2400), .IN1(n2398), .SEL(n2399), .F(n2278) );
  MUX U417 ( .IN0(n125), .IN1(n2602), .SEL(n2603), .F(n2477) );
  IV U418 ( .A(n2604), .Z(n125) );
  MUX U419 ( .IN0(n2596), .IN1(n2594), .SEL(n2595), .F(n2469) );
  MUX U420 ( .IN0(n2557), .IN1(n2555), .SEL(n2556), .F(n2430) );
  MUX U421 ( .IN0(n2539), .IN1(n2537), .SEL(n2538), .F(n126) );
  IV U422 ( .A(n126), .Z(n2409) );
  MUX U423 ( .IN0(n2638), .IN1(n2636), .SEL(n2637), .F(n2512) );
  XNOR U424 ( .A(n2928), .B(n2927), .Z(n3052) );
  MUX U425 ( .IN0(n615), .IN1(n613), .SEL(n614), .F(n569) );
  MUX U426 ( .IN0(n800), .IN1(n798), .SEL(n799), .F(n739) );
  MUX U427 ( .IN0(n971), .IN1(n969), .SEL(n970), .F(n900) );
  MUX U428 ( .IN0(n127), .IN1(n979), .SEL(n980), .F(n910) );
  IV U429 ( .A(n981), .Z(n127) );
  XNOR U430 ( .A(n1100), .B(n1099), .Z(n1171) );
  MUX U431 ( .IN0(n128), .IN1(n1389), .SEL(n1390), .F(n1294) );
  IV U432 ( .A(n1391), .Z(n128) );
  XNOR U433 ( .A(n1717), .B(n1626), .Z(n1627) );
  MUX U434 ( .IN0(n1929), .IN1(n129), .SEL(n1930), .F(n1825) );
  IV U435 ( .A(n1931), .Z(n129) );
  MUX U436 ( .IN0(n2415), .IN1(n2417), .SEL(n2416), .F(n2297) );
  ANDN U437 ( .A(n596), .B(n600), .Z(n599) );
  MUX U438 ( .IN0(n130), .IN1(n830), .SEL(n831), .F(n771) );
  IV U439 ( .A(n832), .Z(n130) );
  ANDN U440 ( .A(n1536), .B(n1538), .Z(n1427) );
  MUX U441 ( .IN0(n178), .IN1(n2177), .SEL(n2176), .F(n2060) );
  NANDN U442 ( .B(n582), .A(n583), .Z(n551) );
  AND U443 ( .A(n631), .B(n633), .Z(n590) );
  NANDN U444 ( .B(n751), .A(n752), .Z(n707) );
  AND U445 ( .A(n949), .B(n951), .Z(n881) );
  MUX U446 ( .IN0(n1442), .IN1(n131), .SEL(n1441), .F(n1340) );
  IV U447 ( .A(n1440), .Z(n131) );
  AND U448 ( .A(n497), .B(n498), .Z(n492) );
  MUX U449 ( .IN0(n553), .IN1(\_MxM/Y0[28] ), .SEL(n554), .F(n524) );
  MUX U450 ( .IN0(n3729), .IN1(n3727), .SEL(n3728), .F(n3685) );
  MUX U451 ( .IN0(n3794), .IN1(n3796), .SEL(n3795), .F(n3791) );
  MUX U452 ( .IN0(n132), .IN1(n5079), .SEL(n5080), .F(n5060) );
  IV U453 ( .A(n5081), .Z(n132) );
  MUX U454 ( .IN0(n133), .IN1(n3752), .SEL(n3753), .F(n3743) );
  IV U455 ( .A(n3754), .Z(n133) );
  MUX U456 ( .IN0(n134), .IN1(n4696), .SEL(n4697), .F(n4684) );
  IV U457 ( .A(n4698), .Z(n134) );
  MUX U458 ( .IN0(n4939), .IN1(n135), .SEL(n4940), .F(n4927) );
  MUX U459 ( .IN0(n136), .IN1(n5065), .SEL(n5066), .F(n5053) );
  IV U460 ( .A(n5067), .Z(n136) );
  XNOR U461 ( .A(n4159), .B(n4158), .Z(n4178) );
  MUX U462 ( .IN0(n1750), .IN1(n1752), .SEL(n1751), .F(n1649) );
  MUX U463 ( .IN0(n1784), .IN1(n137), .SEL(n1785), .F(n1683) );
  IV U464 ( .A(n1786), .Z(n137) );
  MUX U465 ( .IN0(n2232), .IN1(n138), .SEL(n2233), .F(n2113) );
  IV U466 ( .A(n2234), .Z(n138) );
  MUX U467 ( .IN0(n2344), .IN1(n139), .SEL(n2345), .F(n2224) );
  IV U468 ( .A(n2346), .Z(n139) );
  MUX U469 ( .IN0(n2320), .IN1(n2322), .SEL(n2321), .F(n2200) );
  MUX U470 ( .IN0(n2434), .IN1(n2436), .SEL(n2435), .F(n2312) );
  MUX U471 ( .IN0(n2427), .IN1(n140), .SEL(n2428), .F(n2305) );
  IV U472 ( .A(n2429), .Z(n140) );
  MUX U473 ( .IN0(n2583), .IN1(n2585), .SEL(n2584), .F(n2458) );
  MUX U474 ( .IN0(n2517), .IN1(n141), .SEL(n2518), .F(n2395) );
  IV U475 ( .A(n2519), .Z(n141) );
  MUX U476 ( .IN0(n2831), .IN1(n2833), .SEL(n2832), .F(n2699) );
  MUX U477 ( .IN0(n2839), .IN1(n142), .SEL(n2840), .F(n2707) );
  IV U478 ( .A(n2841), .Z(n142) );
  MUX U479 ( .IN0(n2995), .IN1(n143), .SEL(n2996), .F(n2855) );
  IV U480 ( .A(n2997), .Z(n143) );
  MUX U481 ( .IN0(n2956), .IN1(n144), .SEL(n2957), .F(n2816) );
  IV U482 ( .A(n2958), .Z(n144) );
  MUX U483 ( .IN0(n2893), .IN1(n2895), .SEL(n2894), .F(n2755) );
  MUX U484 ( .IN0(n4965), .IN1(n4791), .SEL(n4793), .F(n2982) );
  MUX U485 ( .IN0(n745), .IN1(n747), .SEL(n746), .F(n703) );
  MUX U486 ( .IN0(n1549), .IN1(n1547), .SEL(n1548), .F(n1451) );
  MUX U487 ( .IN0(n1592), .IN1(n1590), .SEL(n1591), .F(n1494) );
  MUX U488 ( .IN0(n145), .IN1(n1598), .SEL(n1599), .F(n1502) );
  IV U489 ( .A(n1600), .Z(n145) );
  MUX U490 ( .IN0(n1986), .IN1(n1984), .SEL(n1985), .F(n1877) );
  MUX U491 ( .IN0(n146), .IN1(n2008), .SEL(n2009), .F(n1901) );
  IV U492 ( .A(n2010), .Z(n146) );
  MUX U493 ( .IN0(n2110), .IN1(n2108), .SEL(n2109), .F(n2000) );
  MUX U494 ( .IN0(n2071), .IN1(n2069), .SEL(n2070), .F(n1961) );
  MUX U495 ( .IN0(n2166), .IN1(n2164), .SEL(n2165), .F(n2050) );
  MUX U496 ( .IN0(n2580), .IN1(n2578), .SEL(n2579), .F(n2453) );
  MUX U497 ( .IN0(n2514), .IN1(n2512), .SEL(n2513), .F(n2390) );
  MUX U498 ( .IN0(n2728), .IN1(n2726), .SEL(n2727), .F(n2594) );
  MUX U499 ( .IN0(n147), .IN1(n2734), .SEL(n2735), .F(n2602) );
  IV U500 ( .A(n2736), .Z(n147) );
  MUX U501 ( .IN0(n2689), .IN1(n2687), .SEL(n2688), .F(n2555) );
  MUX U502 ( .IN0(n2776), .IN1(n2774), .SEL(n2775), .F(n2644) );
  XNOR U503 ( .A(n2904), .B(n2903), .Z(n3027) );
  MUX U504 ( .IN0(n733), .IN1(n731), .SEL(n732), .F(n686) );
  XNOR U505 ( .A(n798), .B(n797), .Z(n855) );
  MUX U506 ( .IN0(n1039), .IN1(n1041), .SEL(n1040), .F(n969) );
  XNOR U507 ( .A(n989), .B(n988), .Z(n1054) );
  XNOR U508 ( .A(n1149), .B(n1148), .Z(n1223) );
  XNOR U509 ( .A(n1178), .B(n1177), .Z(n1253) );
  MUX U510 ( .IN0(n1630), .IN1(n1632), .SEL(n1631), .F(n1529) );
  MUX U511 ( .IN0(n148), .IN1(n1368), .SEL(n1369), .F(n1277) );
  IV U512 ( .A(n1370), .Z(n148) );
  XNOR U513 ( .A(n1718), .B(n1728), .Z(n1828) );
  XOR U514 ( .A(n2146), .B(n2042), .Z(n2043) );
  MUX U515 ( .IN0(n149), .IN1(n2339), .SEL(n2340), .F(n2219) );
  IV U516 ( .A(n2341), .Z(n149) );
  MUX U517 ( .IN0(n2411), .IN1(n150), .SEL(n2410), .F(n2295) );
  IV U518 ( .A(n2409), .Z(n150) );
  MUX U519 ( .IN0(n606), .IN1(n151), .SEL(n605), .F(n578) );
  IV U520 ( .A(n604), .Z(n151) );
  XNOR U521 ( .A(n769), .B(n768), .Z(n822) );
  AND U522 ( .A(n1159), .B(n1161), .Z(n1081) );
  MUX U523 ( .IN0(n152), .IN1(n1267), .SEL(n1268), .F(n1187) );
  IV U524 ( .A(n1269), .Z(n152) );
  MUX U525 ( .IN0(n2421), .IN1(n2423), .SEL(n2422), .F(n2299) );
  NANDN U526 ( .B(n623), .A(n624), .Z(n582) );
  ANDN U527 ( .A(n662), .B(n633), .Z(n622) );
  NANDN U528 ( .B(n810), .A(n811), .Z(n751) );
  NAND U529 ( .A(n1427), .B(n1426), .Z(n1338) );
  MUX U530 ( .IN0(n153), .IN1(n1950), .SEL(n1951), .F(n1842) );
  IV U531 ( .A(n1952), .Z(n153) );
  ANDN U532 ( .A(n1090), .B(n1091), .Z(n1016) );
  MUX U533 ( .IN0(\_MxM/Y0[3] ), .IN1(n2612), .SEL(n2613), .F(n2489) );
  MUX U534 ( .IN0(n489), .IN1(n491), .SEL(n490), .F(n154) );
  IV U535 ( .A(n154), .Z(n488) );
  MUX U536 ( .IN0(n584), .IN1(\_MxM/Y0[27] ), .SEL(n585), .F(n553) );
  MUX U537 ( .IN0(n753), .IN1(\_MxM/Y0[23] ), .SEL(n754), .F(n709) );
  MUX U538 ( .IN0(n1010), .IN1(\_MxM/Y0[19] ), .SEL(n1011), .F(n943) );
  MUX U539 ( .IN0(n1327), .IN1(\_MxM/Y0[15] ), .SEL(n1328), .F(n1243) );
  MUX U540 ( .IN0(n1707), .IN1(\_MxM/Y0[11] ), .SEL(n1708), .F(n1611) );
  MUX U541 ( .IN0(n2129), .IN1(\_MxM/Y0[7] ), .SEL(n2130), .F(n2021) );
  MUX U542 ( .IN0(n4598), .IN1(n4152), .SEL(n4153), .F(n4581) );
  MUX U543 ( .IN0(n155), .IN1(n4129), .SEL(n3694), .F(n4108) );
  IV U544 ( .A(n3692), .Z(n155) );
  MUX U545 ( .IN0(n3568), .IN1(n3566), .SEL(n3567), .F(n3522) );
  MUX U546 ( .IN0(n4289), .IN1(n4287), .SEL(n4288), .F(n4263) );
  XNOR U547 ( .A(n4864), .B(n4863), .Z(n4879) );
  MUX U548 ( .IN0(n4321), .IN1(n4323), .SEL(n4322), .F(n4318) );
  MUX U549 ( .IN0(n156), .IN1(n3757), .SEL(n3758), .F(n3736) );
  IV U550 ( .A(n3759), .Z(n156) );
  NANDN U551 ( .B(n1623), .A(n3009), .Z(n188) );
  MUX U552 ( .IN0(n157), .IN1(n5133), .SEL(n5134), .F(n2987) );
  IV U553 ( .A(n5135), .Z(n157) );
  MUX U554 ( .IN0(n4784), .IN1(n4786), .SEL(n4785), .F(n2971) );
  MUX U555 ( .IN0(n3847), .IN1(n3845), .SEL(n3846), .F(n3059) );
  MUX U556 ( .IN0(n1866), .IN1(n1868), .SEL(n1867), .F(n1758) );
  MUX U557 ( .IN0(n1989), .IN1(n1991), .SEL(n1990), .F(n1882) );
  MUX U558 ( .IN0(n2073), .IN1(n2075), .SEL(n2074), .F(n1965) );
  MUX U559 ( .IN0(n2066), .IN1(n158), .SEL(n2067), .F(n1958) );
  IV U560 ( .A(n2068), .Z(n158) );
  MUX U561 ( .IN0(n2328), .IN1(n159), .SEL(n2329), .F(n2208) );
  IV U562 ( .A(n2330), .Z(n159) );
  MUX U563 ( .IN0(n2442), .IN1(n2444), .SEL(n2443), .F(n2320) );
  MUX U564 ( .IN0(n2458), .IN1(n2460), .SEL(n2459), .F(n2336) );
  MUX U565 ( .IN0(n2591), .IN1(n160), .SEL(n2592), .F(n2466) );
  IV U566 ( .A(n2593), .Z(n160) );
  MUX U567 ( .IN0(n2552), .IN1(n161), .SEL(n2553), .F(n2427) );
  IV U568 ( .A(n2554), .Z(n161) );
  MUX U569 ( .IN0(n2641), .IN1(n162), .SEL(n2642), .F(n2517) );
  IV U570 ( .A(n2643), .Z(n162) );
  MUX U571 ( .IN0(n2731), .IN1(n163), .SEL(n2732), .F(n2599) );
  IV U572 ( .A(n2733), .Z(n163) );
  MUX U573 ( .IN0(n2691), .IN1(n2693), .SEL(n2692), .F(n2559) );
  MUX U574 ( .IN0(g_input[8]), .IN1(n5052), .SEL(g_input[31]), .F(n164) );
  IV U575 ( .A(n164), .Z(n2360) );
  MUX U576 ( .IN0(n2979), .IN1(n165), .SEL(n2980), .F(n2839) );
  IV U577 ( .A(n2981), .Z(n165) );
  MUX U578 ( .IN0(n2932), .IN1(n2934), .SEL(n2933), .F(n2794) );
  MUX U579 ( .IN0(n854), .IN1(n852), .SEL(n853), .F(n790) );
  MUX U580 ( .IN0(n1748), .IN1(n1746), .SEL(n1747), .F(n1645) );
  MUX U581 ( .IN0(n1789), .IN1(n1787), .SEL(n1788), .F(n1686) );
  MUX U582 ( .IN0(n1720), .IN1(n1718), .SEL(n1719), .F(n1626) );
  MUX U583 ( .IN0(n166), .IN1(n1901), .SEL(n1902), .F(n1795) );
  IV U584 ( .A(n1903), .Z(n166) );
  MUX U585 ( .IN0(n2094), .IN1(n2092), .SEL(n2093), .F(n1984) );
  MUX U586 ( .IN0(n2190), .IN1(n2188), .SEL(n2189), .F(n2069) );
  MUX U587 ( .IN0(n2229), .IN1(n2227), .SEL(n2228), .F(n2108) );
  MUX U588 ( .IN0(n2149), .IN1(n2147), .SEL(n2148), .F(n2042) );
  MUX U589 ( .IN0(n2280), .IN1(n2278), .SEL(n2279), .F(n2164) );
  MUX U590 ( .IN0(n167), .IN1(n2355), .SEL(n2356), .F(n2235) );
  IV U591 ( .A(n2357), .Z(n167) );
  MUX U592 ( .IN0(n2658), .IN1(n2656), .SEL(n2657), .F(n2537) );
  MUX U593 ( .IN0(n2712), .IN1(n2710), .SEL(n2711), .F(n2578) );
  MUX U594 ( .IN0(n2821), .IN1(n2819), .SEL(n2820), .F(n2687) );
  MUX U595 ( .IN0(n2860), .IN1(n2858), .SEL(n2859), .F(n2726) );
  MUX U596 ( .IN0(n168), .IN1(n2866), .SEL(n2867), .F(n2734) );
  IV U597 ( .A(n2868), .Z(n168) );
  MUX U598 ( .IN0(n2768), .IN1(n2766), .SEL(n2767), .F(n2636) );
  MUX U599 ( .IN0(n2914), .IN1(n2912), .SEL(n2913), .F(n2774) );
  MUX U600 ( .IN0(n619), .IN1(n621), .SEL(n620), .F(n575) );
  MUX U601 ( .IN0(n741), .IN1(n739), .SEL(n740), .F(n697) );
  XNOR U602 ( .A(n930), .B(n929), .Z(n992) );
  XNOR U603 ( .A(n1141), .B(n1140), .Z(n1213) );
  XNOR U604 ( .A(n1230), .B(n1229), .Z(n1307) );
  XNOR U605 ( .A(n1260), .B(n1259), .Z(n1344) );
  MUX U606 ( .IN0(n169), .IN1(n1486), .SEL(n1487), .F(n1389) );
  IV U607 ( .A(n1488), .Z(n169) );
  XNOR U608 ( .A(n1478), .B(n1477), .Z(n1567) );
  MUX U609 ( .IN0(n2033), .IN1(n170), .SEL(n2034), .F(n1929) );
  IV U610 ( .A(n2035), .Z(n170) );
  MUX U611 ( .IN0(n171), .IN1(n2100), .SEL(n2101), .F(n1992) );
  IV U612 ( .A(n2102), .Z(n171) );
  MUX U613 ( .IN0(n172), .IN1(n2323), .SEL(n2324), .F(n2203) );
  IV U614 ( .A(n2325), .Z(n172) );
  MUX U615 ( .IN0(n173), .IN1(n2586), .SEL(n2587), .F(n2461) );
  IV U616 ( .A(n2588), .Z(n173) );
  MUX U617 ( .IN0(n174), .IN1(n2504), .SEL(n2505), .F(n2380) );
  IV U618 ( .A(n2506), .Z(n174) );
  MUX U619 ( .IN0(n175), .IN1(n566), .SEL(n565), .F(n540) );
  IV U620 ( .A(n564), .Z(n175) );
  AND U621 ( .A(n602), .B(n603), .Z(n598) );
  MUX U622 ( .IN0(n889), .IN1(n887), .SEL(n888), .F(n827) );
  MUX U623 ( .IN0(n176), .IN1(n1034), .SEL(n1035), .F(n966) );
  IV U624 ( .A(n1036), .Z(n176) );
  AND U625 ( .A(n1240), .B(n1242), .Z(n1159) );
  MUX U626 ( .IN0(n1529), .IN1(n1531), .SEL(n1530), .F(n1438) );
  MUX U627 ( .IN0(n177), .IN1(n1753), .SEL(n1754), .F(n1652) );
  IV U628 ( .A(n1755), .Z(n177) );
  ANDN U629 ( .A(n1737), .B(n1739), .Z(n1636) );
  AND U630 ( .A(n2018), .B(n2020), .Z(n1911) );
  MUX U631 ( .IN0(n2301), .IN1(n2299), .SEL(n2300), .F(n178) );
  IV U632 ( .A(n178), .Z(n2175) );
  NANDN U633 ( .B(n663), .A(n664), .Z(n623) );
  MUX U634 ( .IN0(n750), .IN1(n179), .SEL(n749), .F(n706) );
  IV U635 ( .A(n748), .Z(n179) );
  AND U636 ( .A(n818), .B(n820), .Z(n807) );
  NANDN U637 ( .B(n873), .A(n874), .Z(n810) );
  MUX U638 ( .IN0(n180), .IN1(n1533), .SEL(n1534), .F(n1440) );
  IV U639 ( .A(n1535), .Z(n180) );
  MUX U640 ( .IN0(n181), .IN1(n2057), .SEL(n2058), .F(n1950) );
  IV U641 ( .A(n2059), .Z(n181) );
  MUX U642 ( .IN0(n2529), .IN1(n208), .SEL(n2528), .F(n182) );
  IV U643 ( .A(n182), .Z(n2405) );
  AND U644 ( .A(n530), .B(n532), .Z(n507) );
  ANDN U645 ( .A(n1168), .B(n1169), .Z(n1090) );
  NAND U646 ( .A(n478), .B(n480), .Z(n477) );
  MUX U647 ( .IN0(n625), .IN1(\_MxM/Y0[26] ), .SEL(n626), .F(n584) );
  MUX U648 ( .IN0(n812), .IN1(\_MxM/Y0[22] ), .SEL(n813), .F(n753) );
  MUX U649 ( .IN0(n1084), .IN1(\_MxM/Y0[18] ), .SEL(n1085), .F(n1010) );
  MUX U650 ( .IN0(n1418), .IN1(\_MxM/Y0[14] ), .SEL(n1419), .F(n1327) );
  MUX U651 ( .IN0(n1808), .IN1(\_MxM/Y0[10] ), .SEL(n1809), .F(n1707) );
  MUX U652 ( .IN0(n2248), .IN1(\_MxM/Y0[6] ), .SEL(n2249), .F(n2129) );
  MUX U653 ( .IN0(n4143), .IN1(n4141), .SEL(n4142), .F(n4120) );
  MUX U654 ( .IN0(n3718), .IN1(n3716), .SEL(n3717), .F(n183) );
  IV U655 ( .A(n183), .Z(n3674) );
  MUX U656 ( .IN0(n3641), .IN1(n3639), .SEL(n3640), .F(n3593) );
  MUX U657 ( .IN0(n4564), .IN1(n4110), .SEL(n4111), .F(n4547) );
  MUX U658 ( .IN0(n184), .IN1(n4045), .SEL(n3512), .F(n4024) );
  IV U659 ( .A(n3510), .Z(n184) );
  MUX U660 ( .IN0(n4694), .IN1(n4314), .SEL(n4315), .F(n4682) );
  MUX U661 ( .IN0(n4932), .IN1(n4930), .SEL(n4931), .F(n4910) );
  XNOR U662 ( .A(n4263), .B(n4262), .Z(n4280) );
  MUX U663 ( .IN0(n185), .IN1(n3961), .SEL(n3330), .F(n3940) );
  IV U664 ( .A(n3328), .Z(n185) );
  MUX U665 ( .IN0(n4640), .IN1(n4230), .SEL(n4232), .F(n4628) );
  MUX U666 ( .IN0(n5202), .IN1(n5204), .SEL(n5203), .F(n5198) );
  MUX U667 ( .IN0(n4846), .IN1(n4844), .SEL(n4845), .F(n4824) );
  MUX U668 ( .IN0(n186), .IN1(n5158), .SEL(n5159), .F(n5133) );
  IV U669 ( .A(n5160), .Z(n186) );
  MUX U670 ( .IN0(n187), .IN1(n5060), .SEL(n5061), .F(n5046) );
  IV U671 ( .A(n5062), .Z(n187) );
  MUX U672 ( .IN0(n3812), .IN1(n188), .SEL(n3813), .F(n3698) );
  MUX U673 ( .IN0(n189), .IN1(n3878), .SEL(n3157), .F(n3857) );
  IV U674 ( .A(n3155), .Z(n189) );
  MUX U675 ( .IN0(n1882), .IN1(n1884), .SEL(n1883), .F(n1776) );
  MUX U676 ( .IN0(n2855), .IN1(n190), .SEL(n2856), .F(n2723) );
  IV U677 ( .A(n2857), .Z(n190) );
  MUX U678 ( .IN0(g_input[7]), .IN1(n5141), .SEL(g_input[31]), .F(n191) );
  IV U679 ( .A(n191), .Z(n2482) );
  MUX U680 ( .IN0(g_input[11]), .IN1(n5009), .SEL(g_input[31]), .F(n192) );
  IV U681 ( .A(n192), .Z(n2013) );
  MUX U682 ( .IN0(n2916), .IN1(n2918), .SEL(n2917), .F(n2778) );
  MUX U683 ( .IN0(n2909), .IN1(n193), .SEL(n2910), .F(n2771) );
  IV U684 ( .A(n2911), .Z(n193) );
  MUX U685 ( .IN0(n3036), .IN1(n3034), .SEL(n3035), .F(n2904) );
  MUX U686 ( .IN0(n804), .IN1(n806), .SEL(n805), .F(n745) );
  MUX U687 ( .IN0(n1222), .IN1(n1220), .SEL(n1221), .F(n1141) );
  MUX U688 ( .IN0(n1374), .IN1(n1372), .SEL(n1373), .F(n1286) );
  MUX U689 ( .IN0(n1773), .IN1(n1771), .SEL(n1772), .F(n1670) );
  MUX U690 ( .IN0(n2333), .IN1(n2331), .SEL(n2332), .F(n2211) );
  MUX U691 ( .IN0(n2432), .IN1(n2430), .SEL(n2431), .F(n2308) );
  MUX U692 ( .IN0(n2646), .IN1(n2644), .SEL(n2645), .F(n2520) );
  MUX U693 ( .IN0(n2844), .IN1(n2842), .SEL(n2843), .F(n2710) );
  MUX U694 ( .IN0(n194), .IN1(n3006), .SEL(n3007), .F(n2866) );
  IV U695 ( .A(n3008), .Z(n194) );
  MUX U696 ( .IN0(n3000), .IN1(n2998), .SEL(n2999), .F(n2858) );
  MUX U697 ( .IN0(n2961), .IN1(n2959), .SEL(n2960), .F(n2819) );
  XNOR U698 ( .A(n862), .B(n861), .Z(n923) );
  XNOR U699 ( .A(n920), .B(n919), .Z(n982) );
  XNOR U700 ( .A(n1071), .B(n1070), .Z(n1144) );
  MUX U701 ( .IN0(n1200), .IN1(n195), .SEL(n1201), .F(n1121) );
  IV U702 ( .A(n1202), .Z(n195) );
  XNOR U703 ( .A(n1314), .B(n1313), .Z(n1400) );
  XNOR U704 ( .A(n1349), .B(n1348), .Z(n1444) );
  XNOR U705 ( .A(n1494), .B(n1493), .Z(n1585) );
  MUX U706 ( .IN0(n196), .IN1(n1678), .SEL(n1679), .F(n1582) );
  IV U707 ( .A(n1680), .Z(n196) );
  XNOR U708 ( .A(n1598), .B(n1597), .Z(n1689) );
  XNOR U709 ( .A(n1645), .B(n1644), .Z(n1741) );
  MUX U710 ( .IN0(n197), .IN1(n1869), .SEL(n1870), .F(n1761) );
  IV U711 ( .A(n1871), .Z(n197) );
  XNOR U712 ( .A(n1893), .B(n1892), .Z(n1995) );
  XNOR U713 ( .A(n1901), .B(n1900), .Z(n2003) );
  XNOR U714 ( .A(n2050), .B(n2049), .Z(n2159) );
  XNOR U715 ( .A(n2227), .B(n2226), .Z(n2342) );
  XNOR U716 ( .A(n2235), .B(n2234), .Z(n2350) );
  XNOR U717 ( .A(n2270), .B(n2269), .Z(n2383) );
  MUX U718 ( .IN0(n198), .IN1(n2570), .SEL(n2571), .F(n2445) );
  IV U719 ( .A(n2572), .Z(n198) );
  XNOR U720 ( .A(n2656), .B(n2666), .Z(n2785) );
  MUX U721 ( .IN0(n199), .IN1(n2758), .SEL(n2759), .F(n2628) );
  IV U722 ( .A(n2760), .Z(n199) );
  XNOR U723 ( .A(n569), .B(n566), .Z(n607) );
  MUX U724 ( .IN0(n645), .IN1(n643), .SEL(n644), .F(n596) );
  MUX U725 ( .IN0(n200), .IN1(n681), .SEL(n682), .F(n640) );
  IV U726 ( .A(n683), .Z(n200) );
  AND U727 ( .A(n900), .B(n902), .Z(n833) );
  MUX U728 ( .IN0(n201), .IN1(n1109), .SEL(n1110), .F(n1034) );
  IV U729 ( .A(n1111), .Z(n201) );
  MUX U730 ( .IN0(n1525), .IN1(n348), .SEL(n1524), .F(n1437) );
  AND U731 ( .A(n1608), .B(n1610), .Z(n1512) );
  ANDN U732 ( .A(n1845), .B(n1847), .Z(n1737) );
  MUX U733 ( .IN0(n202), .IN1(n1968), .SEL(n1969), .F(n1861) );
  IV U734 ( .A(n1970), .Z(n202) );
  AND U735 ( .A(n2245), .B(n2247), .Z(n2126) );
  MUX U736 ( .IN0(n203), .IN1(n2437), .SEL(n2438), .F(n2315) );
  IV U737 ( .A(n2439), .Z(n203) );
  MUX U738 ( .IN0(n204), .IN1(n2548), .SEL(n2547), .F(n2421) );
  IV U739 ( .A(n2546), .Z(n204) );
  NANDN U740 ( .B(n551), .A(n552), .Z(n522) );
  ANDN U741 ( .A(n706), .B(n673), .Z(n662) );
  NANDN U742 ( .B(n707), .A(n708), .Z(n663) );
  MUX U743 ( .IN0(n829), .IN1(n827), .SEL(n828), .F(n205) );
  IV U744 ( .A(n205), .Z(n767) );
  OR U745 ( .A(n1008), .B(n1009), .Z(n941) );
  MUX U746 ( .IN0(n206), .IN1(n1633), .SEL(n1634), .F(n1533) );
  IV U747 ( .A(n1635), .Z(n206) );
  MUX U748 ( .IN0(n207), .IN1(n2171), .SEL(n2172), .F(n2057) );
  IV U749 ( .A(n2173), .Z(n207) );
  MUX U750 ( .IN0(n2653), .IN1(n241), .SEL(n2652), .F(n208) );
  IV U751 ( .A(n208), .Z(n2527) );
  AND U752 ( .A(n807), .B(n809), .Z(n715) );
  MUX U753 ( .IN0(n209), .IN1(n1249), .SEL(n1250), .F(n1168) );
  IV U754 ( .A(n1251), .Z(n209) );
  ANDN U755 ( .A(n482), .B(n483), .Z(n474) );
  MUX U756 ( .IN0(n665), .IN1(\_MxM/Y0[25] ), .SEL(n666), .F(n625) );
  MUX U757 ( .IN0(n875), .IN1(\_MxM/Y0[21] ), .SEL(n876), .F(n812) );
  MUX U758 ( .IN0(n1162), .IN1(\_MxM/Y0[17] ), .SEL(n1163), .F(n1084) );
  MUX U759 ( .IN0(n1515), .IN1(\_MxM/Y0[13] ), .SEL(n1516), .F(n1418) );
  MUX U760 ( .IN0(n1914), .IN1(\_MxM/Y0[9] ), .SEL(n1915), .F(n1808) );
  MUX U761 ( .IN0(n2368), .IN1(\_MxM/Y0[5] ), .SEL(n2369), .F(n2248) );
  MUX U762 ( .IN0(n501), .IN1(\_MxM/Y0[30] ), .SEL(n502), .F(n467) );
  MUX U763 ( .IN0(n3049), .IN1(n3730), .SEL(n3050), .F(n210) );
  IV U764 ( .A(n210), .Z(n3688) );
  MUX U765 ( .IN0(n211), .IN1(n3674), .SEL(n3675), .F(n3628) );
  IV U766 ( .A(n3676), .Z(n211) );
  MUX U767 ( .IN0(n4080), .IN1(n4078), .SEL(n4079), .F(n4057) );
  MUX U768 ( .IN0(n3595), .IN1(n3593), .SEL(n3594), .F(n3547) );
  MUX U769 ( .IN0(n212), .IN1(n3492), .SEL(n3493), .F(n3446) );
  IV U770 ( .A(n3494), .Z(n212) );
  MUX U771 ( .IN0(n4496), .IN1(n4026), .SEL(n4027), .F(n4479) );
  MUX U772 ( .IN0(n3386), .IN1(n3384), .SEL(n3385), .F(n3340) );
  MUX U773 ( .IN0(n3996), .IN1(n3994), .SEL(n3995), .F(n3973) );
  MUX U774 ( .IN0(n3413), .IN1(n3411), .SEL(n3412), .F(n3365) );
  MUX U775 ( .IN0(n4780), .IN1(n4933), .SEL(n4781), .F(n213) );
  IV U776 ( .A(n213), .Z(n4913) );
  MUX U777 ( .IN0(n214), .IN1(n3310), .SEL(n3311), .F(n3265) );
  IV U778 ( .A(n3312), .Z(n214) );
  MUX U779 ( .IN0(n4428), .IN1(n3942), .SEL(n3943), .F(n4412) );
  MUX U780 ( .IN0(n5013), .IN1(n4871), .SEL(n4873), .F(n5001) );
  MUX U781 ( .IN0(n3210), .IN1(n3208), .SEL(n3209), .F(n3166) );
  MUX U782 ( .IN0(n4751), .IN1(n215), .SEL(n4752), .F(n4740) );
  IV U783 ( .A(n4754), .Z(n215) );
  MUX U784 ( .IN0(n3912), .IN1(n3910), .SEL(n3911), .F(n3890) );
  MUX U785 ( .IN0(n3235), .IN1(n3233), .SEL(n3234), .F(n3190) );
  MUX U786 ( .IN0(n4943), .IN1(n4945), .SEL(n4944), .F(n4939) );
  MUX U787 ( .IN0(n4205), .IN1(n4203), .SEL(n4204), .F(n4183) );
  NANDN U788 ( .B(n5222), .A(n3009), .Z(n250) );
  MUX U789 ( .IN0(n216), .IN1(n3137), .SEL(n3138), .F(n3093) );
  IV U790 ( .A(n3139), .Z(n216) );
  MUX U791 ( .IN0(n2312), .IN1(n2314), .SEL(n2313), .F(n2192) );
  MUX U792 ( .IN0(n2684), .IN1(n217), .SEL(n2685), .F(n2552) );
  IV U793 ( .A(n2686), .Z(n217) );
  MUX U794 ( .IN0(g_input[10]), .IN1(n5023), .SEL(g_input[31]), .F(n218) );
  IV U795 ( .A(n218), .Z(n2121) );
  MUX U796 ( .IN0(g_input[6]), .IN1(n5152), .SEL(g_input[31]), .F(n219) );
  IV U797 ( .A(n219), .Z(n2607) );
  MUX U798 ( .IN0(g_input[5]), .IN1(n5168), .SEL(g_input[31]), .F(n220) );
  IV U799 ( .A(n220), .Z(n2739) );
  MUX U800 ( .IN0(n4362), .IN1(n3859), .SEL(n3860), .F(n4342) );
  XNOR U801 ( .A(n4598), .B(n4596), .Z(n4603) );
  MUX U802 ( .IN0(n3061), .IN1(n3059), .SEL(n3060), .F(n2928) );
  MUX U803 ( .IN0(n736), .IN1(n221), .SEL(n737), .F(n694) );
  IV U804 ( .A(n738), .Z(n221) );
  MUX U805 ( .IN0(n290), .IN1(n1204), .SEL(n1203), .F(n1115) );
  MUX U806 ( .IN0(n1576), .IN1(n1574), .SEL(n1575), .F(n1478) );
  MUX U807 ( .IN0(n222), .IN1(n1795), .SEL(n1796), .F(n1694) );
  IV U808 ( .A(n1797), .Z(n222) );
  MUX U809 ( .IN0(n2455), .IN1(n2453), .SEL(n2454), .F(n2331) );
  MUX U810 ( .IN0(n2392), .IN1(n2390), .SEL(n2391), .F(n2270) );
  MUX U811 ( .IN0(n2522), .IN1(n2520), .SEL(n2521), .F(n2398) );
  MUX U812 ( .IN0(n2984), .IN1(n2982), .SEL(n2983), .F(n2842) );
  MUX U813 ( .IN0(n2906), .IN1(n2904), .SEL(n2905), .F(n2766) );
  XNOR U814 ( .A(n2998), .B(n2997), .Z(n5138) );
  XNOR U815 ( .A(n2959), .B(n2958), .Z(n4768) );
  XNOR U816 ( .A(n2912), .B(n2911), .Z(n3037) );
  MUX U817 ( .IN0(n961), .IN1(n959), .SEL(n960), .F(n887) );
  MUX U818 ( .IN0(n792), .IN1(n790), .SEL(n791), .F(n731) );
  XNOR U819 ( .A(n997), .B(n996), .Z(n1064) );
  MUX U820 ( .IN0(n1123), .IN1(n223), .SEL(n1122), .F(n1039) );
  IV U821 ( .A(n1121), .Z(n223) );
  XNOR U822 ( .A(n1061), .B(n1060), .Z(n1134) );
  XNOR U823 ( .A(n1397), .B(n1396), .Z(n1489) );
  XNOR U824 ( .A(n1405), .B(n1404), .Z(n1497) );
  XNOR U825 ( .A(n1451), .B(n1450), .Z(n1540) );
  MUX U826 ( .IN0(n224), .IN1(n1660), .SEL(n1661), .F(n1564) );
  IV U827 ( .A(n1662), .Z(n224) );
  XNOR U828 ( .A(n1686), .B(n1685), .Z(n1782) );
  MUX U829 ( .IN0(n225), .IN1(n1885), .SEL(n1886), .F(n1779) );
  IV U830 ( .A(n1887), .Z(n225) );
  XNOR U831 ( .A(n1854), .B(n1853), .Z(n1956) );
  XNOR U832 ( .A(n1943), .B(n1942), .Z(n2045) );
  XNOR U833 ( .A(n1984), .B(n1983), .Z(n2087) );
  MUX U834 ( .IN0(n226), .IN1(n2203), .SEL(n2204), .F(n2084) );
  IV U835 ( .A(n2205), .Z(n226) );
  MUX U836 ( .IN0(n227), .IN1(n2260), .SEL(n2261), .F(n2143) );
  IV U837 ( .A(n2262), .Z(n227) );
  XNOR U838 ( .A(n2308), .B(n2307), .Z(n2425) );
  XNOR U839 ( .A(n2347), .B(n2346), .Z(n2464) );
  XNOR U840 ( .A(n2355), .B(n2354), .Z(n2472) );
  XNOR U841 ( .A(n2655), .B(n2537), .Z(n2538) );
  MUX U842 ( .IN0(n228), .IN1(n2834), .SEL(n2835), .F(n2702) );
  IV U843 ( .A(n2836), .Z(n228) );
  MUX U844 ( .IN0(n2852), .IN1(n298), .SEL(n2851), .F(n229) );
  IV U845 ( .A(n229), .Z(n2718) );
  MUX U846 ( .IN0(n230), .IN1(n2810), .SEL(n2811), .F(n2677) );
  IV U847 ( .A(n2812), .Z(n230) );
  MUX U848 ( .IN0(n575), .IN1(n577), .SEL(n576), .F(n545) );
  XNOR U849 ( .A(n613), .B(n612), .Z(n646) );
  MUX U850 ( .IN0(n231), .IN1(n723), .SEL(n724), .F(n681) );
  IV U851 ( .A(n725), .Z(n231) );
  MUX U852 ( .IN0(n232), .IN1(n897), .SEL(n898), .F(n830) );
  IV U853 ( .A(n899), .Z(n232) );
  MUX U854 ( .IN0(n233), .IN1(n1187), .SEL(n1188), .F(n1109) );
  IV U855 ( .A(n1189), .Z(n233) );
  AND U856 ( .A(n1415), .B(n1417), .Z(n1324) );
  MUX U857 ( .IN0(n234), .IN1(n1554), .SEL(n1555), .F(n1458) );
  IV U858 ( .A(n1556), .Z(n234) );
  XNOR U859 ( .A(n1436), .B(n1437), .Z(n1433) );
  AND U860 ( .A(n1636), .B(n1638), .Z(n1536) );
  AND U861 ( .A(n1805), .B(n1807), .Z(n1704) );
  MUX U862 ( .IN0(n235), .IN1(n2076), .SEL(n2077), .F(n1968) );
  IV U863 ( .A(n2078), .Z(n235) );
  AND U864 ( .A(n2365), .B(n2367), .Z(n2245) );
  MUX U865 ( .IN0(n236), .IN1(n2562), .SEL(n2563), .F(n2437) );
  IV U866 ( .A(n2564), .Z(n236) );
  MUX U867 ( .IN0(n237), .IN1(n2674), .SEL(n2675), .F(n2546) );
  IV U868 ( .A(n2676), .Z(n237) );
  NAND U869 ( .A(n540), .B(n539), .Z(n534) );
  XNOR U870 ( .A(n578), .B(n603), .Z(n594) );
  ANDN U871 ( .A(n715), .B(n716), .Z(n671) );
  AND U872 ( .A(n763), .B(n764), .Z(n762) );
  ANDN U873 ( .A(n1016), .B(n1017), .Z(n949) );
  NAND U874 ( .A(n1081), .B(n1083), .Z(n1008) );
  MUX U875 ( .IN0(n238), .IN1(n1842), .SEL(n1843), .F(n1734) );
  IV U876 ( .A(n1844), .Z(n238) );
  MUX U877 ( .IN0(n239), .IN1(n2060), .SEL(n2061), .F(n1953) );
  IV U878 ( .A(n2062), .Z(n239) );
  MUX U879 ( .IN0(n240), .IN1(n2285), .SEL(n2286), .F(n2171) );
  IV U880 ( .A(n2287), .Z(n240) );
  MUX U881 ( .IN0(n2783), .IN1(n272), .SEL(n2782), .F(n241) );
  IV U882 ( .A(n241), .Z(n2651) );
  XNOR U883 ( .A(n551), .B(n556), .Z(n552) );
  XNOR U884 ( .A(n663), .B(n668), .Z(n664) );
  XNOR U885 ( .A(n810), .B(n815), .Z(n811) );
  XOR U886 ( .A(n1249), .B(n1338), .Z(n1333) );
  XNOR U887 ( .A(n2921), .B(n2920), .Z(n2751) );
  MUX U888 ( .IN0(n709), .IN1(\_MxM/Y0[24] ), .SEL(n710), .F(n665) );
  MUX U889 ( .IN0(n943), .IN1(\_MxM/Y0[20] ), .SEL(n944), .F(n875) );
  MUX U890 ( .IN0(n1243), .IN1(\_MxM/Y0[16] ), .SEL(n1244), .F(n1162) );
  MUX U891 ( .IN0(n1611), .IN1(\_MxM/Y0[12] ), .SEL(n1612), .F(n1515) );
  MUX U892 ( .IN0(n2021), .IN1(\_MxM/Y0[8] ), .SEL(n2022), .F(n1914) );
  MUX U893 ( .IN0(\_MxM/Y0[4] ), .IN1(n2489), .SEL(n2490), .F(n2368) );
  XNOR U894 ( .A(n501), .B(n505), .Z(n503) );
  MUX U895 ( .IN0(n3660), .IN1(n3658), .SEL(n3659), .F(n3612) );
  MUX U896 ( .IN0(n4581), .IN1(n4131), .SEL(n4132), .F(n4564) );
  MUX U897 ( .IN0(n242), .IN1(n4108), .SEL(n3648), .F(n4087) );
  IV U898 ( .A(n3646), .Z(n242) );
  MUX U899 ( .IN0(n4059), .IN1(n4057), .SEL(n4058), .F(n4036) );
  MUX U900 ( .IN0(n3549), .IN1(n3547), .SEL(n3548), .F(n3503) );
  MUX U901 ( .IN0(n243), .IN1(n3582), .SEL(n3583), .F(n3536) );
  IV U902 ( .A(n3584), .Z(n243) );
  MUX U903 ( .IN0(n3478), .IN1(n3476), .SEL(n3477), .F(n3430) );
  MUX U904 ( .IN0(n4513), .IN1(n4047), .SEL(n4048), .F(n4496) );
  MUX U905 ( .IN0(n4311), .IN1(n4309), .SEL(n4310), .F(n4287) );
  MUX U906 ( .IN0(n244), .IN1(n4024), .SEL(n3466), .F(n4003) );
  IV U907 ( .A(n3464), .Z(n244) );
  MUX U908 ( .IN0(n4682), .IN1(n4294), .SEL(n4296), .F(n4670) );
  MUX U909 ( .IN0(n3975), .IN1(n3973), .SEL(n3974), .F(n3952) );
  MUX U910 ( .IN0(n3367), .IN1(n3365), .SEL(n3366), .F(n3321) );
  MUX U911 ( .IN0(n245), .IN1(n3400), .SEL(n3401), .F(n3354) );
  IV U912 ( .A(n3402), .Z(n245) );
  MUX U913 ( .IN0(n3296), .IN1(n3294), .SEL(n3295), .F(n3251) );
  MUX U914 ( .IN0(n4445), .IN1(n3963), .SEL(n3964), .F(n4428) );
  MUX U915 ( .IN0(n4748), .IN1(n4334), .SEL(n4335), .F(n246) );
  IV U916 ( .A(n246), .Z(n4734) );
  MUX U917 ( .IN0(n4866), .IN1(n4864), .SEL(n4865), .F(n4844) );
  MUX U918 ( .IN0(n4225), .IN1(n4223), .SEL(n4224), .F(n4203) );
  MUX U919 ( .IN0(n247), .IN1(n3940), .SEL(n3284), .F(n3919) );
  IV U920 ( .A(n3282), .Z(n247) );
  MUX U921 ( .IN0(n5001), .IN1(n4851), .SEL(n4853), .F(n4989) );
  MUX U922 ( .IN0(n3815), .IN1(n3817), .SEL(n3816), .F(n3812) );
  MUX U923 ( .IN0(n4628), .IN1(n4210), .SEL(n4212), .F(n4618) );
  MUX U924 ( .IN0(n3892), .IN1(n3890), .SEL(n3891), .F(n3869) );
  MUX U925 ( .IN0(n3192), .IN1(n3190), .SEL(n3191), .F(n3148) );
  MUX U926 ( .IN0(n248), .IN1(n3222), .SEL(n3223), .F(n3180) );
  IV U927 ( .A(n3224), .Z(n248) );
  MUX U928 ( .IN0(n3123), .IN1(n3121), .SEL(n3122), .F(n3081) );
  MUX U929 ( .IN0(n249), .IN1(n3736), .SEL(n3737), .F(n3711) );
  IV U930 ( .A(n3738), .Z(n249) );
  XNOR U931 ( .A(n5217), .B(g_input[3]), .Z(n5218) );
  XNOR U932 ( .A(n4471), .B(g_input[23]), .Z(n4472) );
  MUX U933 ( .IN0(n4379), .IN1(n3880), .SEL(n3881), .F(n4362) );
  MUX U934 ( .IN0(n5219), .IN1(n250), .SEL(n5220), .F(n3003) );
  MUX U935 ( .IN0(n2097), .IN1(n2099), .SEL(n2098), .F(n1989) );
  MUX U936 ( .IN0(n2352), .IN1(n251), .SEL(n2353), .F(n2232) );
  IV U937 ( .A(n2354), .Z(n251) );
  MUX U938 ( .IN0(n2567), .IN1(n2569), .SEL(n2568), .F(n2442) );
  MUX U939 ( .IN0(n2524), .IN1(n2526), .SEL(n2525), .F(n2402) );
  MUX U940 ( .IN0(n2847), .IN1(n2849), .SEL(n2848), .F(n2715) );
  XNOR U941 ( .A(n5058), .B(n5057), .Z(n5063) );
  XNOR U942 ( .A(n4773), .B(n4772), .Z(n4799) );
  XNOR U943 ( .A(n4141), .B(n4139), .Z(n4154) );
  MUX U944 ( .IN0(n252), .IN1(n3857), .SEL(n3112), .F(n3837) );
  IV U945 ( .A(n3110), .Z(n252) );
  MUX U946 ( .IN0(n922), .IN1(n920), .SEL(n921), .F(n852) );
  MUX U947 ( .IN0(n999), .IN1(n997), .SEL(n998), .F(n930) );
  MUX U948 ( .IN0(n253), .IN1(n5125), .SEL(e_input[31]), .F(n1118) );
  IV U949 ( .A(e_input[19]), .Z(n253) );
  MUX U950 ( .IN0(n254), .IN1(n1405), .SEL(n1406), .F(n1314) );
  IV U951 ( .A(n1407), .Z(n254) );
  MUX U952 ( .IN0(n255), .IN1(n3822), .SEL(e_input[31]), .F(n1623) );
  IV U953 ( .A(e_input[13]), .Z(n255) );
  MUX U954 ( .IN0(n1647), .IN1(n1645), .SEL(n1646), .F(n1547) );
  MUX U955 ( .IN0(n1837), .IN1(n1835), .SEL(n1836), .F(n1718) );
  MUX U956 ( .IN0(n256), .IN1(n2116), .SEL(n2117), .F(n2008) );
  IV U957 ( .A(n2118), .Z(n256) );
  MUX U958 ( .IN0(n2349), .IN1(n2347), .SEL(n2348), .F(n2227) );
  MUX U959 ( .IN0(n2930), .IN1(n2928), .SEL(n2929), .F(n2790) );
  XNOR U960 ( .A(n2982), .B(n2981), .Z(n4958) );
  MUX U961 ( .IN0(n257), .IN1(n3024), .SEL(n3025), .F(n2896) );
  IV U962 ( .A(n3026), .Z(n257) );
  XOR U963 ( .A(n953), .B(n891), .Z(n888) );
  MUX U964 ( .IN0(n258), .IN1(n1051), .SEL(n1052), .F(n979) );
  IV U965 ( .A(n1053), .Z(n258) );
  ANDN U966 ( .A(n1115), .B(n1114), .Z(n1042) );
  XNOR U967 ( .A(n1220), .B(n1219), .Z(n1297) );
  MUX U968 ( .IN0(n1277), .IN1(n259), .SEL(n1278), .F(n1200) );
  IV U969 ( .A(n1279), .Z(n259) );
  XNOR U970 ( .A(n1590), .B(n1589), .Z(n1681) );
  XNOR U971 ( .A(n1574), .B(n1573), .Z(n1663) );
  MUX U972 ( .IN0(n260), .IN1(n1761), .SEL(n1762), .F(n1660) );
  IV U973 ( .A(n1763), .Z(n260) );
  MUX U974 ( .IN0(n261), .IN1(n1779), .SEL(n1780), .F(n1678) );
  IV U975 ( .A(n1781), .Z(n261) );
  XNOR U976 ( .A(n1694), .B(n1693), .Z(n1790) );
  XNOR U977 ( .A(n1877), .B(n1876), .Z(n1979) );
  MUX U978 ( .IN0(n262), .IN1(n2219), .SEL(n2220), .F(n2100) );
  IV U979 ( .A(n2221), .Z(n262) );
  XNOR U980 ( .A(n2147), .B(n2157), .Z(n2263) );
  XNOR U981 ( .A(n2164), .B(n2163), .Z(n2273) );
  XNOR U982 ( .A(n2188), .B(n2187), .Z(n2303) );
  XNOR U983 ( .A(n2211), .B(n2210), .Z(n2326) );
  MUX U984 ( .IN0(n263), .IN1(n2445), .SEL(n2446), .F(n2323) );
  IV U985 ( .A(n2447), .Z(n263) );
  XNOR U986 ( .A(n2520), .B(n2519), .Z(n2639) );
  XNOR U987 ( .A(n2512), .B(n2511), .Z(n2631) );
  XNOR U988 ( .A(n2578), .B(n2577), .Z(n2705) );
  XNOR U989 ( .A(n2687), .B(n2686), .Z(n2814) );
  XNOR U990 ( .A(n2726), .B(n2725), .Z(n2853) );
  XNOR U991 ( .A(n2734), .B(n2733), .Z(n2861) );
  MUX U992 ( .IN0(n580), .IN1(n578), .SEL(n579), .F(n548) );
  NAND U993 ( .A(n691), .B(n690), .Z(n684) );
  XNOR U994 ( .A(n653), .B(n652), .Z(n692) );
  MUX U995 ( .IN0(n264), .IN1(n779), .SEL(n780), .F(n723) );
  IV U996 ( .A(n781), .Z(n264) );
  AND U997 ( .A(n1324), .B(n1326), .Z(n1240) );
  MUX U998 ( .IN0(n265), .IN1(n1358), .SEL(n1359), .F(n1267) );
  IV U999 ( .A(n1360), .Z(n265) );
  MUX U1000 ( .IN0(n266), .IN1(n1861), .SEL(n1862), .F(n1753) );
  IV U1001 ( .A(n1863), .Z(n266) );
  AND U1002 ( .A(n1911), .B(n1913), .Z(n1805) );
  MUX U1003 ( .IN0(n267), .IN1(n2315), .SEL(n2316), .F(n2195) );
  IV U1004 ( .A(n2317), .Z(n267) );
  XNOR U1005 ( .A(n2296), .B(n2295), .Z(n2293) );
  ANDN U1006 ( .A(n2487), .B(n2488), .Z(n2365) );
  MUX U1007 ( .IN0(n2677), .IN1(n2800), .SEL(n2679), .F(n2544) );
  MUX U1008 ( .IN0(n2828), .IN1(n361), .SEL(n2827), .F(n268) );
  IV U1009 ( .A(n268), .Z(n2694) );
  MUX U1010 ( .IN0(n269), .IN1(n2797), .SEL(n2798), .F(n2674) );
  IV U1011 ( .A(n2799), .Z(n269) );
  ANDN U1012 ( .A(n622), .B(n592), .Z(n581) );
  MUX U1013 ( .IN0(n824), .IN1(n826), .SEL(n825), .F(n270) );
  IV U1014 ( .A(n270), .Z(n769) );
  AND U1015 ( .A(n881), .B(n883), .Z(n818) );
  XOR U1016 ( .A(n833), .B(n830), .Z(n884) );
  NANDN U1017 ( .B(n941), .A(n942), .Z(n873) );
  XNOR U1018 ( .A(n1618), .B(n1619), .Z(n1638) );
  MUX U1019 ( .IN0(n271), .IN1(n2405), .SEL(n2406), .F(n2285) );
  IV U1020 ( .A(n2407), .Z(n271) );
  MUX U1021 ( .IN0(n2921), .IN1(n2919), .SEL(n2920), .F(n272) );
  IV U1022 ( .A(n272), .Z(n2781) );
  MUX U1023 ( .IN0(n518), .IN1(n516), .SEL(n517), .F(n273) );
  IV U1024 ( .A(n273), .Z(n495) );
  NANDN U1025 ( .B(n522), .A(n523), .Z(n479) );
  XOR U1026 ( .A(n1111), .B(n1110), .Z(n1091) );
  XOR U1027 ( .A(n1340), .B(n1339), .Z(n1424) );
  XOR U1028 ( .A(n1953), .B(n1950), .Z(n2027) );
  AND U1029 ( .A(n507), .B(n509), .Z(n482) );
  MUX U1030 ( .IN0(n2876), .IN1(\_MxM/Y0[1] ), .SEL(n2877), .F(n2744) );
  XNOR U1031 ( .A(n553), .B(n557), .Z(n555) );
  XNOR U1032 ( .A(n665), .B(n669), .Z(n667) );
  XNOR U1033 ( .A(n812), .B(n816), .Z(n814) );
  XNOR U1034 ( .A(n1010), .B(n1014), .Z(n1012) );
  XNOR U1035 ( .A(n1243), .B(n1247), .Z(n1245) );
  XNOR U1036 ( .A(n1515), .B(n1519), .Z(n1517) );
  XNOR U1037 ( .A(n1808), .B(n1812), .Z(n1810) );
  XNOR U1038 ( .A(n2129), .B(n2133), .Z(n2131) );
  MUX U1039 ( .IN0(n274), .IN1(n4150), .SEL(n3733), .F(n4129) );
  IV U1040 ( .A(n3732), .Z(n274) );
  MUX U1041 ( .IN0(n3614), .IN1(n3612), .SEL(n3613), .F(n3566) );
  MUX U1042 ( .IN0(n4101), .IN1(n4099), .SEL(n4100), .F(n4078) );
  MUX U1043 ( .IN0(n4547), .IN1(n4089), .SEL(n4090), .F(n4530) );
  MUX U1044 ( .IN0(n275), .IN1(n3536), .SEL(n3537), .F(n3492) );
  IV U1045 ( .A(n3538), .Z(n275) );
  MUX U1046 ( .IN0(n276), .IN1(n4066), .SEL(n3556), .F(n4045) );
  IV U1047 ( .A(n3554), .Z(n276) );
  MUX U1048 ( .IN0(n3432), .IN1(n3430), .SEL(n3431), .F(n3384) );
  MUX U1049 ( .IN0(n4017), .IN1(n4015), .SEL(n4016), .F(n3994) );
  MUX U1050 ( .IN0(n3459), .IN1(n3457), .SEL(n3458), .F(n3411) );
  MUX U1051 ( .IN0(n4479), .IN1(n4005), .SEL(n4006), .F(n4462) );
  MUX U1052 ( .IN0(n3828), .IN1(n4312), .SEL(n3829), .F(n277) );
  IV U1053 ( .A(n277), .Z(n4290) );
  MUX U1054 ( .IN0(n4670), .IN1(n4270), .SEL(n4272), .F(n4655) );
  MUX U1055 ( .IN0(n4265), .IN1(n4263), .SEL(n4264), .F(n4243) );
  MUX U1056 ( .IN0(n278), .IN1(n3354), .SEL(n3355), .F(n3310) );
  IV U1057 ( .A(n3356), .Z(n278) );
  MUX U1058 ( .IN0(n279), .IN1(n3982), .SEL(n3374), .F(n3961) );
  IV U1059 ( .A(n3372), .Z(n279) );
  MUX U1060 ( .IN0(n4888), .IN1(n4886), .SEL(n4887), .F(n4864) );
  MUX U1061 ( .IN0(n5027), .IN1(n4893), .SEL(n4895), .F(n5013) );
  MUX U1062 ( .IN0(n3253), .IN1(n3251), .SEL(n3252), .F(n3208) );
  MUX U1063 ( .IN0(n3933), .IN1(n3931), .SEL(n3932), .F(n3910) );
  MUX U1064 ( .IN0(n3277), .IN1(n3275), .SEL(n3276), .F(n3233) );
  MUX U1065 ( .IN0(n4412), .IN1(n3921), .SEL(n3922), .F(n4396) );
  MUX U1066 ( .IN0(g_input[1]), .IN1(n5234), .SEL(g_input[31]), .F(n280) );
  IV U1067 ( .A(n280), .Z(n3802) );
  MUX U1068 ( .IN0(n281), .IN1(n5153), .SEL(n5154), .F(n5142) );
  IV U1069 ( .A(n5155), .Z(n281) );
  MUX U1070 ( .IN0(n4618), .IN1(n4190), .SEL(n4192), .F(n4608) );
  MUX U1071 ( .IN0(n4185), .IN1(n4183), .SEL(n4184), .F(n4159) );
  MUX U1072 ( .IN0(n282), .IN1(n3180), .SEL(n3181), .F(n3137) );
  IV U1073 ( .A(n3182), .Z(n282) );
  MUX U1074 ( .IN0(n283), .IN1(n3899), .SEL(n3199), .F(n3878) );
  IV U1075 ( .A(n3197), .Z(n283) );
  XNOR U1076 ( .A(n5140), .B(g_input[7]), .Z(n5141) );
  XNOR U1077 ( .A(n5008), .B(g_input[11]), .Z(n5009) );
  XNOR U1078 ( .A(n4960), .B(g_input[15]), .Z(n4961) );
  XNOR U1079 ( .A(n4539), .B(g_input[19]), .Z(n4540) );
  MUX U1080 ( .IN0(g_input[2]), .IN1(n5227), .SEL(g_input[31]), .F(n284) );
  IV U1081 ( .A(n284), .Z(n3799) );
  MUX U1082 ( .IN0(n4806), .IN1(n4804), .SEL(n4805), .F(n4773) );
  MUX U1083 ( .IN0(n4977), .IN1(n4811), .SEL(n4813), .F(n4965) );
  MUX U1084 ( .IN0(n3083), .IN1(n3081), .SEL(n3082), .F(n3042) );
  MUX U1085 ( .IN0(n3105), .IN1(n3103), .SEL(n3104), .F(n3034) );
  XNOR U1086 ( .A(n4437), .B(g_input[25]), .Z(n4438) );
  MUX U1087 ( .IN0(n285), .IN1(n3809), .SEL(e_input[31]), .F(n2039) );
  IV U1088 ( .A(e_input[9]), .Z(n285) );
  MUX U1089 ( .IN0(n2559), .IN1(n2561), .SEL(n2560), .F(n2434) );
  MUX U1090 ( .IN0(n2778), .IN1(n2780), .SEL(n2779), .F(n2648) );
  MUX U1091 ( .IN0(g_input[4]), .IN1(n5186), .SEL(g_input[31]), .F(n2737) );
  MUX U1092 ( .IN0(n3003), .IN1(n286), .SEL(n3004), .F(n2863) );
  IV U1093 ( .A(n3005), .Z(n286) );
  MUX U1094 ( .IN0(g_input[9]), .IN1(n5037), .SEL(g_input[31]), .F(n287) );
  IV U1095 ( .A(n287), .Z(n2240) );
  MUX U1096 ( .IN0(n2971), .IN1(n2973), .SEL(n2972), .F(n2831) );
  MUX U1097 ( .IN0(e_input[1]), .IN1(n4766), .SEL(e_input[31]), .F(n288) );
  IV U1098 ( .A(n288), .Z(n4339) );
  XNOR U1099 ( .A(n3727), .B(n3725), .Z(n3741) );
  MUX U1100 ( .IN0(n1063), .IN1(n1061), .SEL(n1062), .F(n989) );
  MUX U1101 ( .IN0(n289), .IN1(n1230), .SEL(n1231), .F(n1149) );
  IV U1102 ( .A(n1232), .Z(n289) );
  MUX U1103 ( .IN0(n1262), .IN1(n1260), .SEL(n1261), .F(n1178) );
  MUX U1104 ( .IN0(n1286), .IN1(n1288), .SEL(n1287), .F(n290) );
  MUX U1105 ( .IN0(n1688), .IN1(n1686), .SEL(n1687), .F(n1590) );
  MUX U1106 ( .IN0(n2272), .IN1(n2270), .SEL(n2271), .F(n2147) );
  MUX U1107 ( .IN0(n2792), .IN1(n2790), .SEL(n2791), .F(n2656) );
  MUX U1108 ( .IN0(n4342), .IN1(n3855), .SEL(n3856), .F(n291) );
  IV U1109 ( .A(n291), .Z(n2949) );
  XNOR U1110 ( .A(n4936), .B(n4933), .Z(n4934) );
  XNOR U1111 ( .A(n5239), .B(e_input[30]), .Z(n5237) );
  MUX U1112 ( .IN0(n292), .IN1(n842), .SEL(n843), .F(n779) );
  IV U1113 ( .A(n844), .Z(n292) );
  XNOR U1114 ( .A(n1304), .B(n1303), .Z(n1392) );
  MUX U1115 ( .IN0(n293), .IN1(n1468), .SEL(n1469), .F(n1368) );
  IV U1116 ( .A(n1470), .Z(n293) );
  MUX U1117 ( .IN0(n294), .IN1(n1582), .SEL(n1583), .F(n1486) );
  IV U1118 ( .A(n1584), .Z(n294) );
  XNOR U1119 ( .A(n1502), .B(n1501), .Z(n1593) );
  XNOR U1120 ( .A(n1547), .B(n1546), .Z(n1640) );
  XNOR U1121 ( .A(n1670), .B(n1669), .Z(n1764) );
  XNOR U1122 ( .A(n1835), .B(n1834), .Z(n1936) );
  XNOR U1123 ( .A(n2000), .B(n1999), .Z(n2103) );
  XNOR U1124 ( .A(n2008), .B(n2007), .Z(n2111) );
  XNOR U1125 ( .A(n1961), .B(n1960), .Z(n2064) );
  MUX U1126 ( .IN0(n295), .IN1(n2084), .SEL(n2085), .F(n1976) );
  IV U1127 ( .A(n2086), .Z(n295) );
  XNOR U1128 ( .A(n2331), .B(n2330), .Z(n2448) );
  MUX U1129 ( .IN0(n296), .IN1(n2461), .SEL(n2462), .F(n2339) );
  IV U1130 ( .A(n2463), .Z(n296) );
  XNOR U1131 ( .A(n2278), .B(n2277), .Z(n2393) );
  MUX U1132 ( .IN0(n297), .IN1(n2380), .SEL(n2381), .F(n2260) );
  IV U1133 ( .A(n2382), .Z(n297) );
  XNOR U1134 ( .A(n2594), .B(n2593), .Z(n2721) );
  XNOR U1135 ( .A(n2602), .B(n2601), .Z(n2729) );
  XNOR U1136 ( .A(n2555), .B(n2554), .Z(n2682) );
  XNOR U1137 ( .A(n2710), .B(n2709), .Z(n2837) );
  XNOR U1138 ( .A(n2644), .B(n2643), .Z(n2769) );
  XNOR U1139 ( .A(n2636), .B(n2635), .Z(n2761) );
  MUX U1140 ( .IN0(n2992), .IN1(n2990), .SEL(n2991), .F(n298) );
  IV U1141 ( .A(n298), .Z(n2850) );
  MUX U1142 ( .IN0(n299), .IN1(n2974), .SEL(n2975), .F(n2834) );
  IV U1143 ( .A(n2976), .Z(n299) );
  MUX U1144 ( .IN0(n300), .IN1(n2896), .SEL(n2897), .F(n2758) );
  IV U1145 ( .A(n2898), .Z(n300) );
  MUX U1146 ( .IN0(n2946), .IN1(n301), .SEL(n2947), .F(n2810) );
  IV U1147 ( .A(n2948), .Z(n301) );
  MUX U1148 ( .IN0(n571), .IN1(n569), .SEL(n570), .F(n536) );
  MUX U1149 ( .IN0(n302), .IN1(n640), .SEL(n641), .F(n604) );
  IV U1150 ( .A(n642), .Z(n302) );
  XNOR U1151 ( .A(n697), .B(n696), .Z(n734) );
  XNOR U1152 ( .A(n731), .B(n729), .Z(n782) );
  AND U1153 ( .A(n833), .B(n834), .Z(n763) );
  MUX U1154 ( .IN0(n303), .IN1(n966), .SEL(n967), .F(n897) );
  IV U1155 ( .A(n968), .Z(n303) );
  XOR U1156 ( .A(n1039), .B(n1043), .Z(n1112) );
  XNOR U1157 ( .A(n1525), .B(n1524), .Z(n1523) );
  MUX U1158 ( .IN0(n304), .IN1(n1652), .SEL(n1653), .F(n1554) );
  IV U1159 ( .A(n1654), .Z(n304) );
  AND U1160 ( .A(n1704), .B(n1706), .Z(n1608) );
  MUX U1161 ( .IN0(n305), .IN1(n1716), .SEL(n1715), .F(n1619) );
  IV U1162 ( .A(n1714), .Z(n305) );
  AND U1163 ( .A(n2126), .B(n2128), .Z(n2018) );
  MUX U1164 ( .IN0(n306), .IN1(n2195), .SEL(n2196), .F(n2076) );
  IV U1165 ( .A(n2197), .Z(n306) );
  MUX U1166 ( .IN0(n307), .IN1(n2694), .SEL(n2695), .F(n2562) );
  IV U1167 ( .A(n2696), .Z(n307) );
  MUX U1168 ( .IN0(n545), .IN1(n547), .SEL(n546), .F(n513) );
  AND U1169 ( .A(n768), .B(n769), .Z(n765) );
  MUX U1170 ( .IN0(n308), .IN1(n1734), .SEL(n1735), .F(n1633) );
  IV U1171 ( .A(n1736), .Z(n308) );
  XOR U1172 ( .A(n2174), .B(n2060), .Z(n2061) );
  XNOR U1173 ( .A(n2421), .B(n2419), .Z(n2530) );
  NANDN U1174 ( .B(n520), .A(n519), .Z(n491) );
  XNOR U1175 ( .A(n522), .B(n527), .Z(n523) );
  XNOR U1176 ( .A(n623), .B(n628), .Z(n624) );
  XNOR U1177 ( .A(n751), .B(n716), .Z(n752) );
  XNOR U1178 ( .A(n941), .B(n946), .Z(n942) );
  XOR U1179 ( .A(n1189), .B(n1188), .Z(n1169) );
  MUX U1180 ( .IN0(\_MxM/Y0[2] ), .IN1(n2744), .SEL(n2745), .F(n2612) );
  XOR U1181 ( .A(n1342), .B(n1341), .Z(n1421) );
  XOR U1182 ( .A(n1952), .B(n1951), .Z(n2024) );
  XOR U1183 ( .A(n2287), .B(n2286), .Z(n2371) );
  XNOR U1184 ( .A(n2617), .B(n2496), .Z(n2497) );
  XOR U1185 ( .A(n2783), .B(n2782), .Z(n2887) );
  XNOR U1186 ( .A(n584), .B(n588), .Z(n586) );
  XNOR U1187 ( .A(n709), .B(n713), .Z(n711) );
  XNOR U1188 ( .A(n875), .B(n879), .Z(n877) );
  XNOR U1189 ( .A(n1084), .B(n1088), .Z(n1086) );
  XNOR U1190 ( .A(n1327), .B(n1331), .Z(n1329) );
  XNOR U1191 ( .A(n1611), .B(n1615), .Z(n1613) );
  XNOR U1192 ( .A(n1914), .B(n1918), .Z(n1916) );
  XNOR U1193 ( .A(n2248), .B(n2252), .Z(n2250) );
  XOR U1194 ( .A(n467), .B(n468), .Z(n365) );
  MUX U1195 ( .IN0(n3704), .IN1(n3702), .SEL(n3703), .F(n3658) );
  MUX U1196 ( .IN0(n3687), .IN1(n3685), .SEL(n3686), .F(n3639) );
  MUX U1197 ( .IN0(n309), .IN1(n3628), .SEL(n3629), .F(n3582) );
  IV U1198 ( .A(n3630), .Z(n309) );
  MUX U1199 ( .IN0(n3524), .IN1(n3522), .SEL(n3523), .F(n3476) );
  MUX U1200 ( .IN0(n310), .IN1(n4087), .SEL(n3602), .F(n4066) );
  IV U1201 ( .A(n3600), .Z(n310) );
  MUX U1202 ( .IN0(n4530), .IN1(n4068), .SEL(n4069), .F(n4513) );
  MUX U1203 ( .IN0(n4038), .IN1(n4036), .SEL(n4037), .F(n4015) );
  MUX U1204 ( .IN0(n3505), .IN1(n3503), .SEL(n3504), .F(n3457) );
  MUX U1205 ( .IN0(n311), .IN1(n3446), .SEL(n3447), .F(n3400) );
  IV U1206 ( .A(n3448), .Z(n311) );
  MUX U1207 ( .IN0(n3342), .IN1(n3340), .SEL(n3341), .F(n3294) );
  MUX U1208 ( .IN0(n312), .IN1(n4003), .SEL(n3420), .F(n3982) );
  IV U1209 ( .A(n3418), .Z(n312) );
  MUX U1210 ( .IN0(n4462), .IN1(n3984), .SEL(n3985), .F(n4445) );
  MUX U1211 ( .IN0(n4912), .IN1(n4910), .SEL(n4911), .F(n4886) );
  MUX U1212 ( .IN0(n5044), .IN1(n4917), .SEL(n4919), .F(n5027) );
  MUX U1213 ( .IN0(n3954), .IN1(n3952), .SEL(n3953), .F(n3931) );
  MUX U1214 ( .IN0(n3323), .IN1(n3321), .SEL(n3322), .F(n3275) );
  MUX U1215 ( .IN0(n4655), .IN1(n4250), .SEL(n4252), .F(n4640) );
  MUX U1216 ( .IN0(n4245), .IN1(n4243), .SEL(n4244), .F(n4223) );
  MUX U1217 ( .IN0(n5112), .IN1(n4956), .SEL(n4957), .F(n313) );
  IV U1218 ( .A(n313), .Z(n5098) );
  MUX U1219 ( .IN0(n3788), .IN1(n3739), .SEL(n3740), .F(n314) );
  IV U1220 ( .A(n314), .Z(n3774) );
  MUX U1221 ( .IN0(n315), .IN1(n3771), .SEL(n3772), .F(n3757) );
  IV U1222 ( .A(n3773), .Z(n315) );
  MUX U1223 ( .IN0(n316), .IN1(n3265), .SEL(n3266), .F(n3222) );
  IV U1224 ( .A(n3267), .Z(n316) );
  MUX U1225 ( .IN0(n5195), .IN1(n5136), .SEL(n5137), .F(n317) );
  IV U1226 ( .A(n317), .Z(n5179) );
  MUX U1227 ( .IN0(n3168), .IN1(n3166), .SEL(n3167), .F(n3121) );
  MUX U1228 ( .IN0(n318), .IN1(n3919), .SEL(n3242), .F(n3899) );
  IV U1229 ( .A(n3240), .Z(n318) );
  MUX U1230 ( .IN0(n4396), .IN1(n3901), .SEL(n3902), .F(n4379) );
  MUX U1231 ( .IN0(n5223), .IN1(n5225), .SEL(n5224), .F(n5219) );
  MUX U1232 ( .IN0(n4826), .IN1(n4824), .SEL(n4825), .F(n4804) );
  MUX U1233 ( .IN0(n4989), .IN1(n4831), .SEL(n4833), .F(n4977) );
  MUX U1234 ( .IN0(n319), .IN1(n3743), .SEL(n3744), .F(n3721) );
  IV U1235 ( .A(n3745), .Z(n319) );
  MUX U1236 ( .IN0(n3871), .IN1(n3869), .SEL(n3870), .F(n3845) );
  MUX U1237 ( .IN0(n3150), .IN1(n3148), .SEL(n3149), .F(n3103) );
  XNOR U1238 ( .A(n5167), .B(g_input[5]), .Z(n5168) );
  XNOR U1239 ( .A(n5036), .B(g_input[9]), .Z(n5037) );
  MUX U1240 ( .IN0(n320), .IN1(n4950), .SEL(e_input[31]), .F(n4942) );
  IV U1241 ( .A(e_input[21]), .Z(n320) );
  XNOR U1242 ( .A(n4984), .B(g_input[13]), .Z(n4985) );
  XNOR U1243 ( .A(n4573), .B(g_input[17]), .Z(n4574) );
  XNOR U1244 ( .A(n4505), .B(g_input[21]), .Z(n4506) );
  AND U1245 ( .A(n5235), .B(g_input[0]), .Z(n3013) );
  MUX U1246 ( .IN0(n4161), .IN1(n4159), .SEL(n4160), .F(n4141) );
  MUX U1247 ( .IN0(n4608), .IN1(n4170), .SEL(n4172), .F(n4598) );
  MUX U1248 ( .IN0(n321), .IN1(n5214), .SEL(e_input[31]), .F(n5201) );
  IV U1249 ( .A(e_input[25]), .Z(n321) );
  MUX U1250 ( .IN0(n322), .IN1(n5232), .SEL(e_input[31]), .F(n5222) );
  IV U1251 ( .A(e_input[29]), .Z(n322) );
  XNOR U1252 ( .A(n4405), .B(g_input[27]), .Z(n4406) );
  MUX U1253 ( .IN0(g_input[3]), .IN1(n5218), .SEL(g_input[31]), .F(n2869) );
  MUX U1254 ( .IN0(n2987), .IN1(n2989), .SEL(n2988), .F(n2847) );
  MUX U1255 ( .IN0(n2963), .IN1(n2965), .SEL(n2964), .F(n2823) );
  MUX U1256 ( .IN0(e_input[20]), .IN1(n323), .SEL(e_input[31]), .F(n1021) );
  IV U1257 ( .A(n4949), .Z(n323) );
  MUX U1258 ( .IN0(e_input[16]), .IN1(n324), .SEL(e_input[31]), .F(n1383) );
  IV U1259 ( .A(n5129), .Z(n324) );
  MUX U1260 ( .IN0(e_input[8]), .IN1(n325), .SEL(e_input[31]), .F(n2158) );
  IV U1261 ( .A(n3808), .Z(n325) );
  MUX U1262 ( .IN0(e_input[12]), .IN1(n326), .SEL(e_input[31]), .F(n1729) );
  IV U1263 ( .A(n3821), .Z(n326) );
  MUX U1264 ( .IN0(e_input[4]), .IN1(n327), .SEL(e_input[31]), .F(n2667) );
  IV U1265 ( .A(n4327), .Z(n327) );
  XNOR U1266 ( .A(n4315), .B(n4312), .Z(n4313) );
  MUX U1267 ( .IN0(n328), .IN1(n3093), .SEL(n3094), .F(n3024) );
  IV U1268 ( .A(n3095), .Z(n328) );
  MUX U1269 ( .IN0(n329), .IN1(n5208), .SEL(e_input[31]), .F(n636) );
  IV U1270 ( .A(e_input[27]), .Z(n329) );
  MUX U1271 ( .IN0(e_input[26]), .IN1(n330), .SEL(e_input[31]), .F(n677) );
  IV U1272 ( .A(n5209), .Z(n330) );
  MUX U1273 ( .IN0(e_input[24]), .IN1(n331), .SEL(e_input[31]), .F(n784) );
  IV U1274 ( .A(n5213), .Z(n331) );
  MUX U1275 ( .IN0(e_input[28]), .IN1(n332), .SEL(e_input[31]), .F(n609) );
  IV U1276 ( .A(n5231), .Z(n332) );
  MUX U1277 ( .IN0(n1102), .IN1(n1100), .SEL(n1101), .F(n1027) );
  MUX U1278 ( .IN0(n333), .IN1(n1149), .SEL(n1150), .F(n1071) );
  IV U1279 ( .A(n1151), .Z(n333) );
  MUX U1280 ( .IN0(n1143), .IN1(n1141), .SEL(n1142), .F(n1061) );
  MUX U1281 ( .IN0(e_input[18]), .IN1(n334), .SEL(e_input[31]), .F(n1199) );
  IV U1282 ( .A(n5124), .Z(n334) );
  MUX U1283 ( .IN0(n335), .IN1(n5130), .SEL(e_input[31]), .F(n1283) );
  IV U1284 ( .A(e_input[17]), .Z(n335) );
  MUX U1285 ( .IN0(n1480), .IN1(n1478), .SEL(n1479), .F(n1372) );
  MUX U1286 ( .IN0(n1453), .IN1(n1451), .SEL(n1452), .F(n1349) );
  MUX U1287 ( .IN0(n1496), .IN1(n1494), .SEL(n1495), .F(n1397) );
  MUX U1288 ( .IN0(n336), .IN1(n1502), .SEL(n1503), .F(n1405) );
  IV U1289 ( .A(n1504), .Z(n336) );
  MUX U1290 ( .IN0(n337), .IN1(n3804), .SEL(e_input[31]), .F(n1822) );
  IV U1291 ( .A(e_input[11]), .Z(n337) );
  MUX U1292 ( .IN0(e_input[10]), .IN1(n338), .SEL(e_input[31]), .F(n1928) );
  IV U1293 ( .A(n3803), .Z(n338) );
  MUX U1294 ( .IN0(n2052), .IN1(n2050), .SEL(n2051), .F(n1943) );
  MUX U1295 ( .IN0(e_input[6]), .IN1(n339), .SEL(e_input[31]), .F(n2418) );
  IV U1296 ( .A(n4332), .Z(n339) );
  MUX U1297 ( .IN0(n340), .IN1(n4328), .SEL(e_input[31]), .F(n2534) );
  IV U1298 ( .A(e_input[5]), .Z(n340) );
  MUX U1299 ( .IN0(n341), .IN1(n4762), .SEL(e_input[31]), .F(n2807) );
  IV U1300 ( .A(e_input[3]), .Z(n341) );
  MUX U1301 ( .IN0(e_input[2]), .IN1(n342), .SEL(e_input[31]), .F(n2945) );
  IV U1302 ( .A(n4761), .Z(n342) );
  MUX U1303 ( .IN0(n3837), .IN1(n343), .SEL(n3074), .F(n2946) );
  IV U1304 ( .A(n3073), .Z(n343) );
  MUX U1305 ( .IN0(e_input[22]), .IN1(n344), .SEL(e_input[31]), .F(n893) );
  IV U1306 ( .A(n4955), .Z(n344) );
  MUX U1307 ( .IN0(n345), .IN1(n4954), .SEL(e_input[31]), .F(n823) );
  IV U1308 ( .A(e_input[23]), .Z(n345) );
  MUX U1309 ( .IN0(n346), .IN1(n910), .SEL(n911), .F(n842) );
  IV U1310 ( .A(n912), .Z(n346) );
  MUX U1311 ( .IN0(n347), .IN1(n1210), .SEL(n1211), .F(n1131) );
  IV U1312 ( .A(n1212), .Z(n347) );
  MUX U1313 ( .IN0(n1628), .IN1(n1626), .SEL(n1627), .F(n348) );
  MUX U1314 ( .IN0(e_input[14]), .IN1(n349), .SEL(e_input[31]), .F(n1532) );
  IV U1315 ( .A(n3826), .Z(n349) );
  MUX U1316 ( .IN0(n350), .IN1(n1564), .SEL(n1565), .F(n1468) );
  IV U1317 ( .A(n1566), .Z(n350) );
  XNOR U1318 ( .A(n1787), .B(n1786), .Z(n1888) );
  XNOR U1319 ( .A(n1795), .B(n1794), .Z(n1896) );
  XNOR U1320 ( .A(n1746), .B(n1745), .Z(n1849) );
  XNOR U1321 ( .A(n1771), .B(n1770), .Z(n1872) );
  MUX U1322 ( .IN0(n351), .IN1(n1976), .SEL(n1977), .F(n1869) );
  IV U1323 ( .A(n1978), .Z(n351) );
  MUX U1324 ( .IN0(n352), .IN1(n1992), .SEL(n1993), .F(n1885) );
  IV U1325 ( .A(n1994), .Z(n352) );
  MUX U1326 ( .IN0(n1932), .IN1(n2036), .SEL(n1934), .F(n1824) );
  XNOR U1327 ( .A(n2092), .B(n2091), .Z(n2206) );
  XNOR U1328 ( .A(n2069), .B(n2068), .Z(n2183) );
  XNOR U1329 ( .A(n2108), .B(n2107), .Z(n2222) );
  XNOR U1330 ( .A(n2116), .B(n2115), .Z(n2230) );
  MUX U1331 ( .IN0(n353), .IN1(n2143), .SEL(n2144), .F(n2033) );
  IV U1332 ( .A(n2145), .Z(n353) );
  MUX U1333 ( .IN0(n354), .IN1(n4333), .SEL(e_input[31]), .F(n2292) );
  IV U1334 ( .A(e_input[7]), .Z(n354) );
  XNOR U1335 ( .A(n2477), .B(n2476), .Z(n2597) );
  XNOR U1336 ( .A(n2469), .B(n2468), .Z(n2589) );
  XNOR U1337 ( .A(n2430), .B(n2429), .Z(n2550) );
  XNOR U1338 ( .A(n2453), .B(n2452), .Z(n2573) );
  XNOR U1339 ( .A(n2390), .B(n2389), .Z(n2507) );
  XNOR U1340 ( .A(n2398), .B(n2397), .Z(n2515) );
  MUX U1341 ( .IN0(n355), .IN1(n2628), .SEL(n2629), .F(n2504) );
  IV U1342 ( .A(n2630), .Z(n355) );
  MUX U1343 ( .IN0(n356), .IN1(n2718), .SEL(n2719), .F(n2586) );
  IV U1344 ( .A(n2720), .Z(n356) );
  MUX U1345 ( .IN0(n357), .IN1(n2702), .SEL(n2703), .F(n2570) );
  IV U1346 ( .A(n2704), .Z(n357) );
  XNOR U1347 ( .A(n2866), .B(n2865), .Z(n3001) );
  XNOR U1348 ( .A(n2858), .B(n2857), .Z(n2993) );
  XNOR U1349 ( .A(n2819), .B(n2818), .Z(n2954) );
  XNOR U1350 ( .A(n2842), .B(n2841), .Z(n2977) );
  XNOR U1351 ( .A(n2766), .B(n2765), .Z(n2899) );
  XNOR U1352 ( .A(n2774), .B(n2773), .Z(n2907) );
  MUX U1353 ( .IN0(n2949), .IN1(n4336), .SEL(n2951), .F(n2809) );
  XNOR U1354 ( .A(n2790), .B(n2789), .Z(n2923) );
  MUX U1355 ( .IN0(e_input[30]), .IN1(n358), .SEL(e_input[31]), .F(n543) );
  IV U1356 ( .A(n5237), .Z(n358) );
  XNOR U1357 ( .A(n686), .B(n690), .Z(n726) );
  NAND U1358 ( .A(n891), .B(n890), .Z(n885) );
  MUX U1359 ( .IN0(n894), .IN1(n896), .SEL(n895), .F(n824) );
  XNOR U1360 ( .A(n739), .B(n738), .Z(n793) );
  NAND U1361 ( .A(n1042), .B(n1043), .Z(n1037) );
  MUX U1362 ( .IN0(n359), .IN1(n1458), .SEL(n1459), .F(n1358) );
  IV U1363 ( .A(n1460), .Z(n359) );
  MUX U1364 ( .IN0(n360), .IN1(n3827), .SEL(e_input[31]), .F(n1431) );
  IV U1365 ( .A(e_input[15]), .Z(n360) );
  AND U1366 ( .A(n1512), .B(n1514), .Z(n1415) );
  ANDN U1367 ( .A(n1953), .B(n1954), .Z(n1845) );
  MUX U1368 ( .IN0(n2968), .IN1(n2966), .SEL(n2967), .F(n361) );
  IV U1369 ( .A(n361), .Z(n2826) );
  MUX U1370 ( .IN0(n362), .IN1(n2935), .SEL(n2936), .F(n2797) );
  IV U1371 ( .A(n2937), .Z(n362) );
  MUX U1372 ( .IN0(n538), .IN1(n536), .SEL(n537), .F(n516) );
  ANDN U1373 ( .A(n548), .B(n549), .Z(n519) );
  MUX U1374 ( .IN0(n363), .IN1(n771), .SEL(n772), .F(n748) );
  IV U1375 ( .A(n773), .Z(n363) );
  XNOR U1376 ( .A(n1433), .B(n1432), .Z(n1426) );
  XNOR U1377 ( .A(n2299), .B(n2294), .Z(n2408) );
  MUX U1378 ( .IN0(n513), .IN1(n515), .SEL(n514), .F(n364) );
  IV U1379 ( .A(n364), .Z(n498) );
  XNOR U1380 ( .A(n582), .B(n587), .Z(n583) );
  XNOR U1381 ( .A(n707), .B(n712), .Z(n708) );
  XNOR U1382 ( .A(n873), .B(n878), .Z(n874) );
  XOR U1383 ( .A(n1036), .B(n1035), .Z(n1017) );
  XOR U1384 ( .A(n1269), .B(n1268), .Z(n1251) );
  XOR U1385 ( .A(n1535), .B(n1534), .Z(n1614) );
  XOR U1386 ( .A(n1736), .B(n1735), .Z(n1811) );
  XOR U1387 ( .A(n1844), .B(n1843), .Z(n1917) );
  XOR U1388 ( .A(n2059), .B(n2058), .Z(n2132) );
  XOR U1389 ( .A(n2173), .B(n2172), .Z(n2251) );
  XOR U1390 ( .A(n2407), .B(n2406), .Z(n2493) );
  XOR U1391 ( .A(n2529), .B(n2528), .Z(n2617) );
  XOR U1392 ( .A(n2653), .B(n2652), .Z(n2747) );
  AND U1393 ( .A(\_MxM/Y0[0] ), .B(n2751), .Z(n2876) );
  XNOR U1394 ( .A(n524), .B(n528), .Z(n526) );
  XNOR U1395 ( .A(n625), .B(n629), .Z(n627) );
  XNOR U1396 ( .A(n753), .B(n756), .Z(n755) );
  XNOR U1397 ( .A(n943), .B(n947), .Z(n945) );
  XNOR U1398 ( .A(n1162), .B(n1166), .Z(n1164) );
  XNOR U1399 ( .A(n1418), .B(n1422), .Z(n1420) );
  XNOR U1400 ( .A(n1707), .B(n1711), .Z(n1709) );
  XNOR U1401 ( .A(n2021), .B(n2025), .Z(n2023) );
  XNOR U1402 ( .A(n2368), .B(n2372), .Z(n2370) );
  MUX U1403 ( .IN0(n365), .IN1(n459), .SEL(n465), .F(n462) );
  NAND U1404 ( .A(n366), .B(n367), .Z(\_MxM/n341 ) );
  NAND U1405 ( .A(n368), .B(n369), .Z(n367) );
  NAND U1406 ( .A(\_MxM/Y0[0] ), .B(rst), .Z(n366) );
  NAND U1407 ( .A(n370), .B(n371), .Z(\_MxM/n340 ) );
  NAND U1408 ( .A(n372), .B(n369), .Z(n371) );
  NAND U1409 ( .A(\_MxM/Y0[1] ), .B(rst), .Z(n370) );
  NAND U1410 ( .A(n373), .B(n374), .Z(\_MxM/n339 ) );
  NAND U1411 ( .A(n375), .B(n369), .Z(n374) );
  NAND U1412 ( .A(\_MxM/Y0[2] ), .B(rst), .Z(n373) );
  NAND U1413 ( .A(n376), .B(n377), .Z(\_MxM/n338 ) );
  NAND U1414 ( .A(n378), .B(n369), .Z(n377) );
  NAND U1415 ( .A(\_MxM/Y0[3] ), .B(rst), .Z(n376) );
  NAND U1416 ( .A(n379), .B(n380), .Z(\_MxM/n337 ) );
  NAND U1417 ( .A(n381), .B(n369), .Z(n380) );
  NAND U1418 ( .A(\_MxM/Y0[4] ), .B(rst), .Z(n379) );
  NAND U1419 ( .A(n382), .B(n383), .Z(\_MxM/n336 ) );
  NAND U1420 ( .A(n384), .B(n369), .Z(n383) );
  NAND U1421 ( .A(rst), .B(\_MxM/Y0[5] ), .Z(n382) );
  NAND U1422 ( .A(n385), .B(n386), .Z(\_MxM/n335 ) );
  NAND U1423 ( .A(n387), .B(n369), .Z(n386) );
  NAND U1424 ( .A(rst), .B(\_MxM/Y0[6] ), .Z(n385) );
  NAND U1425 ( .A(n388), .B(n389), .Z(\_MxM/n334 ) );
  NAND U1426 ( .A(n390), .B(n369), .Z(n389) );
  NAND U1427 ( .A(rst), .B(\_MxM/Y0[7] ), .Z(n388) );
  NAND U1428 ( .A(n391), .B(n392), .Z(\_MxM/n333 ) );
  NAND U1429 ( .A(n393), .B(n369), .Z(n392) );
  NAND U1430 ( .A(rst), .B(\_MxM/Y0[8] ), .Z(n391) );
  NAND U1431 ( .A(n394), .B(n395), .Z(\_MxM/n332 ) );
  NAND U1432 ( .A(n396), .B(n369), .Z(n395) );
  NAND U1433 ( .A(rst), .B(\_MxM/Y0[9] ), .Z(n394) );
  NAND U1434 ( .A(n397), .B(n398), .Z(\_MxM/n331 ) );
  NAND U1435 ( .A(n399), .B(n369), .Z(n398) );
  NAND U1436 ( .A(rst), .B(\_MxM/Y0[10] ), .Z(n397) );
  NAND U1437 ( .A(n400), .B(n401), .Z(\_MxM/n330 ) );
  NAND U1438 ( .A(n402), .B(n369), .Z(n401) );
  NAND U1439 ( .A(rst), .B(\_MxM/Y0[11] ), .Z(n400) );
  NAND U1440 ( .A(n403), .B(n404), .Z(\_MxM/n329 ) );
  NAND U1441 ( .A(n405), .B(n369), .Z(n404) );
  NAND U1442 ( .A(rst), .B(\_MxM/Y0[12] ), .Z(n403) );
  NAND U1443 ( .A(n406), .B(n407), .Z(\_MxM/n328 ) );
  NAND U1444 ( .A(n408), .B(n369), .Z(n407) );
  NAND U1445 ( .A(rst), .B(\_MxM/Y0[13] ), .Z(n406) );
  NAND U1446 ( .A(n409), .B(n410), .Z(\_MxM/n327 ) );
  NAND U1447 ( .A(n411), .B(n369), .Z(n410) );
  NAND U1448 ( .A(rst), .B(\_MxM/Y0[14] ), .Z(n409) );
  NAND U1449 ( .A(n412), .B(n413), .Z(\_MxM/n326 ) );
  NAND U1450 ( .A(n414), .B(n369), .Z(n413) );
  NAND U1451 ( .A(rst), .B(\_MxM/Y0[15] ), .Z(n412) );
  NAND U1452 ( .A(n415), .B(n416), .Z(\_MxM/n325 ) );
  NAND U1453 ( .A(n417), .B(n369), .Z(n416) );
  NAND U1454 ( .A(rst), .B(\_MxM/Y0[16] ), .Z(n415) );
  NAND U1455 ( .A(n418), .B(n419), .Z(\_MxM/n324 ) );
  NAND U1456 ( .A(n420), .B(n369), .Z(n419) );
  NAND U1457 ( .A(rst), .B(\_MxM/Y0[17] ), .Z(n418) );
  NAND U1458 ( .A(n421), .B(n422), .Z(\_MxM/n323 ) );
  NAND U1459 ( .A(n423), .B(n369), .Z(n422) );
  NAND U1460 ( .A(rst), .B(\_MxM/Y0[18] ), .Z(n421) );
  NAND U1461 ( .A(n424), .B(n425), .Z(\_MxM/n322 ) );
  NAND U1462 ( .A(n426), .B(n369), .Z(n425) );
  NAND U1463 ( .A(rst), .B(\_MxM/Y0[19] ), .Z(n424) );
  NAND U1464 ( .A(n427), .B(n428), .Z(\_MxM/n321 ) );
  NAND U1465 ( .A(n429), .B(n369), .Z(n428) );
  NAND U1466 ( .A(rst), .B(\_MxM/Y0[20] ), .Z(n427) );
  NAND U1467 ( .A(n430), .B(n431), .Z(\_MxM/n320 ) );
  NAND U1468 ( .A(n432), .B(n369), .Z(n431) );
  NAND U1469 ( .A(rst), .B(\_MxM/Y0[21] ), .Z(n430) );
  NAND U1470 ( .A(n433), .B(n434), .Z(\_MxM/n319 ) );
  NAND U1471 ( .A(n435), .B(n369), .Z(n434) );
  NAND U1472 ( .A(rst), .B(\_MxM/Y0[22] ), .Z(n433) );
  NAND U1473 ( .A(n436), .B(n437), .Z(\_MxM/n318 ) );
  NAND U1474 ( .A(n438), .B(n369), .Z(n437) );
  NAND U1475 ( .A(rst), .B(\_MxM/Y0[23] ), .Z(n436) );
  NAND U1476 ( .A(n439), .B(n440), .Z(\_MxM/n317 ) );
  NAND U1477 ( .A(n441), .B(n369), .Z(n440) );
  NAND U1478 ( .A(rst), .B(\_MxM/Y0[24] ), .Z(n439) );
  NAND U1479 ( .A(n442), .B(n443), .Z(\_MxM/n316 ) );
  NAND U1480 ( .A(n444), .B(n369), .Z(n443) );
  NAND U1481 ( .A(rst), .B(\_MxM/Y0[25] ), .Z(n442) );
  NAND U1482 ( .A(n445), .B(n446), .Z(\_MxM/n315 ) );
  NAND U1483 ( .A(n447), .B(n369), .Z(n446) );
  NAND U1484 ( .A(rst), .B(\_MxM/Y0[26] ), .Z(n445) );
  NAND U1485 ( .A(n448), .B(n449), .Z(\_MxM/n314 ) );
  NAND U1486 ( .A(n450), .B(n369), .Z(n449) );
  NAND U1487 ( .A(rst), .B(\_MxM/Y0[27] ), .Z(n448) );
  NAND U1488 ( .A(n451), .B(n452), .Z(\_MxM/n313 ) );
  NAND U1489 ( .A(n453), .B(n369), .Z(n452) );
  NAND U1490 ( .A(rst), .B(\_MxM/Y0[28] ), .Z(n451) );
  NAND U1491 ( .A(n454), .B(n455), .Z(\_MxM/n312 ) );
  NAND U1492 ( .A(n456), .B(n369), .Z(n455) );
  NAND U1493 ( .A(rst), .B(\_MxM/Y0[29] ), .Z(n454) );
  NAND U1494 ( .A(n457), .B(n458), .Z(\_MxM/n311 ) );
  NAND U1495 ( .A(n459), .B(n369), .Z(n458) );
  NAND U1496 ( .A(rst), .B(\_MxM/Y0[30] ), .Z(n457) );
  NAND U1497 ( .A(n460), .B(n461), .Z(\_MxM/n310 ) );
  NAND U1498 ( .A(n462), .B(n369), .Z(n461) );
  NOR U1499 ( .A(rst), .B(n463), .Z(n369) );
  NAND U1500 ( .A(\_MxM/Y0[31] ), .B(rst), .Z(n460) );
  MUX U1501 ( .IN0(o[31]), .IN1(n462), .SEL(n464), .F(\_MxM/n309 ) );
  XNOR U1502 ( .A(\_MxM/Y0[31] ), .B(n466), .Z(n465) );
  AND U1503 ( .A(n469), .B(n470), .Z(n468) );
  XNOR U1504 ( .A(\_MxM/Y0[31] ), .B(n471), .Z(n470) );
  MUX U1505 ( .IN0(o[30]), .IN1(n459), .SEL(n464), .F(\_MxM/n308 ) );
  XOR U1506 ( .A(n469), .B(\_MxM/Y0[31] ), .Z(n459) );
  XOR U1507 ( .A(n471), .B(n466), .Z(n469) );
  XOR U1508 ( .A(n472), .B(n473), .Z(n466) );
  XOR U1509 ( .A(n474), .B(n475), .Z(n473) );
  AND U1510 ( .A(n476), .B(n477), .Z(n475) );
  XOR U1511 ( .A(n484), .B(n482), .Z(n472) );
  XOR U1512 ( .A(n485), .B(n486), .Z(n484) );
  XOR U1513 ( .A(n487), .B(n488), .Z(n486) );
  XOR U1514 ( .A(n492), .B(n493), .Z(n487) );
  ANDN U1515 ( .A(n494), .B(n495), .Z(n493) );
  XOR U1516 ( .A(n499), .B(n500), .Z(n485) );
  XOR U1517 ( .A(n489), .B(n491), .Z(n500) );
  XOR U1518 ( .A(n498), .B(n495), .Z(n499) );
  IV U1519 ( .A(n467), .Z(n471) );
  MUX U1520 ( .IN0(o[29]), .IN1(n456), .SEL(n464), .F(\_MxM/n307 ) );
  XOR U1521 ( .A(n502), .B(\_MxM/Y0[30] ), .Z(n456) );
  XNOR U1522 ( .A(n503), .B(n504), .Z(n502) );
  AND U1523 ( .A(n476), .B(n506), .Z(n505) );
  XNOR U1524 ( .A(n480), .B(n504), .Z(n506) );
  XOR U1525 ( .A(n478), .B(n504), .Z(n480) );
  XNOR U1526 ( .A(n483), .B(n481), .Z(n504) );
  IV U1527 ( .A(n482), .Z(n481) );
  XNOR U1528 ( .A(n489), .B(n490), .Z(n483) );
  XNOR U1529 ( .A(n491), .B(n494), .Z(n490) );
  XNOR U1530 ( .A(n495), .B(n510), .Z(n494) );
  XOR U1531 ( .A(n496), .B(n497), .Z(n510) );
  NAND U1532 ( .A(n511), .B(n512), .Z(n497) );
  IV U1533 ( .A(n498), .Z(n496) );
  IV U1534 ( .A(n479), .Z(n478) );
  MUX U1535 ( .IN0(o[28]), .IN1(n453), .SEL(n464), .F(\_MxM/n306 ) );
  XOR U1536 ( .A(n525), .B(\_MxM/Y0[29] ), .Z(n453) );
  XNOR U1537 ( .A(n526), .B(n527), .Z(n525) );
  AND U1538 ( .A(n476), .B(n529), .Z(n528) );
  XNOR U1539 ( .A(n523), .B(n527), .Z(n529) );
  XNOR U1540 ( .A(n509), .B(n508), .Z(n527) );
  IV U1541 ( .A(n507), .Z(n508) );
  XOR U1542 ( .A(n521), .B(n520), .Z(n509) );
  XOR U1543 ( .A(n519), .B(n533), .Z(n520) );
  XNOR U1544 ( .A(n518), .B(n517), .Z(n533) );
  XNOR U1545 ( .A(n534), .B(n535), .Z(n517) );
  IV U1546 ( .A(n516), .Z(n535) );
  XNOR U1547 ( .A(n514), .B(n515), .Z(n518) );
  NAND U1548 ( .A(n541), .B(n512), .Z(n515) );
  XNOR U1549 ( .A(n513), .B(n542), .Z(n514) );
  ANDN U1550 ( .A(n543), .B(n544), .Z(n542) );
  MUX U1551 ( .IN0(o[27]), .IN1(n450), .SEL(n464), .F(\_MxM/n305 ) );
  XOR U1552 ( .A(n554), .B(\_MxM/Y0[28] ), .Z(n450) );
  XNOR U1553 ( .A(n555), .B(n556), .Z(n554) );
  AND U1554 ( .A(n476), .B(n558), .Z(n557) );
  XNOR U1555 ( .A(n552), .B(n556), .Z(n558) );
  XNOR U1556 ( .A(n532), .B(n531), .Z(n556) );
  IV U1557 ( .A(n530), .Z(n531) );
  XOR U1558 ( .A(n550), .B(n549), .Z(n532) );
  XOR U1559 ( .A(n548), .B(n562), .Z(n549) );
  XNOR U1560 ( .A(n538), .B(n537), .Z(n562) );
  XOR U1561 ( .A(n567), .B(n539), .Z(n563) );
  AND U1562 ( .A(n568), .B(n511), .Z(n539) );
  IV U1563 ( .A(n536), .Z(n567) );
  XNOR U1564 ( .A(n546), .B(n547), .Z(n538) );
  NAND U1565 ( .A(n572), .B(n512), .Z(n547) );
  XNOR U1566 ( .A(n545), .B(n573), .Z(n546) );
  ANDN U1567 ( .A(n543), .B(n574), .Z(n573) );
  MUX U1568 ( .IN0(o[26]), .IN1(n447), .SEL(n464), .F(\_MxM/n304 ) );
  XOR U1569 ( .A(n585), .B(\_MxM/Y0[27] ), .Z(n447) );
  XNOR U1570 ( .A(n586), .B(n587), .Z(n585) );
  AND U1571 ( .A(n476), .B(n589), .Z(n588) );
  XNOR U1572 ( .A(n583), .B(n587), .Z(n589) );
  XNOR U1573 ( .A(n561), .B(n560), .Z(n587) );
  IV U1574 ( .A(n559), .Z(n560) );
  XNOR U1575 ( .A(n581), .B(n593), .Z(n561) );
  XOR U1576 ( .A(n580), .B(n579), .Z(n593) );
  XOR U1577 ( .A(n594), .B(n595), .Z(n579) );
  XOR U1578 ( .A(n596), .B(n597), .Z(n595) );
  XOR U1579 ( .A(n598), .B(n599), .Z(n597) );
  XNOR U1580 ( .A(n571), .B(n570), .Z(n580) );
  XOR U1581 ( .A(n607), .B(n565), .Z(n570) );
  XNOR U1582 ( .A(n564), .B(n608), .Z(n565) );
  ANDN U1583 ( .A(n609), .B(n544), .Z(n608) );
  AND U1584 ( .A(n541), .B(n568), .Z(n566) );
  XNOR U1585 ( .A(n576), .B(n577), .Z(n571) );
  NAND U1586 ( .A(n616), .B(n512), .Z(n577) );
  XNOR U1587 ( .A(n575), .B(n617), .Z(n576) );
  ANDN U1588 ( .A(n543), .B(n618), .Z(n617) );
  MUX U1589 ( .IN0(o[25]), .IN1(n444), .SEL(n464), .F(\_MxM/n303 ) );
  XOR U1590 ( .A(n626), .B(\_MxM/Y0[26] ), .Z(n444) );
  XNOR U1591 ( .A(n627), .B(n628), .Z(n626) );
  AND U1592 ( .A(n476), .B(n630), .Z(n629) );
  XNOR U1593 ( .A(n624), .B(n628), .Z(n630) );
  XNOR U1594 ( .A(n592), .B(n591), .Z(n628) );
  IV U1595 ( .A(n590), .Z(n591) );
  XOR U1596 ( .A(n622), .B(n634), .Z(n592) );
  XNOR U1597 ( .A(n606), .B(n605), .Z(n634) );
  XOR U1598 ( .A(n635), .B(n600), .Z(n605) );
  XOR U1599 ( .A(n601), .B(n602), .Z(n600) );
  NANDN U1600 ( .B(n636), .A(n511), .Z(n602) );
  IV U1601 ( .A(n603), .Z(n601) );
  XOR U1602 ( .A(n596), .B(n604), .Z(n635) );
  XNOR U1603 ( .A(n615), .B(n614), .Z(n606) );
  XOR U1604 ( .A(n646), .B(n611), .Z(n614) );
  XNOR U1605 ( .A(n610), .B(n647), .Z(n611) );
  ANDN U1606 ( .A(n609), .B(n574), .Z(n647) );
  XOR U1607 ( .A(n648), .B(n649), .Z(n610) );
  AND U1608 ( .A(n650), .B(n651), .Z(n649) );
  XNOR U1609 ( .A(n652), .B(n648), .Z(n651) );
  AND U1610 ( .A(n572), .B(n568), .Z(n612) );
  XNOR U1611 ( .A(n620), .B(n621), .Z(n615) );
  NAND U1612 ( .A(n656), .B(n512), .Z(n621) );
  XNOR U1613 ( .A(n619), .B(n657), .Z(n620) );
  ANDN U1614 ( .A(n543), .B(n658), .Z(n657) );
  MUX U1615 ( .IN0(o[24]), .IN1(n441), .SEL(n464), .F(\_MxM/n302 ) );
  XOR U1616 ( .A(n666), .B(\_MxM/Y0[25] ), .Z(n441) );
  XNOR U1617 ( .A(n667), .B(n668), .Z(n666) );
  AND U1618 ( .A(n476), .B(n670), .Z(n669) );
  XNOR U1619 ( .A(n664), .B(n668), .Z(n670) );
  XNOR U1620 ( .A(n633), .B(n632), .Z(n668) );
  IV U1621 ( .A(n631), .Z(n632) );
  XOR U1622 ( .A(n662), .B(n674), .Z(n633) );
  XNOR U1623 ( .A(n642), .B(n641), .Z(n674) );
  XOR U1624 ( .A(n675), .B(n645), .Z(n641) );
  XNOR U1625 ( .A(n638), .B(n639), .Z(n645) );
  NANDN U1626 ( .B(n636), .A(n541), .Z(n639) );
  XNOR U1627 ( .A(n637), .B(n676), .Z(n638) );
  ANDN U1628 ( .A(n677), .B(n544), .Z(n676) );
  XNOR U1629 ( .A(n644), .B(n640), .Z(n675) );
  XNOR U1630 ( .A(n684), .B(n685), .Z(n644) );
  IV U1631 ( .A(n643), .Z(n685) );
  XNOR U1632 ( .A(n655), .B(n654), .Z(n642) );
  XOR U1633 ( .A(n692), .B(n650), .Z(n654) );
  XNOR U1634 ( .A(n648), .B(n693), .Z(n650) );
  ANDN U1635 ( .A(n609), .B(n618), .Z(n693) );
  AND U1636 ( .A(n616), .B(n568), .Z(n652) );
  XNOR U1637 ( .A(n660), .B(n661), .Z(n655) );
  NAND U1638 ( .A(n700), .B(n512), .Z(n661) );
  XNOR U1639 ( .A(n659), .B(n701), .Z(n660) );
  ANDN U1640 ( .A(n543), .B(n702), .Z(n701) );
  MUX U1641 ( .IN0(o[23]), .IN1(n438), .SEL(n464), .F(\_MxM/n301 ) );
  XOR U1642 ( .A(n710), .B(\_MxM/Y0[24] ), .Z(n438) );
  XNOR U1643 ( .A(n711), .B(n712), .Z(n710) );
  AND U1644 ( .A(n476), .B(n714), .Z(n713) );
  XNOR U1645 ( .A(n708), .B(n712), .Z(n714) );
  XNOR U1646 ( .A(n673), .B(n672), .Z(n712) );
  IV U1647 ( .A(n671), .Z(n672) );
  XOR U1648 ( .A(n706), .B(n717), .Z(n673) );
  XNOR U1649 ( .A(n683), .B(n682), .Z(n717) );
  XOR U1650 ( .A(n718), .B(n688), .Z(n682) );
  XNOR U1651 ( .A(n679), .B(n680), .Z(n688) );
  NANDN U1652 ( .B(n636), .A(n572), .Z(n680) );
  XNOR U1653 ( .A(n678), .B(n719), .Z(n679) );
  ANDN U1654 ( .A(n677), .B(n574), .Z(n719) );
  XNOR U1655 ( .A(n687), .B(n681), .Z(n718) );
  XNOR U1656 ( .A(n726), .B(n689), .Z(n687) );
  IV U1657 ( .A(n691), .Z(n689) );
  AND U1658 ( .A(n730), .B(n511), .Z(n690) );
  XNOR U1659 ( .A(n699), .B(n698), .Z(n683) );
  XOR U1660 ( .A(n734), .B(n695), .Z(n698) );
  XNOR U1661 ( .A(n694), .B(n735), .Z(n695) );
  ANDN U1662 ( .A(n609), .B(n658), .Z(n735) );
  AND U1663 ( .A(n656), .B(n568), .Z(n696) );
  XNOR U1664 ( .A(n704), .B(n705), .Z(n699) );
  NAND U1665 ( .A(n742), .B(n512), .Z(n705) );
  XNOR U1666 ( .A(n703), .B(n743), .Z(n704) );
  ANDN U1667 ( .A(n543), .B(n744), .Z(n743) );
  MUX U1668 ( .IN0(o[22]), .IN1(n435), .SEL(n464), .F(\_MxM/n300 ) );
  XOR U1669 ( .A(n754), .B(\_MxM/Y0[23] ), .Z(n435) );
  XNOR U1670 ( .A(n755), .B(n716), .Z(n754) );
  AND U1671 ( .A(n476), .B(n757), .Z(n756) );
  XNOR U1672 ( .A(n752), .B(n716), .Z(n757) );
  XOR U1673 ( .A(n715), .B(n758), .Z(n716) );
  XNOR U1674 ( .A(n750), .B(n749), .Z(n758) );
  XOR U1675 ( .A(n759), .B(n760), .Z(n749) );
  XOR U1676 ( .A(n761), .B(n762), .Z(n760) );
  XOR U1677 ( .A(n765), .B(n766), .Z(n761) );
  ANDN U1678 ( .A(n764), .B(n767), .Z(n766) );
  XNOR U1679 ( .A(n770), .B(n748), .Z(n759) );
  XOR U1680 ( .A(n769), .B(n767), .Z(n770) );
  XNOR U1681 ( .A(n725), .B(n724), .Z(n750) );
  XOR U1682 ( .A(n774), .B(n733), .Z(n724) );
  XNOR U1683 ( .A(n721), .B(n722), .Z(n733) );
  NANDN U1684 ( .B(n636), .A(n616), .Z(n722) );
  XNOR U1685 ( .A(n720), .B(n775), .Z(n721) );
  ANDN U1686 ( .A(n677), .B(n618), .Z(n775) );
  XNOR U1687 ( .A(n732), .B(n723), .Z(n774) );
  XOR U1688 ( .A(n782), .B(n728), .Z(n732) );
  XNOR U1689 ( .A(n727), .B(n783), .Z(n728) );
  ANDN U1690 ( .A(n784), .B(n544), .Z(n783) );
  XOR U1691 ( .A(n785), .B(n786), .Z(n727) );
  AND U1692 ( .A(n787), .B(n788), .Z(n786) );
  XNOR U1693 ( .A(n789), .B(n785), .Z(n788) );
  AND U1694 ( .A(n541), .B(n730), .Z(n729) );
  XNOR U1695 ( .A(n741), .B(n740), .Z(n725) );
  XOR U1696 ( .A(n793), .B(n737), .Z(n740) );
  XNOR U1697 ( .A(n736), .B(n794), .Z(n737) );
  ANDN U1698 ( .A(n609), .B(n702), .Z(n794) );
  AND U1699 ( .A(n700), .B(n568), .Z(n738) );
  XNOR U1700 ( .A(n746), .B(n747), .Z(n741) );
  NAND U1701 ( .A(n801), .B(n512), .Z(n747) );
  XNOR U1702 ( .A(n745), .B(n802), .Z(n746) );
  ANDN U1703 ( .A(n543), .B(n803), .Z(n802) );
  MUX U1704 ( .IN0(o[21]), .IN1(n432), .SEL(n464), .F(\_MxM/n299 ) );
  XOR U1705 ( .A(n813), .B(\_MxM/Y0[22] ), .Z(n432) );
  XNOR U1706 ( .A(n814), .B(n815), .Z(n813) );
  AND U1707 ( .A(n476), .B(n817), .Z(n816) );
  XNOR U1708 ( .A(n811), .B(n815), .Z(n817) );
  XNOR U1709 ( .A(n809), .B(n808), .Z(n815) );
  IV U1710 ( .A(n807), .Z(n808) );
  XNOR U1711 ( .A(n773), .B(n772), .Z(n809) );
  XOR U1712 ( .A(n821), .B(n764), .Z(n772) );
  XNOR U1713 ( .A(n767), .B(n822), .Z(n764) );
  NANDN U1714 ( .B(n823), .A(n511), .Z(n768) );
  XOR U1715 ( .A(n763), .B(n771), .Z(n821) );
  XNOR U1716 ( .A(n781), .B(n780), .Z(n773) );
  XOR U1717 ( .A(n835), .B(n792), .Z(n780) );
  XNOR U1718 ( .A(n777), .B(n778), .Z(n792) );
  NANDN U1719 ( .B(n636), .A(n656), .Z(n778) );
  XNOR U1720 ( .A(n776), .B(n836), .Z(n777) );
  ANDN U1721 ( .A(n677), .B(n658), .Z(n836) );
  XOR U1722 ( .A(n837), .B(n838), .Z(n776) );
  AND U1723 ( .A(n839), .B(n840), .Z(n838) );
  XOR U1724 ( .A(n841), .B(n837), .Z(n840) );
  XNOR U1725 ( .A(n791), .B(n779), .Z(n835) );
  XOR U1726 ( .A(n845), .B(n787), .Z(n791) );
  XNOR U1727 ( .A(n785), .B(n846), .Z(n787) );
  ANDN U1728 ( .A(n784), .B(n574), .Z(n846) );
  XOR U1729 ( .A(n847), .B(n848), .Z(n785) );
  AND U1730 ( .A(n849), .B(n850), .Z(n848) );
  XNOR U1731 ( .A(n851), .B(n847), .Z(n850) );
  AND U1732 ( .A(n572), .B(n730), .Z(n789) );
  XNOR U1733 ( .A(n800), .B(n799), .Z(n781) );
  XOR U1734 ( .A(n855), .B(n796), .Z(n799) );
  XNOR U1735 ( .A(n795), .B(n856), .Z(n796) );
  ANDN U1736 ( .A(n609), .B(n744), .Z(n856) );
  XOR U1737 ( .A(n857), .B(n858), .Z(n795) );
  AND U1738 ( .A(n859), .B(n860), .Z(n858) );
  XNOR U1739 ( .A(n861), .B(n857), .Z(n860) );
  AND U1740 ( .A(n742), .B(n568), .Z(n797) );
  XNOR U1741 ( .A(n805), .B(n806), .Z(n800) );
  NAND U1742 ( .A(n865), .B(n512), .Z(n806) );
  XNOR U1743 ( .A(n804), .B(n866), .Z(n805) );
  ANDN U1744 ( .A(n543), .B(n867), .Z(n866) );
  XOR U1745 ( .A(n868), .B(n869), .Z(n804) );
  AND U1746 ( .A(n870), .B(n871), .Z(n869) );
  XOR U1747 ( .A(n872), .B(n868), .Z(n871) );
  MUX U1748 ( .IN0(o[20]), .IN1(n429), .SEL(n464), .F(\_MxM/n298 ) );
  XOR U1749 ( .A(n876), .B(\_MxM/Y0[21] ), .Z(n429) );
  XNOR U1750 ( .A(n877), .B(n878), .Z(n876) );
  AND U1751 ( .A(n476), .B(n880), .Z(n879) );
  XNOR U1752 ( .A(n874), .B(n878), .Z(n880) );
  XNOR U1753 ( .A(n820), .B(n819), .Z(n878) );
  IV U1754 ( .A(n818), .Z(n819) );
  XNOR U1755 ( .A(n832), .B(n831), .Z(n820) );
  XOR U1756 ( .A(n884), .B(n834), .Z(n831) );
  XNOR U1757 ( .A(n829), .B(n828), .Z(n834) );
  XNOR U1758 ( .A(n885), .B(n886), .Z(n828) );
  IV U1759 ( .A(n827), .Z(n886) );
  XNOR U1760 ( .A(n825), .B(n826), .Z(n829) );
  NANDN U1761 ( .B(n823), .A(n541), .Z(n826) );
  XNOR U1762 ( .A(n824), .B(n892), .Z(n825) );
  ANDN U1763 ( .A(n893), .B(n544), .Z(n892) );
  XNOR U1764 ( .A(n844), .B(n843), .Z(n832) );
  XOR U1765 ( .A(n903), .B(n854), .Z(n843) );
  XNOR U1766 ( .A(n839), .B(n841), .Z(n854) );
  NANDN U1767 ( .B(n636), .A(n700), .Z(n841) );
  XNOR U1768 ( .A(n837), .B(n904), .Z(n839) );
  ANDN U1769 ( .A(n677), .B(n702), .Z(n904) );
  XOR U1770 ( .A(n905), .B(n906), .Z(n837) );
  AND U1771 ( .A(n907), .B(n908), .Z(n906) );
  XOR U1772 ( .A(n909), .B(n905), .Z(n908) );
  XNOR U1773 ( .A(n853), .B(n842), .Z(n903) );
  XOR U1774 ( .A(n913), .B(n849), .Z(n853) );
  XNOR U1775 ( .A(n847), .B(n914), .Z(n849) );
  ANDN U1776 ( .A(n784), .B(n618), .Z(n914) );
  XOR U1777 ( .A(n915), .B(n916), .Z(n847) );
  AND U1778 ( .A(n917), .B(n918), .Z(n916) );
  XNOR U1779 ( .A(n919), .B(n915), .Z(n918) );
  AND U1780 ( .A(n616), .B(n730), .Z(n851) );
  XNOR U1781 ( .A(n864), .B(n863), .Z(n844) );
  XOR U1782 ( .A(n923), .B(n859), .Z(n863) );
  XNOR U1783 ( .A(n857), .B(n924), .Z(n859) );
  ANDN U1784 ( .A(n609), .B(n803), .Z(n924) );
  XOR U1785 ( .A(n925), .B(n926), .Z(n857) );
  AND U1786 ( .A(n927), .B(n928), .Z(n926) );
  XNOR U1787 ( .A(n929), .B(n925), .Z(n928) );
  AND U1788 ( .A(n801), .B(n568), .Z(n861) );
  XNOR U1789 ( .A(n870), .B(n872), .Z(n864) );
  NAND U1790 ( .A(n933), .B(n512), .Z(n872) );
  XNOR U1791 ( .A(n868), .B(n934), .Z(n870) );
  ANDN U1792 ( .A(n543), .B(n935), .Z(n934) );
  XOR U1793 ( .A(n936), .B(n937), .Z(n868) );
  AND U1794 ( .A(n938), .B(n939), .Z(n937) );
  XOR U1795 ( .A(n940), .B(n936), .Z(n939) );
  MUX U1796 ( .IN0(o[19]), .IN1(n426), .SEL(n464), .F(\_MxM/n297 ) );
  XOR U1797 ( .A(n944), .B(\_MxM/Y0[20] ), .Z(n426) );
  XNOR U1798 ( .A(n945), .B(n946), .Z(n944) );
  AND U1799 ( .A(n476), .B(n948), .Z(n947) );
  XNOR U1800 ( .A(n942), .B(n946), .Z(n948) );
  XNOR U1801 ( .A(n883), .B(n882), .Z(n946) );
  IV U1802 ( .A(n881), .Z(n882) );
  XNOR U1803 ( .A(n899), .B(n898), .Z(n883) );
  XOR U1804 ( .A(n952), .B(n902), .Z(n898) );
  XNOR U1805 ( .A(n889), .B(n888), .Z(n902) );
  XOR U1806 ( .A(n957), .B(n890), .Z(n953) );
  AND U1807 ( .A(n958), .B(n511), .Z(n890) );
  IV U1808 ( .A(n887), .Z(n957) );
  XNOR U1809 ( .A(n895), .B(n896), .Z(n889) );
  NANDN U1810 ( .B(n823), .A(n572), .Z(n896) );
  XNOR U1811 ( .A(n894), .B(n962), .Z(n895) );
  ANDN U1812 ( .A(n893), .B(n574), .Z(n962) );
  XNOR U1813 ( .A(n901), .B(n897), .Z(n952) );
  IV U1814 ( .A(n900), .Z(n901) );
  XNOR U1815 ( .A(n912), .B(n911), .Z(n899) );
  XOR U1816 ( .A(n972), .B(n922), .Z(n911) );
  XNOR U1817 ( .A(n907), .B(n909), .Z(n922) );
  NANDN U1818 ( .B(n636), .A(n742), .Z(n909) );
  XNOR U1819 ( .A(n905), .B(n973), .Z(n907) );
  ANDN U1820 ( .A(n677), .B(n744), .Z(n973) );
  XOR U1821 ( .A(n974), .B(n975), .Z(n905) );
  AND U1822 ( .A(n976), .B(n977), .Z(n975) );
  XOR U1823 ( .A(n978), .B(n974), .Z(n977) );
  XNOR U1824 ( .A(n921), .B(n910), .Z(n972) );
  XOR U1825 ( .A(n982), .B(n917), .Z(n921) );
  XNOR U1826 ( .A(n915), .B(n983), .Z(n917) );
  ANDN U1827 ( .A(n784), .B(n658), .Z(n983) );
  XOR U1828 ( .A(n984), .B(n985), .Z(n915) );
  AND U1829 ( .A(n986), .B(n987), .Z(n985) );
  XNOR U1830 ( .A(n988), .B(n984), .Z(n987) );
  AND U1831 ( .A(n656), .B(n730), .Z(n919) );
  XNOR U1832 ( .A(n932), .B(n931), .Z(n912) );
  XOR U1833 ( .A(n992), .B(n927), .Z(n931) );
  XNOR U1834 ( .A(n925), .B(n993), .Z(n927) );
  ANDN U1835 ( .A(n609), .B(n867), .Z(n993) );
  AND U1836 ( .A(n865), .B(n568), .Z(n929) );
  XNOR U1837 ( .A(n938), .B(n940), .Z(n932) );
  NAND U1838 ( .A(n1000), .B(n512), .Z(n940) );
  XNOR U1839 ( .A(n936), .B(n1001), .Z(n938) );
  ANDN U1840 ( .A(n543), .B(n1002), .Z(n1001) );
  XOR U1841 ( .A(n1003), .B(n1004), .Z(n936) );
  AND U1842 ( .A(n1005), .B(n1006), .Z(n1004) );
  XOR U1843 ( .A(n1007), .B(n1003), .Z(n1006) );
  MUX U1844 ( .IN0(o[18]), .IN1(n423), .SEL(n464), .F(\_MxM/n296 ) );
  XOR U1845 ( .A(n1011), .B(\_MxM/Y0[19] ), .Z(n423) );
  XNOR U1846 ( .A(n1012), .B(n1013), .Z(n1011) );
  AND U1847 ( .A(n476), .B(n1015), .Z(n1014) );
  XOR U1848 ( .A(n1009), .B(n1013), .Z(n1015) );
  XOR U1849 ( .A(n1008), .B(n1013), .Z(n1009) );
  XNOR U1850 ( .A(n951), .B(n950), .Z(n1013) );
  IV U1851 ( .A(n949), .Z(n950) );
  XNOR U1852 ( .A(n968), .B(n967), .Z(n951) );
  XOR U1853 ( .A(n1018), .B(n971), .Z(n967) );
  XNOR U1854 ( .A(n961), .B(n960), .Z(n971) );
  XOR U1855 ( .A(n1019), .B(n955), .Z(n960) );
  XNOR U1856 ( .A(n954), .B(n1020), .Z(n955) );
  ANDN U1857 ( .A(n1021), .B(n544), .Z(n1020) );
  XOR U1858 ( .A(n1022), .B(n1023), .Z(n954) );
  AND U1859 ( .A(n1024), .B(n1025), .Z(n1023) );
  XNOR U1860 ( .A(n1026), .B(n1022), .Z(n1025) );
  AND U1861 ( .A(n541), .B(n958), .Z(n956) );
  XNOR U1862 ( .A(n964), .B(n965), .Z(n961) );
  NANDN U1863 ( .B(n823), .A(n616), .Z(n965) );
  XNOR U1864 ( .A(n963), .B(n1030), .Z(n964) );
  ANDN U1865 ( .A(n893), .B(n618), .Z(n1030) );
  XNOR U1866 ( .A(n970), .B(n966), .Z(n1018) );
  XNOR U1867 ( .A(n1037), .B(n1038), .Z(n970) );
  IV U1868 ( .A(n969), .Z(n1038) );
  XNOR U1869 ( .A(n981), .B(n980), .Z(n968) );
  XOR U1870 ( .A(n1044), .B(n991), .Z(n980) );
  XNOR U1871 ( .A(n976), .B(n978), .Z(n991) );
  NANDN U1872 ( .B(n636), .A(n801), .Z(n978) );
  XNOR U1873 ( .A(n974), .B(n1045), .Z(n976) );
  ANDN U1874 ( .A(n677), .B(n803), .Z(n1045) );
  XOR U1875 ( .A(n1046), .B(n1047), .Z(n974) );
  AND U1876 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR U1877 ( .A(n1050), .B(n1046), .Z(n1049) );
  XNOR U1878 ( .A(n990), .B(n979), .Z(n1044) );
  XOR U1879 ( .A(n1054), .B(n986), .Z(n990) );
  XNOR U1880 ( .A(n984), .B(n1055), .Z(n986) );
  ANDN U1881 ( .A(n784), .B(n702), .Z(n1055) );
  XOR U1882 ( .A(n1056), .B(n1057), .Z(n984) );
  AND U1883 ( .A(n1058), .B(n1059), .Z(n1057) );
  XNOR U1884 ( .A(n1060), .B(n1056), .Z(n1059) );
  AND U1885 ( .A(n700), .B(n730), .Z(n988) );
  XNOR U1886 ( .A(n999), .B(n998), .Z(n981) );
  XOR U1887 ( .A(n1064), .B(n995), .Z(n998) );
  XNOR U1888 ( .A(n994), .B(n1065), .Z(n995) );
  ANDN U1889 ( .A(n609), .B(n935), .Z(n1065) );
  XOR U1890 ( .A(n1066), .B(n1067), .Z(n994) );
  AND U1891 ( .A(n1068), .B(n1069), .Z(n1067) );
  XNOR U1892 ( .A(n1070), .B(n1066), .Z(n1069) );
  AND U1893 ( .A(n933), .B(n568), .Z(n996) );
  XNOR U1894 ( .A(n1005), .B(n1007), .Z(n999) );
  NAND U1895 ( .A(n1074), .B(n512), .Z(n1007) );
  XNOR U1896 ( .A(n1003), .B(n1075), .Z(n1005) );
  ANDN U1897 ( .A(n543), .B(n1076), .Z(n1075) );
  NANDN U1898 ( .B(n1077), .A(n1078), .Z(n1003) );
  NAND U1899 ( .A(n1079), .B(n1080), .Z(n1078) );
  MUX U1900 ( .IN0(o[17]), .IN1(n420), .SEL(n464), .F(\_MxM/n295 ) );
  XOR U1901 ( .A(n1085), .B(\_MxM/Y0[18] ), .Z(n420) );
  XOR U1902 ( .A(n1086), .B(n1087), .Z(n1085) );
  AND U1903 ( .A(n476), .B(n1089), .Z(n1088) );
  XOR U1904 ( .A(n1083), .B(n1087), .Z(n1089) );
  XOR U1905 ( .A(n1082), .B(n1087), .Z(n1083) );
  XOR U1906 ( .A(n1017), .B(n1016), .Z(n1087) );
  XNOR U1907 ( .A(n1092), .B(n1041), .Z(n1035) );
  XNOR U1908 ( .A(n1029), .B(n1028), .Z(n1041) );
  XOR U1909 ( .A(n1093), .B(n1024), .Z(n1028) );
  XNOR U1910 ( .A(n1022), .B(n1094), .Z(n1024) );
  ANDN U1911 ( .A(n1021), .B(n574), .Z(n1094) );
  XOR U1912 ( .A(n1095), .B(n1096), .Z(n1022) );
  AND U1913 ( .A(n1097), .B(n1098), .Z(n1096) );
  XNOR U1914 ( .A(n1099), .B(n1095), .Z(n1098) );
  AND U1915 ( .A(n572), .B(n958), .Z(n1026) );
  XNOR U1916 ( .A(n1032), .B(n1033), .Z(n1029) );
  NANDN U1917 ( .B(n823), .A(n656), .Z(n1033) );
  XNOR U1918 ( .A(n1031), .B(n1103), .Z(n1032) );
  ANDN U1919 ( .A(n893), .B(n658), .Z(n1103) );
  XOR U1920 ( .A(n1104), .B(n1105), .Z(n1031) );
  AND U1921 ( .A(n1106), .B(n1107), .Z(n1105) );
  XOR U1922 ( .A(n1108), .B(n1104), .Z(n1107) );
  XNOR U1923 ( .A(n1040), .B(n1034), .Z(n1092) );
  XOR U1924 ( .A(n1112), .B(n1042), .Z(n1040) );
  NAND U1925 ( .A(n1116), .B(n1117), .Z(n1043) );
  NANDN U1926 ( .B(n1118), .A(n511), .Z(n1117) );
  NANDN U1927 ( .B(n1119), .A(n1120), .Z(n1116) );
  XNOR U1928 ( .A(n1053), .B(n1052), .Z(n1036) );
  XOR U1929 ( .A(n1124), .B(n1063), .Z(n1052) );
  XNOR U1930 ( .A(n1048), .B(n1050), .Z(n1063) );
  NANDN U1931 ( .B(n636), .A(n865), .Z(n1050) );
  XNOR U1932 ( .A(n1046), .B(n1125), .Z(n1048) );
  ANDN U1933 ( .A(n677), .B(n867), .Z(n1125) );
  XOR U1934 ( .A(n1126), .B(n1127), .Z(n1046) );
  AND U1935 ( .A(n1128), .B(n1129), .Z(n1127) );
  XOR U1936 ( .A(n1130), .B(n1126), .Z(n1129) );
  XNOR U1937 ( .A(n1062), .B(n1051), .Z(n1124) );
  XOR U1938 ( .A(n1134), .B(n1058), .Z(n1062) );
  XNOR U1939 ( .A(n1056), .B(n1135), .Z(n1058) );
  ANDN U1940 ( .A(n784), .B(n744), .Z(n1135) );
  XOR U1941 ( .A(n1136), .B(n1137), .Z(n1056) );
  AND U1942 ( .A(n1138), .B(n1139), .Z(n1137) );
  XNOR U1943 ( .A(n1140), .B(n1136), .Z(n1139) );
  AND U1944 ( .A(n742), .B(n730), .Z(n1060) );
  XOR U1945 ( .A(n1073), .B(n1072), .Z(n1053) );
  XOR U1946 ( .A(n1144), .B(n1068), .Z(n1072) );
  XNOR U1947 ( .A(n1066), .B(n1145), .Z(n1068) );
  ANDN U1948 ( .A(n609), .B(n1002), .Z(n1145) );
  AND U1949 ( .A(n1000), .B(n568), .Z(n1070) );
  XOR U1950 ( .A(n1080), .B(n1079), .Z(n1073) );
  NAND U1951 ( .A(n1152), .B(n512), .Z(n1079) );
  XNOR U1952 ( .A(n1077), .B(n1153), .Z(n1080) );
  ANDN U1953 ( .A(n543), .B(n1154), .Z(n1153) );
  NANDN U1954 ( .B(n1155), .A(n1156), .Z(n1077) );
  NAND U1955 ( .A(n1157), .B(n1158), .Z(n1156) );
  IV U1956 ( .A(n1081), .Z(n1082) );
  MUX U1957 ( .IN0(o[16]), .IN1(n417), .SEL(n464), .F(\_MxM/n294 ) );
  XOR U1958 ( .A(n1163), .B(\_MxM/Y0[17] ), .Z(n417) );
  XOR U1959 ( .A(n1164), .B(n1165), .Z(n1163) );
  AND U1960 ( .A(n476), .B(n1167), .Z(n1166) );
  XOR U1961 ( .A(n1161), .B(n1165), .Z(n1167) );
  XOR U1962 ( .A(n1160), .B(n1165), .Z(n1161) );
  XOR U1963 ( .A(n1091), .B(n1090), .Z(n1165) );
  XNOR U1964 ( .A(n1170), .B(n1123), .Z(n1110) );
  XNOR U1965 ( .A(n1102), .B(n1101), .Z(n1123) );
  XOR U1966 ( .A(n1171), .B(n1097), .Z(n1101) );
  XNOR U1967 ( .A(n1095), .B(n1172), .Z(n1097) );
  ANDN U1968 ( .A(n1021), .B(n618), .Z(n1172) );
  XOR U1969 ( .A(n1173), .B(n1174), .Z(n1095) );
  AND U1970 ( .A(n1175), .B(n1176), .Z(n1174) );
  XNOR U1971 ( .A(n1177), .B(n1173), .Z(n1176) );
  AND U1972 ( .A(n616), .B(n958), .Z(n1099) );
  XNOR U1973 ( .A(n1106), .B(n1108), .Z(n1102) );
  NANDN U1974 ( .B(n823), .A(n700), .Z(n1108) );
  XNOR U1975 ( .A(n1104), .B(n1181), .Z(n1106) );
  ANDN U1976 ( .A(n893), .B(n702), .Z(n1181) );
  XOR U1977 ( .A(n1182), .B(n1183), .Z(n1104) );
  AND U1978 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U1979 ( .A(n1186), .B(n1182), .Z(n1185) );
  XOR U1980 ( .A(n1122), .B(n1109), .Z(n1170) );
  XNOR U1981 ( .A(n1190), .B(n1114), .Z(n1122) );
  XNOR U1982 ( .A(n1191), .B(n1120), .Z(n1114) );
  AND U1983 ( .A(n541), .B(n1192), .Z(n1120) );
  NAND U1984 ( .A(n1193), .B(n1119), .Z(n1191) );
  XOR U1985 ( .A(n1194), .B(n1195), .Z(n1119) );
  AND U1986 ( .A(n1196), .B(n1197), .Z(n1195) );
  XOR U1987 ( .A(n1198), .B(n1194), .Z(n1197) );
  NANDN U1988 ( .B(n544), .A(n1199), .Z(n1193) );
  XNOR U1989 ( .A(n1113), .B(n1121), .Z(n1190) );
  IV U1990 ( .A(n1115), .Z(n1113) );
  XNOR U1991 ( .A(n1133), .B(n1132), .Z(n1111) );
  XOR U1992 ( .A(n1205), .B(n1143), .Z(n1132) );
  XNOR U1993 ( .A(n1128), .B(n1130), .Z(n1143) );
  NANDN U1994 ( .B(n636), .A(n933), .Z(n1130) );
  XNOR U1995 ( .A(n1126), .B(n1206), .Z(n1128) );
  ANDN U1996 ( .A(n677), .B(n935), .Z(n1206) );
  XNOR U1997 ( .A(n1142), .B(n1131), .Z(n1205) );
  XOR U1998 ( .A(n1213), .B(n1138), .Z(n1142) );
  XNOR U1999 ( .A(n1136), .B(n1214), .Z(n1138) );
  ANDN U2000 ( .A(n784), .B(n803), .Z(n1214) );
  XOR U2001 ( .A(n1215), .B(n1216), .Z(n1136) );
  AND U2002 ( .A(n1217), .B(n1218), .Z(n1216) );
  XNOR U2003 ( .A(n1219), .B(n1215), .Z(n1218) );
  AND U2004 ( .A(n801), .B(n730), .Z(n1140) );
  XOR U2005 ( .A(n1151), .B(n1150), .Z(n1133) );
  XOR U2006 ( .A(n1223), .B(n1147), .Z(n1150) );
  XNOR U2007 ( .A(n1146), .B(n1224), .Z(n1147) );
  ANDN U2008 ( .A(n609), .B(n1076), .Z(n1224) );
  XOR U2009 ( .A(n1225), .B(n1226), .Z(n1146) );
  AND U2010 ( .A(n1227), .B(n1228), .Z(n1226) );
  XNOR U2011 ( .A(n1229), .B(n1225), .Z(n1228) );
  AND U2012 ( .A(n1074), .B(n568), .Z(n1148) );
  XOR U2013 ( .A(n1158), .B(n1157), .Z(n1151) );
  NAND U2014 ( .A(n1233), .B(n512), .Z(n1157) );
  XNOR U2015 ( .A(n1155), .B(n1234), .Z(n1158) );
  ANDN U2016 ( .A(n543), .B(n1235), .Z(n1234) );
  NAND U2017 ( .A(n1236), .B(n1237), .Z(n1155) );
  NAND U2018 ( .A(n1238), .B(n1239), .Z(n1236) );
  IV U2019 ( .A(n1159), .Z(n1160) );
  MUX U2020 ( .IN0(o[15]), .IN1(n414), .SEL(n464), .F(\_MxM/n293 ) );
  XOR U2021 ( .A(n1244), .B(\_MxM/Y0[16] ), .Z(n414) );
  XOR U2022 ( .A(n1245), .B(n1246), .Z(n1244) );
  AND U2023 ( .A(n476), .B(n1248), .Z(n1247) );
  XOR U2024 ( .A(n1242), .B(n1246), .Z(n1248) );
  XOR U2025 ( .A(n1241), .B(n1246), .Z(n1242) );
  XOR U2026 ( .A(n1169), .B(n1168), .Z(n1246) );
  XNOR U2027 ( .A(n1252), .B(n1202), .Z(n1188) );
  XNOR U2028 ( .A(n1180), .B(n1179), .Z(n1202) );
  XOR U2029 ( .A(n1253), .B(n1175), .Z(n1179) );
  XNOR U2030 ( .A(n1173), .B(n1254), .Z(n1175) );
  ANDN U2031 ( .A(n1021), .B(n658), .Z(n1254) );
  XOR U2032 ( .A(n1255), .B(n1256), .Z(n1173) );
  AND U2033 ( .A(n1257), .B(n1258), .Z(n1256) );
  XNOR U2034 ( .A(n1259), .B(n1255), .Z(n1258) );
  AND U2035 ( .A(n656), .B(n958), .Z(n1177) );
  XNOR U2036 ( .A(n1184), .B(n1186), .Z(n1180) );
  NANDN U2037 ( .B(n823), .A(n742), .Z(n1186) );
  XNOR U2038 ( .A(n1182), .B(n1263), .Z(n1184) );
  ANDN U2039 ( .A(n893), .B(n744), .Z(n1263) );
  XNOR U2040 ( .A(n1201), .B(n1187), .Z(n1252) );
  XOR U2041 ( .A(n1270), .B(n1204), .Z(n1201) );
  XNOR U2042 ( .A(n1196), .B(n1198), .Z(n1204) );
  NAND U2043 ( .A(n572), .B(n1192), .Z(n1198) );
  XNOR U2044 ( .A(n1194), .B(n1271), .Z(n1196) );
  ANDN U2045 ( .A(n1199), .B(n574), .Z(n1271) );
  XOR U2046 ( .A(n1272), .B(n1273), .Z(n1194) );
  AND U2047 ( .A(n1274), .B(n1275), .Z(n1273) );
  XOR U2048 ( .A(n1276), .B(n1272), .Z(n1275) );
  XNOR U2049 ( .A(n1203), .B(n1200), .Z(n1270) );
  AND U2050 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U2051 ( .B(n1283), .A(n511), .Z(n1282) );
  NANDN U2052 ( .B(n1284), .A(n1285), .Z(n1281) );
  XNOR U2053 ( .A(n1212), .B(n1211), .Z(n1189) );
  XOR U2054 ( .A(n1289), .B(n1222), .Z(n1211) );
  XNOR U2055 ( .A(n1208), .B(n1209), .Z(n1222) );
  NANDN U2056 ( .B(n636), .A(n1000), .Z(n1209) );
  XNOR U2057 ( .A(n1207), .B(n1290), .Z(n1208) );
  ANDN U2058 ( .A(n677), .B(n1002), .Z(n1290) );
  XNOR U2059 ( .A(n1221), .B(n1210), .Z(n1289) );
  XOR U2060 ( .A(n1297), .B(n1217), .Z(n1221) );
  XNOR U2061 ( .A(n1215), .B(n1298), .Z(n1217) );
  ANDN U2062 ( .A(n784), .B(n867), .Z(n1298) );
  XOR U2063 ( .A(n1299), .B(n1300), .Z(n1215) );
  AND U2064 ( .A(n1301), .B(n1302), .Z(n1300) );
  XNOR U2065 ( .A(n1303), .B(n1299), .Z(n1302) );
  AND U2066 ( .A(n865), .B(n730), .Z(n1219) );
  XOR U2067 ( .A(n1232), .B(n1231), .Z(n1212) );
  XOR U2068 ( .A(n1307), .B(n1227), .Z(n1231) );
  XNOR U2069 ( .A(n1225), .B(n1308), .Z(n1227) );
  ANDN U2070 ( .A(n609), .B(n1154), .Z(n1308) );
  XOR U2071 ( .A(n1309), .B(n1310), .Z(n1225) );
  AND U2072 ( .A(n1311), .B(n1312), .Z(n1310) );
  XNOR U2073 ( .A(n1313), .B(n1309), .Z(n1312) );
  AND U2074 ( .A(n1152), .B(n568), .Z(n1229) );
  XOR U2075 ( .A(n1239), .B(n1238), .Z(n1232) );
  NAND U2076 ( .A(n1317), .B(n512), .Z(n1238) );
  XOR U2077 ( .A(n1237), .B(n1318), .Z(n1239) );
  ANDN U2078 ( .A(n543), .B(n1319), .Z(n1318) );
  ANDN U2079 ( .A(n1320), .B(n1321), .Z(n1237) );
  NAND U2080 ( .A(n1322), .B(n1323), .Z(n1320) );
  IV U2081 ( .A(n1240), .Z(n1241) );
  MUX U2082 ( .IN0(o[14]), .IN1(n411), .SEL(n464), .F(\_MxM/n292 ) );
  XOR U2083 ( .A(n1328), .B(\_MxM/Y0[15] ), .Z(n411) );
  XOR U2084 ( .A(n1329), .B(n1330), .Z(n1328) );
  AND U2085 ( .A(n476), .B(n1332), .Z(n1331) );
  XOR U2086 ( .A(n1326), .B(n1330), .Z(n1332) );
  XOR U2087 ( .A(n1325), .B(n1330), .Z(n1326) );
  XNOR U2088 ( .A(n1251), .B(n1250), .Z(n1330) );
  XOR U2089 ( .A(n1333), .B(n1334), .Z(n1250) );
  XOR U2090 ( .A(n1335), .B(n1336), .Z(n1334) );
  XOR U2091 ( .A(n1337), .B(n1335), .Z(n1336) );
  XNOR U2092 ( .A(n1343), .B(n1279), .Z(n1268) );
  XNOR U2093 ( .A(n1262), .B(n1261), .Z(n1279) );
  XOR U2094 ( .A(n1344), .B(n1257), .Z(n1261) );
  XNOR U2095 ( .A(n1255), .B(n1345), .Z(n1257) );
  ANDN U2096 ( .A(n1021), .B(n702), .Z(n1345) );
  AND U2097 ( .A(n700), .B(n958), .Z(n1259) );
  XNOR U2098 ( .A(n1265), .B(n1266), .Z(n1262) );
  NANDN U2099 ( .B(n823), .A(n801), .Z(n1266) );
  XNOR U2100 ( .A(n1264), .B(n1352), .Z(n1265) );
  ANDN U2101 ( .A(n893), .B(n803), .Z(n1352) );
  XOR U2102 ( .A(n1353), .B(n1354), .Z(n1264) );
  AND U2103 ( .A(n1355), .B(n1356), .Z(n1354) );
  XOR U2104 ( .A(n1357), .B(n1353), .Z(n1356) );
  XNOR U2105 ( .A(n1278), .B(n1267), .Z(n1343) );
  XOR U2106 ( .A(n1361), .B(n1288), .Z(n1278) );
  XNOR U2107 ( .A(n1274), .B(n1276), .Z(n1288) );
  NAND U2108 ( .A(n616), .B(n1192), .Z(n1276) );
  XNOR U2109 ( .A(n1272), .B(n1362), .Z(n1274) );
  ANDN U2110 ( .A(n1199), .B(n618), .Z(n1362) );
  XOR U2111 ( .A(n1363), .B(n1364), .Z(n1272) );
  AND U2112 ( .A(n1365), .B(n1366), .Z(n1364) );
  XOR U2113 ( .A(n1367), .B(n1363), .Z(n1366) );
  XNOR U2114 ( .A(n1287), .B(n1277), .Z(n1361) );
  XOR U2115 ( .A(n1375), .B(n1285), .Z(n1371) );
  AND U2116 ( .A(n541), .B(n1376), .Z(n1285) );
  NAND U2117 ( .A(n1377), .B(n1284), .Z(n1375) );
  XOR U2118 ( .A(n1378), .B(n1379), .Z(n1284) );
  AND U2119 ( .A(n1380), .B(n1381), .Z(n1379) );
  XNOR U2120 ( .A(n1382), .B(n1378), .Z(n1381) );
  NANDN U2121 ( .B(n544), .A(n1383), .Z(n1377) );
  XNOR U2122 ( .A(n1296), .B(n1295), .Z(n1269) );
  XOR U2123 ( .A(n1384), .B(n1306), .Z(n1295) );
  XNOR U2124 ( .A(n1292), .B(n1293), .Z(n1306) );
  NANDN U2125 ( .B(n636), .A(n1074), .Z(n1293) );
  XNOR U2126 ( .A(n1291), .B(n1385), .Z(n1292) );
  ANDN U2127 ( .A(n677), .B(n1076), .Z(n1385) );
  XNOR U2128 ( .A(n1305), .B(n1294), .Z(n1384) );
  XOR U2129 ( .A(n1392), .B(n1301), .Z(n1305) );
  XNOR U2130 ( .A(n1299), .B(n1393), .Z(n1301) );
  ANDN U2131 ( .A(n784), .B(n935), .Z(n1393) );
  AND U2132 ( .A(n933), .B(n730), .Z(n1303) );
  XOR U2133 ( .A(n1316), .B(n1315), .Z(n1296) );
  XOR U2134 ( .A(n1400), .B(n1311), .Z(n1315) );
  XNOR U2135 ( .A(n1309), .B(n1401), .Z(n1311) );
  ANDN U2136 ( .A(n609), .B(n1235), .Z(n1401) );
  AND U2137 ( .A(n1233), .B(n568), .Z(n1313) );
  XOR U2138 ( .A(n1323), .B(n1322), .Z(n1316) );
  NAND U2139 ( .A(n1408), .B(n512), .Z(n1322) );
  XNOR U2140 ( .A(n1321), .B(n1409), .Z(n1323) );
  ANDN U2141 ( .A(n543), .B(n1410), .Z(n1409) );
  NAND U2142 ( .A(n1411), .B(n1412), .Z(n1321) );
  NAND U2143 ( .A(n1413), .B(n1414), .Z(n1411) );
  IV U2144 ( .A(n1324), .Z(n1325) );
  MUX U2145 ( .IN0(o[13]), .IN1(n408), .SEL(n464), .F(\_MxM/n291 ) );
  XOR U2146 ( .A(n1419), .B(\_MxM/Y0[14] ), .Z(n408) );
  XOR U2147 ( .A(n1420), .B(n1421), .Z(n1419) );
  AND U2148 ( .A(n476), .B(n1423), .Z(n1422) );
  XOR U2149 ( .A(n1417), .B(n1421), .Z(n1423) );
  XOR U2150 ( .A(n1416), .B(n1421), .Z(n1417) );
  XOR U2151 ( .A(n1424), .B(n1338), .Z(n1341) );
  NAND U2152 ( .A(n1335), .B(n1428), .Z(n1339) );
  AND U2153 ( .A(n1429), .B(n1430), .Z(n1428) );
  NANDN U2154 ( .B(n1431), .A(n511), .Z(n1430) );
  NANDN U2155 ( .B(n1432), .A(n1433), .Z(n1429) );
  AND U2156 ( .A(n1434), .B(n1435), .Z(n1335) );
  NANDN U2157 ( .B(n1436), .A(n1437), .Z(n1435) );
  OR U2158 ( .A(n1438), .B(n1439), .Z(n1434) );
  XNOR U2159 ( .A(n1360), .B(n1359), .Z(n1342) );
  XOR U2160 ( .A(n1443), .B(n1370), .Z(n1359) );
  XNOR U2161 ( .A(n1351), .B(n1350), .Z(n1370) );
  XOR U2162 ( .A(n1444), .B(n1347), .Z(n1350) );
  XNOR U2163 ( .A(n1346), .B(n1445), .Z(n1347) );
  ANDN U2164 ( .A(n1021), .B(n744), .Z(n1445) );
  XOR U2165 ( .A(n1446), .B(n1447), .Z(n1346) );
  AND U2166 ( .A(n1448), .B(n1449), .Z(n1447) );
  XNOR U2167 ( .A(n1450), .B(n1446), .Z(n1449) );
  AND U2168 ( .A(n742), .B(n958), .Z(n1348) );
  XNOR U2169 ( .A(n1355), .B(n1357), .Z(n1351) );
  NANDN U2170 ( .B(n823), .A(n865), .Z(n1357) );
  XNOR U2171 ( .A(n1353), .B(n1454), .Z(n1355) );
  ANDN U2172 ( .A(n893), .B(n867), .Z(n1454) );
  XNOR U2173 ( .A(n1369), .B(n1358), .Z(n1443) );
  XOR U2174 ( .A(n1461), .B(n1374), .Z(n1369) );
  XNOR U2175 ( .A(n1365), .B(n1367), .Z(n1374) );
  NAND U2176 ( .A(n656), .B(n1192), .Z(n1367) );
  XNOR U2177 ( .A(n1363), .B(n1462), .Z(n1365) );
  ANDN U2178 ( .A(n1199), .B(n658), .Z(n1462) );
  XOR U2179 ( .A(n1463), .B(n1464), .Z(n1363) );
  AND U2180 ( .A(n1465), .B(n1466), .Z(n1464) );
  XOR U2181 ( .A(n1467), .B(n1463), .Z(n1466) );
  XNOR U2182 ( .A(n1373), .B(n1368), .Z(n1461) );
  XOR U2183 ( .A(n1471), .B(n1380), .Z(n1373) );
  XNOR U2184 ( .A(n1378), .B(n1472), .Z(n1380) );
  ANDN U2185 ( .A(n1383), .B(n574), .Z(n1472) );
  XOR U2186 ( .A(n1473), .B(n1474), .Z(n1378) );
  AND U2187 ( .A(n1475), .B(n1476), .Z(n1474) );
  XNOR U2188 ( .A(n1477), .B(n1473), .Z(n1476) );
  AND U2189 ( .A(n572), .B(n1376), .Z(n1382) );
  XNOR U2190 ( .A(n1391), .B(n1390), .Z(n1360) );
  XOR U2191 ( .A(n1481), .B(n1399), .Z(n1390) );
  XNOR U2192 ( .A(n1387), .B(n1388), .Z(n1399) );
  NANDN U2193 ( .B(n636), .A(n1152), .Z(n1388) );
  XNOR U2194 ( .A(n1386), .B(n1482), .Z(n1387) );
  ANDN U2195 ( .A(n677), .B(n1154), .Z(n1482) );
  XNOR U2196 ( .A(n1398), .B(n1389), .Z(n1481) );
  XOR U2197 ( .A(n1489), .B(n1395), .Z(n1398) );
  XNOR U2198 ( .A(n1394), .B(n1490), .Z(n1395) );
  ANDN U2199 ( .A(n784), .B(n1002), .Z(n1490) );
  AND U2200 ( .A(n1000), .B(n730), .Z(n1396) );
  XOR U2201 ( .A(n1407), .B(n1406), .Z(n1391) );
  XOR U2202 ( .A(n1497), .B(n1403), .Z(n1406) );
  XNOR U2203 ( .A(n1402), .B(n1498), .Z(n1403) );
  ANDN U2204 ( .A(n609), .B(n1319), .Z(n1498) );
  AND U2205 ( .A(n1317), .B(n568), .Z(n1404) );
  XOR U2206 ( .A(n1414), .B(n1413), .Z(n1407) );
  NAND U2207 ( .A(n1505), .B(n512), .Z(n1413) );
  XOR U2208 ( .A(n1412), .B(n1506), .Z(n1414) );
  ANDN U2209 ( .A(n543), .B(n1507), .Z(n1506) );
  ANDN U2210 ( .A(n1508), .B(n1509), .Z(n1412) );
  NAND U2211 ( .A(n1510), .B(n1511), .Z(n1508) );
  IV U2212 ( .A(n1415), .Z(n1416) );
  MUX U2213 ( .IN0(o[12]), .IN1(n405), .SEL(n464), .F(\_MxM/n290 ) );
  XOR U2214 ( .A(n1516), .B(\_MxM/Y0[13] ), .Z(n405) );
  XNOR U2215 ( .A(n1517), .B(n1518), .Z(n1516) );
  AND U2216 ( .A(n476), .B(n1520), .Z(n1519) );
  XNOR U2217 ( .A(n1514), .B(n1518), .Z(n1520) );
  XNOR U2218 ( .A(n1513), .B(n1518), .Z(n1514) );
  XNOR U2219 ( .A(n1442), .B(n1441), .Z(n1518) );
  XOR U2220 ( .A(n1521), .B(n1426), .Z(n1441) );
  NANDN U2221 ( .B(n1522), .A(n1523), .Z(n1432) );
  XOR U2222 ( .A(n1526), .B(n1439), .Z(n1436) );
  NAND U2223 ( .A(n1527), .B(n541), .Z(n1439) );
  NAND U2224 ( .A(n1528), .B(n1438), .Z(n1526) );
  NANDN U2225 ( .B(n544), .A(n1532), .Z(n1528) );
  XNOR U2226 ( .A(n1425), .B(n1440), .Z(n1521) );
  IV U2227 ( .A(n1427), .Z(n1425) );
  XNOR U2228 ( .A(n1460), .B(n1459), .Z(n1442) );
  XOR U2229 ( .A(n1539), .B(n1470), .Z(n1459) );
  XNOR U2230 ( .A(n1453), .B(n1452), .Z(n1470) );
  XOR U2231 ( .A(n1540), .B(n1448), .Z(n1452) );
  XNOR U2232 ( .A(n1446), .B(n1541), .Z(n1448) );
  ANDN U2233 ( .A(n1021), .B(n803), .Z(n1541) );
  XOR U2234 ( .A(n1542), .B(n1543), .Z(n1446) );
  AND U2235 ( .A(n1544), .B(n1545), .Z(n1543) );
  XNOR U2236 ( .A(n1546), .B(n1542), .Z(n1545) );
  AND U2237 ( .A(n801), .B(n958), .Z(n1450) );
  XNOR U2238 ( .A(n1456), .B(n1457), .Z(n1453) );
  NANDN U2239 ( .B(n823), .A(n933), .Z(n1457) );
  XNOR U2240 ( .A(n1455), .B(n1550), .Z(n1456) );
  ANDN U2241 ( .A(n893), .B(n935), .Z(n1550) );
  XNOR U2242 ( .A(n1469), .B(n1458), .Z(n1539) );
  XOR U2243 ( .A(n1557), .B(n1480), .Z(n1469) );
  XNOR U2244 ( .A(n1465), .B(n1467), .Z(n1480) );
  NAND U2245 ( .A(n700), .B(n1192), .Z(n1467) );
  XNOR U2246 ( .A(n1463), .B(n1558), .Z(n1465) );
  ANDN U2247 ( .A(n1199), .B(n702), .Z(n1558) );
  XOR U2248 ( .A(n1559), .B(n1560), .Z(n1463) );
  AND U2249 ( .A(n1561), .B(n1562), .Z(n1560) );
  XOR U2250 ( .A(n1563), .B(n1559), .Z(n1562) );
  XNOR U2251 ( .A(n1479), .B(n1468), .Z(n1557) );
  XOR U2252 ( .A(n1567), .B(n1475), .Z(n1479) );
  XNOR U2253 ( .A(n1473), .B(n1568), .Z(n1475) );
  ANDN U2254 ( .A(n1383), .B(n618), .Z(n1568) );
  XOR U2255 ( .A(n1569), .B(n1570), .Z(n1473) );
  AND U2256 ( .A(n1571), .B(n1572), .Z(n1570) );
  XNOR U2257 ( .A(n1573), .B(n1569), .Z(n1572) );
  AND U2258 ( .A(n616), .B(n1376), .Z(n1477) );
  XNOR U2259 ( .A(n1488), .B(n1487), .Z(n1460) );
  XOR U2260 ( .A(n1577), .B(n1496), .Z(n1487) );
  XNOR U2261 ( .A(n1484), .B(n1485), .Z(n1496) );
  NANDN U2262 ( .B(n636), .A(n1233), .Z(n1485) );
  XNOR U2263 ( .A(n1483), .B(n1578), .Z(n1484) );
  ANDN U2264 ( .A(n677), .B(n1235), .Z(n1578) );
  XNOR U2265 ( .A(n1495), .B(n1486), .Z(n1577) );
  XOR U2266 ( .A(n1585), .B(n1492), .Z(n1495) );
  XNOR U2267 ( .A(n1491), .B(n1586), .Z(n1492) );
  ANDN U2268 ( .A(n784), .B(n1076), .Z(n1586) );
  AND U2269 ( .A(n1074), .B(n730), .Z(n1493) );
  XOR U2270 ( .A(n1504), .B(n1503), .Z(n1488) );
  XOR U2271 ( .A(n1593), .B(n1500), .Z(n1503) );
  XNOR U2272 ( .A(n1499), .B(n1594), .Z(n1500) );
  ANDN U2273 ( .A(n609), .B(n1410), .Z(n1594) );
  AND U2274 ( .A(n1408), .B(n568), .Z(n1501) );
  XOR U2275 ( .A(n1511), .B(n1510), .Z(n1504) );
  NAND U2276 ( .A(n1601), .B(n512), .Z(n1510) );
  XNOR U2277 ( .A(n1509), .B(n1602), .Z(n1511) );
  ANDN U2278 ( .A(n543), .B(n1603), .Z(n1602) );
  NAND U2279 ( .A(n1604), .B(n1605), .Z(n1509) );
  NAND U2280 ( .A(n1606), .B(n1607), .Z(n1604) );
  IV U2281 ( .A(n1512), .Z(n1513) );
  MUX U2282 ( .IN0(o[11]), .IN1(n402), .SEL(n464), .F(\_MxM/n289 ) );
  XOR U2283 ( .A(n1612), .B(\_MxM/Y0[12] ), .Z(n402) );
  XOR U2284 ( .A(n1613), .B(n1614), .Z(n1612) );
  AND U2285 ( .A(n476), .B(n1616), .Z(n1615) );
  XOR U2286 ( .A(n1610), .B(n1614), .Z(n1616) );
  XOR U2287 ( .A(n1609), .B(n1614), .Z(n1610) );
  XNOR U2288 ( .A(n1617), .B(n1538), .Z(n1534) );
  XOR U2289 ( .A(n1523), .B(n1522), .Z(n1538) );
  NANDN U2290 ( .B(n1618), .A(n1619), .Z(n1522) );
  AND U2291 ( .A(n1621), .B(n1622), .Z(n1620) );
  NANDN U2292 ( .B(n1623), .A(n511), .Z(n1622) );
  NANDN U2293 ( .B(n1624), .A(n1625), .Z(n1621) );
  XNOR U2294 ( .A(n1530), .B(n1531), .Z(n1525) );
  NAND U2295 ( .A(n1527), .B(n572), .Z(n1531) );
  XNOR U2296 ( .A(n1529), .B(n1629), .Z(n1530) );
  ANDN U2297 ( .A(n1532), .B(n574), .Z(n1629) );
  XNOR U2298 ( .A(n1537), .B(n1533), .Z(n1617) );
  IV U2299 ( .A(n1536), .Z(n1537) );
  XNOR U2300 ( .A(n1556), .B(n1555), .Z(n1535) );
  XOR U2301 ( .A(n1639), .B(n1566), .Z(n1555) );
  XNOR U2302 ( .A(n1549), .B(n1548), .Z(n1566) );
  XOR U2303 ( .A(n1640), .B(n1544), .Z(n1548) );
  XNOR U2304 ( .A(n1542), .B(n1641), .Z(n1544) );
  ANDN U2305 ( .A(n1021), .B(n867), .Z(n1641) );
  AND U2306 ( .A(n865), .B(n958), .Z(n1546) );
  XNOR U2307 ( .A(n1552), .B(n1553), .Z(n1549) );
  NANDN U2308 ( .B(n823), .A(n1000), .Z(n1553) );
  XNOR U2309 ( .A(n1551), .B(n1648), .Z(n1552) );
  ANDN U2310 ( .A(n893), .B(n1002), .Z(n1648) );
  XNOR U2311 ( .A(n1565), .B(n1554), .Z(n1639) );
  XOR U2312 ( .A(n1655), .B(n1576), .Z(n1565) );
  XNOR U2313 ( .A(n1561), .B(n1563), .Z(n1576) );
  NAND U2314 ( .A(n742), .B(n1192), .Z(n1563) );
  XNOR U2315 ( .A(n1559), .B(n1656), .Z(n1561) );
  ANDN U2316 ( .A(n1199), .B(n744), .Z(n1656) );
  XNOR U2317 ( .A(n1575), .B(n1564), .Z(n1655) );
  XOR U2318 ( .A(n1663), .B(n1571), .Z(n1575) );
  XNOR U2319 ( .A(n1569), .B(n1664), .Z(n1571) );
  ANDN U2320 ( .A(n1383), .B(n658), .Z(n1664) );
  XOR U2321 ( .A(n1665), .B(n1666), .Z(n1569) );
  AND U2322 ( .A(n1667), .B(n1668), .Z(n1666) );
  XNOR U2323 ( .A(n1669), .B(n1665), .Z(n1668) );
  AND U2324 ( .A(n656), .B(n1376), .Z(n1573) );
  XNOR U2325 ( .A(n1584), .B(n1583), .Z(n1556) );
  XOR U2326 ( .A(n1673), .B(n1592), .Z(n1583) );
  XNOR U2327 ( .A(n1580), .B(n1581), .Z(n1592) );
  NANDN U2328 ( .B(n636), .A(n1317), .Z(n1581) );
  XNOR U2329 ( .A(n1579), .B(n1674), .Z(n1580) );
  ANDN U2330 ( .A(n677), .B(n1319), .Z(n1674) );
  XNOR U2331 ( .A(n1591), .B(n1582), .Z(n1673) );
  XOR U2332 ( .A(n1681), .B(n1588), .Z(n1591) );
  XNOR U2333 ( .A(n1587), .B(n1682), .Z(n1588) );
  ANDN U2334 ( .A(n784), .B(n1154), .Z(n1682) );
  AND U2335 ( .A(n1152), .B(n730), .Z(n1589) );
  XOR U2336 ( .A(n1600), .B(n1599), .Z(n1584) );
  XOR U2337 ( .A(n1689), .B(n1596), .Z(n1599) );
  XNOR U2338 ( .A(n1595), .B(n1690), .Z(n1596) );
  ANDN U2339 ( .A(n609), .B(n1507), .Z(n1690) );
  AND U2340 ( .A(n1505), .B(n568), .Z(n1597) );
  XOR U2341 ( .A(n1607), .B(n1606), .Z(n1600) );
  NAND U2342 ( .A(n1697), .B(n512), .Z(n1606) );
  XOR U2343 ( .A(n1605), .B(n1698), .Z(n1607) );
  ANDN U2344 ( .A(n543), .B(n1699), .Z(n1698) );
  ANDN U2345 ( .A(n1700), .B(n1701), .Z(n1605) );
  NAND U2346 ( .A(n1702), .B(n1703), .Z(n1700) );
  IV U2347 ( .A(n1608), .Z(n1609) );
  MUX U2348 ( .IN0(o[10]), .IN1(n399), .SEL(n464), .F(\_MxM/n288 ) );
  XOR U2349 ( .A(n1708), .B(\_MxM/Y0[11] ), .Z(n399) );
  XNOR U2350 ( .A(n1709), .B(n1710), .Z(n1708) );
  AND U2351 ( .A(n476), .B(n1712), .Z(n1711) );
  XNOR U2352 ( .A(n1706), .B(n1710), .Z(n1712) );
  XNOR U2353 ( .A(n1705), .B(n1710), .Z(n1706) );
  XNOR U2354 ( .A(n1635), .B(n1634), .Z(n1710) );
  XOR U2355 ( .A(n1713), .B(n1638), .Z(n1634) );
  XOR U2356 ( .A(n1628), .B(n1627), .Z(n1618) );
  XOR U2357 ( .A(n1721), .B(n1625), .Z(n1717) );
  AND U2358 ( .A(n1722), .B(n541), .Z(n1625) );
  NAND U2359 ( .A(n1723), .B(n1624), .Z(n1721) );
  XOR U2360 ( .A(n1724), .B(n1725), .Z(n1624) );
  AND U2361 ( .A(n1726), .B(n1727), .Z(n1725) );
  XNOR U2362 ( .A(n1728), .B(n1724), .Z(n1727) );
  NANDN U2363 ( .B(n544), .A(n1729), .Z(n1723) );
  XNOR U2364 ( .A(n1631), .B(n1632), .Z(n1628) );
  NAND U2365 ( .A(n1527), .B(n616), .Z(n1632) );
  XNOR U2366 ( .A(n1630), .B(n1730), .Z(n1631) );
  ANDN U2367 ( .A(n1532), .B(n618), .Z(n1730) );
  XNOR U2368 ( .A(n1637), .B(n1633), .Z(n1713) );
  IV U2369 ( .A(n1636), .Z(n1637) );
  XNOR U2370 ( .A(n1654), .B(n1653), .Z(n1635) );
  XOR U2371 ( .A(n1740), .B(n1662), .Z(n1653) );
  XNOR U2372 ( .A(n1647), .B(n1646), .Z(n1662) );
  XOR U2373 ( .A(n1741), .B(n1643), .Z(n1646) );
  XNOR U2374 ( .A(n1642), .B(n1742), .Z(n1643) );
  ANDN U2375 ( .A(n1021), .B(n935), .Z(n1742) );
  AND U2376 ( .A(n933), .B(n958), .Z(n1644) );
  XNOR U2377 ( .A(n1650), .B(n1651), .Z(n1647) );
  NANDN U2378 ( .B(n823), .A(n1074), .Z(n1651) );
  XNOR U2379 ( .A(n1649), .B(n1749), .Z(n1650) );
  ANDN U2380 ( .A(n893), .B(n1076), .Z(n1749) );
  XNOR U2381 ( .A(n1661), .B(n1652), .Z(n1740) );
  XOR U2382 ( .A(n1756), .B(n1672), .Z(n1661) );
  XNOR U2383 ( .A(n1658), .B(n1659), .Z(n1672) );
  NAND U2384 ( .A(n801), .B(n1192), .Z(n1659) );
  XNOR U2385 ( .A(n1657), .B(n1757), .Z(n1658) );
  ANDN U2386 ( .A(n1199), .B(n803), .Z(n1757) );
  XNOR U2387 ( .A(n1671), .B(n1660), .Z(n1756) );
  XOR U2388 ( .A(n1764), .B(n1667), .Z(n1671) );
  XNOR U2389 ( .A(n1665), .B(n1765), .Z(n1667) );
  ANDN U2390 ( .A(n1383), .B(n702), .Z(n1765) );
  XOR U2391 ( .A(n1766), .B(n1767), .Z(n1665) );
  AND U2392 ( .A(n1768), .B(n1769), .Z(n1767) );
  XNOR U2393 ( .A(n1770), .B(n1766), .Z(n1769) );
  AND U2394 ( .A(n700), .B(n1376), .Z(n1669) );
  XNOR U2395 ( .A(n1680), .B(n1679), .Z(n1654) );
  XOR U2396 ( .A(n1774), .B(n1688), .Z(n1679) );
  XNOR U2397 ( .A(n1676), .B(n1677), .Z(n1688) );
  NANDN U2398 ( .B(n636), .A(n1408), .Z(n1677) );
  XNOR U2399 ( .A(n1675), .B(n1775), .Z(n1676) );
  ANDN U2400 ( .A(n677), .B(n1410), .Z(n1775) );
  XNOR U2401 ( .A(n1687), .B(n1678), .Z(n1774) );
  XOR U2402 ( .A(n1782), .B(n1684), .Z(n1687) );
  XNOR U2403 ( .A(n1683), .B(n1783), .Z(n1684) );
  ANDN U2404 ( .A(n784), .B(n1235), .Z(n1783) );
  AND U2405 ( .A(n1233), .B(n730), .Z(n1685) );
  XOR U2406 ( .A(n1696), .B(n1695), .Z(n1680) );
  XOR U2407 ( .A(n1790), .B(n1692), .Z(n1695) );
  XNOR U2408 ( .A(n1691), .B(n1791), .Z(n1692) );
  ANDN U2409 ( .A(n609), .B(n1603), .Z(n1791) );
  AND U2410 ( .A(n1601), .B(n568), .Z(n1693) );
  XOR U2411 ( .A(n1703), .B(n1702), .Z(n1696) );
  NAND U2412 ( .A(n1798), .B(n512), .Z(n1702) );
  XNOR U2413 ( .A(n1701), .B(n1799), .Z(n1703) );
  ANDN U2414 ( .A(n543), .B(n1800), .Z(n1799) );
  NAND U2415 ( .A(n1801), .B(n1802), .Z(n1701) );
  NAND U2416 ( .A(n1803), .B(n1804), .Z(n1801) );
  IV U2417 ( .A(n1704), .Z(n1705) );
  MUX U2418 ( .IN0(o[9]), .IN1(n396), .SEL(n464), .F(\_MxM/n287 ) );
  XOR U2419 ( .A(n1809), .B(\_MxM/Y0[10] ), .Z(n396) );
  XOR U2420 ( .A(n1810), .B(n1811), .Z(n1809) );
  AND U2421 ( .A(n476), .B(n1813), .Z(n1812) );
  XOR U2422 ( .A(n1807), .B(n1811), .Z(n1813) );
  XOR U2423 ( .A(n1806), .B(n1811), .Z(n1807) );
  XNOR U2424 ( .A(n1814), .B(n1739), .Z(n1735) );
  XNOR U2425 ( .A(n1716), .B(n1715), .Z(n1739) );
  XOR U2426 ( .A(n1714), .B(n1815), .Z(n1715) );
  AND U2427 ( .A(n1816), .B(n1817), .Z(n1815) );
  NANDN U2428 ( .B(n1818), .A(n1819), .Z(n1817) );
  AND U2429 ( .A(n1820), .B(n1821), .Z(n1816) );
  NANDN U2430 ( .B(n1822), .A(n511), .Z(n1821) );
  OR U2431 ( .A(n1823), .B(n1824), .Z(n1820) );
  XNOR U2432 ( .A(n1720), .B(n1719), .Z(n1716) );
  XOR U2433 ( .A(n1828), .B(n1726), .Z(n1719) );
  XNOR U2434 ( .A(n1724), .B(n1829), .Z(n1726) );
  ANDN U2435 ( .A(n1729), .B(n574), .Z(n1829) );
  XOR U2436 ( .A(n1830), .B(n1831), .Z(n1724) );
  AND U2437 ( .A(n1832), .B(n1833), .Z(n1831) );
  XNOR U2438 ( .A(n1834), .B(n1830), .Z(n1833) );
  AND U2439 ( .A(n1722), .B(n572), .Z(n1728) );
  XNOR U2440 ( .A(n1732), .B(n1733), .Z(n1720) );
  NAND U2441 ( .A(n1527), .B(n656), .Z(n1733) );
  XNOR U2442 ( .A(n1731), .B(n1838), .Z(n1732) );
  ANDN U2443 ( .A(n1532), .B(n658), .Z(n1838) );
  XNOR U2444 ( .A(n1738), .B(n1734), .Z(n1814) );
  IV U2445 ( .A(n1737), .Z(n1738) );
  XNOR U2446 ( .A(n1755), .B(n1754), .Z(n1736) );
  XOR U2447 ( .A(n1848), .B(n1763), .Z(n1754) );
  XNOR U2448 ( .A(n1748), .B(n1747), .Z(n1763) );
  XOR U2449 ( .A(n1849), .B(n1744), .Z(n1747) );
  XNOR U2450 ( .A(n1743), .B(n1850), .Z(n1744) );
  ANDN U2451 ( .A(n1021), .B(n1002), .Z(n1850) );
  AND U2452 ( .A(n1000), .B(n958), .Z(n1745) );
  XNOR U2453 ( .A(n1751), .B(n1752), .Z(n1748) );
  NANDN U2454 ( .B(n823), .A(n1152), .Z(n1752) );
  XNOR U2455 ( .A(n1750), .B(n1857), .Z(n1751) );
  ANDN U2456 ( .A(n893), .B(n1154), .Z(n1857) );
  XNOR U2457 ( .A(n1762), .B(n1753), .Z(n1848) );
  XOR U2458 ( .A(n1864), .B(n1773), .Z(n1762) );
  XNOR U2459 ( .A(n1759), .B(n1760), .Z(n1773) );
  NAND U2460 ( .A(n865), .B(n1192), .Z(n1760) );
  XNOR U2461 ( .A(n1758), .B(n1865), .Z(n1759) );
  ANDN U2462 ( .A(n1199), .B(n867), .Z(n1865) );
  XNOR U2463 ( .A(n1772), .B(n1761), .Z(n1864) );
  XOR U2464 ( .A(n1872), .B(n1768), .Z(n1772) );
  XNOR U2465 ( .A(n1766), .B(n1873), .Z(n1768) );
  ANDN U2466 ( .A(n1383), .B(n744), .Z(n1873) );
  AND U2467 ( .A(n742), .B(n1376), .Z(n1770) );
  XNOR U2468 ( .A(n1781), .B(n1780), .Z(n1755) );
  XOR U2469 ( .A(n1880), .B(n1789), .Z(n1780) );
  XNOR U2470 ( .A(n1777), .B(n1778), .Z(n1789) );
  NANDN U2471 ( .B(n636), .A(n1505), .Z(n1778) );
  XNOR U2472 ( .A(n1776), .B(n1881), .Z(n1777) );
  ANDN U2473 ( .A(n677), .B(n1507), .Z(n1881) );
  XNOR U2474 ( .A(n1788), .B(n1779), .Z(n1880) );
  XOR U2475 ( .A(n1888), .B(n1785), .Z(n1788) );
  XNOR U2476 ( .A(n1784), .B(n1889), .Z(n1785) );
  ANDN U2477 ( .A(n784), .B(n1319), .Z(n1889) );
  AND U2478 ( .A(n1317), .B(n730), .Z(n1786) );
  XOR U2479 ( .A(n1797), .B(n1796), .Z(n1781) );
  XOR U2480 ( .A(n1896), .B(n1793), .Z(n1796) );
  XNOR U2481 ( .A(n1792), .B(n1897), .Z(n1793) );
  ANDN U2482 ( .A(n609), .B(n1699), .Z(n1897) );
  AND U2483 ( .A(n1697), .B(n568), .Z(n1794) );
  XOR U2484 ( .A(n1804), .B(n1803), .Z(n1797) );
  NAND U2485 ( .A(n1904), .B(n512), .Z(n1803) );
  XOR U2486 ( .A(n1802), .B(n1905), .Z(n1804) );
  ANDN U2487 ( .A(n543), .B(n1906), .Z(n1905) );
  ANDN U2488 ( .A(n1907), .B(n1908), .Z(n1802) );
  NAND U2489 ( .A(n1909), .B(n1910), .Z(n1907) );
  IV U2490 ( .A(n1805), .Z(n1806) );
  MUX U2491 ( .IN0(o[8]), .IN1(n393), .SEL(n464), .F(\_MxM/n286 ) );
  XOR U2492 ( .A(n1915), .B(\_MxM/Y0[9] ), .Z(n393) );
  XOR U2493 ( .A(n1916), .B(n1917), .Z(n1915) );
  AND U2494 ( .A(n476), .B(n1919), .Z(n1918) );
  XOR U2495 ( .A(n1913), .B(n1917), .Z(n1919) );
  XOR U2496 ( .A(n1912), .B(n1917), .Z(n1913) );
  XNOR U2497 ( .A(n1920), .B(n1847), .Z(n1843) );
  XNOR U2498 ( .A(n1827), .B(n1826), .Z(n1847) );
  XOR U2499 ( .A(n1921), .B(n1823), .Z(n1826) );
  XNOR U2500 ( .A(n1922), .B(n1819), .Z(n1823) );
  AND U2501 ( .A(n1923), .B(n541), .Z(n1819) );
  NAND U2502 ( .A(n1924), .B(n1818), .Z(n1922) );
  NANDN U2503 ( .B(n544), .A(n1928), .Z(n1924) );
  XNOR U2504 ( .A(n1824), .B(n1825), .Z(n1921) );
  XNOR U2505 ( .A(n1932), .B(n1935), .Z(n1934) );
  XNOR U2506 ( .A(n1837), .B(n1836), .Z(n1827) );
  XOR U2507 ( .A(n1936), .B(n1832), .Z(n1836) );
  XNOR U2508 ( .A(n1830), .B(n1937), .Z(n1832) );
  ANDN U2509 ( .A(n1729), .B(n618), .Z(n1937) );
  XOR U2510 ( .A(n1938), .B(n1939), .Z(n1830) );
  AND U2511 ( .A(n1940), .B(n1941), .Z(n1939) );
  XNOR U2512 ( .A(n1942), .B(n1938), .Z(n1941) );
  AND U2513 ( .A(n1722), .B(n616), .Z(n1834) );
  XNOR U2514 ( .A(n1840), .B(n1841), .Z(n1837) );
  NAND U2515 ( .A(n1527), .B(n700), .Z(n1841) );
  XNOR U2516 ( .A(n1839), .B(n1946), .Z(n1840) );
  ANDN U2517 ( .A(n1532), .B(n702), .Z(n1946) );
  XNOR U2518 ( .A(n1846), .B(n1842), .Z(n1920) );
  IV U2519 ( .A(n1845), .Z(n1846) );
  XNOR U2520 ( .A(n1863), .B(n1862), .Z(n1844) );
  XOR U2521 ( .A(n1955), .B(n1871), .Z(n1862) );
  XNOR U2522 ( .A(n1856), .B(n1855), .Z(n1871) );
  XOR U2523 ( .A(n1956), .B(n1852), .Z(n1855) );
  XNOR U2524 ( .A(n1851), .B(n1957), .Z(n1852) );
  ANDN U2525 ( .A(n1021), .B(n1076), .Z(n1957) );
  AND U2526 ( .A(n1074), .B(n958), .Z(n1853) );
  XNOR U2527 ( .A(n1859), .B(n1860), .Z(n1856) );
  NANDN U2528 ( .B(n823), .A(n1233), .Z(n1860) );
  XNOR U2529 ( .A(n1858), .B(n1964), .Z(n1859) );
  ANDN U2530 ( .A(n893), .B(n1235), .Z(n1964) );
  XNOR U2531 ( .A(n1870), .B(n1861), .Z(n1955) );
  XOR U2532 ( .A(n1971), .B(n1879), .Z(n1870) );
  XNOR U2533 ( .A(n1867), .B(n1868), .Z(n1879) );
  NAND U2534 ( .A(n933), .B(n1192), .Z(n1868) );
  XNOR U2535 ( .A(n1866), .B(n1972), .Z(n1867) );
  ANDN U2536 ( .A(n1199), .B(n935), .Z(n1972) );
  XNOR U2537 ( .A(n1878), .B(n1869), .Z(n1971) );
  XOR U2538 ( .A(n1979), .B(n1875), .Z(n1878) );
  XNOR U2539 ( .A(n1874), .B(n1980), .Z(n1875) );
  ANDN U2540 ( .A(n1383), .B(n803), .Z(n1980) );
  AND U2541 ( .A(n801), .B(n1376), .Z(n1876) );
  XNOR U2542 ( .A(n1887), .B(n1886), .Z(n1863) );
  XOR U2543 ( .A(n1987), .B(n1895), .Z(n1886) );
  XNOR U2544 ( .A(n1883), .B(n1884), .Z(n1895) );
  NANDN U2545 ( .B(n636), .A(n1601), .Z(n1884) );
  XNOR U2546 ( .A(n1882), .B(n1988), .Z(n1883) );
  ANDN U2547 ( .A(n677), .B(n1603), .Z(n1988) );
  XNOR U2548 ( .A(n1894), .B(n1885), .Z(n1987) );
  XOR U2549 ( .A(n1995), .B(n1891), .Z(n1894) );
  XNOR U2550 ( .A(n1890), .B(n1996), .Z(n1891) );
  ANDN U2551 ( .A(n784), .B(n1410), .Z(n1996) );
  AND U2552 ( .A(n1408), .B(n730), .Z(n1892) );
  XOR U2553 ( .A(n1903), .B(n1902), .Z(n1887) );
  XOR U2554 ( .A(n2003), .B(n1899), .Z(n1902) );
  XNOR U2555 ( .A(n1898), .B(n2004), .Z(n1899) );
  ANDN U2556 ( .A(n609), .B(n1800), .Z(n2004) );
  AND U2557 ( .A(n1798), .B(n568), .Z(n1900) );
  XOR U2558 ( .A(n1910), .B(n1909), .Z(n1903) );
  NAND U2559 ( .A(n2011), .B(n512), .Z(n1909) );
  XNOR U2560 ( .A(n1908), .B(n2012), .Z(n1910) );
  ANDN U2561 ( .A(n543), .B(n2013), .Z(n2012) );
  NAND U2562 ( .A(n2014), .B(n2015), .Z(n1908) );
  NAND U2563 ( .A(n2016), .B(n2017), .Z(n2014) );
  IV U2564 ( .A(n1911), .Z(n1912) );
  MUX U2565 ( .IN0(o[7]), .IN1(n390), .SEL(n464), .F(\_MxM/n285 ) );
  XOR U2566 ( .A(n2022), .B(\_MxM/Y0[8] ), .Z(n390) );
  XOR U2567 ( .A(n2023), .B(n2024), .Z(n2022) );
  AND U2568 ( .A(n476), .B(n2026), .Z(n2025) );
  XOR U2569 ( .A(n2020), .B(n2024), .Z(n2026) );
  XOR U2570 ( .A(n2019), .B(n2024), .Z(n2020) );
  XNOR U2571 ( .A(n2027), .B(n1954), .Z(n1951) );
  XNOR U2572 ( .A(n1931), .B(n1930), .Z(n1954) );
  XOR U2573 ( .A(n2028), .B(n1935), .Z(n1930) );
  XNOR U2574 ( .A(n1926), .B(n1927), .Z(n1935) );
  NAND U2575 ( .A(n1923), .B(n572), .Z(n1927) );
  XNOR U2576 ( .A(n1925), .B(n2029), .Z(n1926) );
  ANDN U2577 ( .A(n1928), .B(n574), .Z(n2029) );
  XNOR U2578 ( .A(n1933), .B(n1929), .Z(n2028) );
  XOR U2579 ( .A(n1932), .B(n2036), .Z(n1933) );
  AND U2580 ( .A(n2037), .B(n2038), .Z(n2036) );
  NANDN U2581 ( .B(n2039), .A(n511), .Z(n2038) );
  NANDN U2582 ( .B(n2040), .A(n2041), .Z(n2037) );
  XNOR U2583 ( .A(n1945), .B(n1944), .Z(n1931) );
  XOR U2584 ( .A(n2045), .B(n1940), .Z(n1944) );
  XNOR U2585 ( .A(n1938), .B(n2046), .Z(n1940) );
  ANDN U2586 ( .A(n1729), .B(n658), .Z(n2046) );
  AND U2587 ( .A(n1722), .B(n656), .Z(n1942) );
  XNOR U2588 ( .A(n1948), .B(n1949), .Z(n1945) );
  NAND U2589 ( .A(n1527), .B(n742), .Z(n1949) );
  XNOR U2590 ( .A(n1947), .B(n2053), .Z(n1948) );
  ANDN U2591 ( .A(n1532), .B(n744), .Z(n2053) );
  XNOR U2592 ( .A(n1970), .B(n1969), .Z(n1952) );
  XOR U2593 ( .A(n2063), .B(n1978), .Z(n1969) );
  XNOR U2594 ( .A(n1963), .B(n1962), .Z(n1978) );
  XOR U2595 ( .A(n2064), .B(n1959), .Z(n1962) );
  XNOR U2596 ( .A(n1958), .B(n2065), .Z(n1959) );
  ANDN U2597 ( .A(n1021), .B(n1154), .Z(n2065) );
  AND U2598 ( .A(n1152), .B(n958), .Z(n1960) );
  XNOR U2599 ( .A(n1966), .B(n1967), .Z(n1963) );
  NANDN U2600 ( .B(n823), .A(n1317), .Z(n1967) );
  XNOR U2601 ( .A(n1965), .B(n2072), .Z(n1966) );
  ANDN U2602 ( .A(n893), .B(n1319), .Z(n2072) );
  XNOR U2603 ( .A(n1977), .B(n1968), .Z(n2063) );
  XOR U2604 ( .A(n2079), .B(n1986), .Z(n1977) );
  XNOR U2605 ( .A(n1974), .B(n1975), .Z(n1986) );
  NAND U2606 ( .A(n1000), .B(n1192), .Z(n1975) );
  XNOR U2607 ( .A(n1973), .B(n2080), .Z(n1974) );
  ANDN U2608 ( .A(n1199), .B(n1002), .Z(n2080) );
  XNOR U2609 ( .A(n1985), .B(n1976), .Z(n2079) );
  XOR U2610 ( .A(n2087), .B(n1982), .Z(n1985) );
  XNOR U2611 ( .A(n1981), .B(n2088), .Z(n1982) );
  ANDN U2612 ( .A(n1383), .B(n867), .Z(n2088) );
  AND U2613 ( .A(n865), .B(n1376), .Z(n1983) );
  XNOR U2614 ( .A(n1994), .B(n1993), .Z(n1970) );
  XOR U2615 ( .A(n2095), .B(n2002), .Z(n1993) );
  XNOR U2616 ( .A(n1990), .B(n1991), .Z(n2002) );
  NANDN U2617 ( .B(n636), .A(n1697), .Z(n1991) );
  XNOR U2618 ( .A(n1989), .B(n2096), .Z(n1990) );
  ANDN U2619 ( .A(n677), .B(n1699), .Z(n2096) );
  XNOR U2620 ( .A(n2001), .B(n1992), .Z(n2095) );
  XOR U2621 ( .A(n2103), .B(n1998), .Z(n2001) );
  XNOR U2622 ( .A(n1997), .B(n2104), .Z(n1998) );
  ANDN U2623 ( .A(n784), .B(n1507), .Z(n2104) );
  AND U2624 ( .A(n1505), .B(n730), .Z(n1999) );
  XOR U2625 ( .A(n2010), .B(n2009), .Z(n1994) );
  XOR U2626 ( .A(n2111), .B(n2006), .Z(n2009) );
  XNOR U2627 ( .A(n2005), .B(n2112), .Z(n2006) );
  ANDN U2628 ( .A(n609), .B(n1906), .Z(n2112) );
  AND U2629 ( .A(n1904), .B(n568), .Z(n2007) );
  XOR U2630 ( .A(n2017), .B(n2016), .Z(n2010) );
  NAND U2631 ( .A(n2119), .B(n512), .Z(n2016) );
  XOR U2632 ( .A(n2015), .B(n2120), .Z(n2017) );
  ANDN U2633 ( .A(n543), .B(n2121), .Z(n2120) );
  ANDN U2634 ( .A(n2122), .B(n2123), .Z(n2015) );
  NAND U2635 ( .A(n2124), .B(n2125), .Z(n2122) );
  IV U2636 ( .A(n2018), .Z(n2019) );
  MUX U2637 ( .IN0(o[6]), .IN1(n387), .SEL(n464), .F(\_MxM/n284 ) );
  XOR U2638 ( .A(n2130), .B(\_MxM/Y0[7] ), .Z(n387) );
  XOR U2639 ( .A(n2131), .B(n2132), .Z(n2130) );
  AND U2640 ( .A(n476), .B(n2134), .Z(n2133) );
  XOR U2641 ( .A(n2128), .B(n2132), .Z(n2134) );
  XOR U2642 ( .A(n2127), .B(n2132), .Z(n2128) );
  XNOR U2643 ( .A(n2135), .B(n2062), .Z(n2058) );
  XNOR U2644 ( .A(n2035), .B(n2034), .Z(n2062) );
  XOR U2645 ( .A(n2136), .B(n2044), .Z(n2034) );
  XNOR U2646 ( .A(n2031), .B(n2032), .Z(n2044) );
  NAND U2647 ( .A(n1923), .B(n616), .Z(n2032) );
  XNOR U2648 ( .A(n2030), .B(n2137), .Z(n2031) );
  ANDN U2649 ( .A(n1928), .B(n618), .Z(n2137) );
  XOR U2650 ( .A(n2138), .B(n2139), .Z(n2030) );
  AND U2651 ( .A(n2140), .B(n2141), .Z(n2139) );
  XOR U2652 ( .A(n2142), .B(n2138), .Z(n2141) );
  XNOR U2653 ( .A(n2043), .B(n2033), .Z(n2136) );
  XOR U2654 ( .A(n2150), .B(n2041), .Z(n2146) );
  AND U2655 ( .A(n2151), .B(n541), .Z(n2041) );
  NAND U2656 ( .A(n2152), .B(n2040), .Z(n2150) );
  XOR U2657 ( .A(n2153), .B(n2154), .Z(n2040) );
  AND U2658 ( .A(n2155), .B(n2156), .Z(n2154) );
  XNOR U2659 ( .A(n2157), .B(n2153), .Z(n2156) );
  NANDN U2660 ( .B(n544), .A(n2158), .Z(n2152) );
  XNOR U2661 ( .A(n2052), .B(n2051), .Z(n2035) );
  XOR U2662 ( .A(n2159), .B(n2048), .Z(n2051) );
  XNOR U2663 ( .A(n2047), .B(n2160), .Z(n2048) );
  ANDN U2664 ( .A(n1729), .B(n702), .Z(n2160) );
  AND U2665 ( .A(n1722), .B(n700), .Z(n2049) );
  XNOR U2666 ( .A(n2055), .B(n2056), .Z(n2052) );
  NAND U2667 ( .A(n1527), .B(n801), .Z(n2056) );
  XNOR U2668 ( .A(n2054), .B(n2167), .Z(n2055) );
  ANDN U2669 ( .A(n1532), .B(n803), .Z(n2167) );
  XNOR U2670 ( .A(n2061), .B(n2057), .Z(n2135) );
  XOR U2671 ( .A(n2178), .B(n2179), .Z(n2174) );
  NANDN U2672 ( .B(n2180), .A(n2181), .Z(n2178) );
  XNOR U2673 ( .A(n2078), .B(n2077), .Z(n2059) );
  XOR U2674 ( .A(n2182), .B(n2086), .Z(n2077) );
  XNOR U2675 ( .A(n2071), .B(n2070), .Z(n2086) );
  XOR U2676 ( .A(n2183), .B(n2067), .Z(n2070) );
  XNOR U2677 ( .A(n2066), .B(n2184), .Z(n2067) );
  ANDN U2678 ( .A(n1021), .B(n1235), .Z(n2184) );
  AND U2679 ( .A(n1233), .B(n958), .Z(n2068) );
  XNOR U2680 ( .A(n2074), .B(n2075), .Z(n2071) );
  NANDN U2681 ( .B(n823), .A(n1408), .Z(n2075) );
  XNOR U2682 ( .A(n2073), .B(n2191), .Z(n2074) );
  ANDN U2683 ( .A(n893), .B(n1410), .Z(n2191) );
  XNOR U2684 ( .A(n2085), .B(n2076), .Z(n2182) );
  XOR U2685 ( .A(n2198), .B(n2094), .Z(n2085) );
  XNOR U2686 ( .A(n2082), .B(n2083), .Z(n2094) );
  NAND U2687 ( .A(n1074), .B(n1192), .Z(n2083) );
  XNOR U2688 ( .A(n2081), .B(n2199), .Z(n2082) );
  ANDN U2689 ( .A(n1199), .B(n1076), .Z(n2199) );
  XNOR U2690 ( .A(n2093), .B(n2084), .Z(n2198) );
  XOR U2691 ( .A(n2206), .B(n2090), .Z(n2093) );
  XNOR U2692 ( .A(n2089), .B(n2207), .Z(n2090) );
  ANDN U2693 ( .A(n1383), .B(n935), .Z(n2207) );
  AND U2694 ( .A(n933), .B(n1376), .Z(n2091) );
  XNOR U2695 ( .A(n2102), .B(n2101), .Z(n2078) );
  XOR U2696 ( .A(n2214), .B(n2110), .Z(n2101) );
  XNOR U2697 ( .A(n2098), .B(n2099), .Z(n2110) );
  NANDN U2698 ( .B(n636), .A(n1798), .Z(n2099) );
  XNOR U2699 ( .A(n2097), .B(n2215), .Z(n2098) );
  ANDN U2700 ( .A(n677), .B(n1800), .Z(n2215) );
  XNOR U2701 ( .A(n2109), .B(n2100), .Z(n2214) );
  XOR U2702 ( .A(n2222), .B(n2106), .Z(n2109) );
  XNOR U2703 ( .A(n2105), .B(n2223), .Z(n2106) );
  ANDN U2704 ( .A(n784), .B(n1603), .Z(n2223) );
  AND U2705 ( .A(n1601), .B(n730), .Z(n2107) );
  XOR U2706 ( .A(n2118), .B(n2117), .Z(n2102) );
  XOR U2707 ( .A(n2230), .B(n2114), .Z(n2117) );
  XNOR U2708 ( .A(n2113), .B(n2231), .Z(n2114) );
  ANDN U2709 ( .A(n609), .B(n2013), .Z(n2231) );
  AND U2710 ( .A(n2011), .B(n568), .Z(n2115) );
  XOR U2711 ( .A(n2125), .B(n2124), .Z(n2118) );
  NAND U2712 ( .A(n2238), .B(n512), .Z(n2124) );
  XNOR U2713 ( .A(n2123), .B(n2239), .Z(n2125) );
  ANDN U2714 ( .A(n543), .B(n2240), .Z(n2239) );
  NAND U2715 ( .A(n2241), .B(n2242), .Z(n2123) );
  NAND U2716 ( .A(n2243), .B(n2244), .Z(n2241) );
  IV U2717 ( .A(n2126), .Z(n2127) );
  MUX U2718 ( .IN0(o[5]), .IN1(n384), .SEL(n464), .F(\_MxM/n283 ) );
  XOR U2719 ( .A(n2249), .B(\_MxM/Y0[6] ), .Z(n384) );
  XOR U2720 ( .A(n2250), .B(n2251), .Z(n2249) );
  AND U2721 ( .A(n476), .B(n2253), .Z(n2252) );
  XOR U2722 ( .A(n2247), .B(n2251), .Z(n2253) );
  XOR U2723 ( .A(n2246), .B(n2251), .Z(n2247) );
  XNOR U2724 ( .A(n2254), .B(n2177), .Z(n2172) );
  XNOR U2725 ( .A(n2145), .B(n2144), .Z(n2177) );
  XOR U2726 ( .A(n2255), .B(n2149), .Z(n2144) );
  XNOR U2727 ( .A(n2140), .B(n2142), .Z(n2149) );
  NAND U2728 ( .A(n1923), .B(n656), .Z(n2142) );
  XNOR U2729 ( .A(n2138), .B(n2256), .Z(n2140) );
  ANDN U2730 ( .A(n1928), .B(n658), .Z(n2256) );
  XNOR U2731 ( .A(n2148), .B(n2143), .Z(n2255) );
  XOR U2732 ( .A(n2263), .B(n2155), .Z(n2148) );
  XNOR U2733 ( .A(n2153), .B(n2264), .Z(n2155) );
  ANDN U2734 ( .A(n2158), .B(n574), .Z(n2264) );
  XOR U2735 ( .A(n2265), .B(n2266), .Z(n2153) );
  AND U2736 ( .A(n2267), .B(n2268), .Z(n2266) );
  XNOR U2737 ( .A(n2269), .B(n2265), .Z(n2268) );
  AND U2738 ( .A(n2151), .B(n572), .Z(n2157) );
  XNOR U2739 ( .A(n2166), .B(n2165), .Z(n2145) );
  XOR U2740 ( .A(n2273), .B(n2162), .Z(n2165) );
  XNOR U2741 ( .A(n2161), .B(n2274), .Z(n2162) );
  ANDN U2742 ( .A(n1729), .B(n744), .Z(n2274) );
  AND U2743 ( .A(n1722), .B(n742), .Z(n2163) );
  XNOR U2744 ( .A(n2169), .B(n2170), .Z(n2166) );
  NAND U2745 ( .A(n1527), .B(n865), .Z(n2170) );
  XNOR U2746 ( .A(n2168), .B(n2281), .Z(n2169) );
  ANDN U2747 ( .A(n1532), .B(n867), .Z(n2281) );
  XNOR U2748 ( .A(n2176), .B(n2171), .Z(n2254) );
  XOR U2749 ( .A(n2175), .B(n2288), .Z(n2176) );
  AND U2750 ( .A(n2179), .B(n2289), .Z(n2288) );
  AND U2751 ( .A(n2290), .B(n2291), .Z(n2289) );
  NANDN U2752 ( .B(n2292), .A(n511), .Z(n2291) );
  NAND U2753 ( .A(n2293), .B(n2294), .Z(n2290) );
  ANDN U2754 ( .A(n2181), .B(n2180), .Z(n2179) );
  ANDN U2755 ( .A(n2295), .B(n2296), .Z(n2180) );
  OR U2756 ( .A(n2297), .B(n2298), .Z(n2181) );
  XNOR U2757 ( .A(n2197), .B(n2196), .Z(n2173) );
  XOR U2758 ( .A(n2302), .B(n2205), .Z(n2196) );
  XNOR U2759 ( .A(n2190), .B(n2189), .Z(n2205) );
  XOR U2760 ( .A(n2303), .B(n2186), .Z(n2189) );
  XNOR U2761 ( .A(n2185), .B(n2304), .Z(n2186) );
  ANDN U2762 ( .A(n1021), .B(n1319), .Z(n2304) );
  AND U2763 ( .A(n1317), .B(n958), .Z(n2187) );
  XNOR U2764 ( .A(n2193), .B(n2194), .Z(n2190) );
  NANDN U2765 ( .B(n823), .A(n1505), .Z(n2194) );
  XNOR U2766 ( .A(n2192), .B(n2311), .Z(n2193) );
  ANDN U2767 ( .A(n893), .B(n1507), .Z(n2311) );
  XNOR U2768 ( .A(n2204), .B(n2195), .Z(n2302) );
  XOR U2769 ( .A(n2318), .B(n2213), .Z(n2204) );
  XNOR U2770 ( .A(n2201), .B(n2202), .Z(n2213) );
  NAND U2771 ( .A(n1152), .B(n1192), .Z(n2202) );
  XNOR U2772 ( .A(n2200), .B(n2319), .Z(n2201) );
  ANDN U2773 ( .A(n1199), .B(n1154), .Z(n2319) );
  XNOR U2774 ( .A(n2212), .B(n2203), .Z(n2318) );
  XOR U2775 ( .A(n2326), .B(n2209), .Z(n2212) );
  XNOR U2776 ( .A(n2208), .B(n2327), .Z(n2209) );
  ANDN U2777 ( .A(n1383), .B(n1002), .Z(n2327) );
  AND U2778 ( .A(n1000), .B(n1376), .Z(n2210) );
  XNOR U2779 ( .A(n2221), .B(n2220), .Z(n2197) );
  XOR U2780 ( .A(n2334), .B(n2229), .Z(n2220) );
  XNOR U2781 ( .A(n2217), .B(n2218), .Z(n2229) );
  NANDN U2782 ( .B(n636), .A(n1904), .Z(n2218) );
  XNOR U2783 ( .A(n2216), .B(n2335), .Z(n2217) );
  ANDN U2784 ( .A(n677), .B(n1906), .Z(n2335) );
  XNOR U2785 ( .A(n2228), .B(n2219), .Z(n2334) );
  XOR U2786 ( .A(n2342), .B(n2225), .Z(n2228) );
  XNOR U2787 ( .A(n2224), .B(n2343), .Z(n2225) );
  ANDN U2788 ( .A(n784), .B(n1699), .Z(n2343) );
  AND U2789 ( .A(n1697), .B(n730), .Z(n2226) );
  XOR U2790 ( .A(n2237), .B(n2236), .Z(n2221) );
  XOR U2791 ( .A(n2350), .B(n2233), .Z(n2236) );
  XNOR U2792 ( .A(n2232), .B(n2351), .Z(n2233) );
  ANDN U2793 ( .A(n609), .B(n2121), .Z(n2351) );
  AND U2794 ( .A(n2119), .B(n568), .Z(n2234) );
  XOR U2795 ( .A(n2244), .B(n2243), .Z(n2237) );
  NAND U2796 ( .A(n2358), .B(n512), .Z(n2243) );
  XOR U2797 ( .A(n2242), .B(n2359), .Z(n2244) );
  ANDN U2798 ( .A(n543), .B(n2360), .Z(n2359) );
  ANDN U2799 ( .A(n2361), .B(n2362), .Z(n2242) );
  NAND U2800 ( .A(n2363), .B(n2364), .Z(n2361) );
  IV U2801 ( .A(n2245), .Z(n2246) );
  MUX U2802 ( .IN0(o[4]), .IN1(n381), .SEL(n464), .F(\_MxM/n282 ) );
  XOR U2803 ( .A(n2369), .B(\_MxM/Y0[5] ), .Z(n381) );
  XOR U2804 ( .A(n2370), .B(n2371), .Z(n2369) );
  AND U2805 ( .A(n476), .B(n2373), .Z(n2372) );
  XOR U2806 ( .A(n2367), .B(n2371), .Z(n2373) );
  XOR U2807 ( .A(n2366), .B(n2371), .Z(n2367) );
  XNOR U2808 ( .A(n2374), .B(n2301), .Z(n2286) );
  XNOR U2809 ( .A(n2262), .B(n2261), .Z(n2301) );
  XOR U2810 ( .A(n2375), .B(n2272), .Z(n2261) );
  XNOR U2811 ( .A(n2258), .B(n2259), .Z(n2272) );
  NAND U2812 ( .A(n1923), .B(n700), .Z(n2259) );
  XNOR U2813 ( .A(n2257), .B(n2376), .Z(n2258) );
  ANDN U2814 ( .A(n1928), .B(n702), .Z(n2376) );
  XNOR U2815 ( .A(n2271), .B(n2260), .Z(n2375) );
  XOR U2816 ( .A(n2383), .B(n2267), .Z(n2271) );
  XNOR U2817 ( .A(n2265), .B(n2384), .Z(n2267) );
  ANDN U2818 ( .A(n2158), .B(n618), .Z(n2384) );
  XOR U2819 ( .A(n2385), .B(n2386), .Z(n2265) );
  AND U2820 ( .A(n2387), .B(n2388), .Z(n2386) );
  XNOR U2821 ( .A(n2389), .B(n2385), .Z(n2388) );
  AND U2822 ( .A(n2151), .B(n616), .Z(n2269) );
  XNOR U2823 ( .A(n2280), .B(n2279), .Z(n2262) );
  XOR U2824 ( .A(n2393), .B(n2276), .Z(n2279) );
  XNOR U2825 ( .A(n2275), .B(n2394), .Z(n2276) );
  ANDN U2826 ( .A(n1729), .B(n803), .Z(n2394) );
  AND U2827 ( .A(n1722), .B(n801), .Z(n2277) );
  XNOR U2828 ( .A(n2283), .B(n2284), .Z(n2280) );
  NAND U2829 ( .A(n1527), .B(n933), .Z(n2284) );
  XNOR U2830 ( .A(n2282), .B(n2401), .Z(n2283) );
  ANDN U2831 ( .A(n1532), .B(n935), .Z(n2401) );
  XOR U2832 ( .A(n2300), .B(n2285), .Z(n2374) );
  XOR U2833 ( .A(n2408), .B(n2293), .Z(n2300) );
  XOR U2834 ( .A(n2412), .B(n2298), .Z(n2296) );
  NAND U2835 ( .A(n2413), .B(n541), .Z(n2298) );
  NAND U2836 ( .A(n2414), .B(n2297), .Z(n2412) );
  NANDN U2837 ( .B(n544), .A(n2418), .Z(n2414) );
  ANDN U2838 ( .A(n2419), .B(n2420), .Z(n2294) );
  XNOR U2839 ( .A(n2317), .B(n2316), .Z(n2287) );
  XOR U2840 ( .A(n2424), .B(n2325), .Z(n2316) );
  XNOR U2841 ( .A(n2310), .B(n2309), .Z(n2325) );
  XOR U2842 ( .A(n2425), .B(n2306), .Z(n2309) );
  XNOR U2843 ( .A(n2305), .B(n2426), .Z(n2306) );
  ANDN U2844 ( .A(n1021), .B(n1410), .Z(n2426) );
  AND U2845 ( .A(n1408), .B(n958), .Z(n2307) );
  XNOR U2846 ( .A(n2313), .B(n2314), .Z(n2310) );
  NANDN U2847 ( .B(n823), .A(n1601), .Z(n2314) );
  XNOR U2848 ( .A(n2312), .B(n2433), .Z(n2313) );
  ANDN U2849 ( .A(n893), .B(n1603), .Z(n2433) );
  XNOR U2850 ( .A(n2324), .B(n2315), .Z(n2424) );
  XOR U2851 ( .A(n2440), .B(n2333), .Z(n2324) );
  XNOR U2852 ( .A(n2321), .B(n2322), .Z(n2333) );
  NAND U2853 ( .A(n1233), .B(n1192), .Z(n2322) );
  XNOR U2854 ( .A(n2320), .B(n2441), .Z(n2321) );
  ANDN U2855 ( .A(n1199), .B(n1235), .Z(n2441) );
  XNOR U2856 ( .A(n2332), .B(n2323), .Z(n2440) );
  XOR U2857 ( .A(n2448), .B(n2329), .Z(n2332) );
  XNOR U2858 ( .A(n2328), .B(n2449), .Z(n2329) );
  ANDN U2859 ( .A(n1383), .B(n1076), .Z(n2449) );
  AND U2860 ( .A(n1074), .B(n1376), .Z(n2330) );
  XNOR U2861 ( .A(n2341), .B(n2340), .Z(n2317) );
  XOR U2862 ( .A(n2456), .B(n2349), .Z(n2340) );
  XNOR U2863 ( .A(n2337), .B(n2338), .Z(n2349) );
  NANDN U2864 ( .B(n636), .A(n2011), .Z(n2338) );
  XNOR U2865 ( .A(n2336), .B(n2457), .Z(n2337) );
  ANDN U2866 ( .A(n677), .B(n2013), .Z(n2457) );
  XNOR U2867 ( .A(n2348), .B(n2339), .Z(n2456) );
  XOR U2868 ( .A(n2464), .B(n2345), .Z(n2348) );
  XNOR U2869 ( .A(n2344), .B(n2465), .Z(n2345) );
  ANDN U2870 ( .A(n784), .B(n1800), .Z(n2465) );
  AND U2871 ( .A(n1798), .B(n730), .Z(n2346) );
  XOR U2872 ( .A(n2357), .B(n2356), .Z(n2341) );
  XOR U2873 ( .A(n2472), .B(n2353), .Z(n2356) );
  XNOR U2874 ( .A(n2352), .B(n2473), .Z(n2353) );
  ANDN U2875 ( .A(n609), .B(n2240), .Z(n2473) );
  AND U2876 ( .A(n2238), .B(n568), .Z(n2354) );
  XOR U2877 ( .A(n2364), .B(n2363), .Z(n2357) );
  NAND U2878 ( .A(n2480), .B(n512), .Z(n2363) );
  XNOR U2879 ( .A(n2362), .B(n2481), .Z(n2364) );
  ANDN U2880 ( .A(n543), .B(n2482), .Z(n2481) );
  NAND U2881 ( .A(n2483), .B(n2484), .Z(n2362) );
  NAND U2882 ( .A(n2485), .B(n2486), .Z(n2483) );
  IV U2883 ( .A(n2365), .Z(n2366) );
  MUX U2884 ( .IN0(o[3]), .IN1(n378), .SEL(n464), .F(\_MxM/n281 ) );
  XNOR U2885 ( .A(n2490), .B(\_MxM/Y0[4] ), .Z(n378) );
  XNOR U2886 ( .A(n2492), .B(n2493), .Z(n2490) );
  XOR U2887 ( .A(n2491), .B(n2494), .Z(n2492) );
  AND U2888 ( .A(n476), .B(n2495), .Z(n2494) );
  XNOR U2889 ( .A(n2488), .B(n2493), .Z(n2495) );
  XOR U2890 ( .A(n2493), .B(n2487), .Z(n2488) );
  NOR U2891 ( .A(n2496), .B(n2497), .Z(n2487) );
  XNOR U2892 ( .A(n2498), .B(n2423), .Z(n2406) );
  XNOR U2893 ( .A(n2382), .B(n2381), .Z(n2423) );
  XOR U2894 ( .A(n2499), .B(n2392), .Z(n2381) );
  XNOR U2895 ( .A(n2378), .B(n2379), .Z(n2392) );
  NAND U2896 ( .A(n1923), .B(n742), .Z(n2379) );
  XNOR U2897 ( .A(n2377), .B(n2500), .Z(n2378) );
  ANDN U2898 ( .A(n1928), .B(n744), .Z(n2500) );
  XNOR U2899 ( .A(n2391), .B(n2380), .Z(n2499) );
  XOR U2900 ( .A(n2507), .B(n2387), .Z(n2391) );
  XNOR U2901 ( .A(n2385), .B(n2508), .Z(n2387) );
  ANDN U2902 ( .A(n2158), .B(n658), .Z(n2508) );
  AND U2903 ( .A(n2151), .B(n656), .Z(n2389) );
  XNOR U2904 ( .A(n2400), .B(n2399), .Z(n2382) );
  XOR U2905 ( .A(n2515), .B(n2396), .Z(n2399) );
  XNOR U2906 ( .A(n2395), .B(n2516), .Z(n2396) );
  ANDN U2907 ( .A(n1729), .B(n867), .Z(n2516) );
  AND U2908 ( .A(n1722), .B(n865), .Z(n2397) );
  XNOR U2909 ( .A(n2403), .B(n2404), .Z(n2400) );
  NAND U2910 ( .A(n1527), .B(n1000), .Z(n2404) );
  XNOR U2911 ( .A(n2402), .B(n2523), .Z(n2403) );
  ANDN U2912 ( .A(n1532), .B(n1002), .Z(n2523) );
  XNOR U2913 ( .A(n2422), .B(n2405), .Z(n2498) );
  XOR U2914 ( .A(n2530), .B(n2420), .Z(n2422) );
  XOR U2915 ( .A(n2411), .B(n2410), .Z(n2420) );
  XNOR U2916 ( .A(n2409), .B(n2531), .Z(n2410) );
  AND U2917 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2918 ( .B(n2534), .A(n511), .Z(n2533) );
  NANDN U2919 ( .B(n2535), .A(n2536), .Z(n2532) );
  XNOR U2920 ( .A(n2416), .B(n2417), .Z(n2411) );
  NAND U2921 ( .A(n2413), .B(n572), .Z(n2417) );
  XNOR U2922 ( .A(n2415), .B(n2540), .Z(n2416) );
  ANDN U2923 ( .A(n2418), .B(n574), .Z(n2540) );
  NOR U2924 ( .A(n2544), .B(n2545), .Z(n2419) );
  XNOR U2925 ( .A(n2439), .B(n2438), .Z(n2407) );
  XOR U2926 ( .A(n2549), .B(n2447), .Z(n2438) );
  XNOR U2927 ( .A(n2432), .B(n2431), .Z(n2447) );
  XOR U2928 ( .A(n2550), .B(n2428), .Z(n2431) );
  XNOR U2929 ( .A(n2427), .B(n2551), .Z(n2428) );
  ANDN U2930 ( .A(n1021), .B(n1507), .Z(n2551) );
  AND U2931 ( .A(n1505), .B(n958), .Z(n2429) );
  XNOR U2932 ( .A(n2435), .B(n2436), .Z(n2432) );
  NANDN U2933 ( .B(n823), .A(n1697), .Z(n2436) );
  XNOR U2934 ( .A(n2434), .B(n2558), .Z(n2435) );
  ANDN U2935 ( .A(n893), .B(n1699), .Z(n2558) );
  XNOR U2936 ( .A(n2446), .B(n2437), .Z(n2549) );
  XOR U2937 ( .A(n2565), .B(n2455), .Z(n2446) );
  XNOR U2938 ( .A(n2443), .B(n2444), .Z(n2455) );
  NAND U2939 ( .A(n1317), .B(n1192), .Z(n2444) );
  XNOR U2940 ( .A(n2442), .B(n2566), .Z(n2443) );
  ANDN U2941 ( .A(n1199), .B(n1319), .Z(n2566) );
  XNOR U2942 ( .A(n2454), .B(n2445), .Z(n2565) );
  XOR U2943 ( .A(n2573), .B(n2451), .Z(n2454) );
  XNOR U2944 ( .A(n2450), .B(n2574), .Z(n2451) );
  ANDN U2945 ( .A(n1383), .B(n1154), .Z(n2574) );
  AND U2946 ( .A(n1152), .B(n1376), .Z(n2452) );
  XNOR U2947 ( .A(n2463), .B(n2462), .Z(n2439) );
  XOR U2948 ( .A(n2581), .B(n2471), .Z(n2462) );
  XNOR U2949 ( .A(n2459), .B(n2460), .Z(n2471) );
  NANDN U2950 ( .B(n636), .A(n2119), .Z(n2460) );
  XNOR U2951 ( .A(n2458), .B(n2582), .Z(n2459) );
  ANDN U2952 ( .A(n677), .B(n2121), .Z(n2582) );
  XNOR U2953 ( .A(n2470), .B(n2461), .Z(n2581) );
  XOR U2954 ( .A(n2589), .B(n2467), .Z(n2470) );
  XNOR U2955 ( .A(n2466), .B(n2590), .Z(n2467) );
  ANDN U2956 ( .A(n784), .B(n1906), .Z(n2590) );
  AND U2957 ( .A(n1904), .B(n730), .Z(n2468) );
  XOR U2958 ( .A(n2479), .B(n2478), .Z(n2463) );
  XOR U2959 ( .A(n2597), .B(n2475), .Z(n2478) );
  XNOR U2960 ( .A(n2474), .B(n2598), .Z(n2475) );
  ANDN U2961 ( .A(n609), .B(n2360), .Z(n2598) );
  AND U2962 ( .A(n2358), .B(n568), .Z(n2476) );
  XOR U2963 ( .A(n2486), .B(n2485), .Z(n2479) );
  NAND U2964 ( .A(n2605), .B(n512), .Z(n2485) );
  XOR U2965 ( .A(n2484), .B(n2606), .Z(n2486) );
  ANDN U2966 ( .A(n543), .B(n2607), .Z(n2606) );
  ANDN U2967 ( .A(n2608), .B(n2609), .Z(n2484) );
  NAND U2968 ( .A(n2610), .B(n2611), .Z(n2608) );
  IV U2969 ( .A(n2489), .Z(n2491) );
  MUX U2970 ( .IN0(o[2]), .IN1(n375), .SEL(n464), .F(\_MxM/n280 ) );
  IV U2971 ( .A(n2615), .Z(n464) );
  XNOR U2972 ( .A(n2613), .B(\_MxM/Y0[3] ), .Z(n375) );
  XNOR U2973 ( .A(n2616), .B(n2617), .Z(n2613) );
  XOR U2974 ( .A(n2614), .B(n2618), .Z(n2616) );
  AND U2975 ( .A(n476), .B(n2619), .Z(n2618) );
  XNOR U2976 ( .A(n2497), .B(n2617), .Z(n2619) );
  NANDN U2977 ( .B(n2620), .A(n2621), .Z(n2496) );
  XNOR U2978 ( .A(n2622), .B(n2548), .Z(n2528) );
  XNOR U2979 ( .A(n2506), .B(n2505), .Z(n2548) );
  XOR U2980 ( .A(n2623), .B(n2514), .Z(n2505) );
  XNOR U2981 ( .A(n2502), .B(n2503), .Z(n2514) );
  NAND U2982 ( .A(n1923), .B(n801), .Z(n2503) );
  XNOR U2983 ( .A(n2501), .B(n2624), .Z(n2502) );
  ANDN U2984 ( .A(n1928), .B(n803), .Z(n2624) );
  XNOR U2985 ( .A(n2513), .B(n2504), .Z(n2623) );
  XOR U2986 ( .A(n2631), .B(n2510), .Z(n2513) );
  XNOR U2987 ( .A(n2509), .B(n2632), .Z(n2510) );
  ANDN U2988 ( .A(n2158), .B(n702), .Z(n2632) );
  AND U2989 ( .A(n2151), .B(n700), .Z(n2511) );
  XNOR U2990 ( .A(n2522), .B(n2521), .Z(n2506) );
  XOR U2991 ( .A(n2639), .B(n2518), .Z(n2521) );
  XNOR U2992 ( .A(n2517), .B(n2640), .Z(n2518) );
  ANDN U2993 ( .A(n1729), .B(n935), .Z(n2640) );
  AND U2994 ( .A(n1722), .B(n933), .Z(n2519) );
  XNOR U2995 ( .A(n2525), .B(n2526), .Z(n2522) );
  NAND U2996 ( .A(n1527), .B(n1074), .Z(n2526) );
  XNOR U2997 ( .A(n2524), .B(n2647), .Z(n2525) );
  ANDN U2998 ( .A(n1532), .B(n1076), .Z(n2647) );
  XNOR U2999 ( .A(n2547), .B(n2527), .Z(n2622) );
  XOR U3000 ( .A(n2654), .B(n2545), .Z(n2547) );
  XOR U3001 ( .A(n2539), .B(n2538), .Z(n2545) );
  XOR U3002 ( .A(n2659), .B(n2536), .Z(n2655) );
  AND U3003 ( .A(n2660), .B(n541), .Z(n2536) );
  NAND U3004 ( .A(n2661), .B(n2535), .Z(n2659) );
  XOR U3005 ( .A(n2662), .B(n2663), .Z(n2535) );
  AND U3006 ( .A(n2664), .B(n2665), .Z(n2663) );
  XNOR U3007 ( .A(n2666), .B(n2662), .Z(n2665) );
  NANDN U3008 ( .B(n544), .A(n2667), .Z(n2661) );
  XNOR U3009 ( .A(n2542), .B(n2543), .Z(n2539) );
  NAND U3010 ( .A(n2413), .B(n616), .Z(n2543) );
  XNOR U3011 ( .A(n2541), .B(n2668), .Z(n2542) );
  ANDN U3012 ( .A(n2418), .B(n618), .Z(n2668) );
  XOR U3013 ( .A(n2669), .B(n2670), .Z(n2541) );
  AND U3014 ( .A(n2671), .B(n2672), .Z(n2670) );
  XOR U3015 ( .A(n2673), .B(n2669), .Z(n2672) );
  XNOR U3016 ( .A(n2544), .B(n2546), .Z(n2654) );
  XNOR U3017 ( .A(n2677), .B(n2680), .Z(n2679) );
  XNOR U3018 ( .A(n2564), .B(n2563), .Z(n2529) );
  XOR U3019 ( .A(n2681), .B(n2572), .Z(n2563) );
  XNOR U3020 ( .A(n2557), .B(n2556), .Z(n2572) );
  XOR U3021 ( .A(n2682), .B(n2553), .Z(n2556) );
  XNOR U3022 ( .A(n2552), .B(n2683), .Z(n2553) );
  ANDN U3023 ( .A(n1021), .B(n1603), .Z(n2683) );
  AND U3024 ( .A(n1601), .B(n958), .Z(n2554) );
  XNOR U3025 ( .A(n2560), .B(n2561), .Z(n2557) );
  NANDN U3026 ( .B(n823), .A(n1798), .Z(n2561) );
  XNOR U3027 ( .A(n2559), .B(n2690), .Z(n2560) );
  ANDN U3028 ( .A(n893), .B(n1800), .Z(n2690) );
  XNOR U3029 ( .A(n2571), .B(n2562), .Z(n2681) );
  XOR U3030 ( .A(n2697), .B(n2580), .Z(n2571) );
  XNOR U3031 ( .A(n2568), .B(n2569), .Z(n2580) );
  NAND U3032 ( .A(n1408), .B(n1192), .Z(n2569) );
  XNOR U3033 ( .A(n2567), .B(n2698), .Z(n2568) );
  ANDN U3034 ( .A(n1199), .B(n1410), .Z(n2698) );
  XNOR U3035 ( .A(n2579), .B(n2570), .Z(n2697) );
  XOR U3036 ( .A(n2705), .B(n2576), .Z(n2579) );
  XNOR U3037 ( .A(n2575), .B(n2706), .Z(n2576) );
  ANDN U3038 ( .A(n1383), .B(n1235), .Z(n2706) );
  AND U3039 ( .A(n1233), .B(n1376), .Z(n2577) );
  XNOR U3040 ( .A(n2588), .B(n2587), .Z(n2564) );
  XOR U3041 ( .A(n2713), .B(n2596), .Z(n2587) );
  XNOR U3042 ( .A(n2584), .B(n2585), .Z(n2596) );
  NANDN U3043 ( .B(n636), .A(n2238), .Z(n2585) );
  XNOR U3044 ( .A(n2583), .B(n2714), .Z(n2584) );
  ANDN U3045 ( .A(n677), .B(n2240), .Z(n2714) );
  XNOR U3046 ( .A(n2595), .B(n2586), .Z(n2713) );
  XOR U3047 ( .A(n2721), .B(n2592), .Z(n2595) );
  XNOR U3048 ( .A(n2591), .B(n2722), .Z(n2592) );
  ANDN U3049 ( .A(n784), .B(n2013), .Z(n2722) );
  AND U3050 ( .A(n2011), .B(n730), .Z(n2593) );
  XOR U3051 ( .A(n2604), .B(n2603), .Z(n2588) );
  XOR U3052 ( .A(n2729), .B(n2600), .Z(n2603) );
  XNOR U3053 ( .A(n2599), .B(n2730), .Z(n2600) );
  ANDN U3054 ( .A(n609), .B(n2482), .Z(n2730) );
  AND U3055 ( .A(n2480), .B(n568), .Z(n2601) );
  XOR U3056 ( .A(n2611), .B(n2610), .Z(n2604) );
  NAND U3057 ( .A(n2737), .B(n512), .Z(n2610) );
  XNOR U3058 ( .A(n2609), .B(n2738), .Z(n2611) );
  ANDN U3059 ( .A(n543), .B(n2739), .Z(n2738) );
  NAND U3060 ( .A(n2740), .B(n2741), .Z(n2609) );
  NAND U3061 ( .A(n2742), .B(n2743), .Z(n2740) );
  IV U3062 ( .A(n2612), .Z(n2614) );
  MUX U3063 ( .IN0(n372), .IN1(o[1]), .SEL(n2615), .F(\_MxM/n279 ) );
  XNOR U3064 ( .A(n2745), .B(\_MxM/Y0[2] ), .Z(n372) );
  XNOR U3065 ( .A(n2746), .B(n2747), .Z(n2745) );
  XNOR U3066 ( .A(n2744), .B(n2748), .Z(n2746) );
  AND U3067 ( .A(n476), .B(n2749), .Z(n2748) );
  XNOR U3068 ( .A(n2620), .B(n2747), .Z(n2749) );
  XOR U3069 ( .A(n2747), .B(n2621), .Z(n2620) );
  ANDN U3070 ( .A(n2750), .B(n2751), .Z(n2621) );
  XNOR U3071 ( .A(n2752), .B(n2676), .Z(n2652) );
  XNOR U3072 ( .A(n2630), .B(n2629), .Z(n2676) );
  XOR U3073 ( .A(n2753), .B(n2638), .Z(n2629) );
  XNOR U3074 ( .A(n2626), .B(n2627), .Z(n2638) );
  NAND U3075 ( .A(n1923), .B(n865), .Z(n2627) );
  XNOR U3076 ( .A(n2625), .B(n2754), .Z(n2626) );
  ANDN U3077 ( .A(n1928), .B(n867), .Z(n2754) );
  XNOR U3078 ( .A(n2637), .B(n2628), .Z(n2753) );
  XOR U3079 ( .A(n2761), .B(n2634), .Z(n2637) );
  XNOR U3080 ( .A(n2633), .B(n2762), .Z(n2634) );
  ANDN U3081 ( .A(n2158), .B(n744), .Z(n2762) );
  AND U3082 ( .A(n2151), .B(n742), .Z(n2635) );
  XNOR U3083 ( .A(n2646), .B(n2645), .Z(n2630) );
  XOR U3084 ( .A(n2769), .B(n2642), .Z(n2645) );
  XNOR U3085 ( .A(n2641), .B(n2770), .Z(n2642) );
  ANDN U3086 ( .A(n1729), .B(n1002), .Z(n2770) );
  AND U3087 ( .A(n1722), .B(n1000), .Z(n2643) );
  XNOR U3088 ( .A(n2649), .B(n2650), .Z(n2646) );
  NAND U3089 ( .A(n1527), .B(n1152), .Z(n2650) );
  XNOR U3090 ( .A(n2648), .B(n2777), .Z(n2649) );
  ANDN U3091 ( .A(n1532), .B(n1154), .Z(n2777) );
  XOR U3092 ( .A(n2675), .B(n2651), .Z(n2752) );
  XNOR U3093 ( .A(n2784), .B(n2680), .Z(n2675) );
  XNOR U3094 ( .A(n2658), .B(n2657), .Z(n2680) );
  XOR U3095 ( .A(n2785), .B(n2664), .Z(n2657) );
  XNOR U3096 ( .A(n2662), .B(n2786), .Z(n2664) );
  ANDN U3097 ( .A(n2667), .B(n574), .Z(n2786) );
  AND U3098 ( .A(n2660), .B(n572), .Z(n2666) );
  XNOR U3099 ( .A(n2671), .B(n2673), .Z(n2658) );
  NAND U3100 ( .A(n2413), .B(n656), .Z(n2673) );
  XNOR U3101 ( .A(n2669), .B(n2793), .Z(n2671) );
  ANDN U3102 ( .A(n2418), .B(n658), .Z(n2793) );
  XNOR U3103 ( .A(n2678), .B(n2674), .Z(n2784) );
  XOR U3104 ( .A(n2677), .B(n2800), .Z(n2678) );
  AND U3105 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U3106 ( .B(n2803), .A(n2804), .Z(n2802) );
  AND U3107 ( .A(n2805), .B(n2806), .Z(n2801) );
  NANDN U3108 ( .B(n2807), .A(n511), .Z(n2806) );
  OR U3109 ( .A(n2808), .B(n2809), .Z(n2805) );
  XNOR U3110 ( .A(n2696), .B(n2695), .Z(n2653) );
  XOR U3111 ( .A(n2813), .B(n2704), .Z(n2695) );
  XNOR U3112 ( .A(n2689), .B(n2688), .Z(n2704) );
  XOR U3113 ( .A(n2814), .B(n2685), .Z(n2688) );
  XNOR U3114 ( .A(n2684), .B(n2815), .Z(n2685) );
  ANDN U3115 ( .A(n1021), .B(n1699), .Z(n2815) );
  AND U3116 ( .A(n1697), .B(n958), .Z(n2686) );
  XNOR U3117 ( .A(n2692), .B(n2693), .Z(n2689) );
  NANDN U3118 ( .B(n823), .A(n1904), .Z(n2693) );
  XNOR U3119 ( .A(n2691), .B(n2822), .Z(n2692) );
  ANDN U3120 ( .A(n893), .B(n1906), .Z(n2822) );
  XNOR U3121 ( .A(n2703), .B(n2694), .Z(n2813) );
  XOR U3122 ( .A(n2829), .B(n2712), .Z(n2703) );
  XNOR U3123 ( .A(n2700), .B(n2701), .Z(n2712) );
  NAND U3124 ( .A(n1505), .B(n1192), .Z(n2701) );
  XNOR U3125 ( .A(n2699), .B(n2830), .Z(n2700) );
  ANDN U3126 ( .A(n1199), .B(n1507), .Z(n2830) );
  XNOR U3127 ( .A(n2711), .B(n2702), .Z(n2829) );
  XOR U3128 ( .A(n2837), .B(n2708), .Z(n2711) );
  XNOR U3129 ( .A(n2707), .B(n2838), .Z(n2708) );
  ANDN U3130 ( .A(n1383), .B(n1319), .Z(n2838) );
  AND U3131 ( .A(n1317), .B(n1376), .Z(n2709) );
  XNOR U3132 ( .A(n2720), .B(n2719), .Z(n2696) );
  XOR U3133 ( .A(n2845), .B(n2728), .Z(n2719) );
  XNOR U3134 ( .A(n2716), .B(n2717), .Z(n2728) );
  NANDN U3135 ( .B(n636), .A(n2358), .Z(n2717) );
  XNOR U3136 ( .A(n2715), .B(n2846), .Z(n2716) );
  ANDN U3137 ( .A(n677), .B(n2360), .Z(n2846) );
  XNOR U3138 ( .A(n2727), .B(n2718), .Z(n2845) );
  XOR U3139 ( .A(n2853), .B(n2724), .Z(n2727) );
  XNOR U3140 ( .A(n2723), .B(n2854), .Z(n2724) );
  ANDN U3141 ( .A(n784), .B(n2121), .Z(n2854) );
  AND U3142 ( .A(n2119), .B(n730), .Z(n2725) );
  XOR U3143 ( .A(n2736), .B(n2735), .Z(n2720) );
  XOR U3144 ( .A(n2861), .B(n2732), .Z(n2735) );
  XNOR U3145 ( .A(n2731), .B(n2862), .Z(n2732) );
  ANDN U3146 ( .A(n609), .B(n2607), .Z(n2862) );
  AND U3147 ( .A(n2605), .B(n568), .Z(n2733) );
  XOR U3148 ( .A(n2743), .B(n2742), .Z(n2736) );
  NAND U3149 ( .A(n2869), .B(n512), .Z(n2742) );
  XOR U3150 ( .A(n2741), .B(n2870), .Z(n2743) );
  ANDN U3151 ( .A(n543), .B(n2871), .Z(n2870) );
  ANDN U3152 ( .A(n2872), .B(n2873), .Z(n2741) );
  NAND U3153 ( .A(n2874), .B(n2875), .Z(n2872) );
  MUX U3154 ( .IN0(n368), .IN1(o[0]), .SEL(n2615), .F(\_MxM/n278 ) );
  NANDN U3155 ( .B(rst), .A(n463), .Z(n2615) );
  AND U3156 ( .A(n2878), .B(n2879), .Z(n463) );
  AND U3157 ( .A(n2880), .B(n2881), .Z(n2879) );
  ANDN U3158 ( .A(n2882), .B(\_MxM/n[7] ), .Z(n2881) );
  NOR U3159 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n2882) );
  NOR U3160 ( .A(\_MxM/n[5] ), .B(\_MxM/n[6] ), .Z(n2880) );
  AND U3161 ( .A(n2883), .B(n2884), .Z(n2878) );
  NOR U3162 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n2884) );
  NOR U3163 ( .A(\_MxM/n[0] ), .B(n2885), .Z(n2883) );
  XOR U3164 ( .A(n2877), .B(\_MxM/Y0[1] ), .Z(n368) );
  XOR U3165 ( .A(n2886), .B(n2887), .Z(n2877) );
  XOR U3166 ( .A(n2888), .B(n2876), .Z(n2886) );
  NAND U3167 ( .A(n2889), .B(n476), .Z(n2888) );
  XOR U3168 ( .A(e_input[31]), .B(g_input[31]), .Z(n476) );
  XOR U3169 ( .A(n2750), .B(n2887), .Z(n2889) );
  XOR U3170 ( .A(n2751), .B(n2887), .Z(n2750) );
  XNOR U3171 ( .A(n2890), .B(n2799), .Z(n2782) );
  XNOR U3172 ( .A(n2760), .B(n2759), .Z(n2799) );
  XOR U3173 ( .A(n2891), .B(n2768), .Z(n2759) );
  XNOR U3174 ( .A(n2756), .B(n2757), .Z(n2768) );
  NAND U3175 ( .A(n1923), .B(n933), .Z(n2757) );
  XNOR U3176 ( .A(n2755), .B(n2892), .Z(n2756) );
  ANDN U3177 ( .A(n1928), .B(n935), .Z(n2892) );
  XNOR U3178 ( .A(n2767), .B(n2758), .Z(n2891) );
  XOR U3179 ( .A(n2899), .B(n2764), .Z(n2767) );
  XNOR U3180 ( .A(n2763), .B(n2900), .Z(n2764) );
  ANDN U3181 ( .A(n2158), .B(n803), .Z(n2900) );
  AND U3182 ( .A(n2151), .B(n801), .Z(n2765) );
  XNOR U3183 ( .A(n2776), .B(n2775), .Z(n2760) );
  XOR U3184 ( .A(n2907), .B(n2772), .Z(n2775) );
  XNOR U3185 ( .A(n2771), .B(n2908), .Z(n2772) );
  ANDN U3186 ( .A(n1729), .B(n1076), .Z(n2908) );
  AND U3187 ( .A(n1722), .B(n1074), .Z(n2773) );
  XNOR U3188 ( .A(n2779), .B(n2780), .Z(n2776) );
  NAND U3189 ( .A(n1527), .B(n1233), .Z(n2780) );
  XNOR U3190 ( .A(n2778), .B(n2915), .Z(n2779) );
  ANDN U3191 ( .A(n1532), .B(n1235), .Z(n2915) );
  XOR U3192 ( .A(n2798), .B(n2781), .Z(n2890) );
  XNOR U3193 ( .A(n2922), .B(n2812), .Z(n2798) );
  XNOR U3194 ( .A(n2792), .B(n2791), .Z(n2812) );
  XOR U3195 ( .A(n2923), .B(n2788), .Z(n2791) );
  XNOR U3196 ( .A(n2787), .B(n2924), .Z(n2788) );
  ANDN U3197 ( .A(n2667), .B(n618), .Z(n2924) );
  AND U3198 ( .A(n2660), .B(n616), .Z(n2789) );
  XNOR U3199 ( .A(n2795), .B(n2796), .Z(n2792) );
  NAND U3200 ( .A(n2413), .B(n700), .Z(n2796) );
  XNOR U3201 ( .A(n2794), .B(n2931), .Z(n2795) );
  ANDN U3202 ( .A(n2418), .B(n702), .Z(n2931) );
  XOR U3203 ( .A(n2811), .B(n2797), .Z(n2922) );
  XNOR U3204 ( .A(n2938), .B(n2808), .Z(n2811) );
  XNOR U3205 ( .A(n2939), .B(n2804), .Z(n2808) );
  AND U3206 ( .A(n2940), .B(n541), .Z(n2804) );
  NAND U3207 ( .A(n2941), .B(n2803), .Z(n2939) );
  NANDN U3208 ( .B(n544), .A(n2945), .Z(n2941) );
  XNOR U3209 ( .A(n2809), .B(n2810), .Z(n2938) );
  XNOR U3210 ( .A(n2949), .B(n2952), .Z(n2951) );
  XNOR U3211 ( .A(n2828), .B(n2827), .Z(n2783) );
  XOR U3212 ( .A(n2953), .B(n2836), .Z(n2827) );
  XNOR U3213 ( .A(n2821), .B(n2820), .Z(n2836) );
  XOR U3214 ( .A(n2954), .B(n2817), .Z(n2820) );
  XNOR U3215 ( .A(n2816), .B(n2955), .Z(n2817) );
  ANDN U3216 ( .A(n1021), .B(n1800), .Z(n2955) );
  AND U3217 ( .A(n1798), .B(n958), .Z(n2818) );
  XNOR U3218 ( .A(n2824), .B(n2825), .Z(n2821) );
  NANDN U3219 ( .B(n823), .A(n2011), .Z(n2825) );
  XNOR U3220 ( .A(n2823), .B(n2962), .Z(n2824) );
  ANDN U3221 ( .A(n893), .B(n2013), .Z(n2962) );
  XNOR U3222 ( .A(n2835), .B(n2826), .Z(n2953) );
  XOR U3223 ( .A(n2969), .B(n2844), .Z(n2835) );
  XNOR U3224 ( .A(n2832), .B(n2833), .Z(n2844) );
  NAND U3225 ( .A(n1601), .B(n1192), .Z(n2833) );
  XNOR U3226 ( .A(n2831), .B(n2970), .Z(n2832) );
  ANDN U3227 ( .A(n1199), .B(n1603), .Z(n2970) );
  XNOR U3228 ( .A(n2843), .B(n2834), .Z(n2969) );
  XOR U3229 ( .A(n2977), .B(n2840), .Z(n2843) );
  XNOR U3230 ( .A(n2839), .B(n2978), .Z(n2840) );
  ANDN U3231 ( .A(n1383), .B(n1410), .Z(n2978) );
  AND U3232 ( .A(n1408), .B(n1376), .Z(n2841) );
  XNOR U3233 ( .A(n2852), .B(n2851), .Z(n2828) );
  XOR U3234 ( .A(n2985), .B(n2860), .Z(n2851) );
  XNOR U3235 ( .A(n2848), .B(n2849), .Z(n2860) );
  NANDN U3236 ( .B(n636), .A(n2480), .Z(n2849) );
  XNOR U3237 ( .A(n2847), .B(n2986), .Z(n2848) );
  ANDN U3238 ( .A(n677), .B(n2482), .Z(n2986) );
  XNOR U3239 ( .A(n2859), .B(n2850), .Z(n2985) );
  XOR U3240 ( .A(n2993), .B(n2856), .Z(n2859) );
  XNOR U3241 ( .A(n2855), .B(n2994), .Z(n2856) );
  ANDN U3242 ( .A(n784), .B(n2240), .Z(n2994) );
  AND U3243 ( .A(n2238), .B(n730), .Z(n2857) );
  XOR U3244 ( .A(n2868), .B(n2867), .Z(n2852) );
  XOR U3245 ( .A(n3001), .B(n2864), .Z(n2867) );
  XNOR U3246 ( .A(n2863), .B(n3002), .Z(n2864) );
  ANDN U3247 ( .A(n609), .B(n2739), .Z(n3002) );
  AND U3248 ( .A(n2737), .B(n568), .Z(n2865) );
  XOR U3249 ( .A(n2875), .B(n2874), .Z(n2868) );
  NAND U3250 ( .A(n3009), .B(n512), .Z(n2874) );
  XNOR U3251 ( .A(n2873), .B(n3010), .Z(n2875) );
  ANDN U3252 ( .A(n543), .B(n3011), .Z(n3010) );
  NAND U3253 ( .A(n3012), .B(n3013), .Z(n2873) );
  NAND U3254 ( .A(n3014), .B(n3015), .Z(n3012) );
  XNOR U3255 ( .A(n3016), .B(n2937), .Z(n2920) );
  XNOR U3256 ( .A(n2898), .B(n2897), .Z(n2937) );
  XOR U3257 ( .A(n3017), .B(n2906), .Z(n2897) );
  XNOR U3258 ( .A(n2894), .B(n2895), .Z(n2906) );
  NAND U3259 ( .A(n1923), .B(n1000), .Z(n2895) );
  XNOR U3260 ( .A(n2893), .B(n3018), .Z(n2894) );
  ANDN U3261 ( .A(n1928), .B(n1002), .Z(n3018) );
  XOR U3262 ( .A(n3019), .B(n3020), .Z(n2893) );
  AND U3263 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR U3264 ( .A(n3023), .B(n3019), .Z(n3022) );
  XNOR U3265 ( .A(n2905), .B(n2896), .Z(n3017) );
  XOR U3266 ( .A(n3027), .B(n2902), .Z(n2905) );
  XNOR U3267 ( .A(n2901), .B(n3028), .Z(n2902) );
  ANDN U3268 ( .A(n2158), .B(n867), .Z(n3028) );
  XOR U3269 ( .A(n3029), .B(n3030), .Z(n2901) );
  AND U3270 ( .A(n3031), .B(n3032), .Z(n3030) );
  XNOR U3271 ( .A(n3033), .B(n3029), .Z(n3032) );
  AND U3272 ( .A(n2151), .B(n865), .Z(n2903) );
  XNOR U3273 ( .A(n2914), .B(n2913), .Z(n2898) );
  XOR U3274 ( .A(n3037), .B(n2910), .Z(n2913) );
  XNOR U3275 ( .A(n2909), .B(n3038), .Z(n2910) );
  ANDN U3276 ( .A(n1729), .B(n1154), .Z(n3038) );
  AND U3277 ( .A(n1722), .B(n1152), .Z(n2911) );
  XNOR U3278 ( .A(n2917), .B(n2918), .Z(n2914) );
  NAND U3279 ( .A(n1527), .B(n1317), .Z(n2918) );
  XNOR U3280 ( .A(n2916), .B(n3045), .Z(n2917) );
  ANDN U3281 ( .A(n1532), .B(n1319), .Z(n3045) );
  XNOR U3282 ( .A(n2936), .B(n2919), .Z(n3016) );
  XNOR U3283 ( .A(n3049), .B(n3050), .Z(n2919) );
  XNOR U3284 ( .A(n3051), .B(n2948), .Z(n2936) );
  XNOR U3285 ( .A(n2930), .B(n2929), .Z(n2948) );
  XOR U3286 ( .A(n3052), .B(n2926), .Z(n2929) );
  XNOR U3287 ( .A(n2925), .B(n3053), .Z(n2926) );
  ANDN U3288 ( .A(n2667), .B(n658), .Z(n3053) );
  XOR U3289 ( .A(n3054), .B(n3055), .Z(n2925) );
  AND U3290 ( .A(n3056), .B(n3057), .Z(n3055) );
  XNOR U3291 ( .A(n3058), .B(n3054), .Z(n3057) );
  AND U3292 ( .A(n2660), .B(n656), .Z(n2927) );
  XNOR U3293 ( .A(n2933), .B(n2934), .Z(n2930) );
  NAND U3294 ( .A(n2413), .B(n742), .Z(n2934) );
  XNOR U3295 ( .A(n2932), .B(n3062), .Z(n2933) );
  ANDN U3296 ( .A(n2418), .B(n744), .Z(n3062) );
  XOR U3297 ( .A(n3063), .B(n3064), .Z(n2932) );
  AND U3298 ( .A(n3065), .B(n3066), .Z(n3064) );
  XOR U3299 ( .A(n3067), .B(n3063), .Z(n3066) );
  XNOR U3300 ( .A(n2947), .B(n2935), .Z(n3051) );
  XOR U3301 ( .A(n3068), .B(n3069), .Z(n2935) );
  AND U3302 ( .A(n3070), .B(n3071), .Z(n3069) );
  XOR U3303 ( .A(n3072), .B(n3073), .Z(n3071) );
  XNOR U3304 ( .A(n3074), .B(n3068), .Z(n3072) );
  XNOR U3305 ( .A(n3025), .B(n3075), .Z(n3070) );
  XNOR U3306 ( .A(n3068), .B(n3026), .Z(n3075) );
  XNOR U3307 ( .A(n3044), .B(n3043), .Z(n3026) );
  XOR U3308 ( .A(n3076), .B(n3040), .Z(n3043) );
  XNOR U3309 ( .A(n3039), .B(n3077), .Z(n3040) );
  ANDN U3310 ( .A(n1729), .B(n1235), .Z(n3077) );
  AND U3311 ( .A(n1722), .B(n1233), .Z(n3041) );
  XNOR U3312 ( .A(n3047), .B(n3048), .Z(n3044) );
  NAND U3313 ( .A(n1408), .B(n1527), .Z(n3048) );
  XNOR U3314 ( .A(n3046), .B(n3084), .Z(n3047) );
  ANDN U3315 ( .A(n1532), .B(n1410), .Z(n3084) );
  XOR U3316 ( .A(n3088), .B(n3036), .Z(n3025) );
  XNOR U3317 ( .A(n3021), .B(n3023), .Z(n3036) );
  NAND U3318 ( .A(n1923), .B(n1074), .Z(n3023) );
  XNOR U3319 ( .A(n3019), .B(n3089), .Z(n3021) );
  ANDN U3320 ( .A(n1928), .B(n1076), .Z(n3089) );
  XNOR U3321 ( .A(n3035), .B(n3024), .Z(n3088) );
  XOR U3322 ( .A(n3096), .B(n3031), .Z(n3035) );
  XNOR U3323 ( .A(n3029), .B(n3097), .Z(n3031) );
  ANDN U3324 ( .A(n2158), .B(n935), .Z(n3097) );
  XOR U3325 ( .A(n3098), .B(n3099), .Z(n3029) );
  AND U3326 ( .A(n3100), .B(n3101), .Z(n3099) );
  XNOR U3327 ( .A(n3102), .B(n3098), .Z(n3101) );
  AND U3328 ( .A(n2151), .B(n933), .Z(n3033) );
  XOR U3329 ( .A(n3106), .B(n3107), .Z(n3068) );
  AND U3330 ( .A(n3108), .B(n3109), .Z(n3107) );
  XOR U3331 ( .A(n3110), .B(n3111), .Z(n3109) );
  XOR U3332 ( .A(n3106), .B(n3112), .Z(n3111) );
  XNOR U3333 ( .A(n3094), .B(n3113), .Z(n3108) );
  XNOR U3334 ( .A(n3106), .B(n3095), .Z(n3113) );
  XNOR U3335 ( .A(n3083), .B(n3082), .Z(n3095) );
  XOR U3336 ( .A(n3114), .B(n3079), .Z(n3082) );
  XNOR U3337 ( .A(n3078), .B(n3115), .Z(n3079) );
  ANDN U3338 ( .A(n1729), .B(n1319), .Z(n3115) );
  XOR U3339 ( .A(n3116), .B(n3117), .Z(n3078) );
  AND U3340 ( .A(n3118), .B(n3119), .Z(n3117) );
  XNOR U3341 ( .A(n3120), .B(n3116), .Z(n3119) );
  AND U3342 ( .A(n1722), .B(n1317), .Z(n3080) );
  XNOR U3343 ( .A(n3086), .B(n3087), .Z(n3083) );
  NAND U3344 ( .A(n1505), .B(n1527), .Z(n3087) );
  XNOR U3345 ( .A(n3085), .B(n3124), .Z(n3086) );
  ANDN U3346 ( .A(n1532), .B(n1507), .Z(n3124) );
  XOR U3347 ( .A(n3125), .B(n3126), .Z(n3085) );
  AND U3348 ( .A(n3127), .B(n3128), .Z(n3126) );
  XOR U3349 ( .A(n3129), .B(n3125), .Z(n3128) );
  XOR U3350 ( .A(n3130), .B(n3105), .Z(n3094) );
  XNOR U3351 ( .A(n3091), .B(n3092), .Z(n3105) );
  NAND U3352 ( .A(n1923), .B(n1152), .Z(n3092) );
  XNOR U3353 ( .A(n3090), .B(n3131), .Z(n3091) );
  ANDN U3354 ( .A(n1928), .B(n1154), .Z(n3131) );
  XOR U3355 ( .A(n3132), .B(n3133), .Z(n3090) );
  AND U3356 ( .A(n3134), .B(n3135), .Z(n3133) );
  XOR U3357 ( .A(n3136), .B(n3132), .Z(n3135) );
  XNOR U3358 ( .A(n3104), .B(n3093), .Z(n3130) );
  XOR U3359 ( .A(n3140), .B(n3100), .Z(n3104) );
  XNOR U3360 ( .A(n3098), .B(n3141), .Z(n3100) );
  ANDN U3361 ( .A(n2158), .B(n1002), .Z(n3141) );
  XOR U3362 ( .A(n3142), .B(n3143), .Z(n3098) );
  AND U3363 ( .A(n3144), .B(n3145), .Z(n3143) );
  XNOR U3364 ( .A(n3146), .B(n3142), .Z(n3145) );
  XOR U3365 ( .A(n3147), .B(n3102), .Z(n3140) );
  AND U3366 ( .A(n2151), .B(n1000), .Z(n3102) );
  IV U3367 ( .A(n3103), .Z(n3147) );
  XOR U3368 ( .A(n3151), .B(n3152), .Z(n3106) );
  AND U3369 ( .A(n3153), .B(n3154), .Z(n3152) );
  XOR U3370 ( .A(n3155), .B(n3156), .Z(n3154) );
  XOR U3371 ( .A(n3151), .B(n3157), .Z(n3156) );
  XNOR U3372 ( .A(n3138), .B(n3158), .Z(n3153) );
  XNOR U3373 ( .A(n3151), .B(n3139), .Z(n3158) );
  XNOR U3374 ( .A(n3123), .B(n3122), .Z(n3139) );
  XOR U3375 ( .A(n3159), .B(n3118), .Z(n3122) );
  XNOR U3376 ( .A(n3116), .B(n3160), .Z(n3118) );
  ANDN U3377 ( .A(n1729), .B(n1410), .Z(n3160) );
  XOR U3378 ( .A(n3161), .B(n3162), .Z(n3116) );
  AND U3379 ( .A(n3163), .B(n3164), .Z(n3162) );
  XNOR U3380 ( .A(n3165), .B(n3161), .Z(n3164) );
  AND U3381 ( .A(n1408), .B(n1722), .Z(n3120) );
  XNOR U3382 ( .A(n3127), .B(n3129), .Z(n3123) );
  NAND U3383 ( .A(n1601), .B(n1527), .Z(n3129) );
  XNOR U3384 ( .A(n3125), .B(n3169), .Z(n3127) );
  ANDN U3385 ( .A(n1532), .B(n1603), .Z(n3169) );
  XOR U3386 ( .A(n3173), .B(n3150), .Z(n3138) );
  XNOR U3387 ( .A(n3134), .B(n3136), .Z(n3150) );
  NAND U3388 ( .A(n1923), .B(n1233), .Z(n3136) );
  XNOR U3389 ( .A(n3132), .B(n3174), .Z(n3134) );
  ANDN U3390 ( .A(n1928), .B(n1235), .Z(n3174) );
  XOR U3391 ( .A(n3175), .B(n3176), .Z(n3132) );
  AND U3392 ( .A(n3177), .B(n3178), .Z(n3176) );
  XOR U3393 ( .A(n3179), .B(n3175), .Z(n3178) );
  XNOR U3394 ( .A(n3149), .B(n3137), .Z(n3173) );
  XOR U3395 ( .A(n3183), .B(n3144), .Z(n3149) );
  XNOR U3396 ( .A(n3142), .B(n3184), .Z(n3144) );
  ANDN U3397 ( .A(n2158), .B(n1076), .Z(n3184) );
  XOR U3398 ( .A(n3185), .B(n3186), .Z(n3142) );
  AND U3399 ( .A(n3187), .B(n3188), .Z(n3186) );
  XNOR U3400 ( .A(n3189), .B(n3185), .Z(n3188) );
  AND U3401 ( .A(n2151), .B(n1074), .Z(n3146) );
  XOR U3402 ( .A(n3193), .B(n3194), .Z(n3151) );
  AND U3403 ( .A(n3195), .B(n3196), .Z(n3194) );
  XOR U3404 ( .A(n3197), .B(n3198), .Z(n3196) );
  XOR U3405 ( .A(n3193), .B(n3199), .Z(n3198) );
  XNOR U3406 ( .A(n3181), .B(n3200), .Z(n3195) );
  XNOR U3407 ( .A(n3193), .B(n3182), .Z(n3200) );
  XNOR U3408 ( .A(n3168), .B(n3167), .Z(n3182) );
  XOR U3409 ( .A(n3201), .B(n3163), .Z(n3167) );
  XNOR U3410 ( .A(n3161), .B(n3202), .Z(n3163) );
  ANDN U3411 ( .A(n1729), .B(n1507), .Z(n3202) );
  XOR U3412 ( .A(n3203), .B(n3204), .Z(n3161) );
  AND U3413 ( .A(n3205), .B(n3206), .Z(n3204) );
  XNOR U3414 ( .A(n3207), .B(n3203), .Z(n3206) );
  AND U3415 ( .A(n1505), .B(n1722), .Z(n3165) );
  XNOR U3416 ( .A(n3171), .B(n3172), .Z(n3168) );
  NAND U3417 ( .A(n1697), .B(n1527), .Z(n3172) );
  XNOR U3418 ( .A(n3170), .B(n3211), .Z(n3171) );
  ANDN U3419 ( .A(n1532), .B(n1699), .Z(n3211) );
  XOR U3420 ( .A(n3212), .B(n3213), .Z(n3170) );
  AND U3421 ( .A(n3214), .B(n3215), .Z(n3213) );
  XOR U3422 ( .A(n3216), .B(n3212), .Z(n3215) );
  XOR U3423 ( .A(n3217), .B(n3192), .Z(n3181) );
  XNOR U3424 ( .A(n3177), .B(n3179), .Z(n3192) );
  NAND U3425 ( .A(n1923), .B(n1317), .Z(n3179) );
  XNOR U3426 ( .A(n3175), .B(n3218), .Z(n3177) );
  ANDN U3427 ( .A(n1928), .B(n1319), .Z(n3218) );
  XNOR U3428 ( .A(n3191), .B(n3180), .Z(n3217) );
  XOR U3429 ( .A(n3225), .B(n3187), .Z(n3191) );
  XNOR U3430 ( .A(n3185), .B(n3226), .Z(n3187) );
  ANDN U3431 ( .A(n2158), .B(n1154), .Z(n3226) );
  XOR U3432 ( .A(n3227), .B(n3228), .Z(n3185) );
  AND U3433 ( .A(n3229), .B(n3230), .Z(n3228) );
  XNOR U3434 ( .A(n3231), .B(n3227), .Z(n3230) );
  XOR U3435 ( .A(n3232), .B(n3189), .Z(n3225) );
  AND U3436 ( .A(n2151), .B(n1152), .Z(n3189) );
  IV U3437 ( .A(n3190), .Z(n3232) );
  XOR U3438 ( .A(n3236), .B(n3237), .Z(n3193) );
  AND U3439 ( .A(n3238), .B(n3239), .Z(n3237) );
  XOR U3440 ( .A(n3240), .B(n3241), .Z(n3239) );
  XOR U3441 ( .A(n3236), .B(n3242), .Z(n3241) );
  XNOR U3442 ( .A(n3223), .B(n3243), .Z(n3238) );
  XNOR U3443 ( .A(n3236), .B(n3224), .Z(n3243) );
  XNOR U3444 ( .A(n3210), .B(n3209), .Z(n3224) );
  XOR U3445 ( .A(n3244), .B(n3205), .Z(n3209) );
  XNOR U3446 ( .A(n3203), .B(n3245), .Z(n3205) );
  ANDN U3447 ( .A(n1729), .B(n1603), .Z(n3245) );
  XOR U3448 ( .A(n3246), .B(n3247), .Z(n3203) );
  AND U3449 ( .A(n3248), .B(n3249), .Z(n3247) );
  XNOR U3450 ( .A(n3250), .B(n3246), .Z(n3249) );
  AND U3451 ( .A(n1601), .B(n1722), .Z(n3207) );
  XNOR U3452 ( .A(n3214), .B(n3216), .Z(n3210) );
  NAND U3453 ( .A(n1798), .B(n1527), .Z(n3216) );
  XNOR U3454 ( .A(n3212), .B(n3254), .Z(n3214) );
  ANDN U3455 ( .A(n1532), .B(n1800), .Z(n3254) );
  XOR U3456 ( .A(n3258), .B(n3235), .Z(n3223) );
  XNOR U3457 ( .A(n3220), .B(n3221), .Z(n3235) );
  NAND U3458 ( .A(n1408), .B(n1923), .Z(n3221) );
  XNOR U3459 ( .A(n3219), .B(n3259), .Z(n3220) );
  ANDN U3460 ( .A(n1928), .B(n1410), .Z(n3259) );
  XOR U3461 ( .A(n3260), .B(n3261), .Z(n3219) );
  AND U3462 ( .A(n3262), .B(n3263), .Z(n3261) );
  XOR U3463 ( .A(n3264), .B(n3260), .Z(n3263) );
  XNOR U3464 ( .A(n3234), .B(n3222), .Z(n3258) );
  XOR U3465 ( .A(n3268), .B(n3229), .Z(n3234) );
  XNOR U3466 ( .A(n3227), .B(n3269), .Z(n3229) );
  ANDN U3467 ( .A(n2158), .B(n1235), .Z(n3269) );
  XOR U3468 ( .A(n3270), .B(n3271), .Z(n3227) );
  AND U3469 ( .A(n3272), .B(n3273), .Z(n3271) );
  XNOR U3470 ( .A(n3274), .B(n3270), .Z(n3273) );
  AND U3471 ( .A(n2151), .B(n1233), .Z(n3231) );
  XOR U3472 ( .A(n3278), .B(n3279), .Z(n3236) );
  AND U3473 ( .A(n3280), .B(n3281), .Z(n3279) );
  XOR U3474 ( .A(n3282), .B(n3283), .Z(n3281) );
  XOR U3475 ( .A(n3278), .B(n3284), .Z(n3283) );
  XNOR U3476 ( .A(n3266), .B(n3285), .Z(n3280) );
  XNOR U3477 ( .A(n3278), .B(n3267), .Z(n3285) );
  XNOR U3478 ( .A(n3253), .B(n3252), .Z(n3267) );
  XOR U3479 ( .A(n3286), .B(n3248), .Z(n3252) );
  XNOR U3480 ( .A(n3246), .B(n3287), .Z(n3248) );
  ANDN U3481 ( .A(n1729), .B(n1699), .Z(n3287) );
  XOR U3482 ( .A(n3288), .B(n3289), .Z(n3246) );
  AND U3483 ( .A(n3290), .B(n3291), .Z(n3289) );
  XNOR U3484 ( .A(n3292), .B(n3288), .Z(n3291) );
  XOR U3485 ( .A(n3293), .B(n3250), .Z(n3286) );
  AND U3486 ( .A(n1697), .B(n1722), .Z(n3250) );
  IV U3487 ( .A(n3251), .Z(n3293) );
  XNOR U3488 ( .A(n3256), .B(n3257), .Z(n3253) );
  NAND U3489 ( .A(n1904), .B(n1527), .Z(n3257) );
  XNOR U3490 ( .A(n3255), .B(n3297), .Z(n3256) );
  ANDN U3491 ( .A(n1532), .B(n1906), .Z(n3297) );
  XOR U3492 ( .A(n3298), .B(n3299), .Z(n3255) );
  AND U3493 ( .A(n3300), .B(n3301), .Z(n3299) );
  XOR U3494 ( .A(n3302), .B(n3298), .Z(n3301) );
  XOR U3495 ( .A(n3303), .B(n3277), .Z(n3266) );
  XNOR U3496 ( .A(n3262), .B(n3264), .Z(n3277) );
  NAND U3497 ( .A(n1505), .B(n1923), .Z(n3264) );
  XNOR U3498 ( .A(n3260), .B(n3304), .Z(n3262) );
  ANDN U3499 ( .A(n1928), .B(n1507), .Z(n3304) );
  XOR U3500 ( .A(n3305), .B(n3306), .Z(n3260) );
  AND U3501 ( .A(n3307), .B(n3308), .Z(n3306) );
  XOR U3502 ( .A(n3309), .B(n3305), .Z(n3308) );
  XNOR U3503 ( .A(n3276), .B(n3265), .Z(n3303) );
  XOR U3504 ( .A(n3313), .B(n3272), .Z(n3276) );
  XNOR U3505 ( .A(n3270), .B(n3314), .Z(n3272) );
  ANDN U3506 ( .A(n2158), .B(n1319), .Z(n3314) );
  XOR U3507 ( .A(n3315), .B(n3316), .Z(n3270) );
  AND U3508 ( .A(n3317), .B(n3318), .Z(n3316) );
  XNOR U3509 ( .A(n3319), .B(n3315), .Z(n3318) );
  XOR U3510 ( .A(n3320), .B(n3274), .Z(n3313) );
  AND U3511 ( .A(n2151), .B(n1317), .Z(n3274) );
  IV U3512 ( .A(n3275), .Z(n3320) );
  XOR U3513 ( .A(n3324), .B(n3325), .Z(n3278) );
  AND U3514 ( .A(n3326), .B(n3327), .Z(n3325) );
  XOR U3515 ( .A(n3328), .B(n3329), .Z(n3327) );
  XOR U3516 ( .A(n3324), .B(n3330), .Z(n3329) );
  XNOR U3517 ( .A(n3311), .B(n3331), .Z(n3326) );
  XNOR U3518 ( .A(n3324), .B(n3312), .Z(n3331) );
  XNOR U3519 ( .A(n3296), .B(n3295), .Z(n3312) );
  XOR U3520 ( .A(n3332), .B(n3290), .Z(n3295) );
  XNOR U3521 ( .A(n3288), .B(n3333), .Z(n3290) );
  ANDN U3522 ( .A(n1729), .B(n1800), .Z(n3333) );
  XOR U3523 ( .A(n3334), .B(n3335), .Z(n3288) );
  AND U3524 ( .A(n3336), .B(n3337), .Z(n3335) );
  XNOR U3525 ( .A(n3338), .B(n3334), .Z(n3337) );
  XOR U3526 ( .A(n3339), .B(n3292), .Z(n3332) );
  AND U3527 ( .A(n1798), .B(n1722), .Z(n3292) );
  IV U3528 ( .A(n3294), .Z(n3339) );
  XNOR U3529 ( .A(n3300), .B(n3302), .Z(n3296) );
  NAND U3530 ( .A(n2011), .B(n1527), .Z(n3302) );
  XNOR U3531 ( .A(n3298), .B(n3343), .Z(n3300) );
  ANDN U3532 ( .A(n1532), .B(n2013), .Z(n3343) );
  XOR U3533 ( .A(n3344), .B(n3345), .Z(n3298) );
  AND U3534 ( .A(n3346), .B(n3347), .Z(n3345) );
  XOR U3535 ( .A(n3348), .B(n3344), .Z(n3347) );
  XOR U3536 ( .A(n3349), .B(n3323), .Z(n3311) );
  XNOR U3537 ( .A(n3307), .B(n3309), .Z(n3323) );
  NAND U3538 ( .A(n1601), .B(n1923), .Z(n3309) );
  XNOR U3539 ( .A(n3305), .B(n3350), .Z(n3307) );
  ANDN U3540 ( .A(n1928), .B(n1603), .Z(n3350) );
  XNOR U3541 ( .A(n3322), .B(n3310), .Z(n3349) );
  XOR U3542 ( .A(n3357), .B(n3317), .Z(n3322) );
  XNOR U3543 ( .A(n3315), .B(n3358), .Z(n3317) );
  ANDN U3544 ( .A(n2158), .B(n1410), .Z(n3358) );
  XOR U3545 ( .A(n3359), .B(n3360), .Z(n3315) );
  AND U3546 ( .A(n3361), .B(n3362), .Z(n3360) );
  XNOR U3547 ( .A(n3363), .B(n3359), .Z(n3362) );
  XOR U3548 ( .A(n3364), .B(n3319), .Z(n3357) );
  AND U3549 ( .A(n1408), .B(n2151), .Z(n3319) );
  IV U3550 ( .A(n3321), .Z(n3364) );
  XOR U3551 ( .A(n3368), .B(n3369), .Z(n3324) );
  AND U3552 ( .A(n3370), .B(n3371), .Z(n3369) );
  XOR U3553 ( .A(n3372), .B(n3373), .Z(n3371) );
  XOR U3554 ( .A(n3368), .B(n3374), .Z(n3373) );
  XNOR U3555 ( .A(n3355), .B(n3375), .Z(n3370) );
  XNOR U3556 ( .A(n3368), .B(n3356), .Z(n3375) );
  XNOR U3557 ( .A(n3342), .B(n3341), .Z(n3356) );
  XOR U3558 ( .A(n3376), .B(n3336), .Z(n3341) );
  XNOR U3559 ( .A(n3334), .B(n3377), .Z(n3336) );
  ANDN U3560 ( .A(n1729), .B(n1906), .Z(n3377) );
  XOR U3561 ( .A(n3378), .B(n3379), .Z(n3334) );
  AND U3562 ( .A(n3380), .B(n3381), .Z(n3379) );
  XNOR U3563 ( .A(n3382), .B(n3378), .Z(n3381) );
  XOR U3564 ( .A(n3383), .B(n3338), .Z(n3376) );
  AND U3565 ( .A(n1904), .B(n1722), .Z(n3338) );
  IV U3566 ( .A(n3340), .Z(n3383) );
  XNOR U3567 ( .A(n3346), .B(n3348), .Z(n3342) );
  NAND U3568 ( .A(n2119), .B(n1527), .Z(n3348) );
  XNOR U3569 ( .A(n3344), .B(n3387), .Z(n3346) );
  ANDN U3570 ( .A(n1532), .B(n2121), .Z(n3387) );
  XOR U3571 ( .A(n3388), .B(n3389), .Z(n3344) );
  AND U3572 ( .A(n3390), .B(n3391), .Z(n3389) );
  XOR U3573 ( .A(n3392), .B(n3388), .Z(n3391) );
  XOR U3574 ( .A(n3393), .B(n3367), .Z(n3355) );
  XNOR U3575 ( .A(n3352), .B(n3353), .Z(n3367) );
  NAND U3576 ( .A(n1697), .B(n1923), .Z(n3353) );
  XNOR U3577 ( .A(n3351), .B(n3394), .Z(n3352) );
  ANDN U3578 ( .A(n1928), .B(n1699), .Z(n3394) );
  XOR U3579 ( .A(n3395), .B(n3396), .Z(n3351) );
  AND U3580 ( .A(n3397), .B(n3398), .Z(n3396) );
  XOR U3581 ( .A(n3399), .B(n3395), .Z(n3398) );
  XNOR U3582 ( .A(n3366), .B(n3354), .Z(n3393) );
  XOR U3583 ( .A(n3403), .B(n3361), .Z(n3366) );
  XNOR U3584 ( .A(n3359), .B(n3404), .Z(n3361) );
  ANDN U3585 ( .A(n2158), .B(n1507), .Z(n3404) );
  XOR U3586 ( .A(n3405), .B(n3406), .Z(n3359) );
  AND U3587 ( .A(n3407), .B(n3408), .Z(n3406) );
  XNOR U3588 ( .A(n3409), .B(n3405), .Z(n3408) );
  XOR U3589 ( .A(n3410), .B(n3363), .Z(n3403) );
  AND U3590 ( .A(n1505), .B(n2151), .Z(n3363) );
  IV U3591 ( .A(n3365), .Z(n3410) );
  XOR U3592 ( .A(n3414), .B(n3415), .Z(n3368) );
  AND U3593 ( .A(n3416), .B(n3417), .Z(n3415) );
  XOR U3594 ( .A(n3418), .B(n3419), .Z(n3417) );
  XOR U3595 ( .A(n3414), .B(n3420), .Z(n3419) );
  XNOR U3596 ( .A(n3401), .B(n3421), .Z(n3416) );
  XNOR U3597 ( .A(n3414), .B(n3402), .Z(n3421) );
  XNOR U3598 ( .A(n3386), .B(n3385), .Z(n3402) );
  XOR U3599 ( .A(n3422), .B(n3380), .Z(n3385) );
  XNOR U3600 ( .A(n3378), .B(n3423), .Z(n3380) );
  ANDN U3601 ( .A(n1729), .B(n2013), .Z(n3423) );
  XOR U3602 ( .A(n3424), .B(n3425), .Z(n3378) );
  AND U3603 ( .A(n3426), .B(n3427), .Z(n3425) );
  XNOR U3604 ( .A(n3428), .B(n3424), .Z(n3427) );
  XOR U3605 ( .A(n3429), .B(n3382), .Z(n3422) );
  AND U3606 ( .A(n2011), .B(n1722), .Z(n3382) );
  IV U3607 ( .A(n3384), .Z(n3429) );
  XNOR U3608 ( .A(n3390), .B(n3392), .Z(n3386) );
  NAND U3609 ( .A(n2238), .B(n1527), .Z(n3392) );
  XNOR U3610 ( .A(n3388), .B(n3433), .Z(n3390) );
  ANDN U3611 ( .A(n1532), .B(n2240), .Z(n3433) );
  XOR U3612 ( .A(n3434), .B(n3435), .Z(n3388) );
  AND U3613 ( .A(n3436), .B(n3437), .Z(n3435) );
  XOR U3614 ( .A(n3438), .B(n3434), .Z(n3437) );
  XOR U3615 ( .A(n3439), .B(n3413), .Z(n3401) );
  XNOR U3616 ( .A(n3397), .B(n3399), .Z(n3413) );
  NAND U3617 ( .A(n1798), .B(n1923), .Z(n3399) );
  XNOR U3618 ( .A(n3395), .B(n3440), .Z(n3397) );
  ANDN U3619 ( .A(n1928), .B(n1800), .Z(n3440) );
  XOR U3620 ( .A(n3441), .B(n3442), .Z(n3395) );
  AND U3621 ( .A(n3443), .B(n3444), .Z(n3442) );
  XOR U3622 ( .A(n3445), .B(n3441), .Z(n3444) );
  XNOR U3623 ( .A(n3412), .B(n3400), .Z(n3439) );
  XOR U3624 ( .A(n3449), .B(n3407), .Z(n3412) );
  XNOR U3625 ( .A(n3405), .B(n3450), .Z(n3407) );
  ANDN U3626 ( .A(n2158), .B(n1603), .Z(n3450) );
  XOR U3627 ( .A(n3451), .B(n3452), .Z(n3405) );
  AND U3628 ( .A(n3453), .B(n3454), .Z(n3452) );
  XNOR U3629 ( .A(n3455), .B(n3451), .Z(n3454) );
  XOR U3630 ( .A(n3456), .B(n3409), .Z(n3449) );
  AND U3631 ( .A(n1601), .B(n2151), .Z(n3409) );
  IV U3632 ( .A(n3411), .Z(n3456) );
  XOR U3633 ( .A(n3460), .B(n3461), .Z(n3414) );
  AND U3634 ( .A(n3462), .B(n3463), .Z(n3461) );
  XOR U3635 ( .A(n3464), .B(n3465), .Z(n3463) );
  XOR U3636 ( .A(n3460), .B(n3466), .Z(n3465) );
  XNOR U3637 ( .A(n3447), .B(n3467), .Z(n3462) );
  XNOR U3638 ( .A(n3460), .B(n3448), .Z(n3467) );
  XNOR U3639 ( .A(n3432), .B(n3431), .Z(n3448) );
  XOR U3640 ( .A(n3468), .B(n3426), .Z(n3431) );
  XNOR U3641 ( .A(n3424), .B(n3469), .Z(n3426) );
  ANDN U3642 ( .A(n1729), .B(n2121), .Z(n3469) );
  XOR U3643 ( .A(n3470), .B(n3471), .Z(n3424) );
  AND U3644 ( .A(n3472), .B(n3473), .Z(n3471) );
  XNOR U3645 ( .A(n3474), .B(n3470), .Z(n3473) );
  XOR U3646 ( .A(n3475), .B(n3428), .Z(n3468) );
  AND U3647 ( .A(n2119), .B(n1722), .Z(n3428) );
  IV U3648 ( .A(n3430), .Z(n3475) );
  XNOR U3649 ( .A(n3436), .B(n3438), .Z(n3432) );
  NAND U3650 ( .A(n2358), .B(n1527), .Z(n3438) );
  XNOR U3651 ( .A(n3434), .B(n3479), .Z(n3436) );
  ANDN U3652 ( .A(n1532), .B(n2360), .Z(n3479) );
  XOR U3653 ( .A(n3480), .B(n3481), .Z(n3434) );
  AND U3654 ( .A(n3482), .B(n3483), .Z(n3481) );
  XOR U3655 ( .A(n3484), .B(n3480), .Z(n3483) );
  XOR U3656 ( .A(n3485), .B(n3459), .Z(n3447) );
  XNOR U3657 ( .A(n3443), .B(n3445), .Z(n3459) );
  NAND U3658 ( .A(n1904), .B(n1923), .Z(n3445) );
  XNOR U3659 ( .A(n3441), .B(n3486), .Z(n3443) );
  ANDN U3660 ( .A(n1928), .B(n1906), .Z(n3486) );
  XOR U3661 ( .A(n3487), .B(n3488), .Z(n3441) );
  AND U3662 ( .A(n3489), .B(n3490), .Z(n3488) );
  XOR U3663 ( .A(n3491), .B(n3487), .Z(n3490) );
  XNOR U3664 ( .A(n3458), .B(n3446), .Z(n3485) );
  XOR U3665 ( .A(n3495), .B(n3453), .Z(n3458) );
  XNOR U3666 ( .A(n3451), .B(n3496), .Z(n3453) );
  ANDN U3667 ( .A(n2158), .B(n1699), .Z(n3496) );
  XOR U3668 ( .A(n3497), .B(n3498), .Z(n3451) );
  AND U3669 ( .A(n3499), .B(n3500), .Z(n3498) );
  XNOR U3670 ( .A(n3501), .B(n3497), .Z(n3500) );
  XOR U3671 ( .A(n3502), .B(n3455), .Z(n3495) );
  AND U3672 ( .A(n1697), .B(n2151), .Z(n3455) );
  IV U3673 ( .A(n3457), .Z(n3502) );
  XOR U3674 ( .A(n3506), .B(n3507), .Z(n3460) );
  AND U3675 ( .A(n3508), .B(n3509), .Z(n3507) );
  XOR U3676 ( .A(n3510), .B(n3511), .Z(n3509) );
  XOR U3677 ( .A(n3506), .B(n3512), .Z(n3511) );
  XNOR U3678 ( .A(n3493), .B(n3513), .Z(n3508) );
  XNOR U3679 ( .A(n3506), .B(n3494), .Z(n3513) );
  XNOR U3680 ( .A(n3478), .B(n3477), .Z(n3494) );
  XOR U3681 ( .A(n3514), .B(n3472), .Z(n3477) );
  XNOR U3682 ( .A(n3470), .B(n3515), .Z(n3472) );
  ANDN U3683 ( .A(n1729), .B(n2240), .Z(n3515) );
  XOR U3684 ( .A(n3516), .B(n3517), .Z(n3470) );
  AND U3685 ( .A(n3518), .B(n3519), .Z(n3517) );
  XNOR U3686 ( .A(n3520), .B(n3516), .Z(n3519) );
  XOR U3687 ( .A(n3521), .B(n3474), .Z(n3514) );
  AND U3688 ( .A(n2238), .B(n1722), .Z(n3474) );
  IV U3689 ( .A(n3476), .Z(n3521) );
  XNOR U3690 ( .A(n3482), .B(n3484), .Z(n3478) );
  NAND U3691 ( .A(n2480), .B(n1527), .Z(n3484) );
  XNOR U3692 ( .A(n3480), .B(n3525), .Z(n3482) );
  ANDN U3693 ( .A(n1532), .B(n2482), .Z(n3525) );
  XOR U3694 ( .A(n3529), .B(n3505), .Z(n3493) );
  XNOR U3695 ( .A(n3489), .B(n3491), .Z(n3505) );
  NAND U3696 ( .A(n2011), .B(n1923), .Z(n3491) );
  XNOR U3697 ( .A(n3487), .B(n3530), .Z(n3489) );
  ANDN U3698 ( .A(n1928), .B(n2013), .Z(n3530) );
  XOR U3699 ( .A(n3531), .B(n3532), .Z(n3487) );
  AND U3700 ( .A(n3533), .B(n3534), .Z(n3532) );
  XOR U3701 ( .A(n3535), .B(n3531), .Z(n3534) );
  XNOR U3702 ( .A(n3504), .B(n3492), .Z(n3529) );
  XOR U3703 ( .A(n3539), .B(n3499), .Z(n3504) );
  XNOR U3704 ( .A(n3497), .B(n3540), .Z(n3499) );
  ANDN U3705 ( .A(n2158), .B(n1800), .Z(n3540) );
  XOR U3706 ( .A(n3541), .B(n3542), .Z(n3497) );
  AND U3707 ( .A(n3543), .B(n3544), .Z(n3542) );
  XNOR U3708 ( .A(n3545), .B(n3541), .Z(n3544) );
  XOR U3709 ( .A(n3546), .B(n3501), .Z(n3539) );
  AND U3710 ( .A(n1798), .B(n2151), .Z(n3501) );
  IV U3711 ( .A(n3503), .Z(n3546) );
  XOR U3712 ( .A(n3550), .B(n3551), .Z(n3506) );
  AND U3713 ( .A(n3552), .B(n3553), .Z(n3551) );
  XOR U3714 ( .A(n3554), .B(n3555), .Z(n3553) );
  XOR U3715 ( .A(n3550), .B(n3556), .Z(n3555) );
  XNOR U3716 ( .A(n3537), .B(n3557), .Z(n3552) );
  XNOR U3717 ( .A(n3550), .B(n3538), .Z(n3557) );
  XNOR U3718 ( .A(n3524), .B(n3523), .Z(n3538) );
  XOR U3719 ( .A(n3558), .B(n3518), .Z(n3523) );
  XNOR U3720 ( .A(n3516), .B(n3559), .Z(n3518) );
  ANDN U3721 ( .A(n1729), .B(n2360), .Z(n3559) );
  XOR U3722 ( .A(n3560), .B(n3561), .Z(n3516) );
  AND U3723 ( .A(n3562), .B(n3563), .Z(n3561) );
  XNOR U3724 ( .A(n3564), .B(n3560), .Z(n3563) );
  XOR U3725 ( .A(n3565), .B(n3520), .Z(n3558) );
  AND U3726 ( .A(n2358), .B(n1722), .Z(n3520) );
  IV U3727 ( .A(n3522), .Z(n3565) );
  XNOR U3728 ( .A(n3527), .B(n3528), .Z(n3524) );
  NAND U3729 ( .A(n2605), .B(n1527), .Z(n3528) );
  XNOR U3730 ( .A(n3526), .B(n3569), .Z(n3527) );
  ANDN U3731 ( .A(n1532), .B(n2607), .Z(n3569) );
  XOR U3732 ( .A(n3570), .B(n3571), .Z(n3526) );
  AND U3733 ( .A(n3572), .B(n3573), .Z(n3571) );
  XOR U3734 ( .A(n3574), .B(n3570), .Z(n3573) );
  XOR U3735 ( .A(n3575), .B(n3549), .Z(n3537) );
  XNOR U3736 ( .A(n3533), .B(n3535), .Z(n3549) );
  NAND U3737 ( .A(n2119), .B(n1923), .Z(n3535) );
  XNOR U3738 ( .A(n3531), .B(n3576), .Z(n3533) );
  ANDN U3739 ( .A(n1928), .B(n2121), .Z(n3576) );
  XOR U3740 ( .A(n3577), .B(n3578), .Z(n3531) );
  AND U3741 ( .A(n3579), .B(n3580), .Z(n3578) );
  XOR U3742 ( .A(n3581), .B(n3577), .Z(n3580) );
  XNOR U3743 ( .A(n3548), .B(n3536), .Z(n3575) );
  XOR U3744 ( .A(n3585), .B(n3543), .Z(n3548) );
  XNOR U3745 ( .A(n3541), .B(n3586), .Z(n3543) );
  ANDN U3746 ( .A(n2158), .B(n1906), .Z(n3586) );
  XOR U3747 ( .A(n3587), .B(n3588), .Z(n3541) );
  AND U3748 ( .A(n3589), .B(n3590), .Z(n3588) );
  XNOR U3749 ( .A(n3591), .B(n3587), .Z(n3590) );
  XOR U3750 ( .A(n3592), .B(n3545), .Z(n3585) );
  AND U3751 ( .A(n1904), .B(n2151), .Z(n3545) );
  IV U3752 ( .A(n3547), .Z(n3592) );
  XOR U3753 ( .A(n3596), .B(n3597), .Z(n3550) );
  AND U3754 ( .A(n3598), .B(n3599), .Z(n3597) );
  XOR U3755 ( .A(n3600), .B(n3601), .Z(n3599) );
  XOR U3756 ( .A(n3596), .B(n3602), .Z(n3601) );
  XNOR U3757 ( .A(n3583), .B(n3603), .Z(n3598) );
  XNOR U3758 ( .A(n3596), .B(n3584), .Z(n3603) );
  XNOR U3759 ( .A(n3568), .B(n3567), .Z(n3584) );
  XOR U3760 ( .A(n3604), .B(n3562), .Z(n3567) );
  XNOR U3761 ( .A(n3560), .B(n3605), .Z(n3562) );
  ANDN U3762 ( .A(n1729), .B(n2482), .Z(n3605) );
  XOR U3763 ( .A(n3606), .B(n3607), .Z(n3560) );
  AND U3764 ( .A(n3608), .B(n3609), .Z(n3607) );
  XNOR U3765 ( .A(n3610), .B(n3606), .Z(n3609) );
  XOR U3766 ( .A(n3611), .B(n3564), .Z(n3604) );
  AND U3767 ( .A(n2480), .B(n1722), .Z(n3564) );
  IV U3768 ( .A(n3566), .Z(n3611) );
  XNOR U3769 ( .A(n3572), .B(n3574), .Z(n3568) );
  NAND U3770 ( .A(n2737), .B(n1527), .Z(n3574) );
  XNOR U3771 ( .A(n3570), .B(n3615), .Z(n3572) );
  ANDN U3772 ( .A(n1532), .B(n2739), .Z(n3615) );
  XOR U3773 ( .A(n3616), .B(n3617), .Z(n3570) );
  AND U3774 ( .A(n3618), .B(n3619), .Z(n3617) );
  XOR U3775 ( .A(n3620), .B(n3616), .Z(n3619) );
  XOR U3776 ( .A(n3621), .B(n3595), .Z(n3583) );
  XNOR U3777 ( .A(n3579), .B(n3581), .Z(n3595) );
  NAND U3778 ( .A(n2238), .B(n1923), .Z(n3581) );
  XNOR U3779 ( .A(n3577), .B(n3622), .Z(n3579) );
  ANDN U3780 ( .A(n1928), .B(n2240), .Z(n3622) );
  XOR U3781 ( .A(n3623), .B(n3624), .Z(n3577) );
  AND U3782 ( .A(n3625), .B(n3626), .Z(n3624) );
  XOR U3783 ( .A(n3627), .B(n3623), .Z(n3626) );
  XNOR U3784 ( .A(n3594), .B(n3582), .Z(n3621) );
  XOR U3785 ( .A(n3631), .B(n3589), .Z(n3594) );
  XNOR U3786 ( .A(n3587), .B(n3632), .Z(n3589) );
  ANDN U3787 ( .A(n2158), .B(n2013), .Z(n3632) );
  XOR U3788 ( .A(n3633), .B(n3634), .Z(n3587) );
  AND U3789 ( .A(n3635), .B(n3636), .Z(n3634) );
  XNOR U3790 ( .A(n3637), .B(n3633), .Z(n3636) );
  XOR U3791 ( .A(n3638), .B(n3591), .Z(n3631) );
  AND U3792 ( .A(n2011), .B(n2151), .Z(n3591) );
  IV U3793 ( .A(n3593), .Z(n3638) );
  XOR U3794 ( .A(n3642), .B(n3643), .Z(n3596) );
  AND U3795 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U3796 ( .A(n3646), .B(n3647), .Z(n3645) );
  XOR U3797 ( .A(n3642), .B(n3648), .Z(n3647) );
  XNOR U3798 ( .A(n3629), .B(n3649), .Z(n3644) );
  XNOR U3799 ( .A(n3642), .B(n3630), .Z(n3649) );
  XNOR U3800 ( .A(n3614), .B(n3613), .Z(n3630) );
  XOR U3801 ( .A(n3650), .B(n3608), .Z(n3613) );
  XNOR U3802 ( .A(n3606), .B(n3651), .Z(n3608) );
  ANDN U3803 ( .A(n1729), .B(n2607), .Z(n3651) );
  XOR U3804 ( .A(n3652), .B(n3653), .Z(n3606) );
  AND U3805 ( .A(n3654), .B(n3655), .Z(n3653) );
  XNOR U3806 ( .A(n3656), .B(n3652), .Z(n3655) );
  XOR U3807 ( .A(n3657), .B(n3610), .Z(n3650) );
  AND U3808 ( .A(n2605), .B(n1722), .Z(n3610) );
  IV U3809 ( .A(n3612), .Z(n3657) );
  XNOR U3810 ( .A(n3618), .B(n3620), .Z(n3614) );
  NAND U3811 ( .A(n2869), .B(n1527), .Z(n3620) );
  XNOR U3812 ( .A(n3616), .B(n3661), .Z(n3618) );
  ANDN U3813 ( .A(n1532), .B(n2871), .Z(n3661) );
  XOR U3814 ( .A(n3662), .B(n3663), .Z(n3616) );
  AND U3815 ( .A(n3664), .B(n3665), .Z(n3663) );
  XOR U3816 ( .A(n3666), .B(n3662), .Z(n3665) );
  XOR U3817 ( .A(n3667), .B(n3641), .Z(n3629) );
  XNOR U3818 ( .A(n3625), .B(n3627), .Z(n3641) );
  NAND U3819 ( .A(n2358), .B(n1923), .Z(n3627) );
  XNOR U3820 ( .A(n3623), .B(n3668), .Z(n3625) );
  ANDN U3821 ( .A(n1928), .B(n2360), .Z(n3668) );
  XOR U3822 ( .A(n3669), .B(n3670), .Z(n3623) );
  AND U3823 ( .A(n3671), .B(n3672), .Z(n3670) );
  XOR U3824 ( .A(n3673), .B(n3669), .Z(n3672) );
  XNOR U3825 ( .A(n3640), .B(n3628), .Z(n3667) );
  XOR U3826 ( .A(n3677), .B(n3635), .Z(n3640) );
  XNOR U3827 ( .A(n3633), .B(n3678), .Z(n3635) );
  ANDN U3828 ( .A(n2158), .B(n2121), .Z(n3678) );
  XOR U3829 ( .A(n3679), .B(n3680), .Z(n3633) );
  AND U3830 ( .A(n3681), .B(n3682), .Z(n3680) );
  XNOR U3831 ( .A(n3683), .B(n3679), .Z(n3682) );
  XOR U3832 ( .A(n3684), .B(n3637), .Z(n3677) );
  AND U3833 ( .A(n2119), .B(n2151), .Z(n3637) );
  IV U3834 ( .A(n3639), .Z(n3684) );
  XOR U3835 ( .A(n3688), .B(n3689), .Z(n3642) );
  AND U3836 ( .A(n3690), .B(n3691), .Z(n3689) );
  XOR U3837 ( .A(n3692), .B(n3693), .Z(n3691) );
  XOR U3838 ( .A(n3688), .B(n3694), .Z(n3693) );
  XNOR U3839 ( .A(n3675), .B(n3695), .Z(n3690) );
  XNOR U3840 ( .A(n3688), .B(n3676), .Z(n3695) );
  XNOR U3841 ( .A(n3660), .B(n3659), .Z(n3676) );
  XOR U3842 ( .A(n3696), .B(n3654), .Z(n3659) );
  XNOR U3843 ( .A(n3652), .B(n3697), .Z(n3654) );
  ANDN U3844 ( .A(n1729), .B(n2739), .Z(n3697) );
  XOR U3845 ( .A(n3701), .B(n3656), .Z(n3696) );
  AND U3846 ( .A(n2737), .B(n1722), .Z(n3656) );
  IV U3847 ( .A(n3658), .Z(n3701) );
  XNOR U3848 ( .A(n3664), .B(n3666), .Z(n3660) );
  NAND U3849 ( .A(n3009), .B(n1527), .Z(n3666) );
  XNOR U3850 ( .A(n3662), .B(n3705), .Z(n3664) );
  ANDN U3851 ( .A(n1532), .B(n3011), .Z(n3705) );
  XOR U3852 ( .A(n3709), .B(n3687), .Z(n3675) );
  XNOR U3853 ( .A(n3671), .B(n3673), .Z(n3687) );
  NAND U3854 ( .A(n2480), .B(n1923), .Z(n3673) );
  XNOR U3855 ( .A(n3669), .B(n3710), .Z(n3671) );
  ANDN U3856 ( .A(n1928), .B(n2482), .Z(n3710) );
  XOR U3857 ( .A(n3711), .B(n3712), .Z(n3669) );
  AND U3858 ( .A(n3713), .B(n3714), .Z(n3712) );
  XOR U3859 ( .A(n3715), .B(n3711), .Z(n3714) );
  XNOR U3860 ( .A(n3686), .B(n3674), .Z(n3709) );
  XOR U3861 ( .A(n3719), .B(n3681), .Z(n3686) );
  XNOR U3862 ( .A(n3679), .B(n3720), .Z(n3681) );
  ANDN U3863 ( .A(n2158), .B(n2240), .Z(n3720) );
  XOR U3864 ( .A(n3721), .B(n3722), .Z(n3679) );
  AND U3865 ( .A(n3723), .B(n3724), .Z(n3722) );
  XNOR U3866 ( .A(n3725), .B(n3721), .Z(n3724) );
  XOR U3867 ( .A(n3726), .B(n3683), .Z(n3719) );
  AND U3868 ( .A(n2238), .B(n2151), .Z(n3683) );
  IV U3869 ( .A(n3685), .Z(n3726) );
  XOR U3870 ( .A(n3731), .B(n3732), .Z(n3050) );
  XOR U3871 ( .A(n3733), .B(n3730), .Z(n3731) );
  XNOR U3872 ( .A(n3718), .B(n3717), .Z(n3049) );
  XOR U3873 ( .A(n3734), .B(n3729), .Z(n3717) );
  XNOR U3874 ( .A(n3713), .B(n3715), .Z(n3729) );
  NAND U3875 ( .A(n2605), .B(n1923), .Z(n3715) );
  XNOR U3876 ( .A(n3711), .B(n3735), .Z(n3713) );
  ANDN U3877 ( .A(n1928), .B(n2607), .Z(n3735) );
  XOR U3878 ( .A(n3728), .B(n3716), .Z(n3734) );
  XOR U3879 ( .A(n3739), .B(n3740), .Z(n3716) );
  XOR U3880 ( .A(n3741), .B(n3723), .Z(n3728) );
  XNOR U3881 ( .A(n3721), .B(n3742), .Z(n3723) );
  ANDN U3882 ( .A(n2158), .B(n2360), .Z(n3742) );
  AND U3883 ( .A(n2358), .B(n2151), .Z(n3725) );
  XNOR U3884 ( .A(n3746), .B(n3747), .Z(n3727) );
  AND U3885 ( .A(n3748), .B(n3749), .Z(n3747) );
  XNOR U3886 ( .A(n3744), .B(n3750), .Z(n3749) );
  XNOR U3887 ( .A(n3745), .B(n3746), .Z(n3750) );
  AND U3888 ( .A(n2480), .B(n2151), .Z(n3745) );
  XOR U3889 ( .A(n3743), .B(n3751), .Z(n3744) );
  ANDN U3890 ( .A(n2158), .B(n2482), .Z(n3751) );
  XNOR U3891 ( .A(n3737), .B(n3755), .Z(n3748) );
  XNOR U3892 ( .A(n3738), .B(n3746), .Z(n3755) );
  AND U3893 ( .A(n2737), .B(n1923), .Z(n3738) );
  XOR U3894 ( .A(n3736), .B(n3756), .Z(n3737) );
  ANDN U3895 ( .A(n1928), .B(n2739), .Z(n3756) );
  XOR U3896 ( .A(n3760), .B(n3761), .Z(n3746) );
  AND U3897 ( .A(n3762), .B(n3763), .Z(n3761) );
  XNOR U3898 ( .A(n3753), .B(n3764), .Z(n3763) );
  XNOR U3899 ( .A(n3754), .B(n3760), .Z(n3764) );
  AND U3900 ( .A(n2605), .B(n2151), .Z(n3754) );
  XOR U3901 ( .A(n3752), .B(n3765), .Z(n3753) );
  ANDN U3902 ( .A(n2158), .B(n2607), .Z(n3765) );
  XNOR U3903 ( .A(n3758), .B(n3769), .Z(n3762) );
  XNOR U3904 ( .A(n3759), .B(n3760), .Z(n3769) );
  AND U3905 ( .A(n2869), .B(n1923), .Z(n3759) );
  XOR U3906 ( .A(n3757), .B(n3770), .Z(n3758) );
  ANDN U3907 ( .A(n1928), .B(n2871), .Z(n3770) );
  XOR U3908 ( .A(n3774), .B(n3775), .Z(n3760) );
  AND U3909 ( .A(n3776), .B(n3777), .Z(n3775) );
  XNOR U3910 ( .A(n3767), .B(n3778), .Z(n3777) );
  XNOR U3911 ( .A(n3768), .B(n3774), .Z(n3778) );
  AND U3912 ( .A(n2737), .B(n2151), .Z(n3768) );
  XOR U3913 ( .A(n3766), .B(n3779), .Z(n3767) );
  ANDN U3914 ( .A(n2158), .B(n2739), .Z(n3779) );
  XNOR U3915 ( .A(n3772), .B(n3783), .Z(n3776) );
  XNOR U3916 ( .A(n3773), .B(n3774), .Z(n3783) );
  AND U3917 ( .A(n3009), .B(n1923), .Z(n3773) );
  XOR U3918 ( .A(n3771), .B(n3784), .Z(n3772) );
  ANDN U3919 ( .A(n1928), .B(n3011), .Z(n3784) );
  XNOR U3920 ( .A(n3789), .B(n3781), .Z(n3740) );
  XNOR U3921 ( .A(n3780), .B(n3790), .Z(n3781) );
  ANDN U3922 ( .A(n2158), .B(n2871), .Z(n3790) );
  XNOR U3923 ( .A(n3793), .B(n3791), .Z(n3792) );
  ANDN U3924 ( .A(n2158), .B(n3011), .Z(n3793) );
  XNOR U3925 ( .A(n3788), .B(n3782), .Z(n3789) );
  AND U3926 ( .A(n2869), .B(n2151), .Z(n3782) );
  XNOR U3927 ( .A(n3786), .B(n3787), .Z(n3739) );
  NAND U3928 ( .A(n3797), .B(n1923), .Z(n3787) );
  XNOR U3929 ( .A(n3785), .B(n3798), .Z(n3786) );
  ANDN U3930 ( .A(n1928), .B(n3799), .Z(n3798) );
  NAND U3931 ( .A(g_input[0]), .B(n3800), .Z(n3785) );
  NANDN U3932 ( .B(n1923), .A(n3801), .Z(n3800) );
  NANDN U3933 ( .B(n3802), .A(n1928), .Z(n3801) );
  IV U3934 ( .A(n1822), .Z(n1923) );
  XNOR U3935 ( .A(n3795), .B(n3796), .Z(n3788) );
  NAND U3936 ( .A(n3797), .B(n2151), .Z(n3796) );
  XNOR U3937 ( .A(n3794), .B(n3805), .Z(n3795) );
  ANDN U3938 ( .A(n2158), .B(n3799), .Z(n3805) );
  NAND U3939 ( .A(g_input[0]), .B(n3806), .Z(n3794) );
  NANDN U3940 ( .B(n2151), .A(n3807), .Z(n3806) );
  NANDN U3941 ( .B(n3802), .A(n2158), .Z(n3807) );
  IV U3942 ( .A(n2039), .Z(n2151) );
  XNOR U3943 ( .A(n3704), .B(n3703), .Z(n3718) );
  XOR U3944 ( .A(n3810), .B(n3699), .Z(n3703) );
  XNOR U3945 ( .A(n3698), .B(n3811), .Z(n3699) );
  ANDN U3946 ( .A(n1729), .B(n2871), .Z(n3811) );
  XNOR U3947 ( .A(n3814), .B(n3812), .Z(n3813) );
  ANDN U3948 ( .A(n1729), .B(n3011), .Z(n3814) );
  XNOR U3949 ( .A(n3702), .B(n3700), .Z(n3810) );
  AND U3950 ( .A(n2869), .B(n1722), .Z(n3700) );
  XNOR U3951 ( .A(n3816), .B(n3817), .Z(n3702) );
  NAND U3952 ( .A(n3797), .B(n1722), .Z(n3817) );
  XNOR U3953 ( .A(n3815), .B(n3818), .Z(n3816) );
  ANDN U3954 ( .A(n1729), .B(n3799), .Z(n3818) );
  NAND U3955 ( .A(g_input[0]), .B(n3819), .Z(n3815) );
  NANDN U3956 ( .B(n1722), .A(n3820), .Z(n3819) );
  NANDN U3957 ( .B(n3802), .A(n1729), .Z(n3820) );
  IV U3958 ( .A(n1623), .Z(n1722) );
  XNOR U3959 ( .A(n3707), .B(n3708), .Z(n3704) );
  NAND U3960 ( .A(n3797), .B(n1527), .Z(n3708) );
  XNOR U3961 ( .A(n3706), .B(n3823), .Z(n3707) );
  ANDN U3962 ( .A(n1532), .B(n3799), .Z(n3823) );
  NAND U3963 ( .A(g_input[0]), .B(n3824), .Z(n3706) );
  NANDN U3964 ( .B(n1527), .A(n3825), .Z(n3824) );
  NANDN U3965 ( .B(n3802), .A(n1532), .Z(n3825) );
  IV U3966 ( .A(n1431), .Z(n1527) );
  XNOR U3967 ( .A(n3828), .B(n3829), .Z(n3730) );
  XOR U3968 ( .A(n3830), .B(n2952), .Z(n2947) );
  XNOR U3969 ( .A(n2943), .B(n2944), .Z(n2952) );
  NAND U3970 ( .A(n2940), .B(n572), .Z(n2944) );
  XNOR U3971 ( .A(n2942), .B(n3831), .Z(n2943) );
  ANDN U3972 ( .A(n2945), .B(n574), .Z(n3831) );
  XOR U3973 ( .A(n3832), .B(n3833), .Z(n2942) );
  AND U3974 ( .A(n3834), .B(n3835), .Z(n3833) );
  XOR U3975 ( .A(n3836), .B(n3832), .Z(n3835) );
  XNOR U3976 ( .A(n2950), .B(n2946), .Z(n3830) );
  XNOR U3977 ( .A(n3061), .B(n3060), .Z(n3073) );
  XOR U3978 ( .A(n3838), .B(n3056), .Z(n3060) );
  XNOR U3979 ( .A(n3054), .B(n3839), .Z(n3056) );
  ANDN U3980 ( .A(n2667), .B(n702), .Z(n3839) );
  XOR U3981 ( .A(n3840), .B(n3841), .Z(n3054) );
  AND U3982 ( .A(n3842), .B(n3843), .Z(n3841) );
  XNOR U3983 ( .A(n3844), .B(n3840), .Z(n3843) );
  AND U3984 ( .A(n2660), .B(n700), .Z(n3058) );
  XNOR U3985 ( .A(n3065), .B(n3067), .Z(n3061) );
  NAND U3986 ( .A(n2413), .B(n801), .Z(n3067) );
  XNOR U3987 ( .A(n3063), .B(n3848), .Z(n3065) );
  ANDN U3988 ( .A(n2418), .B(n803), .Z(n3848) );
  XOR U3989 ( .A(n3849), .B(n3850), .Z(n3063) );
  AND U3990 ( .A(n3851), .B(n3852), .Z(n3850) );
  XOR U3991 ( .A(n3853), .B(n3849), .Z(n3852) );
  XOR U3992 ( .A(n3854), .B(n3855), .Z(n3074) );
  XNOR U3993 ( .A(n3856), .B(n3837), .Z(n3854) );
  XOR U3994 ( .A(n3858), .B(n3859), .Z(n3112) );
  XOR U3995 ( .A(n3860), .B(n3857), .Z(n3858) );
  XNOR U3996 ( .A(n3847), .B(n3846), .Z(n3110) );
  XOR U3997 ( .A(n3861), .B(n3842), .Z(n3846) );
  XNOR U3998 ( .A(n3840), .B(n3862), .Z(n3842) );
  ANDN U3999 ( .A(n2667), .B(n744), .Z(n3862) );
  XOR U4000 ( .A(n3863), .B(n3864), .Z(n3840) );
  AND U4001 ( .A(n3865), .B(n3866), .Z(n3864) );
  XNOR U4002 ( .A(n3867), .B(n3863), .Z(n3866) );
  XOR U4003 ( .A(n3868), .B(n3844), .Z(n3861) );
  AND U4004 ( .A(n2660), .B(n742), .Z(n3844) );
  IV U4005 ( .A(n3845), .Z(n3868) );
  XNOR U4006 ( .A(n3851), .B(n3853), .Z(n3847) );
  NAND U4007 ( .A(n2413), .B(n865), .Z(n3853) );
  XNOR U4008 ( .A(n3849), .B(n3872), .Z(n3851) );
  ANDN U4009 ( .A(n2418), .B(n867), .Z(n3872) );
  XOR U4010 ( .A(n3873), .B(n3874), .Z(n3849) );
  AND U4011 ( .A(n3875), .B(n3876), .Z(n3874) );
  XOR U4012 ( .A(n3877), .B(n3873), .Z(n3876) );
  XOR U4013 ( .A(n3879), .B(n3880), .Z(n3157) );
  XOR U4014 ( .A(n3881), .B(n3878), .Z(n3879) );
  XNOR U4015 ( .A(n3871), .B(n3870), .Z(n3155) );
  XOR U4016 ( .A(n3882), .B(n3865), .Z(n3870) );
  XNOR U4017 ( .A(n3863), .B(n3883), .Z(n3865) );
  ANDN U4018 ( .A(n2667), .B(n803), .Z(n3883) );
  XOR U4019 ( .A(n3884), .B(n3885), .Z(n3863) );
  AND U4020 ( .A(n3886), .B(n3887), .Z(n3885) );
  XNOR U4021 ( .A(n3888), .B(n3884), .Z(n3887) );
  XOR U4022 ( .A(n3889), .B(n3867), .Z(n3882) );
  AND U4023 ( .A(n2660), .B(n801), .Z(n3867) );
  IV U4024 ( .A(n3869), .Z(n3889) );
  XNOR U4025 ( .A(n3875), .B(n3877), .Z(n3871) );
  NAND U4026 ( .A(n2413), .B(n933), .Z(n3877) );
  XNOR U4027 ( .A(n3873), .B(n3893), .Z(n3875) );
  ANDN U4028 ( .A(n2418), .B(n935), .Z(n3893) );
  XOR U4029 ( .A(n3894), .B(n3895), .Z(n3873) );
  AND U4030 ( .A(n3896), .B(n3897), .Z(n3895) );
  XOR U4031 ( .A(n3898), .B(n3894), .Z(n3897) );
  XOR U4032 ( .A(n3900), .B(n3901), .Z(n3199) );
  XOR U4033 ( .A(n3902), .B(n3899), .Z(n3900) );
  XNOR U4034 ( .A(n3892), .B(n3891), .Z(n3197) );
  XOR U4035 ( .A(n3903), .B(n3886), .Z(n3891) );
  XNOR U4036 ( .A(n3884), .B(n3904), .Z(n3886) );
  ANDN U4037 ( .A(n2667), .B(n867), .Z(n3904) );
  XOR U4038 ( .A(n3905), .B(n3906), .Z(n3884) );
  AND U4039 ( .A(n3907), .B(n3908), .Z(n3906) );
  XNOR U4040 ( .A(n3909), .B(n3905), .Z(n3908) );
  AND U4041 ( .A(n2660), .B(n865), .Z(n3888) );
  XNOR U4042 ( .A(n3896), .B(n3898), .Z(n3892) );
  NAND U4043 ( .A(n2413), .B(n1000), .Z(n3898) );
  XNOR U4044 ( .A(n3894), .B(n3913), .Z(n3896) );
  ANDN U4045 ( .A(n2418), .B(n1002), .Z(n3913) );
  XOR U4046 ( .A(n3914), .B(n3915), .Z(n3894) );
  AND U4047 ( .A(n3916), .B(n3917), .Z(n3915) );
  XOR U4048 ( .A(n3918), .B(n3914), .Z(n3917) );
  XOR U4049 ( .A(n3920), .B(n3921), .Z(n3242) );
  XOR U4050 ( .A(n3922), .B(n3919), .Z(n3920) );
  XNOR U4051 ( .A(n3912), .B(n3911), .Z(n3240) );
  XOR U4052 ( .A(n3923), .B(n3907), .Z(n3911) );
  XNOR U4053 ( .A(n3905), .B(n3924), .Z(n3907) );
  ANDN U4054 ( .A(n2667), .B(n935), .Z(n3924) );
  XOR U4055 ( .A(n3925), .B(n3926), .Z(n3905) );
  AND U4056 ( .A(n3927), .B(n3928), .Z(n3926) );
  XNOR U4057 ( .A(n3929), .B(n3925), .Z(n3928) );
  XOR U4058 ( .A(n3930), .B(n3909), .Z(n3923) );
  AND U4059 ( .A(n2660), .B(n933), .Z(n3909) );
  IV U4060 ( .A(n3910), .Z(n3930) );
  XNOR U4061 ( .A(n3916), .B(n3918), .Z(n3912) );
  NAND U4062 ( .A(n2413), .B(n1074), .Z(n3918) );
  XNOR U4063 ( .A(n3914), .B(n3934), .Z(n3916) );
  ANDN U4064 ( .A(n2418), .B(n1076), .Z(n3934) );
  XOR U4065 ( .A(n3935), .B(n3936), .Z(n3914) );
  AND U4066 ( .A(n3937), .B(n3938), .Z(n3936) );
  XOR U4067 ( .A(n3939), .B(n3935), .Z(n3938) );
  XOR U4068 ( .A(n3941), .B(n3942), .Z(n3284) );
  XOR U4069 ( .A(n3943), .B(n3940), .Z(n3941) );
  XNOR U4070 ( .A(n3933), .B(n3932), .Z(n3282) );
  XOR U4071 ( .A(n3944), .B(n3927), .Z(n3932) );
  XNOR U4072 ( .A(n3925), .B(n3945), .Z(n3927) );
  ANDN U4073 ( .A(n2667), .B(n1002), .Z(n3945) );
  XOR U4074 ( .A(n3946), .B(n3947), .Z(n3925) );
  AND U4075 ( .A(n3948), .B(n3949), .Z(n3947) );
  XNOR U4076 ( .A(n3950), .B(n3946), .Z(n3949) );
  XOR U4077 ( .A(n3951), .B(n3929), .Z(n3944) );
  AND U4078 ( .A(n2660), .B(n1000), .Z(n3929) );
  IV U4079 ( .A(n3931), .Z(n3951) );
  XNOR U4080 ( .A(n3937), .B(n3939), .Z(n3933) );
  NAND U4081 ( .A(n2413), .B(n1152), .Z(n3939) );
  XNOR U4082 ( .A(n3935), .B(n3955), .Z(n3937) );
  ANDN U4083 ( .A(n2418), .B(n1154), .Z(n3955) );
  XOR U4084 ( .A(n3956), .B(n3957), .Z(n3935) );
  AND U4085 ( .A(n3958), .B(n3959), .Z(n3957) );
  XOR U4086 ( .A(n3960), .B(n3956), .Z(n3959) );
  XOR U4087 ( .A(n3962), .B(n3963), .Z(n3330) );
  XOR U4088 ( .A(n3964), .B(n3961), .Z(n3962) );
  XNOR U4089 ( .A(n3954), .B(n3953), .Z(n3328) );
  XOR U4090 ( .A(n3965), .B(n3948), .Z(n3953) );
  XNOR U4091 ( .A(n3946), .B(n3966), .Z(n3948) );
  ANDN U4092 ( .A(n2667), .B(n1076), .Z(n3966) );
  XOR U4093 ( .A(n3967), .B(n3968), .Z(n3946) );
  AND U4094 ( .A(n3969), .B(n3970), .Z(n3968) );
  XNOR U4095 ( .A(n3971), .B(n3967), .Z(n3970) );
  XOR U4096 ( .A(n3972), .B(n3950), .Z(n3965) );
  AND U4097 ( .A(n2660), .B(n1074), .Z(n3950) );
  IV U4098 ( .A(n3952), .Z(n3972) );
  XNOR U4099 ( .A(n3958), .B(n3960), .Z(n3954) );
  NAND U4100 ( .A(n2413), .B(n1233), .Z(n3960) );
  XNOR U4101 ( .A(n3956), .B(n3976), .Z(n3958) );
  ANDN U4102 ( .A(n2418), .B(n1235), .Z(n3976) );
  XOR U4103 ( .A(n3977), .B(n3978), .Z(n3956) );
  AND U4104 ( .A(n3979), .B(n3980), .Z(n3978) );
  XOR U4105 ( .A(n3981), .B(n3977), .Z(n3980) );
  XOR U4106 ( .A(n3983), .B(n3984), .Z(n3374) );
  XOR U4107 ( .A(n3985), .B(n3982), .Z(n3983) );
  XNOR U4108 ( .A(n3975), .B(n3974), .Z(n3372) );
  XOR U4109 ( .A(n3986), .B(n3969), .Z(n3974) );
  XNOR U4110 ( .A(n3967), .B(n3987), .Z(n3969) );
  ANDN U4111 ( .A(n2667), .B(n1154), .Z(n3987) );
  XOR U4112 ( .A(n3988), .B(n3989), .Z(n3967) );
  AND U4113 ( .A(n3990), .B(n3991), .Z(n3989) );
  XNOR U4114 ( .A(n3992), .B(n3988), .Z(n3991) );
  XOR U4115 ( .A(n3993), .B(n3971), .Z(n3986) );
  AND U4116 ( .A(n2660), .B(n1152), .Z(n3971) );
  IV U4117 ( .A(n3973), .Z(n3993) );
  XNOR U4118 ( .A(n3979), .B(n3981), .Z(n3975) );
  NAND U4119 ( .A(n2413), .B(n1317), .Z(n3981) );
  XNOR U4120 ( .A(n3977), .B(n3997), .Z(n3979) );
  ANDN U4121 ( .A(n2418), .B(n1319), .Z(n3997) );
  XOR U4122 ( .A(n3998), .B(n3999), .Z(n3977) );
  AND U4123 ( .A(n4000), .B(n4001), .Z(n3999) );
  XOR U4124 ( .A(n4002), .B(n3998), .Z(n4001) );
  XOR U4125 ( .A(n4004), .B(n4005), .Z(n3420) );
  XOR U4126 ( .A(n4006), .B(n4003), .Z(n4004) );
  XNOR U4127 ( .A(n3996), .B(n3995), .Z(n3418) );
  XOR U4128 ( .A(n4007), .B(n3990), .Z(n3995) );
  XNOR U4129 ( .A(n3988), .B(n4008), .Z(n3990) );
  ANDN U4130 ( .A(n2667), .B(n1235), .Z(n4008) );
  XOR U4131 ( .A(n4009), .B(n4010), .Z(n3988) );
  AND U4132 ( .A(n4011), .B(n4012), .Z(n4010) );
  XNOR U4133 ( .A(n4013), .B(n4009), .Z(n4012) );
  XOR U4134 ( .A(n4014), .B(n3992), .Z(n4007) );
  AND U4135 ( .A(n2660), .B(n1233), .Z(n3992) );
  IV U4136 ( .A(n3994), .Z(n4014) );
  XNOR U4137 ( .A(n4000), .B(n4002), .Z(n3996) );
  NAND U4138 ( .A(n2413), .B(n1408), .Z(n4002) );
  XNOR U4139 ( .A(n3998), .B(n4018), .Z(n4000) );
  ANDN U4140 ( .A(n2418), .B(n1410), .Z(n4018) );
  XOR U4141 ( .A(n4019), .B(n4020), .Z(n3998) );
  AND U4142 ( .A(n4021), .B(n4022), .Z(n4020) );
  XOR U4143 ( .A(n4023), .B(n4019), .Z(n4022) );
  XOR U4144 ( .A(n4025), .B(n4026), .Z(n3466) );
  XOR U4145 ( .A(n4027), .B(n4024), .Z(n4025) );
  XNOR U4146 ( .A(n4017), .B(n4016), .Z(n3464) );
  XOR U4147 ( .A(n4028), .B(n4011), .Z(n4016) );
  XNOR U4148 ( .A(n4009), .B(n4029), .Z(n4011) );
  ANDN U4149 ( .A(n2667), .B(n1319), .Z(n4029) );
  XOR U4150 ( .A(n4030), .B(n4031), .Z(n4009) );
  AND U4151 ( .A(n4032), .B(n4033), .Z(n4031) );
  XNOR U4152 ( .A(n4034), .B(n4030), .Z(n4033) );
  XOR U4153 ( .A(n4035), .B(n4013), .Z(n4028) );
  AND U4154 ( .A(n2660), .B(n1317), .Z(n4013) );
  IV U4155 ( .A(n4015), .Z(n4035) );
  XNOR U4156 ( .A(n4021), .B(n4023), .Z(n4017) );
  NAND U4157 ( .A(n2413), .B(n1505), .Z(n4023) );
  XNOR U4158 ( .A(n4019), .B(n4039), .Z(n4021) );
  ANDN U4159 ( .A(n2418), .B(n1507), .Z(n4039) );
  XOR U4160 ( .A(n4040), .B(n4041), .Z(n4019) );
  AND U4161 ( .A(n4042), .B(n4043), .Z(n4041) );
  XOR U4162 ( .A(n4044), .B(n4040), .Z(n4043) );
  XOR U4163 ( .A(n4046), .B(n4047), .Z(n3512) );
  XOR U4164 ( .A(n4048), .B(n4045), .Z(n4046) );
  XNOR U4165 ( .A(n4038), .B(n4037), .Z(n3510) );
  XOR U4166 ( .A(n4049), .B(n4032), .Z(n4037) );
  XNOR U4167 ( .A(n4030), .B(n4050), .Z(n4032) );
  ANDN U4168 ( .A(n2667), .B(n1410), .Z(n4050) );
  XOR U4169 ( .A(n4051), .B(n4052), .Z(n4030) );
  AND U4170 ( .A(n4053), .B(n4054), .Z(n4052) );
  XNOR U4171 ( .A(n4055), .B(n4051), .Z(n4054) );
  XOR U4172 ( .A(n4056), .B(n4034), .Z(n4049) );
  AND U4173 ( .A(n2660), .B(n1408), .Z(n4034) );
  IV U4174 ( .A(n4036), .Z(n4056) );
  XNOR U4175 ( .A(n4042), .B(n4044), .Z(n4038) );
  NAND U4176 ( .A(n2413), .B(n1601), .Z(n4044) );
  XNOR U4177 ( .A(n4040), .B(n4060), .Z(n4042) );
  ANDN U4178 ( .A(n2418), .B(n1603), .Z(n4060) );
  XOR U4179 ( .A(n4061), .B(n4062), .Z(n4040) );
  AND U4180 ( .A(n4063), .B(n4064), .Z(n4062) );
  XOR U4181 ( .A(n4065), .B(n4061), .Z(n4064) );
  XOR U4182 ( .A(n4067), .B(n4068), .Z(n3556) );
  XOR U4183 ( .A(n4069), .B(n4066), .Z(n4067) );
  XNOR U4184 ( .A(n4059), .B(n4058), .Z(n3554) );
  XOR U4185 ( .A(n4070), .B(n4053), .Z(n4058) );
  XNOR U4186 ( .A(n4051), .B(n4071), .Z(n4053) );
  ANDN U4187 ( .A(n2667), .B(n1507), .Z(n4071) );
  XOR U4188 ( .A(n4072), .B(n4073), .Z(n4051) );
  AND U4189 ( .A(n4074), .B(n4075), .Z(n4073) );
  XNOR U4190 ( .A(n4076), .B(n4072), .Z(n4075) );
  XOR U4191 ( .A(n4077), .B(n4055), .Z(n4070) );
  AND U4192 ( .A(n2660), .B(n1505), .Z(n4055) );
  IV U4193 ( .A(n4057), .Z(n4077) );
  XNOR U4194 ( .A(n4063), .B(n4065), .Z(n4059) );
  NAND U4195 ( .A(n2413), .B(n1697), .Z(n4065) );
  XNOR U4196 ( .A(n4061), .B(n4081), .Z(n4063) );
  ANDN U4197 ( .A(n2418), .B(n1699), .Z(n4081) );
  XOR U4198 ( .A(n4082), .B(n4083), .Z(n4061) );
  AND U4199 ( .A(n4084), .B(n4085), .Z(n4083) );
  XOR U4200 ( .A(n4086), .B(n4082), .Z(n4085) );
  XOR U4201 ( .A(n4088), .B(n4089), .Z(n3602) );
  XOR U4202 ( .A(n4090), .B(n4087), .Z(n4088) );
  XNOR U4203 ( .A(n4080), .B(n4079), .Z(n3600) );
  XOR U4204 ( .A(n4091), .B(n4074), .Z(n4079) );
  XNOR U4205 ( .A(n4072), .B(n4092), .Z(n4074) );
  ANDN U4206 ( .A(n2667), .B(n1603), .Z(n4092) );
  XOR U4207 ( .A(n4093), .B(n4094), .Z(n4072) );
  AND U4208 ( .A(n4095), .B(n4096), .Z(n4094) );
  XNOR U4209 ( .A(n4097), .B(n4093), .Z(n4096) );
  XOR U4210 ( .A(n4098), .B(n4076), .Z(n4091) );
  AND U4211 ( .A(n2660), .B(n1601), .Z(n4076) );
  IV U4212 ( .A(n4078), .Z(n4098) );
  XNOR U4213 ( .A(n4084), .B(n4086), .Z(n4080) );
  NAND U4214 ( .A(n2413), .B(n1798), .Z(n4086) );
  XNOR U4215 ( .A(n4082), .B(n4102), .Z(n4084) );
  ANDN U4216 ( .A(n2418), .B(n1800), .Z(n4102) );
  XOR U4217 ( .A(n4103), .B(n4104), .Z(n4082) );
  AND U4218 ( .A(n4105), .B(n4106), .Z(n4104) );
  XOR U4219 ( .A(n4107), .B(n4103), .Z(n4106) );
  XOR U4220 ( .A(n4109), .B(n4110), .Z(n3648) );
  XOR U4221 ( .A(n4111), .B(n4108), .Z(n4109) );
  XNOR U4222 ( .A(n4101), .B(n4100), .Z(n3646) );
  XOR U4223 ( .A(n4112), .B(n4095), .Z(n4100) );
  XNOR U4224 ( .A(n4093), .B(n4113), .Z(n4095) );
  ANDN U4225 ( .A(n2667), .B(n1699), .Z(n4113) );
  XOR U4226 ( .A(n4114), .B(n4115), .Z(n4093) );
  AND U4227 ( .A(n4116), .B(n4117), .Z(n4115) );
  XNOR U4228 ( .A(n4118), .B(n4114), .Z(n4117) );
  XOR U4229 ( .A(n4119), .B(n4097), .Z(n4112) );
  AND U4230 ( .A(n2660), .B(n1697), .Z(n4097) );
  IV U4231 ( .A(n4099), .Z(n4119) );
  XNOR U4232 ( .A(n4105), .B(n4107), .Z(n4101) );
  NAND U4233 ( .A(n2413), .B(n1904), .Z(n4107) );
  XNOR U4234 ( .A(n4103), .B(n4123), .Z(n4105) );
  ANDN U4235 ( .A(n2418), .B(n1906), .Z(n4123) );
  XOR U4236 ( .A(n4124), .B(n4125), .Z(n4103) );
  AND U4237 ( .A(n4126), .B(n4127), .Z(n4125) );
  XOR U4238 ( .A(n4128), .B(n4124), .Z(n4127) );
  XOR U4239 ( .A(n4130), .B(n4131), .Z(n3694) );
  XOR U4240 ( .A(n4132), .B(n4129), .Z(n4130) );
  XNOR U4241 ( .A(n4122), .B(n4121), .Z(n3692) );
  XOR U4242 ( .A(n4133), .B(n4116), .Z(n4121) );
  XNOR U4243 ( .A(n4114), .B(n4134), .Z(n4116) );
  ANDN U4244 ( .A(n2667), .B(n1800), .Z(n4134) );
  XOR U4245 ( .A(n4135), .B(n4136), .Z(n4114) );
  AND U4246 ( .A(n4137), .B(n4138), .Z(n4136) );
  XNOR U4247 ( .A(n4139), .B(n4135), .Z(n4138) );
  XOR U4248 ( .A(n4140), .B(n4118), .Z(n4133) );
  AND U4249 ( .A(n2660), .B(n1798), .Z(n4118) );
  IV U4250 ( .A(n4120), .Z(n4140) );
  XNOR U4251 ( .A(n4126), .B(n4128), .Z(n4122) );
  NAND U4252 ( .A(n2413), .B(n2011), .Z(n4128) );
  XNOR U4253 ( .A(n4124), .B(n4144), .Z(n4126) );
  ANDN U4254 ( .A(n2418), .B(n2013), .Z(n4144) );
  XOR U4255 ( .A(n4145), .B(n4146), .Z(n4124) );
  AND U4256 ( .A(n4147), .B(n4148), .Z(n4146) );
  XOR U4257 ( .A(n4149), .B(n4145), .Z(n4148) );
  XOR U4258 ( .A(n4151), .B(n4152), .Z(n3733) );
  XOR U4259 ( .A(n4153), .B(n4150), .Z(n4151) );
  XNOR U4260 ( .A(n4143), .B(n4142), .Z(n3732) );
  XOR U4261 ( .A(n4154), .B(n4137), .Z(n4142) );
  XNOR U4262 ( .A(n4135), .B(n4155), .Z(n4137) );
  ANDN U4263 ( .A(n2667), .B(n1906), .Z(n4155) );
  AND U4264 ( .A(n2660), .B(n1904), .Z(n4139) );
  XNOR U4265 ( .A(n4147), .B(n4149), .Z(n4143) );
  NAND U4266 ( .A(n2413), .B(n2119), .Z(n4149) );
  XNOR U4267 ( .A(n4145), .B(n4162), .Z(n4147) );
  ANDN U4268 ( .A(n2418), .B(n2121), .Z(n4162) );
  XOR U4269 ( .A(n4166), .B(n4167), .Z(n4150) );
  AND U4270 ( .A(n4168), .B(n4169), .Z(n4167) );
  XOR U4271 ( .A(n4170), .B(n4171), .Z(n4169) );
  XNOR U4272 ( .A(n4166), .B(n4172), .Z(n4171) );
  XNOR U4273 ( .A(n4160), .B(n4173), .Z(n4168) );
  XNOR U4274 ( .A(n4166), .B(n4161), .Z(n4173) );
  XNOR U4275 ( .A(n4164), .B(n4165), .Z(n4161) );
  NAND U4276 ( .A(n2238), .B(n2413), .Z(n4165) );
  XNOR U4277 ( .A(n4163), .B(n4174), .Z(n4164) );
  ANDN U4278 ( .A(n2418), .B(n2240), .Z(n4174) );
  XOR U4279 ( .A(n4178), .B(n4157), .Z(n4160) );
  XNOR U4280 ( .A(n4156), .B(n4179), .Z(n4157) );
  ANDN U4281 ( .A(n2667), .B(n2013), .Z(n4179) );
  AND U4282 ( .A(n2660), .B(n2011), .Z(n4158) );
  XOR U4283 ( .A(n4186), .B(n4187), .Z(n4166) );
  AND U4284 ( .A(n4188), .B(n4189), .Z(n4187) );
  XOR U4285 ( .A(n4190), .B(n4191), .Z(n4189) );
  XNOR U4286 ( .A(n4186), .B(n4192), .Z(n4191) );
  XNOR U4287 ( .A(n4184), .B(n4193), .Z(n4188) );
  XNOR U4288 ( .A(n4186), .B(n4185), .Z(n4193) );
  XNOR U4289 ( .A(n4176), .B(n4177), .Z(n4185) );
  NAND U4290 ( .A(n2358), .B(n2413), .Z(n4177) );
  XNOR U4291 ( .A(n4175), .B(n4194), .Z(n4176) );
  ANDN U4292 ( .A(n2418), .B(n2360), .Z(n4194) );
  XOR U4293 ( .A(n4198), .B(n4181), .Z(n4184) );
  XNOR U4294 ( .A(n4180), .B(n4199), .Z(n4181) );
  ANDN U4295 ( .A(n2667), .B(n2121), .Z(n4199) );
  AND U4296 ( .A(n2660), .B(n2119), .Z(n4182) );
  XOR U4297 ( .A(n4206), .B(n4207), .Z(n4186) );
  AND U4298 ( .A(n4208), .B(n4209), .Z(n4207) );
  XOR U4299 ( .A(n4210), .B(n4211), .Z(n4209) );
  XNOR U4300 ( .A(n4206), .B(n4212), .Z(n4211) );
  XNOR U4301 ( .A(n4204), .B(n4213), .Z(n4208) );
  XNOR U4302 ( .A(n4206), .B(n4205), .Z(n4213) );
  XNOR U4303 ( .A(n4196), .B(n4197), .Z(n4205) );
  NAND U4304 ( .A(n2480), .B(n2413), .Z(n4197) );
  XNOR U4305 ( .A(n4195), .B(n4214), .Z(n4196) );
  ANDN U4306 ( .A(n2418), .B(n2482), .Z(n4214) );
  XOR U4307 ( .A(n4218), .B(n4201), .Z(n4204) );
  XNOR U4308 ( .A(n4200), .B(n4219), .Z(n4201) );
  ANDN U4309 ( .A(n2667), .B(n2240), .Z(n4219) );
  AND U4310 ( .A(n2238), .B(n2660), .Z(n4202) );
  XOR U4311 ( .A(n4226), .B(n4227), .Z(n4206) );
  AND U4312 ( .A(n4228), .B(n4229), .Z(n4227) );
  XOR U4313 ( .A(n4230), .B(n4231), .Z(n4229) );
  XNOR U4314 ( .A(n4226), .B(n4232), .Z(n4231) );
  XNOR U4315 ( .A(n4224), .B(n4233), .Z(n4228) );
  XNOR U4316 ( .A(n4226), .B(n4225), .Z(n4233) );
  XNOR U4317 ( .A(n4216), .B(n4217), .Z(n4225) );
  NAND U4318 ( .A(n2605), .B(n2413), .Z(n4217) );
  XNOR U4319 ( .A(n4215), .B(n4234), .Z(n4216) );
  ANDN U4320 ( .A(n2418), .B(n2607), .Z(n4234) );
  XOR U4321 ( .A(n4238), .B(n4221), .Z(n4224) );
  XNOR U4322 ( .A(n4220), .B(n4239), .Z(n4221) );
  ANDN U4323 ( .A(n2667), .B(n2360), .Z(n4239) );
  AND U4324 ( .A(n2358), .B(n2660), .Z(n4222) );
  XOR U4325 ( .A(n4246), .B(n4247), .Z(n4226) );
  AND U4326 ( .A(n4248), .B(n4249), .Z(n4247) );
  XOR U4327 ( .A(n4250), .B(n4251), .Z(n4249) );
  XNOR U4328 ( .A(n4246), .B(n4252), .Z(n4251) );
  XNOR U4329 ( .A(n4244), .B(n4253), .Z(n4248) );
  XNOR U4330 ( .A(n4246), .B(n4245), .Z(n4253) );
  XNOR U4331 ( .A(n4236), .B(n4237), .Z(n4245) );
  NAND U4332 ( .A(n2737), .B(n2413), .Z(n4237) );
  XNOR U4333 ( .A(n4235), .B(n4254), .Z(n4236) );
  ANDN U4334 ( .A(n2418), .B(n2739), .Z(n4254) );
  XOR U4335 ( .A(n4258), .B(n4241), .Z(n4244) );
  XNOR U4336 ( .A(n4240), .B(n4259), .Z(n4241) );
  ANDN U4337 ( .A(n2667), .B(n2482), .Z(n4259) );
  AND U4338 ( .A(n2480), .B(n2660), .Z(n4242) );
  XOR U4339 ( .A(n4266), .B(n4267), .Z(n4246) );
  AND U4340 ( .A(n4268), .B(n4269), .Z(n4267) );
  XOR U4341 ( .A(n4270), .B(n4271), .Z(n4269) );
  XNOR U4342 ( .A(n4266), .B(n4272), .Z(n4271) );
  XNOR U4343 ( .A(n4264), .B(n4273), .Z(n4268) );
  XNOR U4344 ( .A(n4266), .B(n4265), .Z(n4273) );
  XNOR U4345 ( .A(n4256), .B(n4257), .Z(n4265) );
  NAND U4346 ( .A(n2869), .B(n2413), .Z(n4257) );
  XNOR U4347 ( .A(n4255), .B(n4274), .Z(n4256) );
  ANDN U4348 ( .A(n2418), .B(n2871), .Z(n4274) );
  XOR U4349 ( .A(n4275), .B(n4276), .Z(n4255) );
  AND U4350 ( .A(n4277), .B(n4278), .Z(n4276) );
  XOR U4351 ( .A(n4279), .B(n4275), .Z(n4278) );
  XOR U4352 ( .A(n4280), .B(n4261), .Z(n4264) );
  XNOR U4353 ( .A(n4260), .B(n4281), .Z(n4261) );
  ANDN U4354 ( .A(n2667), .B(n2607), .Z(n4281) );
  XOR U4355 ( .A(n4282), .B(n4283), .Z(n4260) );
  AND U4356 ( .A(n4284), .B(n4285), .Z(n4283) );
  XNOR U4357 ( .A(n4286), .B(n4282), .Z(n4285) );
  AND U4358 ( .A(n2605), .B(n2660), .Z(n4262) );
  XOR U4359 ( .A(n4290), .B(n4291), .Z(n4266) );
  AND U4360 ( .A(n4292), .B(n4293), .Z(n4291) );
  XOR U4361 ( .A(n4294), .B(n4295), .Z(n4293) );
  XNOR U4362 ( .A(n4290), .B(n4296), .Z(n4295) );
  XNOR U4363 ( .A(n4288), .B(n4297), .Z(n4292) );
  XNOR U4364 ( .A(n4290), .B(n4289), .Z(n4297) );
  XNOR U4365 ( .A(n4277), .B(n4279), .Z(n4289) );
  NAND U4366 ( .A(n3009), .B(n2413), .Z(n4279) );
  XNOR U4367 ( .A(n4275), .B(n4298), .Z(n4277) );
  ANDN U4368 ( .A(n2418), .B(n3011), .Z(n4298) );
  XOR U4369 ( .A(n4302), .B(n4284), .Z(n4288) );
  XNOR U4370 ( .A(n4282), .B(n4303), .Z(n4284) );
  ANDN U4371 ( .A(n2667), .B(n2739), .Z(n4303) );
  XOR U4372 ( .A(n4304), .B(n4305), .Z(n4282) );
  AND U4373 ( .A(n4306), .B(n4307), .Z(n4305) );
  XNOR U4374 ( .A(n4308), .B(n4304), .Z(n4307) );
  AND U4375 ( .A(n2737), .B(n2660), .Z(n4286) );
  XOR U4376 ( .A(n4313), .B(n4314), .Z(n3829) );
  XNOR U4377 ( .A(n4311), .B(n4310), .Z(n3828) );
  XOR U4378 ( .A(n4316), .B(n4306), .Z(n4310) );
  XNOR U4379 ( .A(n4304), .B(n4317), .Z(n4306) );
  ANDN U4380 ( .A(n2667), .B(n2871), .Z(n4317) );
  XNOR U4381 ( .A(n4320), .B(n4318), .Z(n4319) );
  ANDN U4382 ( .A(n2667), .B(n3011), .Z(n4320) );
  XNOR U4383 ( .A(n4309), .B(n4308), .Z(n4316) );
  AND U4384 ( .A(n2869), .B(n2660), .Z(n4308) );
  XNOR U4385 ( .A(n4322), .B(n4323), .Z(n4309) );
  NAND U4386 ( .A(n3797), .B(n2660), .Z(n4323) );
  XNOR U4387 ( .A(n4321), .B(n4324), .Z(n4322) );
  ANDN U4388 ( .A(n2667), .B(n3799), .Z(n4324) );
  NAND U4389 ( .A(g_input[0]), .B(n4325), .Z(n4321) );
  NANDN U4390 ( .B(n2660), .A(n4326), .Z(n4325) );
  NANDN U4391 ( .B(n3802), .A(n2667), .Z(n4326) );
  IV U4392 ( .A(n2534), .Z(n2660) );
  XNOR U4393 ( .A(n4300), .B(n4301), .Z(n4311) );
  NAND U4394 ( .A(n3797), .B(n2413), .Z(n4301) );
  XNOR U4395 ( .A(n4299), .B(n4329), .Z(n4300) );
  ANDN U4396 ( .A(n2418), .B(n3799), .Z(n4329) );
  NAND U4397 ( .A(g_input[0]), .B(n4330), .Z(n4299) );
  NANDN U4398 ( .B(n2413), .A(n4331), .Z(n4330) );
  NANDN U4399 ( .B(n3802), .A(n2418), .Z(n4331) );
  IV U4400 ( .A(n2292), .Z(n2413) );
  XOR U4401 ( .A(n4334), .B(n4335), .Z(n4312) );
  XOR U4402 ( .A(n2949), .B(n4336), .Z(n2950) );
  AND U4403 ( .A(n4337), .B(n4338), .Z(n4336) );
  NANDN U4404 ( .B(n4339), .A(n511), .Z(n4338) );
  NANDN U4405 ( .B(n4340), .A(n4341), .Z(n4337) );
  XNOR U4406 ( .A(n3834), .B(n3836), .Z(n3855) );
  NAND U4407 ( .A(n2940), .B(n616), .Z(n3836) );
  XNOR U4408 ( .A(n3832), .B(n4343), .Z(n3834) );
  ANDN U4409 ( .A(n2945), .B(n618), .Z(n4343) );
  XOR U4410 ( .A(n4344), .B(n4345), .Z(n3832) );
  AND U4411 ( .A(n4346), .B(n4347), .Z(n4345) );
  XOR U4412 ( .A(n4348), .B(n4344), .Z(n4347) );
  XNOR U4413 ( .A(n4349), .B(n4350), .Z(n3856) );
  IV U4414 ( .A(n4342), .Z(n4350) );
  XOR U4415 ( .A(n4351), .B(n4341), .Z(n4349) );
  AND U4416 ( .A(n4352), .B(n541), .Z(n4341) );
  IV U4417 ( .A(n574), .Z(n541) );
  NAND U4418 ( .A(n4353), .B(n4340), .Z(n4351) );
  XOR U4419 ( .A(n4354), .B(n4355), .Z(n4340) );
  AND U4420 ( .A(n4356), .B(n4357), .Z(n4355) );
  XNOR U4421 ( .A(n4358), .B(n4354), .Z(n4357) );
  NANDN U4422 ( .B(n544), .A(e_input[0]), .Z(n4353) );
  IV U4423 ( .A(n511), .Z(n544) );
  AND U4424 ( .A(n4359), .B(n4360), .Z(n511) );
  ANDN U4425 ( .A(g_input[31]), .B(n4361), .Z(n4359) );
  XNOR U4426 ( .A(n4346), .B(n4348), .Z(n3859) );
  NAND U4427 ( .A(n2940), .B(n656), .Z(n4348) );
  XNOR U4428 ( .A(n4344), .B(n4363), .Z(n4346) );
  ANDN U4429 ( .A(n2945), .B(n658), .Z(n4363) );
  XOR U4430 ( .A(n4364), .B(n4365), .Z(n4344) );
  AND U4431 ( .A(n4366), .B(n4367), .Z(n4365) );
  XOR U4432 ( .A(n4368), .B(n4364), .Z(n4367) );
  XNOR U4433 ( .A(n4369), .B(n4356), .Z(n3860) );
  XNOR U4434 ( .A(n4354), .B(n4370), .Z(n4356) );
  ANDN U4435 ( .A(e_input[0]), .B(n574), .Z(n4370) );
  XNOR U4436 ( .A(n4361), .B(g_input[30]), .Z(n4360) );
  NANDN U4437 ( .B(n4371), .A(n4372), .Z(n4361) );
  XOR U4438 ( .A(n4373), .B(n4374), .Z(n4354) );
  AND U4439 ( .A(n4375), .B(n4376), .Z(n4374) );
  XNOR U4440 ( .A(n4377), .B(n4373), .Z(n4376) );
  XOR U4441 ( .A(n4378), .B(n4358), .Z(n4369) );
  AND U4442 ( .A(n4352), .B(n572), .Z(n4358) );
  IV U4443 ( .A(n618), .Z(n572) );
  IV U4444 ( .A(n4362), .Z(n4378) );
  XNOR U4445 ( .A(n4366), .B(n4368), .Z(n3880) );
  NAND U4446 ( .A(n2940), .B(n700), .Z(n4368) );
  XNOR U4447 ( .A(n4364), .B(n4380), .Z(n4366) );
  ANDN U4448 ( .A(n2945), .B(n702), .Z(n4380) );
  XOR U4449 ( .A(n4381), .B(n4382), .Z(n4364) );
  AND U4450 ( .A(n4383), .B(n4384), .Z(n4382) );
  XOR U4451 ( .A(n4385), .B(n4381), .Z(n4384) );
  XNOR U4452 ( .A(n4386), .B(n4375), .Z(n3881) );
  XNOR U4453 ( .A(n4373), .B(n4387), .Z(n4375) );
  ANDN U4454 ( .A(e_input[0]), .B(n618), .Z(n4387) );
  XNOR U4455 ( .A(n4372), .B(g_input[29]), .Z(n4371) );
  ANDN U4456 ( .A(n4388), .B(n4389), .Z(n4372) );
  XOR U4457 ( .A(n4390), .B(n4391), .Z(n4373) );
  AND U4458 ( .A(n4392), .B(n4393), .Z(n4391) );
  XNOR U4459 ( .A(n4394), .B(n4390), .Z(n4393) );
  XOR U4460 ( .A(n4395), .B(n4377), .Z(n4386) );
  AND U4461 ( .A(n4352), .B(n616), .Z(n4377) );
  IV U4462 ( .A(n658), .Z(n616) );
  IV U4463 ( .A(n4379), .Z(n4395) );
  XNOR U4464 ( .A(n4383), .B(n4385), .Z(n3901) );
  NAND U4465 ( .A(n2940), .B(n742), .Z(n4385) );
  XNOR U4466 ( .A(n4381), .B(n4397), .Z(n4383) );
  ANDN U4467 ( .A(n2945), .B(n744), .Z(n4397) );
  XOR U4468 ( .A(n4398), .B(n4399), .Z(n4381) );
  AND U4469 ( .A(n4400), .B(n4401), .Z(n4399) );
  XOR U4470 ( .A(n4402), .B(n4398), .Z(n4401) );
  XNOR U4471 ( .A(n4403), .B(n4392), .Z(n3902) );
  XNOR U4472 ( .A(n4390), .B(n4404), .Z(n4392) );
  ANDN U4473 ( .A(e_input[0]), .B(n658), .Z(n4404) );
  XNOR U4474 ( .A(n4388), .B(g_input[28]), .Z(n4389) );
  ANDN U4475 ( .A(n4405), .B(n4406), .Z(n4388) );
  XOR U4476 ( .A(n4407), .B(n4408), .Z(n4390) );
  AND U4477 ( .A(n4409), .B(n4410), .Z(n4408) );
  XNOR U4478 ( .A(n4411), .B(n4407), .Z(n4410) );
  AND U4479 ( .A(n4352), .B(n656), .Z(n4394) );
  IV U4480 ( .A(n702), .Z(n656) );
  XNOR U4481 ( .A(n4400), .B(n4402), .Z(n3921) );
  NAND U4482 ( .A(n2940), .B(n801), .Z(n4402) );
  XNOR U4483 ( .A(n4398), .B(n4413), .Z(n4400) );
  ANDN U4484 ( .A(n2945), .B(n803), .Z(n4413) );
  XOR U4485 ( .A(n4414), .B(n4415), .Z(n4398) );
  AND U4486 ( .A(n4416), .B(n4417), .Z(n4415) );
  XOR U4487 ( .A(n4418), .B(n4414), .Z(n4417) );
  XNOR U4488 ( .A(n4419), .B(n4409), .Z(n3922) );
  XNOR U4489 ( .A(n4407), .B(n4420), .Z(n4409) );
  ANDN U4490 ( .A(e_input[0]), .B(n702), .Z(n4420) );
  ANDN U4491 ( .A(n4421), .B(n4422), .Z(n4405) );
  XOR U4492 ( .A(n4423), .B(n4424), .Z(n4407) );
  AND U4493 ( .A(n4425), .B(n4426), .Z(n4424) );
  XNOR U4494 ( .A(n4427), .B(n4423), .Z(n4426) );
  AND U4495 ( .A(n4352), .B(n700), .Z(n4411) );
  IV U4496 ( .A(n744), .Z(n700) );
  XNOR U4497 ( .A(n4416), .B(n4418), .Z(n3942) );
  NAND U4498 ( .A(n2940), .B(n865), .Z(n4418) );
  XNOR U4499 ( .A(n4414), .B(n4429), .Z(n4416) );
  ANDN U4500 ( .A(n2945), .B(n867), .Z(n4429) );
  XOR U4501 ( .A(n4430), .B(n4431), .Z(n4414) );
  AND U4502 ( .A(n4432), .B(n4433), .Z(n4431) );
  XOR U4503 ( .A(n4434), .B(n4430), .Z(n4433) );
  XNOR U4504 ( .A(n4435), .B(n4425), .Z(n3943) );
  XNOR U4505 ( .A(n4423), .B(n4436), .Z(n4425) );
  ANDN U4506 ( .A(e_input[0]), .B(n744), .Z(n4436) );
  XNOR U4507 ( .A(n4421), .B(g_input[26]), .Z(n4422) );
  ANDN U4508 ( .A(n4437), .B(n4438), .Z(n4421) );
  XOR U4509 ( .A(n4439), .B(n4440), .Z(n4423) );
  AND U4510 ( .A(n4441), .B(n4442), .Z(n4440) );
  XNOR U4511 ( .A(n4443), .B(n4439), .Z(n4442) );
  XOR U4512 ( .A(n4444), .B(n4427), .Z(n4435) );
  AND U4513 ( .A(n4352), .B(n742), .Z(n4427) );
  IV U4514 ( .A(n803), .Z(n742) );
  IV U4515 ( .A(n4428), .Z(n4444) );
  XNOR U4516 ( .A(n4432), .B(n4434), .Z(n3963) );
  NAND U4517 ( .A(n2940), .B(n933), .Z(n4434) );
  XNOR U4518 ( .A(n4430), .B(n4446), .Z(n4432) );
  ANDN U4519 ( .A(n2945), .B(n935), .Z(n4446) );
  XOR U4520 ( .A(n4447), .B(n4448), .Z(n4430) );
  AND U4521 ( .A(n4449), .B(n4450), .Z(n4448) );
  XOR U4522 ( .A(n4451), .B(n4447), .Z(n4450) );
  XNOR U4523 ( .A(n4452), .B(n4441), .Z(n3964) );
  XNOR U4524 ( .A(n4439), .B(n4453), .Z(n4441) );
  ANDN U4525 ( .A(e_input[0]), .B(n803), .Z(n4453) );
  ANDN U4526 ( .A(n4454), .B(n4455), .Z(n4437) );
  XOR U4527 ( .A(n4456), .B(n4457), .Z(n4439) );
  AND U4528 ( .A(n4458), .B(n4459), .Z(n4457) );
  XNOR U4529 ( .A(n4460), .B(n4456), .Z(n4459) );
  XOR U4530 ( .A(n4461), .B(n4443), .Z(n4452) );
  AND U4531 ( .A(n4352), .B(n801), .Z(n4443) );
  IV U4532 ( .A(n867), .Z(n801) );
  IV U4533 ( .A(n4445), .Z(n4461) );
  XNOR U4534 ( .A(n4449), .B(n4451), .Z(n3984) );
  NAND U4535 ( .A(n2940), .B(n1000), .Z(n4451) );
  XNOR U4536 ( .A(n4447), .B(n4463), .Z(n4449) );
  ANDN U4537 ( .A(n2945), .B(n1002), .Z(n4463) );
  XOR U4538 ( .A(n4464), .B(n4465), .Z(n4447) );
  AND U4539 ( .A(n4466), .B(n4467), .Z(n4465) );
  XOR U4540 ( .A(n4468), .B(n4464), .Z(n4467) );
  XNOR U4541 ( .A(n4469), .B(n4458), .Z(n3985) );
  XNOR U4542 ( .A(n4456), .B(n4470), .Z(n4458) );
  ANDN U4543 ( .A(e_input[0]), .B(n867), .Z(n4470) );
  XNOR U4544 ( .A(n4454), .B(g_input[24]), .Z(n4455) );
  ANDN U4545 ( .A(n4471), .B(n4472), .Z(n4454) );
  XOR U4546 ( .A(n4473), .B(n4474), .Z(n4456) );
  AND U4547 ( .A(n4475), .B(n4476), .Z(n4474) );
  XNOR U4548 ( .A(n4477), .B(n4473), .Z(n4476) );
  XOR U4549 ( .A(n4478), .B(n4460), .Z(n4469) );
  AND U4550 ( .A(n4352), .B(n865), .Z(n4460) );
  IV U4551 ( .A(n935), .Z(n865) );
  IV U4552 ( .A(n4462), .Z(n4478) );
  XNOR U4553 ( .A(n4466), .B(n4468), .Z(n4005) );
  NAND U4554 ( .A(n2940), .B(n1074), .Z(n4468) );
  XNOR U4555 ( .A(n4464), .B(n4480), .Z(n4466) );
  ANDN U4556 ( .A(n2945), .B(n1076), .Z(n4480) );
  XOR U4557 ( .A(n4481), .B(n4482), .Z(n4464) );
  AND U4558 ( .A(n4483), .B(n4484), .Z(n4482) );
  XOR U4559 ( .A(n4485), .B(n4481), .Z(n4484) );
  XNOR U4560 ( .A(n4486), .B(n4475), .Z(n4006) );
  XNOR U4561 ( .A(n4473), .B(n4487), .Z(n4475) );
  ANDN U4562 ( .A(e_input[0]), .B(n935), .Z(n4487) );
  ANDN U4563 ( .A(n4488), .B(n4489), .Z(n4471) );
  XOR U4564 ( .A(n4490), .B(n4491), .Z(n4473) );
  AND U4565 ( .A(n4492), .B(n4493), .Z(n4491) );
  XNOR U4566 ( .A(n4494), .B(n4490), .Z(n4493) );
  XOR U4567 ( .A(n4495), .B(n4477), .Z(n4486) );
  AND U4568 ( .A(n4352), .B(n933), .Z(n4477) );
  IV U4569 ( .A(n1002), .Z(n933) );
  IV U4570 ( .A(n4479), .Z(n4495) );
  XNOR U4571 ( .A(n4483), .B(n4485), .Z(n4026) );
  NAND U4572 ( .A(n2940), .B(n1152), .Z(n4485) );
  XNOR U4573 ( .A(n4481), .B(n4497), .Z(n4483) );
  ANDN U4574 ( .A(n2945), .B(n1154), .Z(n4497) );
  XOR U4575 ( .A(n4498), .B(n4499), .Z(n4481) );
  AND U4576 ( .A(n4500), .B(n4501), .Z(n4499) );
  XOR U4577 ( .A(n4502), .B(n4498), .Z(n4501) );
  XNOR U4578 ( .A(n4503), .B(n4492), .Z(n4027) );
  XNOR U4579 ( .A(n4490), .B(n4504), .Z(n4492) );
  ANDN U4580 ( .A(e_input[0]), .B(n1002), .Z(n4504) );
  XNOR U4581 ( .A(n4488), .B(g_input[22]), .Z(n4489) );
  ANDN U4582 ( .A(n4505), .B(n4506), .Z(n4488) );
  XOR U4583 ( .A(n4507), .B(n4508), .Z(n4490) );
  AND U4584 ( .A(n4509), .B(n4510), .Z(n4508) );
  XNOR U4585 ( .A(n4511), .B(n4507), .Z(n4510) );
  XOR U4586 ( .A(n4512), .B(n4494), .Z(n4503) );
  AND U4587 ( .A(n4352), .B(n1000), .Z(n4494) );
  IV U4588 ( .A(n1076), .Z(n1000) );
  IV U4589 ( .A(n4496), .Z(n4512) );
  XNOR U4590 ( .A(n4500), .B(n4502), .Z(n4047) );
  NAND U4591 ( .A(n2940), .B(n1233), .Z(n4502) );
  XNOR U4592 ( .A(n4498), .B(n4514), .Z(n4500) );
  ANDN U4593 ( .A(n2945), .B(n1235), .Z(n4514) );
  XOR U4594 ( .A(n4515), .B(n4516), .Z(n4498) );
  AND U4595 ( .A(n4517), .B(n4518), .Z(n4516) );
  XOR U4596 ( .A(n4519), .B(n4515), .Z(n4518) );
  XNOR U4597 ( .A(n4520), .B(n4509), .Z(n4048) );
  XNOR U4598 ( .A(n4507), .B(n4521), .Z(n4509) );
  ANDN U4599 ( .A(e_input[0]), .B(n1076), .Z(n4521) );
  ANDN U4600 ( .A(n4522), .B(n4523), .Z(n4505) );
  XOR U4601 ( .A(n4524), .B(n4525), .Z(n4507) );
  AND U4602 ( .A(n4526), .B(n4527), .Z(n4525) );
  XNOR U4603 ( .A(n4528), .B(n4524), .Z(n4527) );
  XOR U4604 ( .A(n4529), .B(n4511), .Z(n4520) );
  AND U4605 ( .A(n4352), .B(n1074), .Z(n4511) );
  IV U4606 ( .A(n1154), .Z(n1074) );
  IV U4607 ( .A(n4513), .Z(n4529) );
  XNOR U4608 ( .A(n4517), .B(n4519), .Z(n4068) );
  NAND U4609 ( .A(n2940), .B(n1317), .Z(n4519) );
  XNOR U4610 ( .A(n4515), .B(n4531), .Z(n4517) );
  ANDN U4611 ( .A(n2945), .B(n1319), .Z(n4531) );
  XOR U4612 ( .A(n4532), .B(n4533), .Z(n4515) );
  AND U4613 ( .A(n4534), .B(n4535), .Z(n4533) );
  XOR U4614 ( .A(n4536), .B(n4532), .Z(n4535) );
  XNOR U4615 ( .A(n4537), .B(n4526), .Z(n4069) );
  XNOR U4616 ( .A(n4524), .B(n4538), .Z(n4526) );
  ANDN U4617 ( .A(e_input[0]), .B(n1154), .Z(n4538) );
  XNOR U4618 ( .A(n4522), .B(g_input[20]), .Z(n4523) );
  ANDN U4619 ( .A(n4539), .B(n4540), .Z(n4522) );
  XOR U4620 ( .A(n4541), .B(n4542), .Z(n4524) );
  AND U4621 ( .A(n4543), .B(n4544), .Z(n4542) );
  XNOR U4622 ( .A(n4545), .B(n4541), .Z(n4544) );
  XOR U4623 ( .A(n4546), .B(n4528), .Z(n4537) );
  AND U4624 ( .A(n4352), .B(n1152), .Z(n4528) );
  IV U4625 ( .A(n1235), .Z(n1152) );
  IV U4626 ( .A(n4530), .Z(n4546) );
  XNOR U4627 ( .A(n4534), .B(n4536), .Z(n4089) );
  NAND U4628 ( .A(n2940), .B(n1408), .Z(n4536) );
  XNOR U4629 ( .A(n4532), .B(n4548), .Z(n4534) );
  ANDN U4630 ( .A(n2945), .B(n1410), .Z(n4548) );
  XOR U4631 ( .A(n4549), .B(n4550), .Z(n4532) );
  AND U4632 ( .A(n4551), .B(n4552), .Z(n4550) );
  XOR U4633 ( .A(n4553), .B(n4549), .Z(n4552) );
  XNOR U4634 ( .A(n4554), .B(n4543), .Z(n4090) );
  XNOR U4635 ( .A(n4541), .B(n4555), .Z(n4543) );
  ANDN U4636 ( .A(e_input[0]), .B(n1235), .Z(n4555) );
  ANDN U4637 ( .A(n4556), .B(n4557), .Z(n4539) );
  XOR U4638 ( .A(n4558), .B(n4559), .Z(n4541) );
  AND U4639 ( .A(n4560), .B(n4561), .Z(n4559) );
  XNOR U4640 ( .A(n4562), .B(n4558), .Z(n4561) );
  XOR U4641 ( .A(n4563), .B(n4545), .Z(n4554) );
  AND U4642 ( .A(n4352), .B(n1233), .Z(n4545) );
  IV U4643 ( .A(n1319), .Z(n1233) );
  IV U4644 ( .A(n4547), .Z(n4563) );
  XNOR U4645 ( .A(n4551), .B(n4553), .Z(n4110) );
  NAND U4646 ( .A(n2940), .B(n1505), .Z(n4553) );
  XNOR U4647 ( .A(n4549), .B(n4565), .Z(n4551) );
  ANDN U4648 ( .A(n2945), .B(n1507), .Z(n4565) );
  XOR U4649 ( .A(n4566), .B(n4567), .Z(n4549) );
  AND U4650 ( .A(n4568), .B(n4569), .Z(n4567) );
  XOR U4651 ( .A(n4570), .B(n4566), .Z(n4569) );
  XNOR U4652 ( .A(n4571), .B(n4560), .Z(n4111) );
  XNOR U4653 ( .A(n4558), .B(n4572), .Z(n4560) );
  ANDN U4654 ( .A(e_input[0]), .B(n1319), .Z(n4572) );
  XNOR U4655 ( .A(n4556), .B(g_input[18]), .Z(n4557) );
  ANDN U4656 ( .A(n4573), .B(n4574), .Z(n4556) );
  XOR U4657 ( .A(n4575), .B(n4576), .Z(n4558) );
  AND U4658 ( .A(n4577), .B(n4578), .Z(n4576) );
  XNOR U4659 ( .A(n4579), .B(n4575), .Z(n4578) );
  XOR U4660 ( .A(n4580), .B(n4562), .Z(n4571) );
  AND U4661 ( .A(n4352), .B(n1317), .Z(n4562) );
  IV U4662 ( .A(n1410), .Z(n1317) );
  IV U4663 ( .A(n4564), .Z(n4580) );
  XNOR U4664 ( .A(n4568), .B(n4570), .Z(n4131) );
  NAND U4665 ( .A(n2940), .B(n1601), .Z(n4570) );
  XNOR U4666 ( .A(n4566), .B(n4582), .Z(n4568) );
  ANDN U4667 ( .A(n2945), .B(n1603), .Z(n4582) );
  XOR U4668 ( .A(n4583), .B(n4584), .Z(n4566) );
  AND U4669 ( .A(n4585), .B(n4586), .Z(n4584) );
  XOR U4670 ( .A(n4587), .B(n4583), .Z(n4586) );
  XNOR U4671 ( .A(n4588), .B(n4577), .Z(n4132) );
  XNOR U4672 ( .A(n4575), .B(n4589), .Z(n4577) );
  ANDN U4673 ( .A(e_input[0]), .B(n1410), .Z(n4589) );
  ANDN U4674 ( .A(n4590), .B(n4591), .Z(n4573) );
  XOR U4675 ( .A(n4592), .B(n4593), .Z(n4575) );
  AND U4676 ( .A(n4594), .B(n4595), .Z(n4593) );
  XNOR U4677 ( .A(n4596), .B(n4592), .Z(n4595) );
  XOR U4678 ( .A(n4597), .B(n4579), .Z(n4588) );
  AND U4679 ( .A(n4352), .B(n1408), .Z(n4579) );
  IV U4680 ( .A(n1507), .Z(n1408) );
  IV U4681 ( .A(n4581), .Z(n4597) );
  XNOR U4682 ( .A(n4585), .B(n4587), .Z(n4152) );
  NAND U4683 ( .A(n2940), .B(n1697), .Z(n4587) );
  XNOR U4684 ( .A(n4583), .B(n4599), .Z(n4585) );
  ANDN U4685 ( .A(n2945), .B(n1699), .Z(n4599) );
  XNOR U4686 ( .A(n4603), .B(n4594), .Z(n4153) );
  XNOR U4687 ( .A(n4592), .B(n4604), .Z(n4594) );
  ANDN U4688 ( .A(e_input[0]), .B(n1507), .Z(n4604) );
  AND U4689 ( .A(n4352), .B(n1505), .Z(n4596) );
  XNOR U4690 ( .A(n4601), .B(n4602), .Z(n4170) );
  NAND U4691 ( .A(n2940), .B(n1798), .Z(n4602) );
  XNOR U4692 ( .A(n4600), .B(n4609), .Z(n4601) );
  ANDN U4693 ( .A(n2945), .B(n1800), .Z(n4609) );
  XNOR U4694 ( .A(n4613), .B(n4606), .Z(n4172) );
  XNOR U4695 ( .A(n4605), .B(n4614), .Z(n4606) );
  ANDN U4696 ( .A(e_input[0]), .B(n1603), .Z(n4614) );
  AND U4697 ( .A(n4352), .B(n1601), .Z(n4607) );
  XNOR U4698 ( .A(n4611), .B(n4612), .Z(n4190) );
  NAND U4699 ( .A(n2940), .B(n1904), .Z(n4612) );
  XNOR U4700 ( .A(n4610), .B(n4619), .Z(n4611) );
  ANDN U4701 ( .A(n2945), .B(n1906), .Z(n4619) );
  XNOR U4702 ( .A(n4623), .B(n4616), .Z(n4192) );
  XNOR U4703 ( .A(n4615), .B(n4624), .Z(n4616) );
  ANDN U4704 ( .A(e_input[0]), .B(n1699), .Z(n4624) );
  AND U4705 ( .A(n4352), .B(n1697), .Z(n4617) );
  XNOR U4706 ( .A(n4621), .B(n4622), .Z(n4210) );
  NAND U4707 ( .A(n2940), .B(n2011), .Z(n4622) );
  XNOR U4708 ( .A(n4620), .B(n4629), .Z(n4621) );
  ANDN U4709 ( .A(n2945), .B(n2013), .Z(n4629) );
  XNOR U4710 ( .A(n4633), .B(n4626), .Z(n4212) );
  XNOR U4711 ( .A(n4625), .B(n4634), .Z(n4626) );
  ANDN U4712 ( .A(e_input[0]), .B(n1800), .Z(n4634) );
  XOR U4713 ( .A(n4635), .B(n4636), .Z(n4625) );
  AND U4714 ( .A(n4637), .B(n4638), .Z(n4636) );
  XNOR U4715 ( .A(n4639), .B(n4635), .Z(n4638) );
  AND U4716 ( .A(n4352), .B(n1798), .Z(n4627) );
  XNOR U4717 ( .A(n4631), .B(n4632), .Z(n4230) );
  NAND U4718 ( .A(n2940), .B(n2119), .Z(n4632) );
  XNOR U4719 ( .A(n4630), .B(n4641), .Z(n4631) );
  ANDN U4720 ( .A(n2945), .B(n2121), .Z(n4641) );
  XOR U4721 ( .A(n4642), .B(n4643), .Z(n4630) );
  AND U4722 ( .A(n4644), .B(n4645), .Z(n4643) );
  XOR U4723 ( .A(n4646), .B(n4642), .Z(n4645) );
  XNOR U4724 ( .A(n4647), .B(n4637), .Z(n4232) );
  XNOR U4725 ( .A(n4635), .B(n4648), .Z(n4637) );
  ANDN U4726 ( .A(e_input[0]), .B(n1906), .Z(n4648) );
  XOR U4727 ( .A(n4649), .B(n4650), .Z(n4635) );
  AND U4728 ( .A(n4651), .B(n4652), .Z(n4650) );
  XNOR U4729 ( .A(n4653), .B(n4649), .Z(n4652) );
  XOR U4730 ( .A(n4654), .B(n4639), .Z(n4647) );
  AND U4731 ( .A(n4352), .B(n1904), .Z(n4639) );
  IV U4732 ( .A(n4640), .Z(n4654) );
  XNOR U4733 ( .A(n4644), .B(n4646), .Z(n4250) );
  NAND U4734 ( .A(n2940), .B(n2238), .Z(n4646) );
  XNOR U4735 ( .A(n4642), .B(n4656), .Z(n4644) );
  ANDN U4736 ( .A(n2945), .B(n2240), .Z(n4656) );
  XOR U4737 ( .A(n4657), .B(n4658), .Z(n4642) );
  AND U4738 ( .A(n4659), .B(n4660), .Z(n4658) );
  XOR U4739 ( .A(n4661), .B(n4657), .Z(n4660) );
  XNOR U4740 ( .A(n4662), .B(n4651), .Z(n4252) );
  XNOR U4741 ( .A(n4649), .B(n4663), .Z(n4651) );
  ANDN U4742 ( .A(e_input[0]), .B(n2013), .Z(n4663) );
  XOR U4743 ( .A(n4664), .B(n4665), .Z(n4649) );
  AND U4744 ( .A(n4666), .B(n4667), .Z(n4665) );
  XNOR U4745 ( .A(n4668), .B(n4664), .Z(n4667) );
  XOR U4746 ( .A(n4669), .B(n4653), .Z(n4662) );
  AND U4747 ( .A(n4352), .B(n2011), .Z(n4653) );
  IV U4748 ( .A(n4655), .Z(n4669) );
  XNOR U4749 ( .A(n4659), .B(n4661), .Z(n4270) );
  NAND U4750 ( .A(n2940), .B(n2358), .Z(n4661) );
  XNOR U4751 ( .A(n4657), .B(n4671), .Z(n4659) );
  ANDN U4752 ( .A(n2945), .B(n2360), .Z(n4671) );
  XNOR U4753 ( .A(n4675), .B(n4666), .Z(n4272) );
  XNOR U4754 ( .A(n4664), .B(n4676), .Z(n4666) );
  ANDN U4755 ( .A(e_input[0]), .B(n2121), .Z(n4676) );
  XOR U4756 ( .A(n4677), .B(n4678), .Z(n4664) );
  AND U4757 ( .A(n4679), .B(n4680), .Z(n4678) );
  XNOR U4758 ( .A(n4681), .B(n4677), .Z(n4680) );
  AND U4759 ( .A(n4352), .B(n2119), .Z(n4668) );
  XNOR U4760 ( .A(n4673), .B(n4674), .Z(n4294) );
  NAND U4761 ( .A(n2940), .B(n2480), .Z(n4674) );
  XNOR U4762 ( .A(n4672), .B(n4683), .Z(n4673) );
  ANDN U4763 ( .A(n2945), .B(n2482), .Z(n4683) );
  XNOR U4764 ( .A(n4687), .B(n4679), .Z(n4296) );
  XNOR U4765 ( .A(n4677), .B(n4688), .Z(n4679) );
  ANDN U4766 ( .A(e_input[0]), .B(n2240), .Z(n4688) );
  XOR U4767 ( .A(n4689), .B(n4690), .Z(n4677) );
  AND U4768 ( .A(n4691), .B(n4692), .Z(n4690) );
  XNOR U4769 ( .A(n4693), .B(n4689), .Z(n4692) );
  AND U4770 ( .A(n4352), .B(n2238), .Z(n4681) );
  XNOR U4771 ( .A(n4685), .B(n4686), .Z(n4314) );
  NAND U4772 ( .A(n2940), .B(n2605), .Z(n4686) );
  XNOR U4773 ( .A(n4684), .B(n4695), .Z(n4685) );
  ANDN U4774 ( .A(n2945), .B(n2607), .Z(n4695) );
  XNOR U4775 ( .A(n4699), .B(n4691), .Z(n4315) );
  XNOR U4776 ( .A(n4689), .B(n4700), .Z(n4691) );
  ANDN U4777 ( .A(e_input[0]), .B(n2360), .Z(n4700) );
  AND U4778 ( .A(n4352), .B(n2358), .Z(n4693) );
  XNOR U4779 ( .A(n4704), .B(n4705), .Z(n4694) );
  AND U4780 ( .A(n4706), .B(n4707), .Z(n4705) );
  XNOR U4781 ( .A(n4702), .B(n4708), .Z(n4707) );
  XNOR U4782 ( .A(n4703), .B(n4704), .Z(n4708) );
  AND U4783 ( .A(n4352), .B(n2480), .Z(n4703) );
  XOR U4784 ( .A(n4701), .B(n4709), .Z(n4702) );
  ANDN U4785 ( .A(e_input[0]), .B(n2482), .Z(n4709) );
  XNOR U4786 ( .A(n4697), .B(n4713), .Z(n4706) );
  XNOR U4787 ( .A(n4698), .B(n4704), .Z(n4713) );
  AND U4788 ( .A(n2737), .B(n2940), .Z(n4698) );
  XOR U4789 ( .A(n4696), .B(n4714), .Z(n4697) );
  ANDN U4790 ( .A(n2945), .B(n2739), .Z(n4714) );
  XOR U4791 ( .A(n4718), .B(n4719), .Z(n4704) );
  AND U4792 ( .A(n4720), .B(n4721), .Z(n4719) );
  XNOR U4793 ( .A(n4711), .B(n4722), .Z(n4721) );
  XNOR U4794 ( .A(n4712), .B(n4718), .Z(n4722) );
  AND U4795 ( .A(n4352), .B(n2605), .Z(n4712) );
  XOR U4796 ( .A(n4710), .B(n4723), .Z(n4711) );
  ANDN U4797 ( .A(e_input[0]), .B(n2607), .Z(n4723) );
  XNOR U4798 ( .A(n4716), .B(n4727), .Z(n4720) );
  XNOR U4799 ( .A(n4717), .B(n4718), .Z(n4727) );
  AND U4800 ( .A(n2869), .B(n2940), .Z(n4717) );
  XOR U4801 ( .A(n4715), .B(n4728), .Z(n4716) );
  ANDN U4802 ( .A(n2945), .B(n2871), .Z(n4728) );
  XOR U4803 ( .A(n4729), .B(n4730), .Z(n4715) );
  ANDN U4804 ( .A(n4731), .B(n4732), .Z(n4730) );
  XNOR U4805 ( .A(n4733), .B(n4729), .Z(n4731) );
  XOR U4806 ( .A(n4734), .B(n4735), .Z(n4718) );
  AND U4807 ( .A(n4736), .B(n4737), .Z(n4735) );
  XNOR U4808 ( .A(n4725), .B(n4738), .Z(n4737) );
  XNOR U4809 ( .A(n4726), .B(n4734), .Z(n4738) );
  AND U4810 ( .A(n4352), .B(n2737), .Z(n4726) );
  XOR U4811 ( .A(n4724), .B(n4739), .Z(n4725) );
  ANDN U4812 ( .A(e_input[0]), .B(n2739), .Z(n4739) );
  XNOR U4813 ( .A(n4732), .B(n4743), .Z(n4736) );
  XNOR U4814 ( .A(n4733), .B(n4734), .Z(n4743) );
  AND U4815 ( .A(n3009), .B(n2940), .Z(n4733) );
  XOR U4816 ( .A(n4729), .B(n4744), .Z(n4732) );
  ANDN U4817 ( .A(n2945), .B(n3011), .Z(n4744) );
  XNOR U4818 ( .A(n4749), .B(n4741), .Z(n4335) );
  XNOR U4819 ( .A(n4740), .B(n4750), .Z(n4741) );
  ANDN U4820 ( .A(e_input[0]), .B(n2871), .Z(n4750) );
  XNOR U4821 ( .A(n4753), .B(n4751), .Z(n4752) );
  ANDN U4822 ( .A(e_input[0]), .B(n3011), .Z(n4753) );
  ANDN U4823 ( .A(n4352), .B(n3799), .Z(n4754) );
  XNOR U4824 ( .A(n4748), .B(n4742), .Z(n4749) );
  AND U4825 ( .A(n4352), .B(n2869), .Z(n4742) );
  XNOR U4826 ( .A(n4746), .B(n4747), .Z(n4334) );
  NAND U4827 ( .A(n3797), .B(n2940), .Z(n4747) );
  XNOR U4828 ( .A(n4745), .B(n4758), .Z(n4746) );
  ANDN U4829 ( .A(n2945), .B(n3799), .Z(n4758) );
  NAND U4830 ( .A(g_input[0]), .B(n4759), .Z(n4745) );
  NANDN U4831 ( .B(n2940), .A(n4760), .Z(n4759) );
  NANDN U4832 ( .B(n3802), .A(n2945), .Z(n4760) );
  IV U4833 ( .A(n2807), .Z(n2940) );
  XNOR U4834 ( .A(n4756), .B(n4757), .Z(n4748) );
  NAND U4835 ( .A(n3797), .B(n4352), .Z(n4757) );
  XNOR U4836 ( .A(n4755), .B(n4763), .Z(n4756) );
  ANDN U4837 ( .A(e_input[0]), .B(n3799), .Z(n4763) );
  NAND U4838 ( .A(g_input[0]), .B(n4764), .Z(n4755) );
  NANDN U4839 ( .B(n4352), .A(n4765), .Z(n4764) );
  NANDN U4840 ( .B(n3802), .A(e_input[0]), .Z(n4765) );
  IV U4841 ( .A(n4339), .Z(n4352) );
  XNOR U4842 ( .A(n2968), .B(n2967), .Z(n2921) );
  XOR U4843 ( .A(n4767), .B(n2976), .Z(n2967) );
  XNOR U4844 ( .A(n2961), .B(n2960), .Z(n2976) );
  XOR U4845 ( .A(n4768), .B(n2957), .Z(n2960) );
  XNOR U4846 ( .A(n2956), .B(n4769), .Z(n2957) );
  ANDN U4847 ( .A(n1021), .B(n1906), .Z(n4769) );
  AND U4848 ( .A(n1904), .B(n958), .Z(n2958) );
  XNOR U4849 ( .A(n2964), .B(n2965), .Z(n2961) );
  NANDN U4850 ( .B(n823), .A(n2119), .Z(n2965) );
  XNOR U4851 ( .A(n2963), .B(n4776), .Z(n2964) );
  ANDN U4852 ( .A(n893), .B(n2121), .Z(n4776) );
  XOR U4853 ( .A(n2975), .B(n2966), .Z(n4767) );
  XNOR U4854 ( .A(n4780), .B(n4781), .Z(n2966) );
  XOR U4855 ( .A(n4782), .B(n2984), .Z(n2975) );
  XNOR U4856 ( .A(n2972), .B(n2973), .Z(n2984) );
  NAND U4857 ( .A(n1697), .B(n1192), .Z(n2973) );
  XNOR U4858 ( .A(n2971), .B(n4783), .Z(n2972) );
  ANDN U4859 ( .A(n1199), .B(n1699), .Z(n4783) );
  XNOR U4860 ( .A(n2983), .B(n2974), .Z(n4782) );
  XOR U4861 ( .A(n4787), .B(n4788), .Z(n2974) );
  AND U4862 ( .A(n4789), .B(n4790), .Z(n4788) );
  XOR U4863 ( .A(n4791), .B(n4792), .Z(n4790) );
  XNOR U4864 ( .A(n4787), .B(n4793), .Z(n4792) );
  XNOR U4865 ( .A(n4774), .B(n4794), .Z(n4789) );
  XNOR U4866 ( .A(n4787), .B(n4775), .Z(n4794) );
  XNOR U4867 ( .A(n4778), .B(n4779), .Z(n4775) );
  NANDN U4868 ( .B(n823), .A(n2238), .Z(n4779) );
  XNOR U4869 ( .A(n4777), .B(n4795), .Z(n4778) );
  ANDN U4870 ( .A(n893), .B(n2240), .Z(n4795) );
  XOR U4871 ( .A(n4799), .B(n4771), .Z(n4774) );
  XNOR U4872 ( .A(n4770), .B(n4800), .Z(n4771) );
  ANDN U4873 ( .A(n1021), .B(n2013), .Z(n4800) );
  AND U4874 ( .A(n2011), .B(n958), .Z(n4772) );
  XOR U4875 ( .A(n4807), .B(n4808), .Z(n4787) );
  AND U4876 ( .A(n4809), .B(n4810), .Z(n4808) );
  XOR U4877 ( .A(n4811), .B(n4812), .Z(n4810) );
  XNOR U4878 ( .A(n4807), .B(n4813), .Z(n4812) );
  XNOR U4879 ( .A(n4805), .B(n4814), .Z(n4809) );
  XNOR U4880 ( .A(n4807), .B(n4806), .Z(n4814) );
  XNOR U4881 ( .A(n4797), .B(n4798), .Z(n4806) );
  NANDN U4882 ( .B(n823), .A(n2358), .Z(n4798) );
  XNOR U4883 ( .A(n4796), .B(n4815), .Z(n4797) );
  ANDN U4884 ( .A(n893), .B(n2360), .Z(n4815) );
  XOR U4885 ( .A(n4819), .B(n4802), .Z(n4805) );
  XNOR U4886 ( .A(n4801), .B(n4820), .Z(n4802) );
  ANDN U4887 ( .A(n1021), .B(n2121), .Z(n4820) );
  AND U4888 ( .A(n2119), .B(n958), .Z(n4803) );
  XOR U4889 ( .A(n4827), .B(n4828), .Z(n4807) );
  AND U4890 ( .A(n4829), .B(n4830), .Z(n4828) );
  XOR U4891 ( .A(n4831), .B(n4832), .Z(n4830) );
  XNOR U4892 ( .A(n4827), .B(n4833), .Z(n4832) );
  XNOR U4893 ( .A(n4825), .B(n4834), .Z(n4829) );
  XNOR U4894 ( .A(n4827), .B(n4826), .Z(n4834) );
  XNOR U4895 ( .A(n4817), .B(n4818), .Z(n4826) );
  NANDN U4896 ( .B(n823), .A(n2480), .Z(n4818) );
  XNOR U4897 ( .A(n4816), .B(n4835), .Z(n4817) );
  ANDN U4898 ( .A(n893), .B(n2482), .Z(n4835) );
  XOR U4899 ( .A(n4839), .B(n4822), .Z(n4825) );
  XNOR U4900 ( .A(n4821), .B(n4840), .Z(n4822) );
  ANDN U4901 ( .A(n1021), .B(n2240), .Z(n4840) );
  AND U4902 ( .A(n2238), .B(n958), .Z(n4823) );
  XOR U4903 ( .A(n4847), .B(n4848), .Z(n4827) );
  AND U4904 ( .A(n4849), .B(n4850), .Z(n4848) );
  XOR U4905 ( .A(n4851), .B(n4852), .Z(n4850) );
  XNOR U4906 ( .A(n4847), .B(n4853), .Z(n4852) );
  XNOR U4907 ( .A(n4845), .B(n4854), .Z(n4849) );
  XNOR U4908 ( .A(n4847), .B(n4846), .Z(n4854) );
  XNOR U4909 ( .A(n4837), .B(n4838), .Z(n4846) );
  NANDN U4910 ( .B(n823), .A(n2605), .Z(n4838) );
  XNOR U4911 ( .A(n4836), .B(n4855), .Z(n4837) );
  ANDN U4912 ( .A(n893), .B(n2607), .Z(n4855) );
  XOR U4913 ( .A(n4859), .B(n4842), .Z(n4845) );
  XNOR U4914 ( .A(n4841), .B(n4860), .Z(n4842) );
  ANDN U4915 ( .A(n1021), .B(n2360), .Z(n4860) );
  AND U4916 ( .A(n2358), .B(n958), .Z(n4843) );
  XOR U4917 ( .A(n4867), .B(n4868), .Z(n4847) );
  AND U4918 ( .A(n4869), .B(n4870), .Z(n4868) );
  XOR U4919 ( .A(n4871), .B(n4872), .Z(n4870) );
  XNOR U4920 ( .A(n4867), .B(n4873), .Z(n4872) );
  XNOR U4921 ( .A(n4865), .B(n4874), .Z(n4869) );
  XNOR U4922 ( .A(n4867), .B(n4866), .Z(n4874) );
  XNOR U4923 ( .A(n4857), .B(n4858), .Z(n4866) );
  NANDN U4924 ( .B(n823), .A(n2737), .Z(n4858) );
  XNOR U4925 ( .A(n4856), .B(n4875), .Z(n4857) );
  ANDN U4926 ( .A(n893), .B(n2739), .Z(n4875) );
  XOR U4927 ( .A(n4879), .B(n4862), .Z(n4865) );
  XNOR U4928 ( .A(n4861), .B(n4880), .Z(n4862) );
  ANDN U4929 ( .A(n1021), .B(n2482), .Z(n4880) );
  XOR U4930 ( .A(n4881), .B(n4882), .Z(n4861) );
  AND U4931 ( .A(n4883), .B(n4884), .Z(n4882) );
  XNOR U4932 ( .A(n4885), .B(n4881), .Z(n4884) );
  AND U4933 ( .A(n2480), .B(n958), .Z(n4863) );
  XOR U4934 ( .A(n4889), .B(n4890), .Z(n4867) );
  AND U4935 ( .A(n4891), .B(n4892), .Z(n4890) );
  XOR U4936 ( .A(n4893), .B(n4894), .Z(n4892) );
  XNOR U4937 ( .A(n4889), .B(n4895), .Z(n4894) );
  XNOR U4938 ( .A(n4887), .B(n4896), .Z(n4891) );
  XNOR U4939 ( .A(n4889), .B(n4888), .Z(n4896) );
  XNOR U4940 ( .A(n4877), .B(n4878), .Z(n4888) );
  NANDN U4941 ( .B(n823), .A(n2869), .Z(n4878) );
  XNOR U4942 ( .A(n4876), .B(n4897), .Z(n4877) );
  ANDN U4943 ( .A(n893), .B(n2871), .Z(n4897) );
  XOR U4944 ( .A(n4898), .B(n4899), .Z(n4876) );
  AND U4945 ( .A(n4900), .B(n4901), .Z(n4899) );
  XOR U4946 ( .A(n4902), .B(n4898), .Z(n4901) );
  XOR U4947 ( .A(n4903), .B(n4883), .Z(n4887) );
  XNOR U4948 ( .A(n4881), .B(n4904), .Z(n4883) );
  ANDN U4949 ( .A(n1021), .B(n2607), .Z(n4904) );
  XOR U4950 ( .A(n4905), .B(n4906), .Z(n4881) );
  AND U4951 ( .A(n4907), .B(n4908), .Z(n4906) );
  XNOR U4952 ( .A(n4909), .B(n4905), .Z(n4908) );
  AND U4953 ( .A(n2605), .B(n958), .Z(n4885) );
  XOR U4954 ( .A(n4913), .B(n4914), .Z(n4889) );
  AND U4955 ( .A(n4915), .B(n4916), .Z(n4914) );
  XOR U4956 ( .A(n4917), .B(n4918), .Z(n4916) );
  XNOR U4957 ( .A(n4913), .B(n4919), .Z(n4918) );
  XNOR U4958 ( .A(n4911), .B(n4920), .Z(n4915) );
  XNOR U4959 ( .A(n4913), .B(n4912), .Z(n4920) );
  XNOR U4960 ( .A(n4900), .B(n4902), .Z(n4912) );
  NANDN U4961 ( .B(n823), .A(n3009), .Z(n4902) );
  XNOR U4962 ( .A(n4898), .B(n4921), .Z(n4900) );
  ANDN U4963 ( .A(n893), .B(n3011), .Z(n4921) );
  XOR U4964 ( .A(n4925), .B(n4907), .Z(n4911) );
  XNOR U4965 ( .A(n4905), .B(n4926), .Z(n4907) );
  ANDN U4966 ( .A(n1021), .B(n2739), .Z(n4926) );
  AND U4967 ( .A(n2737), .B(n958), .Z(n4909) );
  XOR U4968 ( .A(n4934), .B(n4935), .Z(n4781) );
  XNOR U4969 ( .A(n4932), .B(n4931), .Z(n4780) );
  XOR U4970 ( .A(n4937), .B(n4928), .Z(n4931) );
  XNOR U4971 ( .A(n4927), .B(n4938), .Z(n4928) );
  ANDN U4972 ( .A(n1021), .B(n2871), .Z(n4938) );
  XNOR U4973 ( .A(n4941), .B(n4939), .Z(n4940) );
  ANDN U4974 ( .A(n1021), .B(n3011), .Z(n4941) );
  XNOR U4975 ( .A(n4930), .B(n4929), .Z(n4937) );
  AND U4976 ( .A(n2869), .B(n958), .Z(n4929) );
  XNOR U4977 ( .A(n4944), .B(n4945), .Z(n4930) );
  NAND U4978 ( .A(n3797), .B(n958), .Z(n4945) );
  XNOR U4979 ( .A(n4943), .B(n4946), .Z(n4944) );
  ANDN U4980 ( .A(n1021), .B(n3799), .Z(n4946) );
  NAND U4981 ( .A(g_input[0]), .B(n4947), .Z(n4943) );
  NANDN U4982 ( .B(n958), .A(n4948), .Z(n4947) );
  NANDN U4983 ( .B(n3802), .A(n1021), .Z(n4948) );
  IV U4984 ( .A(n4942), .Z(n958) );
  XNOR U4985 ( .A(n4923), .B(n4924), .Z(n4932) );
  NANDN U4986 ( .B(n823), .A(n3797), .Z(n4924) );
  XNOR U4987 ( .A(n4922), .B(n4951), .Z(n4923) );
  ANDN U4988 ( .A(n893), .B(n3799), .Z(n4951) );
  NAND U4989 ( .A(g_input[0]), .B(n4952), .Z(n4922) );
  NAND U4990 ( .A(n4953), .B(n823), .Z(n4952) );
  NANDN U4991 ( .B(n3802), .A(n893), .Z(n4953) );
  XOR U4992 ( .A(n4956), .B(n4957), .Z(n4933) );
  XOR U4993 ( .A(n4958), .B(n2980), .Z(n2983) );
  XNOR U4994 ( .A(n2979), .B(n4959), .Z(n2980) );
  ANDN U4995 ( .A(n1383), .B(n1507), .Z(n4959) );
  XNOR U4996 ( .A(n4590), .B(g_input[16]), .Z(n4591) );
  ANDN U4997 ( .A(n4960), .B(n4961), .Z(n4590) );
  AND U4998 ( .A(n1505), .B(n1376), .Z(n2981) );
  IV U4999 ( .A(n1603), .Z(n1505) );
  XNOR U5000 ( .A(n4785), .B(n4786), .Z(n4791) );
  NAND U5001 ( .A(n1798), .B(n1192), .Z(n4786) );
  XNOR U5002 ( .A(n4784), .B(n4966), .Z(n4785) );
  ANDN U5003 ( .A(n1199), .B(n1800), .Z(n4966) );
  XNOR U5004 ( .A(n4970), .B(n4963), .Z(n4793) );
  XNOR U5005 ( .A(n4962), .B(n4971), .Z(n4963) );
  ANDN U5006 ( .A(n1383), .B(n1603), .Z(n4971) );
  ANDN U5007 ( .A(n4972), .B(n4973), .Z(n4960) );
  AND U5008 ( .A(n1601), .B(n1376), .Z(n4964) );
  IV U5009 ( .A(n1699), .Z(n1601) );
  XNOR U5010 ( .A(n4968), .B(n4969), .Z(n4811) );
  NAND U5011 ( .A(n1904), .B(n1192), .Z(n4969) );
  XNOR U5012 ( .A(n4967), .B(n4978), .Z(n4968) );
  ANDN U5013 ( .A(n1199), .B(n1906), .Z(n4978) );
  XNOR U5014 ( .A(n4982), .B(n4975), .Z(n4813) );
  XNOR U5015 ( .A(n4974), .B(n4983), .Z(n4975) );
  ANDN U5016 ( .A(n1383), .B(n1699), .Z(n4983) );
  XNOR U5017 ( .A(n4972), .B(g_input[14]), .Z(n4973) );
  ANDN U5018 ( .A(n4984), .B(n4985), .Z(n4972) );
  AND U5019 ( .A(n1697), .B(n1376), .Z(n4976) );
  IV U5020 ( .A(n1800), .Z(n1697) );
  XNOR U5021 ( .A(n4980), .B(n4981), .Z(n4831) );
  NAND U5022 ( .A(n2011), .B(n1192), .Z(n4981) );
  XNOR U5023 ( .A(n4979), .B(n4990), .Z(n4980) );
  ANDN U5024 ( .A(n1199), .B(n2013), .Z(n4990) );
  XNOR U5025 ( .A(n4994), .B(n4987), .Z(n4833) );
  XNOR U5026 ( .A(n4986), .B(n4995), .Z(n4987) );
  ANDN U5027 ( .A(n1383), .B(n1800), .Z(n4995) );
  ANDN U5028 ( .A(n4996), .B(n4997), .Z(n4984) );
  AND U5029 ( .A(n1798), .B(n1376), .Z(n4988) );
  IV U5030 ( .A(n1906), .Z(n1798) );
  XNOR U5031 ( .A(n4992), .B(n4993), .Z(n4851) );
  NAND U5032 ( .A(n2119), .B(n1192), .Z(n4993) );
  XNOR U5033 ( .A(n4991), .B(n5002), .Z(n4992) );
  ANDN U5034 ( .A(n1199), .B(n2121), .Z(n5002) );
  XNOR U5035 ( .A(n5006), .B(n4999), .Z(n4853) );
  XNOR U5036 ( .A(n4998), .B(n5007), .Z(n4999) );
  ANDN U5037 ( .A(n1383), .B(n1906), .Z(n5007) );
  XNOR U5038 ( .A(n4996), .B(g_input[12]), .Z(n4997) );
  ANDN U5039 ( .A(n5008), .B(n5009), .Z(n4996) );
  AND U5040 ( .A(n1904), .B(n1376), .Z(n5000) );
  IV U5041 ( .A(n2013), .Z(n1904) );
  XNOR U5042 ( .A(n5004), .B(n5005), .Z(n4871) );
  NAND U5043 ( .A(n2238), .B(n1192), .Z(n5005) );
  XNOR U5044 ( .A(n5003), .B(n5014), .Z(n5004) );
  ANDN U5045 ( .A(n1199), .B(n2240), .Z(n5014) );
  XOR U5046 ( .A(n5015), .B(n5016), .Z(n5003) );
  AND U5047 ( .A(n5017), .B(n5018), .Z(n5016) );
  XOR U5048 ( .A(n5019), .B(n5015), .Z(n5018) );
  XNOR U5049 ( .A(n5020), .B(n5011), .Z(n4873) );
  XNOR U5050 ( .A(n5010), .B(n5021), .Z(n5011) );
  ANDN U5051 ( .A(n1383), .B(n2013), .Z(n5021) );
  ANDN U5052 ( .A(n5022), .B(n5023), .Z(n5008) );
  AND U5053 ( .A(n2011), .B(n1376), .Z(n5012) );
  IV U5054 ( .A(n2121), .Z(n2011) );
  XNOR U5055 ( .A(n5017), .B(n5019), .Z(n4893) );
  NAND U5056 ( .A(n2358), .B(n1192), .Z(n5019) );
  XNOR U5057 ( .A(n5015), .B(n5028), .Z(n5017) );
  ANDN U5058 ( .A(n1199), .B(n2360), .Z(n5028) );
  XOR U5059 ( .A(n5029), .B(n5030), .Z(n5015) );
  AND U5060 ( .A(n5031), .B(n5032), .Z(n5030) );
  XOR U5061 ( .A(n5033), .B(n5029), .Z(n5032) );
  XNOR U5062 ( .A(n5034), .B(n5025), .Z(n4895) );
  XNOR U5063 ( .A(n5024), .B(n5035), .Z(n5025) );
  ANDN U5064 ( .A(n1383), .B(n2121), .Z(n5035) );
  XNOR U5065 ( .A(n5022), .B(g_input[10]), .Z(n5023) );
  ANDN U5066 ( .A(n5036), .B(n5037), .Z(n5022) );
  XOR U5067 ( .A(n5038), .B(n5039), .Z(n5024) );
  AND U5068 ( .A(n5040), .B(n5041), .Z(n5039) );
  XNOR U5069 ( .A(n5042), .B(n5038), .Z(n5041) );
  XOR U5070 ( .A(n5043), .B(n5026), .Z(n5034) );
  AND U5071 ( .A(n2119), .B(n1376), .Z(n5026) );
  IV U5072 ( .A(n2240), .Z(n2119) );
  IV U5073 ( .A(n5027), .Z(n5043) );
  XNOR U5074 ( .A(n5031), .B(n5033), .Z(n4917) );
  NAND U5075 ( .A(n2480), .B(n1192), .Z(n5033) );
  XNOR U5076 ( .A(n5029), .B(n5045), .Z(n5031) );
  ANDN U5077 ( .A(n1199), .B(n2482), .Z(n5045) );
  XNOR U5078 ( .A(n5049), .B(n5040), .Z(n4919) );
  XNOR U5079 ( .A(n5038), .B(n5050), .Z(n5040) );
  ANDN U5080 ( .A(n1383), .B(n2240), .Z(n5050) );
  ANDN U5081 ( .A(n5051), .B(n5052), .Z(n5036) );
  XOR U5082 ( .A(n5053), .B(n5054), .Z(n5038) );
  AND U5083 ( .A(n5055), .B(n5056), .Z(n5054) );
  XNOR U5084 ( .A(n5057), .B(n5053), .Z(n5056) );
  AND U5085 ( .A(n2238), .B(n1376), .Z(n5042) );
  IV U5086 ( .A(n2360), .Z(n2238) );
  XNOR U5087 ( .A(n5047), .B(n5048), .Z(n4935) );
  NAND U5088 ( .A(n2605), .B(n1192), .Z(n5048) );
  XNOR U5089 ( .A(n5046), .B(n5059), .Z(n5047) );
  ANDN U5090 ( .A(n1199), .B(n2607), .Z(n5059) );
  XNOR U5091 ( .A(n5063), .B(n5055), .Z(n4936) );
  XNOR U5092 ( .A(n5053), .B(n5064), .Z(n5055) );
  ANDN U5093 ( .A(n1383), .B(n2360), .Z(n5064) );
  AND U5094 ( .A(n2358), .B(n1376), .Z(n5057) );
  XNOR U5095 ( .A(n5068), .B(n5069), .Z(n5058) );
  AND U5096 ( .A(n5070), .B(n5071), .Z(n5069) );
  XNOR U5097 ( .A(n5066), .B(n5072), .Z(n5071) );
  XNOR U5098 ( .A(n5067), .B(n5068), .Z(n5072) );
  AND U5099 ( .A(n2480), .B(n1376), .Z(n5067) );
  XOR U5100 ( .A(n5065), .B(n5073), .Z(n5066) );
  ANDN U5101 ( .A(n1383), .B(n2482), .Z(n5073) );
  XNOR U5102 ( .A(n5061), .B(n5077), .Z(n5070) );
  XNOR U5103 ( .A(n5062), .B(n5068), .Z(n5077) );
  AND U5104 ( .A(n2737), .B(n1192), .Z(n5062) );
  XOR U5105 ( .A(n5060), .B(n5078), .Z(n5061) );
  ANDN U5106 ( .A(n1199), .B(n2739), .Z(n5078) );
  XOR U5107 ( .A(n5082), .B(n5083), .Z(n5068) );
  AND U5108 ( .A(n5084), .B(n5085), .Z(n5083) );
  XNOR U5109 ( .A(n5075), .B(n5086), .Z(n5085) );
  XNOR U5110 ( .A(n5076), .B(n5082), .Z(n5086) );
  AND U5111 ( .A(n2605), .B(n1376), .Z(n5076) );
  XOR U5112 ( .A(n5074), .B(n5087), .Z(n5075) );
  ANDN U5113 ( .A(n1383), .B(n2607), .Z(n5087) );
  XNOR U5114 ( .A(n5080), .B(n5091), .Z(n5084) );
  XNOR U5115 ( .A(n5081), .B(n5082), .Z(n5091) );
  AND U5116 ( .A(n2869), .B(n1192), .Z(n5081) );
  XOR U5117 ( .A(n5079), .B(n5092), .Z(n5080) );
  ANDN U5118 ( .A(n1199), .B(n2871), .Z(n5092) );
  XOR U5119 ( .A(n5093), .B(n5094), .Z(n5079) );
  ANDN U5120 ( .A(n5095), .B(n5096), .Z(n5094) );
  XNOR U5121 ( .A(n5097), .B(n5093), .Z(n5095) );
  XOR U5122 ( .A(n5098), .B(n5099), .Z(n5082) );
  AND U5123 ( .A(n5100), .B(n5101), .Z(n5099) );
  XNOR U5124 ( .A(n5089), .B(n5102), .Z(n5101) );
  XNOR U5125 ( .A(n5090), .B(n5098), .Z(n5102) );
  AND U5126 ( .A(n2737), .B(n1376), .Z(n5090) );
  XOR U5127 ( .A(n5088), .B(n5103), .Z(n5089) );
  ANDN U5128 ( .A(n1383), .B(n2739), .Z(n5103) );
  XNOR U5129 ( .A(n5096), .B(n5107), .Z(n5100) );
  XNOR U5130 ( .A(n5097), .B(n5098), .Z(n5107) );
  AND U5131 ( .A(n3009), .B(n1192), .Z(n5097) );
  XOR U5132 ( .A(n5093), .B(n5108), .Z(n5096) );
  ANDN U5133 ( .A(n1199), .B(n3011), .Z(n5108) );
  XNOR U5134 ( .A(n5113), .B(n5105), .Z(n4957) );
  XNOR U5135 ( .A(n5104), .B(n5114), .Z(n5105) );
  ANDN U5136 ( .A(n1383), .B(n2871), .Z(n5114) );
  XNOR U5137 ( .A(n5117), .B(n5115), .Z(n5116) );
  ANDN U5138 ( .A(n1383), .B(n3011), .Z(n5117) );
  XNOR U5139 ( .A(n5112), .B(n5106), .Z(n5113) );
  AND U5140 ( .A(n2869), .B(n1376), .Z(n5106) );
  XNOR U5141 ( .A(n5110), .B(n5111), .Z(n4956) );
  NAND U5142 ( .A(n3797), .B(n1192), .Z(n5111) );
  XNOR U5143 ( .A(n5109), .B(n5121), .Z(n5110) );
  ANDN U5144 ( .A(n1199), .B(n3799), .Z(n5121) );
  NAND U5145 ( .A(g_input[0]), .B(n5122), .Z(n5109) );
  NANDN U5146 ( .B(n1192), .A(n5123), .Z(n5122) );
  NANDN U5147 ( .B(n3802), .A(n1199), .Z(n5123) );
  IV U5148 ( .A(n1118), .Z(n1192) );
  XNOR U5149 ( .A(n5119), .B(n5120), .Z(n5112) );
  NAND U5150 ( .A(n3797), .B(n1376), .Z(n5120) );
  XNOR U5151 ( .A(n5118), .B(n5126), .Z(n5119) );
  ANDN U5152 ( .A(n1383), .B(n3799), .Z(n5126) );
  NAND U5153 ( .A(g_input[0]), .B(n5127), .Z(n5118) );
  NANDN U5154 ( .B(n1376), .A(n5128), .Z(n5127) );
  NANDN U5155 ( .B(n3802), .A(n1383), .Z(n5128) );
  IV U5156 ( .A(n1283), .Z(n1376) );
  XNOR U5157 ( .A(n2992), .B(n2991), .Z(n2968) );
  XOR U5158 ( .A(n5131), .B(n3000), .Z(n2991) );
  XNOR U5159 ( .A(n2988), .B(n2989), .Z(n3000) );
  NANDN U5160 ( .B(n636), .A(n2605), .Z(n2989) );
  XNOR U5161 ( .A(n2987), .B(n5132), .Z(n2988) );
  ANDN U5162 ( .A(n677), .B(n2607), .Z(n5132) );
  XOR U5163 ( .A(n2999), .B(n2990), .Z(n5131) );
  XOR U5164 ( .A(n5136), .B(n5137), .Z(n2990) );
  XOR U5165 ( .A(n5138), .B(n2996), .Z(n2999) );
  XNOR U5166 ( .A(n2995), .B(n5139), .Z(n2996) );
  ANDN U5167 ( .A(n784), .B(n2360), .Z(n5139) );
  XNOR U5168 ( .A(n5051), .B(g_input[8]), .Z(n5052) );
  ANDN U5169 ( .A(n5140), .B(n5141), .Z(n5051) );
  AND U5170 ( .A(n2358), .B(n730), .Z(n2997) );
  IV U5171 ( .A(n2482), .Z(n2358) );
  XNOR U5172 ( .A(n5145), .B(n5146), .Z(n2998) );
  AND U5173 ( .A(n5147), .B(n5148), .Z(n5146) );
  XNOR U5174 ( .A(n5143), .B(n5149), .Z(n5148) );
  XNOR U5175 ( .A(n5144), .B(n5145), .Z(n5149) );
  AND U5176 ( .A(n2480), .B(n730), .Z(n5144) );
  IV U5177 ( .A(n2607), .Z(n2480) );
  XOR U5178 ( .A(n5142), .B(n5150), .Z(n5143) );
  ANDN U5179 ( .A(n784), .B(n2482), .Z(n5150) );
  ANDN U5180 ( .A(n5151), .B(n5152), .Z(n5140) );
  XNOR U5181 ( .A(n5134), .B(n5156), .Z(n5147) );
  XNOR U5182 ( .A(n5135), .B(n5145), .Z(n5156) );
  ANDN U5183 ( .A(n2737), .B(n636), .Z(n5135) );
  XOR U5184 ( .A(n5133), .B(n5157), .Z(n5134) );
  ANDN U5185 ( .A(n677), .B(n2739), .Z(n5157) );
  XOR U5186 ( .A(n5161), .B(n5162), .Z(n5145) );
  AND U5187 ( .A(n5163), .B(n5164), .Z(n5162) );
  XNOR U5188 ( .A(n5154), .B(n5165), .Z(n5164) );
  XNOR U5189 ( .A(n5155), .B(n5161), .Z(n5165) );
  AND U5190 ( .A(n2605), .B(n730), .Z(n5155) );
  IV U5191 ( .A(n2739), .Z(n2605) );
  XOR U5192 ( .A(n5153), .B(n5166), .Z(n5154) );
  ANDN U5193 ( .A(n784), .B(n2607), .Z(n5166) );
  XNOR U5194 ( .A(n5151), .B(g_input[6]), .Z(n5152) );
  ANDN U5195 ( .A(n5167), .B(n5168), .Z(n5151) );
  XNOR U5196 ( .A(n5159), .B(n5172), .Z(n5163) );
  XNOR U5197 ( .A(n5160), .B(n5161), .Z(n5172) );
  ANDN U5198 ( .A(n2869), .B(n636), .Z(n5160) );
  XOR U5199 ( .A(n5158), .B(n5173), .Z(n5159) );
  ANDN U5200 ( .A(n677), .B(n2871), .Z(n5173) );
  XOR U5201 ( .A(n5174), .B(n5175), .Z(n5158) );
  ANDN U5202 ( .A(n5176), .B(n5177), .Z(n5175) );
  XNOR U5203 ( .A(n5178), .B(n5174), .Z(n5176) );
  XOR U5204 ( .A(n5179), .B(n5180), .Z(n5161) );
  AND U5205 ( .A(n5181), .B(n5182), .Z(n5180) );
  XNOR U5206 ( .A(n5170), .B(n5183), .Z(n5182) );
  XNOR U5207 ( .A(n5171), .B(n5179), .Z(n5183) );
  AND U5208 ( .A(n2737), .B(n730), .Z(n5171) );
  XOR U5209 ( .A(n5169), .B(n5184), .Z(n5170) );
  ANDN U5210 ( .A(n784), .B(n2739), .Z(n5184) );
  ANDN U5211 ( .A(n5185), .B(n5186), .Z(n5167) );
  XNOR U5212 ( .A(n5177), .B(n5190), .Z(n5181) );
  XNOR U5213 ( .A(n5178), .B(n5179), .Z(n5190) );
  ANDN U5214 ( .A(n3009), .B(n636), .Z(n5178) );
  XOR U5215 ( .A(n5174), .B(n5191), .Z(n5177) );
  ANDN U5216 ( .A(n677), .B(n3011), .Z(n5191) );
  XNOR U5217 ( .A(n5196), .B(n5188), .Z(n5137) );
  XNOR U5218 ( .A(n5187), .B(n5197), .Z(n5188) );
  ANDN U5219 ( .A(n784), .B(n2871), .Z(n5197) );
  XNOR U5220 ( .A(n5200), .B(n5198), .Z(n5199) );
  ANDN U5221 ( .A(n784), .B(n3011), .Z(n5200) );
  XNOR U5222 ( .A(n5195), .B(n5189), .Z(n5196) );
  AND U5223 ( .A(n2869), .B(n730), .Z(n5189) );
  XNOR U5224 ( .A(n5193), .B(n5194), .Z(n5136) );
  NANDN U5225 ( .B(n636), .A(n3797), .Z(n5194) );
  XNOR U5226 ( .A(n5192), .B(n5205), .Z(n5193) );
  ANDN U5227 ( .A(n677), .B(n3799), .Z(n5205) );
  NAND U5228 ( .A(g_input[0]), .B(n5206), .Z(n5192) );
  NAND U5229 ( .A(n5207), .B(n636), .Z(n5206) );
  NANDN U5230 ( .B(n3802), .A(n677), .Z(n5207) );
  XNOR U5231 ( .A(n5203), .B(n5204), .Z(n5195) );
  NAND U5232 ( .A(n3797), .B(n730), .Z(n5204) );
  XNOR U5233 ( .A(n5202), .B(n5210), .Z(n5203) );
  ANDN U5234 ( .A(n784), .B(n3799), .Z(n5210) );
  NAND U5235 ( .A(g_input[0]), .B(n5211), .Z(n5202) );
  NANDN U5236 ( .B(n730), .A(n5212), .Z(n5211) );
  NANDN U5237 ( .B(n3802), .A(n784), .Z(n5212) );
  IV U5238 ( .A(n5201), .Z(n730) );
  XOR U5239 ( .A(n3008), .B(n3007), .Z(n2992) );
  XOR U5240 ( .A(n5215), .B(n3004), .Z(n3007) );
  XNOR U5241 ( .A(n3003), .B(n5216), .Z(n3004) );
  ANDN U5242 ( .A(n609), .B(n2871), .Z(n5216) );
  IV U5243 ( .A(n2737), .Z(n2871) );
  XNOR U5244 ( .A(n5185), .B(g_input[4]), .Z(n5186) );
  ANDN U5245 ( .A(n5217), .B(n5218), .Z(n5185) );
  XNOR U5246 ( .A(n5221), .B(n5219), .Z(n5220) );
  ANDN U5247 ( .A(n609), .B(n3011), .Z(n5221) );
  IV U5248 ( .A(n2869), .Z(n3011) );
  IV U5249 ( .A(n3799), .Z(n3009) );
  XNOR U5250 ( .A(n3006), .B(n3005), .Z(n5215) );
  AND U5251 ( .A(n2869), .B(n568), .Z(n3005) );
  ANDN U5252 ( .A(n5226), .B(n5227), .Z(n5217) );
  XNOR U5253 ( .A(n5224), .B(n5225), .Z(n3006) );
  NAND U5254 ( .A(n3797), .B(n568), .Z(n5225) );
  XNOR U5255 ( .A(n5223), .B(n5228), .Z(n5224) );
  ANDN U5256 ( .A(n609), .B(n3799), .Z(n5228) );
  NAND U5257 ( .A(g_input[0]), .B(n5229), .Z(n5223) );
  NANDN U5258 ( .B(n568), .A(n5230), .Z(n5229) );
  NANDN U5259 ( .B(n3802), .A(n609), .Z(n5230) );
  IV U5260 ( .A(n5222), .Z(n568) );
  XOR U5261 ( .A(n3015), .B(n3014), .Z(n3008) );
  NAND U5262 ( .A(n3797), .B(n512), .Z(n3014) );
  IV U5263 ( .A(n3802), .Z(n3797) );
  XOR U5264 ( .A(n3013), .B(n5233), .Z(n3015) );
  ANDN U5265 ( .A(n543), .B(n3799), .Z(n5233) );
  XNOR U5266 ( .A(n5226), .B(g_input[2]), .Z(n5227) );
  NOR U5267 ( .A(g_input[0]), .B(n5234), .Z(n5226) );
  NANDN U5268 ( .B(n512), .A(n5236), .Z(n5235) );
  NANDN U5269 ( .B(n3802), .A(n543), .Z(n5236) );
  XOR U5270 ( .A(g_input[0]), .B(g_input[1]), .Z(n5234) );
  AND U5271 ( .A(n5238), .B(n5237), .Z(n512) );
  ANDN U5272 ( .A(e_input[31]), .B(n5239), .Z(n5238) );
  NANDN U5273 ( .B(n5240), .A(n5232), .Z(n5239) );
  XNOR U5274 ( .A(n5240), .B(e_input[29]), .Z(n5232) );
  NAND U5275 ( .A(n5231), .B(n5241), .Z(n5240) );
  XOR U5276 ( .A(n5241), .B(e_input[28]), .Z(n5231) );
  ANDN U5277 ( .A(n5208), .B(n5242), .Z(n5241) );
  XNOR U5278 ( .A(n5242), .B(e_input[27]), .Z(n5208) );
  NAND U5279 ( .A(n5209), .B(n5243), .Z(n5242) );
  XOR U5280 ( .A(n5243), .B(e_input[26]), .Z(n5209) );
  ANDN U5281 ( .A(n5214), .B(n5244), .Z(n5243) );
  XNOR U5282 ( .A(n5244), .B(e_input[25]), .Z(n5214) );
  NAND U5283 ( .A(n5213), .B(n5245), .Z(n5244) );
  XOR U5284 ( .A(n5245), .B(e_input[24]), .Z(n5213) );
  ANDN U5285 ( .A(n4954), .B(n5246), .Z(n5245) );
  XNOR U5286 ( .A(n5246), .B(e_input[23]), .Z(n4954) );
  NAND U5287 ( .A(n4955), .B(n5247), .Z(n5246) );
  XOR U5288 ( .A(n5247), .B(e_input[22]), .Z(n4955) );
  ANDN U5289 ( .A(n4950), .B(n5248), .Z(n5247) );
  XNOR U5290 ( .A(n5248), .B(e_input[21]), .Z(n4950) );
  NAND U5291 ( .A(n4949), .B(n5249), .Z(n5248) );
  XOR U5292 ( .A(n5249), .B(e_input[20]), .Z(n4949) );
  ANDN U5293 ( .A(n5125), .B(n5250), .Z(n5249) );
  XNOR U5294 ( .A(n5250), .B(e_input[19]), .Z(n5125) );
  NAND U5295 ( .A(n5124), .B(n5251), .Z(n5250) );
  XOR U5296 ( .A(n5251), .B(e_input[18]), .Z(n5124) );
  ANDN U5297 ( .A(n5130), .B(n5252), .Z(n5251) );
  XNOR U5298 ( .A(n5252), .B(e_input[17]), .Z(n5130) );
  NAND U5299 ( .A(n5129), .B(n5253), .Z(n5252) );
  XOR U5300 ( .A(n5253), .B(e_input[16]), .Z(n5129) );
  ANDN U5301 ( .A(n3827), .B(n5254), .Z(n5253) );
  XNOR U5302 ( .A(n5254), .B(e_input[15]), .Z(n3827) );
  NAND U5303 ( .A(n3826), .B(n5255), .Z(n5254) );
  XOR U5304 ( .A(n5255), .B(e_input[14]), .Z(n3826) );
  ANDN U5305 ( .A(n3822), .B(n5256), .Z(n5255) );
  XNOR U5306 ( .A(n5256), .B(e_input[13]), .Z(n3822) );
  NAND U5307 ( .A(n3821), .B(n5257), .Z(n5256) );
  XOR U5308 ( .A(n5257), .B(e_input[12]), .Z(n3821) );
  ANDN U5309 ( .A(n3804), .B(n5258), .Z(n5257) );
  XNOR U5310 ( .A(n5258), .B(e_input[11]), .Z(n3804) );
  NAND U5311 ( .A(n3803), .B(n5259), .Z(n5258) );
  XOR U5312 ( .A(n5259), .B(e_input[10]), .Z(n3803) );
  ANDN U5313 ( .A(n3809), .B(n5260), .Z(n5259) );
  XNOR U5314 ( .A(n5260), .B(e_input[9]), .Z(n3809) );
  NAND U5315 ( .A(n3808), .B(n5261), .Z(n5260) );
  XOR U5316 ( .A(n5261), .B(e_input[8]), .Z(n3808) );
  ANDN U5317 ( .A(n4333), .B(n5262), .Z(n5261) );
  XNOR U5318 ( .A(n5262), .B(e_input[7]), .Z(n4333) );
  NAND U5319 ( .A(n4332), .B(n5263), .Z(n5262) );
  XOR U5320 ( .A(n5263), .B(e_input[6]), .Z(n4332) );
  ANDN U5321 ( .A(n4328), .B(n5264), .Z(n5263) );
  XNOR U5322 ( .A(n5264), .B(e_input[5]), .Z(n4328) );
  NAND U5323 ( .A(n4327), .B(n5265), .Z(n5264) );
  XOR U5324 ( .A(n5265), .B(e_input[4]), .Z(n4327) );
  ANDN U5325 ( .A(n4762), .B(n5266), .Z(n5265) );
  XNOR U5326 ( .A(n5266), .B(e_input[3]), .Z(n4762) );
  NAND U5327 ( .A(n4761), .B(n5267), .Z(n5266) );
  XOR U5328 ( .A(n5267), .B(e_input[2]), .Z(n4761) );
  NOR U5329 ( .A(n4766), .B(e_input[0]), .Z(n5267) );
  XOR U5330 ( .A(e_input[0]), .B(e_input[1]), .Z(n4766) );
  AND U5331 ( .A(n5268), .B(n5269), .Z(\_MxM/N24 ) );
  XOR U5332 ( .A(\_MxM/n[9] ), .B(\_MxM/add_39/carry[9] ), .Z(n5269) );
  AND U5333 ( .A(\_MxM/N13 ), .B(n5268), .Z(\_MxM/N23 ) );
  AND U5334 ( .A(\_MxM/N12 ), .B(n5268), .Z(\_MxM/N22 ) );
  AND U5335 ( .A(\_MxM/N11 ), .B(n5268), .Z(\_MxM/N21 ) );
  AND U5336 ( .A(\_MxM/N10 ), .B(n5268), .Z(\_MxM/N20 ) );
  AND U5337 ( .A(\_MxM/N9 ), .B(n5268), .Z(\_MxM/N19 ) );
  AND U5338 ( .A(\_MxM/N8 ), .B(n5268), .Z(\_MxM/N18 ) );
  AND U5339 ( .A(\_MxM/N7 ), .B(n5268), .Z(\_MxM/N17 ) );
  AND U5340 ( .A(\_MxM/N6 ), .B(n5268), .Z(\_MxM/N16 ) );
  NAND U5341 ( .A(n5270), .B(n5271), .Z(n5268) );
  AND U5342 ( .A(n5272), .B(n5273), .Z(n5271) );
  AND U5343 ( .A(\_MxM/n[1] ), .B(n5274), .Z(n5273) );
  NOR U5344 ( .A(\_MxM/N15 ), .B(n2885), .Z(n5274) );
  OR U5345 ( .A(\_MxM/n[3] ), .B(\_MxM/n[4] ), .Z(n2885) );
  AND U5346 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n5272) );
  AND U5347 ( .A(n5275), .B(n5276), .Z(n5270) );
  AND U5348 ( .A(\_MxM/n[6] ), .B(\_MxM/n[7] ), .Z(n5276) );
  AND U5349 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n5275) );
  IV U5350 ( .A(\_MxM/n[0] ), .Z(\_MxM/N15 ) );
endmodule

