
module MxM_W32_N10000 ( clk, rst, A, X, Y );
  input [31:0] A;
  input [31:0] X;
  output [31:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         \add_25/carry[13] , \add_25/carry[12] , \add_25/carry[11] ,
         \add_25/carry[10] , \add_25/carry[9] , \add_25/carry[8] ,
         \add_25/carry[7] , \add_25/carry[6] , \add_25/carry[5] ,
         \add_25/carry[4] , \add_25/carry[3] , \add_25/carry[2] , n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673;
  wire   [31:0] Y0;
  wire   [13:0] n;

  DFF \n_reg[0]  ( .D(n390), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n389), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n388), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n387), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n386), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n385), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n384), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \n_reg[7]  ( .D(n383), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[7]) );
  DFF \n_reg[8]  ( .D(n382), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[8]) );
  DFF \n_reg[9]  ( .D(n381), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[9]) );
  DFF \n_reg[10]  ( .D(n380), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[10]) );
  DFF \n_reg[11]  ( .D(n379), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[11]) );
  DFF \n_reg[12]  ( .D(n378), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[12]) );
  DFF \n_reg[13]  ( .D(n377), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[13]) );
  DFF \Y0_reg[0]  ( .D(n376), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n375), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n374), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n373), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n372), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n371), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n370), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n369), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y0_reg[8]  ( .D(n368), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[8]) );
  DFF \Y0_reg[9]  ( .D(n367), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[9]) );
  DFF \Y0_reg[10]  ( .D(n366), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[10]) );
  DFF \Y0_reg[11]  ( .D(n365), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[11]) );
  DFF \Y0_reg[12]  ( .D(n364), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[12]) );
  DFF \Y0_reg[13]  ( .D(n363), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[13]) );
  DFF \Y0_reg[14]  ( .D(n362), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[14]) );
  DFF \Y0_reg[15]  ( .D(n361), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[15]) );
  DFF \Y0_reg[16]  ( .D(n360), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[16]) );
  DFF \Y0_reg[17]  ( .D(n359), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[17]) );
  DFF \Y0_reg[18]  ( .D(n358), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[18]) );
  DFF \Y0_reg[19]  ( .D(n357), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[19]) );
  DFF \Y0_reg[20]  ( .D(n356), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[20]) );
  DFF \Y0_reg[21]  ( .D(n355), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[21]) );
  DFF \Y0_reg[22]  ( .D(n354), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[22]) );
  DFF \Y0_reg[23]  ( .D(n353), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[23]) );
  DFF \Y0_reg[24]  ( .D(n352), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[24]) );
  DFF \Y0_reg[25]  ( .D(n351), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[25]) );
  DFF \Y0_reg[26]  ( .D(n350), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[26]) );
  DFF \Y0_reg[27]  ( .D(n349), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[27]) );
  DFF \Y0_reg[28]  ( .D(n348), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[28]) );
  DFF \Y0_reg[29]  ( .D(n347), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[29]) );
  DFF \Y0_reg[30]  ( .D(n346), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[30]) );
  DFF \Y0_reg[31]  ( .D(n345), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[31]) );
  DFF \Y_reg[31]  ( .D(n344), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[31]) );
  DFF \Y_reg[30]  ( .D(n343), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[30]) );
  DFF \Y_reg[29]  ( .D(n342), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[29]) );
  DFF \Y_reg[28]  ( .D(n341), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[28]) );
  DFF \Y_reg[27]  ( .D(n340), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[27]) );
  DFF \Y_reg[26]  ( .D(n339), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[26]) );
  DFF \Y_reg[25]  ( .D(n338), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[25]) );
  DFF \Y_reg[24]  ( .D(n337), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[24]) );
  DFF \Y_reg[23]  ( .D(n336), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[23]) );
  DFF \Y_reg[22]  ( .D(n335), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[22]) );
  DFF \Y_reg[21]  ( .D(n334), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[21]) );
  DFF \Y_reg[20]  ( .D(n333), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[20]) );
  DFF \Y_reg[19]  ( .D(n332), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[19]) );
  DFF \Y_reg[18]  ( .D(n331), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[18]) );
  DFF \Y_reg[17]  ( .D(n330), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[17]) );
  DFF \Y_reg[16]  ( .D(n329), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[16]) );
  DFF \Y_reg[15]  ( .D(n328), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[15]) );
  DFF \Y_reg[14]  ( .D(n327), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[14]) );
  DFF \Y_reg[13]  ( .D(n326), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[13]) );
  DFF \Y_reg[12]  ( .D(n325), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[12]) );
  DFF \Y_reg[11]  ( .D(n324), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[11]) );
  DFF \Y_reg[10]  ( .D(n323), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[10]) );
  DFF \Y_reg[9]  ( .D(n322), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[9]) );
  DFF \Y_reg[8]  ( .D(n321), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[8]) );
  DFF \Y_reg[7]  ( .D(n320), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n319), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n318), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n317), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n316), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n315), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n314), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n313), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  HADDER \add_25/U1_1_6  ( .IN0(n[6]), .IN1(\add_25/carry[6] ), .COUT(
        \add_25/carry[7] ), .SUM(N13) );
  HADDER \add_25/U1_1_7  ( .IN0(n[7]), .IN1(\add_25/carry[7] ), .COUT(
        \add_25/carry[8] ), .SUM(N14) );
  HADDER \add_25/U1_1_8  ( .IN0(n[8]), .IN1(\add_25/carry[8] ), .COUT(
        \add_25/carry[9] ), .SUM(N15) );
  HADDER \add_25/U1_1_9  ( .IN0(n[9]), .IN1(\add_25/carry[9] ), .COUT(
        \add_25/carry[10] ), .SUM(N16) );
  HADDER \add_25/U1_1_10  ( .IN0(n[10]), .IN1(\add_25/carry[10] ), .COUT(
        \add_25/carry[11] ), .SUM(N17) );
  HADDER \add_25/U1_1_11  ( .IN0(n[11]), .IN1(\add_25/carry[11] ), .COUT(
        \add_25/carry[12] ), .SUM(N18) );
  HADDER \add_25/U1_1_12  ( .IN0(n[12]), .IN1(\add_25/carry[12] ), .COUT(
        \add_25/carry[13] ), .SUM(N19) );
  MUX U393 ( .IN0(n4104), .IN1(n391), .SEL(n4105), .F(n4058) );
  IV U394 ( .A(n4106), .Z(n391) );
  MUX U395 ( .IN0(n3932), .IN1(n3934), .SEL(n3933), .F(n3886) );
  MUX U396 ( .IN0(n4705), .IN1(n4707), .SEL(n4706), .F(n4681) );
  MUX U397 ( .IN0(n3757), .IN1(n3759), .SEL(n3758), .F(n3711) );
  XNOR U398 ( .A(n4693), .B(n4692), .Z(n4708) );
  XNOR U399 ( .A(n5076), .B(n5074), .Z(n5081) );
  MUX U400 ( .IN0(n3661), .IN1(n3663), .SEL(n3662), .F(n3618) );
  MUX U401 ( .IN0(n5409), .IN1(n5411), .SEL(n5410), .F(n5397) );
  MUX U402 ( .IN0(n5267), .IN1(n392), .SEL(n5268), .F(n5247) );
  IV U403 ( .A(n5269), .Z(n392) );
  MUX U404 ( .IN0(n5416), .IN1(n393), .SEL(n5417), .F(n5404) );
  IV U405 ( .A(n5418), .Z(n393) );
  MUX U406 ( .IN0(n4626), .IN1(n394), .SEL(n4627), .F(n4606) );
  IV U407 ( .A(n4628), .Z(n394) );
  XNOR U408 ( .A(n3614), .B(n3613), .Z(n3650) );
  MUX U409 ( .IN0(n5031), .IN1(n395), .SEL(n5032), .F(n5021) );
  IV U410 ( .A(n5033), .Z(n395) );
  XNOR U411 ( .A(n3639), .B(n3637), .Z(n3674) );
  XNOR U412 ( .A(n4802), .B(n4800), .Z(n4809) );
  NANDN U413 ( .B(n1688), .A(n3415), .Z(n408) );
  MUX U414 ( .IN0(n3491), .IN1(n3493), .SEL(n3492), .F(n3452) );
  MUX U415 ( .IN0(n3484), .IN1(n396), .SEL(n3485), .F(n3445) );
  IV U416 ( .A(n3486), .Z(n396) );
  MUX U417 ( .IN0(n3496), .IN1(n3498), .SEL(n3497), .F(n3425) );
  MUX U418 ( .IN0(n1399), .IN1(n397), .SEL(n1400), .F(n1330) );
  IV U419 ( .A(n1401), .Z(n397) );
  MUX U420 ( .IN0(n1696), .IN1(n1698), .SEL(n1697), .F(n1612) );
  MUX U421 ( .IN0(n1751), .IN1(n398), .SEL(n1752), .F(n1660) );
  IV U422 ( .A(n1753), .Z(n398) );
  MUX U423 ( .IN0(n1799), .IN1(n399), .SEL(n1800), .F(n1704) );
  IV U424 ( .A(n1801), .Z(n399) );
  MUX U425 ( .IN0(n1904), .IN1(n400), .SEL(n1905), .F(n1807) );
  IV U426 ( .A(n1906), .Z(n400) );
  MUX U427 ( .IN0(n2163), .IN1(n2165), .SEL(n2164), .F(n2062) );
  MUX U428 ( .IN0(n2279), .IN1(n401), .SEL(n2280), .F(n2171) );
  IV U429 ( .A(n2281), .Z(n401) );
  MUX U430 ( .IN0(n2452), .IN1(n402), .SEL(n2453), .F(n2343) );
  IV U431 ( .A(n2454), .Z(n402) );
  MUX U432 ( .IN0(A[29]), .IN1(n4778), .SEL(A[31]), .F(n403) );
  IV U433 ( .A(n403), .Z(n1023) );
  MUX U434 ( .IN0(n404), .IN1(n4766), .SEL(A[31]), .F(n979) );
  IV U435 ( .A(A[30]), .Z(n404) );
  MUX U436 ( .IN0(n5328), .IN1(n5330), .SEL(n5329), .F(n5304) );
  MUX U437 ( .IN0(n5078), .IN1(n5080), .SEL(n5079), .F(n5063) );
  XNOR U438 ( .A(n5450), .B(n5448), .Z(n5455) );
  MUX U439 ( .IN0(n4661), .IN1(n4663), .SEL(n4662), .F(n4641) );
  MUX U440 ( .IN0(n4666), .IN1(n405), .SEL(n4667), .F(n4646) );
  IV U441 ( .A(n4668), .Z(n405) );
  XNOR U442 ( .A(n5316), .B(n5315), .Z(n5331) );
  MUX U443 ( .IN0(n5397), .IN1(n5399), .SEL(n5398), .F(n5385) );
  MUX U444 ( .IN0(n5247), .IN1(n406), .SEL(n5248), .F(n5227) );
  IV U445 ( .A(n5249), .Z(n406) );
  MUX U446 ( .IN0(n5404), .IN1(n407), .SEL(n5405), .F(n5392) );
  IV U447 ( .A(n5406), .Z(n407) );
  MUX U448 ( .IN0(n3576), .IN1(n3578), .SEL(n3577), .F(n3531) );
  XNOR U449 ( .A(n5034), .B(n5033), .Z(n5039) );
  MUX U450 ( .IN0(n5026), .IN1(n5028), .SEL(n5027), .F(n5016) );
  MUX U451 ( .IN0(n5521), .IN1(n408), .SEL(n5522), .F(n5510) );
  XNOR U452 ( .A(n3527), .B(n3526), .Z(n3565) );
  MUX U453 ( .IN0(n5011), .IN1(n409), .SEL(n5012), .F(n4998) );
  IV U454 ( .A(n5013), .Z(n409) );
  MUX U455 ( .IN0(n3445), .IN1(n410), .SEL(n3446), .F(n3315) );
  IV U456 ( .A(n3447), .Z(n410) );
  MUX U457 ( .IN0(n1551), .IN1(n411), .SEL(n1552), .F(n1471) );
  IV U458 ( .A(n1553), .Z(n411) );
  MUX U459 ( .IN0(n1612), .IN1(n1614), .SEL(n1613), .F(n1531) );
  MUX U460 ( .IN0(n1669), .IN1(n1671), .SEL(n1670), .F(n1587) );
  MUX U461 ( .IN0(n1984), .IN1(n1986), .SEL(n1985), .F(n1888) );
  MUX U462 ( .IN0(n1992), .IN1(n412), .SEL(n1993), .F(n1896) );
  IV U463 ( .A(n1994), .Z(n412) );
  MUX U464 ( .IN0(n2000), .IN1(n413), .SEL(n2001), .F(n1904) );
  IV U465 ( .A(n2002), .Z(n413) );
  MUX U466 ( .IN0(n2047), .IN1(n414), .SEL(n2048), .F(n1947) );
  IV U467 ( .A(n2049), .Z(n414) );
  MUX U468 ( .IN0(n2244), .IN1(n2246), .SEL(n2245), .F(n2136) );
  MUX U469 ( .IN0(n2386), .IN1(n415), .SEL(n2387), .F(n2279) );
  IV U470 ( .A(n2388), .Z(n415) );
  MUX U471 ( .IN0(n2566), .IN1(n416), .SEL(n2567), .F(n2452) );
  IV U472 ( .A(n2568), .Z(n416) );
  MUX U473 ( .IN0(n3192), .IN1(n417), .SEL(n3193), .F(n3067) );
  IV U474 ( .A(n3194), .Z(n417) );
  MUX U475 ( .IN0(n1099), .IN1(n418), .SEL(n1100), .F(n1053) );
  IV U476 ( .A(n1101), .Z(n418) );
  MUX U477 ( .IN0(n3348), .IN1(n3350), .SEL(n3349), .F(n3208) );
  MUX U478 ( .IN0(n419), .IN1(n1134), .SEL(n1133), .F(n1096) );
  IV U479 ( .A(n1132), .Z(n419) );
  MUX U480 ( .IN0(n4112), .IN1(n4114), .SEL(n4113), .F(n4068) );
  MUX U481 ( .IN0(n5090), .IN1(n5092), .SEL(n5091), .F(n5078) );
  XNOR U482 ( .A(n5088), .B(n5087), .Z(n5093) );
  MUX U483 ( .IN0(n5282), .IN1(n5284), .SEL(n5283), .F(n5262) );
  MUX U484 ( .IN0(n5430), .IN1(n420), .SEL(n5431), .F(n5416) );
  IV U485 ( .A(n5432), .Z(n420) );
  MUX U486 ( .IN0(n4641), .IN1(n4643), .SEL(n4642), .F(n4621) );
  MUX U487 ( .IN0(n4646), .IN1(n421), .SEL(n4647), .F(n4626) );
  IV U488 ( .A(n4648), .Z(n421) );
  MUX U489 ( .IN0(n3625), .IN1(n3627), .SEL(n3626), .F(n3581) );
  XNOR U490 ( .A(n5250), .B(n5249), .Z(n5265) );
  MUX U491 ( .IN0(n5385), .IN1(n5387), .SEL(n5386), .F(n5373) );
  XNOR U492 ( .A(n5395), .B(n5394), .Z(n5400) );
  NANDN U493 ( .B(n2444), .A(n3415), .Z(n434) );
  MUX U494 ( .IN0(n5021), .IN1(n422), .SEL(n5022), .F(n5011) );
  IV U495 ( .A(n5023), .Z(n422) );
  MUX U496 ( .IN0(n5016), .IN1(n5018), .SEL(n5017), .F(n5006) );
  XNOR U497 ( .A(n3487), .B(n3486), .Z(n3520) );
  MUX U498 ( .IN0(n1791), .IN1(n1793), .SEL(n1792), .F(n1696) );
  MUX U499 ( .IN0(n2088), .IN1(n423), .SEL(n2089), .F(n1992) );
  IV U500 ( .A(n2090), .Z(n423) );
  MUX U501 ( .IN0(n2096), .IN1(n424), .SEL(n2097), .F(n2000) );
  IV U502 ( .A(n2098), .Z(n424) );
  MUX U503 ( .IN0(n2054), .IN1(n2056), .SEL(n2055), .F(n1956) );
  MUX U504 ( .IN0(n2062), .IN1(n2064), .SEL(n2063), .F(n1964) );
  MUX U505 ( .IN0(n2148), .IN1(n425), .SEL(n2149), .F(n2047) );
  IV U506 ( .A(n2150), .Z(n425) );
  MUX U507 ( .IN0(n2181), .IN1(n2183), .SEL(n2182), .F(n2080) );
  MUX U508 ( .IN0(n2352), .IN1(n2354), .SEL(n2353), .F(n2244) );
  MUX U509 ( .IN0(n2494), .IN1(n426), .SEL(n2495), .F(n2386) );
  IV U510 ( .A(n2496), .Z(n426) );
  MUX U511 ( .IN0(n2662), .IN1(n2664), .SEL(n2663), .F(n2543) );
  MUX U512 ( .IN0(n2800), .IN1(n427), .SEL(n2801), .F(n2680) );
  IV U513 ( .A(n2802), .Z(n427) );
  MUX U514 ( .IN0(n3331), .IN1(n428), .SEL(n3332), .F(n3192) );
  IV U515 ( .A(n3333), .Z(n428) );
  MUX U516 ( .IN0(n1125), .IN1(n1127), .SEL(n1126), .F(n1083) );
  MUX U517 ( .IN0(n1015), .IN1(n429), .SEL(n1016), .F(n969) );
  IV U518 ( .A(n1017), .Z(n429) );
  MUX U519 ( .IN0(n430), .IN1(n1361), .SEL(n1360), .F(n1296) );
  IV U520 ( .A(n1359), .Z(n430) );
  MUX U521 ( .IN0(n5452), .IN1(n5454), .SEL(n5453), .F(n5435) );
  MUX U522 ( .IN0(n5333), .IN1(n431), .SEL(n5334), .F(n5311) );
  IV U523 ( .A(n5335), .Z(n431) );
  MUX U524 ( .IN0(n5151), .IN1(n5153), .SEL(n5152), .F(n5135) );
  MUX U525 ( .IN0(n5262), .IN1(n5264), .SEL(n5263), .F(n5242) );
  MUX U526 ( .IN0(n5036), .IN1(n5038), .SEL(n5037), .F(n5026) );
  XNOR U527 ( .A(n4818), .B(n4817), .Z(n4825) );
  MUX U528 ( .IN0(n4601), .IN1(n4603), .SEL(n4602), .F(n4581) );
  XNOR U529 ( .A(n4629), .B(n4628), .Z(n4644) );
  MUX U530 ( .IN0(n5227), .IN1(n432), .SEL(n5228), .F(n5207) );
  IV U531 ( .A(n5229), .Z(n432) );
  MUX U532 ( .IN0(n5392), .IN1(n433), .SEL(n5393), .F(n5380) );
  IV U533 ( .A(n5394), .Z(n433) );
  MUX U534 ( .IN0(n4197), .IN1(n434), .SEL(n4198), .F(n4186) );
  MUX U535 ( .IN0(n5373), .IN1(n5375), .SEL(n5374), .F(n5190) );
  MUX U536 ( .IN0(n4562), .IN1(n435), .SEL(n4563), .F(n4541) );
  IV U537 ( .A(n4564), .Z(n435) );
  XNOR U538 ( .A(n5014), .B(n5013), .Z(n5019) );
  MUX U539 ( .IN0(n3452), .IN1(n3454), .SEL(n3453), .F(n3322) );
  MUX U540 ( .IN0(n1860), .IN1(n1862), .SEL(n1861), .F(n1758) );
  MUX U541 ( .IN0(n1896), .IN1(n436), .SEL(n1897), .F(n1799) );
  IV U542 ( .A(n1898), .Z(n436) );
  MUX U543 ( .IN0(n1888), .IN1(n1890), .SEL(n1889), .F(n1791) );
  MUX U544 ( .IN0(n2197), .IN1(n437), .SEL(n2198), .F(n2096) );
  IV U545 ( .A(n2199), .Z(n437) );
  MUX U546 ( .IN0(n2370), .IN1(n2372), .SEL(n2371), .F(n2263) );
  MUX U547 ( .IN0(n2363), .IN1(n438), .SEL(n2364), .F(n2256) );
  IV U548 ( .A(n2365), .Z(n438) );
  MUX U549 ( .IN0(n2402), .IN1(n439), .SEL(n2403), .F(n2295) );
  IV U550 ( .A(n2404), .Z(n439) );
  MUX U551 ( .IN0(n2459), .IN1(n2461), .SEL(n2460), .F(n2352) );
  MUX U552 ( .IN0(n2613), .IN1(n440), .SEL(n2614), .F(n2494) );
  IV U553 ( .A(n2615), .Z(n440) );
  MUX U554 ( .IN0(n3030), .IN1(n3032), .SEL(n3031), .F(n2906) );
  MUX U555 ( .IN0(n3038), .IN1(n441), .SEL(n3039), .F(n2914) );
  IV U556 ( .A(n3040), .Z(n441) );
  MUX U557 ( .IN0(A[28]), .IN1(n4795), .SEL(A[31]), .F(n442) );
  IV U558 ( .A(n442), .Z(n1063) );
  MUX U559 ( .IN0(n1083), .IN1(n1085), .SEL(n1084), .F(n1042) );
  XNOR U560 ( .A(n1364), .B(n1361), .Z(n1424) );
  MUX U561 ( .IN0(n5515), .IN1(n5517), .SEL(n5516), .F(n5499) );
  MUX U562 ( .IN0(n443), .IN1(n5130), .SEL(n5131), .F(n5116) );
  IV U563 ( .A(n5132), .Z(n443) );
  XNOR U564 ( .A(n4649), .B(n4648), .Z(n4664) );
  MUX U565 ( .IN0(n5593), .IN1(n444), .SEL(n5594), .F(n5575) );
  IV U566 ( .A(n5595), .Z(n444) );
  MUX U567 ( .IN0(n5242), .IN1(n5244), .SEL(n5243), .F(n5222) );
  MUX U568 ( .IN0(n4581), .IN1(n4583), .SEL(n4582), .F(n4569) );
  NANDN U569 ( .B(n2939), .A(n3415), .Z(n457) );
  MUX U570 ( .IN0(n4586), .IN1(n445), .SEL(n4587), .F(n4562) );
  IV U571 ( .A(n4588), .Z(n445) );
  XNOR U572 ( .A(n4296), .B(n4294), .Z(n4309) );
  XNOR U573 ( .A(n5230), .B(n5229), .Z(n5245) );
  MUX U574 ( .IN0(n5380), .IN1(n446), .SEL(n5381), .F(n5368) );
  IV U575 ( .A(n5382), .Z(n446) );
  MUX U576 ( .IN0(n5006), .IN1(n5008), .SEL(n5007), .F(n4989) );
  MUX U577 ( .IN0(n5176), .IN1(n447), .SEL(n5177), .F(n3362) );
  IV U578 ( .A(n5178), .Z(n447) );
  MUX U579 ( .IN0(n1807), .IN1(n448), .SEL(n1808), .F(n1714) );
  IV U580 ( .A(n1809), .Z(n448) );
  MUX U581 ( .IN0(n1956), .IN1(n1958), .SEL(n1957), .F(n1860) );
  MUX U582 ( .IN0(n2080), .IN1(n2082), .SEL(n2081), .F(n1984) );
  MUX U583 ( .IN0(n2256), .IN1(n449), .SEL(n2257), .F(n2148) );
  IV U584 ( .A(n2258), .Z(n449) );
  MUX U585 ( .IN0(n2410), .IN1(n450), .SEL(n2411), .F(n2303) );
  IV U586 ( .A(n2412), .Z(n450) );
  MUX U587 ( .IN0(n2510), .IN1(n451), .SEL(n2511), .F(n2402) );
  IV U588 ( .A(n2512), .Z(n451) );
  MUX U589 ( .IN0(n2605), .IN1(n2607), .SEL(n2606), .F(n2486) );
  MUX U590 ( .IN0(n2597), .IN1(n2599), .SEL(n2598), .F(n2478) );
  MUX U591 ( .IN0(n2687), .IN1(n2689), .SEL(n2688), .F(n2573) );
  MUX U592 ( .IN0(n2980), .IN1(n452), .SEL(n2981), .F(n2855) );
  IV U593 ( .A(n2982), .Z(n452) );
  MUX U594 ( .IN0(n1064), .IN1(n1066), .SEL(n1065), .F(n1024) );
  MUX U595 ( .IN0(n1436), .IN1(n1438), .SEL(n1437), .F(n1368) );
  MUX U596 ( .IN0(A[25]), .IN1(n4844), .SEL(A[31]), .F(n453) );
  IV U597 ( .A(n453), .Z(n1208) );
  MUX U598 ( .IN0(n2435), .IN1(n2437), .SEL(n2436), .F(n2330) );
  XNOR U599 ( .A(n1195), .B(n1194), .Z(n1250) );
  XNOR U600 ( .A(n680), .B(n1685), .Z(n1608) );
  AND U601 ( .A(n964), .B(n966), .Z(n935) );
  MUX U602 ( .IN0(n5146), .IN1(n454), .SEL(n5147), .F(n5130) );
  IV U603 ( .A(n5148), .Z(n454) );
  XNOR U604 ( .A(n5292), .B(n5291), .Z(n5309) );
  MUX U605 ( .IN0(n4191), .IN1(n4193), .SEL(n4192), .F(n4177) );
  MUX U606 ( .IN0(n4606), .IN1(n455), .SEL(n4607), .F(n4586) );
  IV U607 ( .A(n4608), .Z(n455) );
  XNOR U608 ( .A(n3572), .B(n3571), .Z(n3607) );
  MUX U609 ( .IN0(n456), .IN1(n5575), .SEL(n5576), .F(n5559) );
  IV U610 ( .A(n5577), .Z(n456) );
  MUX U611 ( .IN0(n5222), .IN1(n5224), .SEL(n5223), .F(n5202) );
  MUX U612 ( .IN0(n4724), .IN1(n457), .SEL(n4725), .F(n4710) );
  XNOR U613 ( .A(n5024), .B(n5023), .Z(n5029) );
  MUX U614 ( .IN0(n5207), .IN1(n458), .SEL(n5208), .F(n5176) );
  IV U615 ( .A(n5209), .Z(n458) );
  XNOR U616 ( .A(n3554), .B(n3552), .Z(n3589) );
  MUX U617 ( .IN0(n5368), .IN1(n459), .SEL(n5369), .F(n3385) );
  IV U618 ( .A(n5370), .Z(n459) );
  MUX U619 ( .IN0(n2303), .IN1(n460), .SEL(n2304), .F(n2197) );
  IV U620 ( .A(n2305), .Z(n460) );
  MUX U621 ( .IN0(n2741), .IN1(n2743), .SEL(n2742), .F(n2621) );
  MUX U622 ( .IN0(n2871), .IN1(n461), .SEL(n2872), .F(n2749) );
  IV U623 ( .A(n2873), .Z(n461) );
  MUX U624 ( .IN0(n2879), .IN1(n462), .SEL(n2880), .F(n2757) );
  IV U625 ( .A(n2881), .Z(n462) );
  MUX U626 ( .IN0(A[22]), .IN1(n4895), .SEL(A[31]), .F(n463) );
  IV U627 ( .A(n463), .Z(n1407) );
  MUX U628 ( .IN0(A[24]), .IN1(n4861), .SEL(A[31]), .F(n464) );
  IV U629 ( .A(n464), .Z(n1272) );
  MUX U630 ( .IN0(A[17]), .IN1(n4980), .SEL(A[31]), .F(n465) );
  IV U631 ( .A(n465), .Z(n1815) );
  MUX U632 ( .IN0(A[19]), .IN1(n4946), .SEL(A[31]), .F(n466) );
  IV U633 ( .A(n466), .Z(n1640) );
  MUX U634 ( .IN0(A[26]), .IN1(n4828), .SEL(A[31]), .F(n467) );
  IV U635 ( .A(n467), .Z(n1149) );
  MUX U636 ( .IN0(A[27]), .IN1(n4812), .SEL(A[31]), .F(n468) );
  IV U637 ( .A(n468), .Z(n1107) );
  MUX U638 ( .IN0(n1269), .IN1(n1267), .SEL(n1268), .F(n1203) );
  MUX U639 ( .IN0(n2946), .IN1(n2948), .SEL(n2947), .F(n2820) );
  XNOR U640 ( .A(n1432), .B(n1431), .Z(n1498) );
  XOR U641 ( .A(n1776), .B(n1691), .Z(n1692) );
  ANDN U642 ( .A(n986), .B(n966), .Z(n955) );
  XNOR U643 ( .A(n5419), .B(n5418), .Z(n5426) );
  MUX U644 ( .IN0(n4186), .IN1(n469), .SEL(n4187), .F(n4172) );
  IV U645 ( .A(n4188), .Z(n469) );
  MUX U646 ( .IN0(n5161), .IN1(n5163), .SEL(n5162), .F(n5157) );
  MUX U647 ( .IN0(n470), .IN1(n5494), .SEL(n5495), .F(n5480) );
  IV U648 ( .A(n5496), .Z(n470) );
  MUX U649 ( .IN0(n471), .IN1(n5116), .SEL(n5117), .F(n5107) );
  IV U650 ( .A(n5118), .Z(n471) );
  XNOR U651 ( .A(n4609), .B(n4608), .Z(n4624) );
  NANDN U652 ( .B(n5607), .A(n3415), .Z(n487) );
  MUX U653 ( .IN0(n5202), .IN1(n5204), .SEL(n5203), .F(n5183) );
  XNOR U654 ( .A(n5383), .B(n5382), .Z(n5388) );
  XNOR U655 ( .A(n5210), .B(n5209), .Z(n5225) );
  XNOR U656 ( .A(n3448), .B(n3447), .Z(n3482) );
  MUX U657 ( .IN0(n2295), .IN1(n472), .SEL(n2296), .F(n2189) );
  IV U658 ( .A(n2297), .Z(n472) );
  MUX U659 ( .IN0(n2590), .IN1(n473), .SEL(n2591), .F(n2471) );
  IV U660 ( .A(n2592), .Z(n473) );
  MUX U661 ( .IN0(n2782), .IN1(n2784), .SEL(n2783), .F(n2662) );
  MUX U662 ( .IN0(n3004), .IN1(n474), .SEL(n3005), .F(n2879) );
  IV U663 ( .A(n3006), .Z(n474) );
  MUX U664 ( .IN0(A[12]), .IN1(n5403), .SEL(A[31]), .F(n475) );
  IV U665 ( .A(n475), .Z(n2311) );
  MUX U666 ( .IN0(n3199), .IN1(n3201), .SEL(n3200), .F(n3074) );
  MUX U667 ( .IN0(A[20]), .IN1(n4929), .SEL(A[31]), .F(n476) );
  IV U668 ( .A(n476), .Z(n1559) );
  MUX U669 ( .IN0(n3168), .IN1(n477), .SEL(n3169), .F(n3038) );
  IV U670 ( .A(n3170), .Z(n477) );
  MUX U671 ( .IN0(A[15]), .IN1(n5367), .SEL(A[31]), .F(n478) );
  IV U672 ( .A(n478), .Z(n2008) );
  MUX U673 ( .IN0(A[23]), .IN1(n4878), .SEL(A[31]), .F(n479) );
  IV U674 ( .A(n479), .Z(n1340) );
  MUX U675 ( .IN0(A[21]), .IN1(n4912), .SEL(A[31]), .F(n480) );
  IV U676 ( .A(n480), .Z(n1481) );
  MUX U677 ( .IN0(n1181), .IN1(n1183), .SEL(n1182), .F(n1125) );
  MUX U678 ( .IN0(n1337), .IN1(n1335), .SEL(n1336), .F(n1267) );
  MUX U679 ( .IN0(n1396), .IN1(n1394), .SEL(n1395), .F(n1325) );
  MUX U680 ( .IN0(n1585), .IN1(n1583), .SEL(n1584), .F(n1505) );
  MUX U681 ( .IN0(n481), .IN1(n1719), .SEL(n1720), .F(n1635) );
  IV U682 ( .A(n1721), .Z(n481) );
  MUX U683 ( .IN0(n2350), .IN1(n2348), .SEL(n2349), .F(n2240) );
  MUX U684 ( .IN0(n482), .IN1(n2640), .SEL(n2641), .F(n2521) );
  IV U685 ( .A(n2642), .Z(n482) );
  MUX U686 ( .IN0(n1060), .IN1(n1058), .SEL(n1059), .F(n1018) );
  MUX U687 ( .IN0(n1368), .IN1(n1370), .SEL(n1369), .F(n1299) );
  MUX U688 ( .IN0(n483), .IN1(n1536), .SEL(n1537), .F(n1456) );
  IV U689 ( .A(n1538), .Z(n483) );
  XOR U690 ( .A(n738), .B(n2025), .Z(n1929) );
  MUX U691 ( .IN0(n2330), .IN1(n2332), .SEL(n2331), .F(n2223) );
  ANDN U692 ( .A(n955), .B(n937), .Z(n926) );
  AND U693 ( .A(n995), .B(n997), .Z(n964) );
  MUX U694 ( .IN0(n1747), .IN1(n1745), .SEL(n1746), .F(n1654) );
  MUX U695 ( .IN0(n5510), .IN1(n484), .SEL(n5511), .F(n5494) );
  IV U696 ( .A(n5512), .Z(n484) );
  MUX U697 ( .IN0(n4621), .IN1(n4623), .SEL(n4622), .F(n4601) );
  MUX U698 ( .IN0(n5598), .IN1(n5600), .SEL(n5599), .F(n5580) );
  XNOR U699 ( .A(n5407), .B(n5406), .Z(n5412) );
  MUX U700 ( .IN0(n485), .IN1(n4172), .SEL(n4173), .F(n4158) );
  IV U701 ( .A(n4174), .Z(n485) );
  MUX U702 ( .IN0(n486), .IN1(n5107), .SEL(n5108), .F(n5095) );
  IV U703 ( .A(n5109), .Z(n486) );
  MUX U704 ( .IN0(n5604), .IN1(n487), .SEL(n5605), .F(n5593) );
  MUX U705 ( .IN0(n5183), .IN1(n5185), .SEL(n5184), .F(n3369) );
  MUX U706 ( .IN0(n2518), .IN1(n488), .SEL(n2519), .F(n2410) );
  IV U707 ( .A(n2520), .Z(n488) );
  MUX U708 ( .IN0(n2486), .IN1(n2488), .SEL(n2487), .F(n2378) );
  MUX U709 ( .IN0(n2680), .IN1(n489), .SEL(n2681), .F(n2566) );
  IV U710 ( .A(n2682), .Z(n489) );
  MUX U711 ( .IN0(n2855), .IN1(n490), .SEL(n2856), .F(n2733) );
  IV U712 ( .A(n2857), .Z(n490) );
  MUX U713 ( .IN0(n2807), .IN1(n2809), .SEL(n2808), .F(n2687) );
  MUX U714 ( .IN0(n3120), .IN1(n3122), .SEL(n3121), .F(n2988) );
  MUX U715 ( .IN0(n3128), .IN1(n491), .SEL(n3129), .F(n2996) );
  IV U716 ( .A(n3130), .Z(n491) );
  MUX U717 ( .IN0(A[16]), .IN1(n4997), .SEL(A[31]), .F(n492) );
  IV U718 ( .A(n492), .Z(n1912) );
  MUX U719 ( .IN0(A[18]), .IN1(n4963), .SEL(A[31]), .F(n493) );
  IV U720 ( .A(n493), .Z(n1724) );
  MUX U721 ( .IN0(A[14]), .IN1(n5379), .SEL(A[31]), .F(n494) );
  IV U722 ( .A(n494), .Z(n2104) );
  MUX U723 ( .IN0(n3160), .IN1(n3162), .SEL(n3161), .F(n3030) );
  MUX U724 ( .IN0(A[13]), .IN1(n5391), .SEL(A[31]), .F(n495) );
  IV U725 ( .A(n495), .Z(n2205) );
  MUX U726 ( .IN0(n3307), .IN1(n496), .SEL(n3308), .F(n3168) );
  IV U727 ( .A(n3309), .Z(n496) );
  XNOR U728 ( .A(n3465), .B(n3464), .Z(n4244) );
  MUX U729 ( .IN0(n1200), .IN1(n497), .SEL(n1201), .F(n1141) );
  IV U730 ( .A(n1202), .Z(n497) );
  MUX U731 ( .IN0(n1434), .IN1(n1432), .SEL(n1433), .F(n1364) );
  MUX U732 ( .IN0(n498), .IN1(n1476), .SEL(n1477), .F(n1402) );
  IV U733 ( .A(n1478), .Z(n498) );
  MUX U734 ( .IN0(n2136), .IN1(n2138), .SEL(n2137), .F(n2035) );
  MUX U735 ( .IN0(n1756), .IN1(n1754), .SEL(n1755), .F(n1665) );
  MUX U736 ( .IN0(n1804), .IN1(n1802), .SEL(n1803), .F(n1709) );
  MUX U737 ( .IN0(n2300), .IN1(n2298), .SEL(n2299), .F(n2192) );
  MUX U738 ( .IN0(n2261), .IN1(n2259), .SEL(n2260), .F(n2151) );
  MUX U739 ( .IN0(n2284), .IN1(n2282), .SEL(n2283), .F(n2176) );
  MUX U740 ( .IN0(n2715), .IN1(n2713), .SEL(n2714), .F(n2593) );
  MUX U741 ( .IN0(n2876), .IN1(n2874), .SEL(n2875), .F(n2752) );
  MUX U742 ( .IN0(n499), .IN1(n2882), .SEL(n2883), .F(n2760) );
  IV U743 ( .A(n2884), .Z(n499) );
  MUX U744 ( .IN0(n1093), .IN1(n1091), .SEL(n1092), .F(n1048) );
  MUX U745 ( .IN0(n1104), .IN1(n1102), .SEL(n1103), .F(n1058) );
  XNOR U746 ( .A(n1257), .B(n1256), .Z(n1318) );
  MUX U747 ( .IN0(n500), .IN1(n1699), .SEL(n1700), .F(n1615) );
  IV U748 ( .A(n1701), .Z(n500) );
  XNOR U749 ( .A(n1777), .B(n1787), .Z(n1876) );
  MUX U750 ( .IN0(n2230), .IN1(n501), .SEL(n2231), .F(n2119) );
  IV U751 ( .A(n2232), .Z(n501) );
  XOR U752 ( .A(n968), .B(n945), .Z(n942) );
  MUX U753 ( .IN0(n1042), .IN1(n1044), .SEL(n1043), .F(n502) );
  IV U754 ( .A(n502), .Z(n1008) );
  AND U755 ( .A(n1076), .B(n1078), .Z(n1036) );
  NOR U756 ( .A(n1743), .B(n1744), .Z(n1742) );
  NANDN U757 ( .B(n914), .A(n926), .Z(n894) );
  MUX U758 ( .IN0(n929), .IN1(Y0[29]), .SEL(n930), .F(n906) );
  MUX U759 ( .IN0(n4528), .IN1(n4526), .SEL(n4527), .F(n4505) );
  MUX U760 ( .IN0(n5464), .IN1(n5341), .SEL(n5342), .F(n5450) );
  MUX U761 ( .IN0(n5524), .IN1(n5526), .SEL(n5525), .F(n5521) );
  MUX U762 ( .IN0(n503), .IN1(n5121), .SEL(n5122), .F(n5102) );
  IV U763 ( .A(n5123), .Z(n503) );
  MUX U764 ( .IN0(n504), .IN1(n5480), .SEL(n5481), .F(n5471) );
  IV U765 ( .A(n5482), .Z(n504) );
  NANDN U766 ( .B(n5348), .A(n3415), .Z(n525) );
  MUX U767 ( .IN0(n4569), .IN1(n4571), .SEL(n4570), .F(n4551) );
  XNOR U768 ( .A(n4589), .B(n4588), .Z(n4604) );
  MUX U769 ( .IN0(n505), .IN1(n5548), .SEL(n5549), .F(n3401) );
  IV U770 ( .A(n5550), .Z(n505) );
  XNOR U771 ( .A(n5371), .B(n5370), .Z(n5376) );
  XNOR U772 ( .A(n5100), .B(n5099), .Z(n5105) );
  MUX U773 ( .IN0(n2263), .IN1(n2265), .SEL(n2264), .F(n2155) );
  MUX U774 ( .IN0(n2378), .IN1(n2380), .SEL(n2379), .F(n2271) );
  MUX U775 ( .IN0(n2621), .IN1(n2623), .SEL(n2622), .F(n2502) );
  MUX U776 ( .IN0(n2629), .IN1(n506), .SEL(n2630), .F(n2510) );
  IV U777 ( .A(n2631), .Z(n506) );
  MUX U778 ( .IN0(n2573), .IN1(n2575), .SEL(n2574), .F(n2459) );
  MUX U779 ( .IN0(n2710), .IN1(n507), .SEL(n2711), .F(n2590) );
  IV U780 ( .A(n2712), .Z(n507) );
  MUX U781 ( .IN0(n2906), .IN1(n2908), .SEL(n2907), .F(n2782) );
  MUX U782 ( .IN0(n2914), .IN1(n508), .SEL(n2915), .F(n2790) );
  IV U783 ( .A(n2916), .Z(n508) );
  MUX U784 ( .IN0(n3053), .IN1(n3055), .SEL(n3054), .F(n2929) );
  MUX U785 ( .IN0(n3104), .IN1(n3106), .SEL(n3105), .F(n2972) );
  MUX U786 ( .IN0(n3112), .IN1(n509), .SEL(n3113), .F(n2980) );
  IV U787 ( .A(n3114), .Z(n509) );
  MUX U788 ( .IN0(n3228), .IN1(n3230), .SEL(n3229), .F(n3096) );
  MUX U789 ( .IN0(n3221), .IN1(n510), .SEL(n3222), .F(n3089) );
  IV U790 ( .A(n3223), .Z(n510) );
  MUX U791 ( .IN0(n3268), .IN1(n511), .SEL(n3269), .F(n3136) );
  IV U792 ( .A(n3270), .Z(n511) );
  MUX U793 ( .IN0(n3176), .IN1(n512), .SEL(n3177), .F(n3046) );
  IV U794 ( .A(n3178), .Z(n512) );
  MUX U795 ( .IN0(n5181), .IN1(n5179), .SEL(n5180), .F(n3365) );
  MUX U796 ( .IN0(n3450), .IN1(n3448), .SEL(n3449), .F(n3318) );
  XNOR U797 ( .A(n3440), .B(n3439), .Z(n3502) );
  MUX U798 ( .IN0(n1108), .IN1(n1110), .SEL(n1109), .F(n1064) );
  MUX U799 ( .IN0(n1711), .IN1(n1709), .SEL(n1710), .F(n1625) );
  MUX U800 ( .IN0(n513), .IN1(n2099), .SEL(n2100), .F(n2003) );
  IV U801 ( .A(n2101), .Z(n513) );
  MUX U802 ( .IN0(n2077), .IN1(n2075), .SEL(n2076), .F(n1979) );
  MUX U803 ( .IN0(n2368), .IN1(n2366), .SEL(n2367), .F(n2259) );
  MUX U804 ( .IN0(n2407), .IN1(n2405), .SEL(n2406), .F(n2298) );
  MUX U805 ( .IN0(n2447), .IN1(n2449), .SEL(n2448), .F(n514) );
  IV U806 ( .A(n514), .Z(n2337) );
  MUX U807 ( .IN0(n2618), .IN1(n2616), .SEL(n2617), .F(n2497) );
  MUX U808 ( .IN0(n2805), .IN1(n2803), .SEL(n2804), .F(n2683) );
  MUX U809 ( .IN0(n515), .IN1(n3007), .SEL(n3008), .F(n2882) );
  IV U810 ( .A(n3009), .Z(n515) );
  MUX U811 ( .IN0(n3001), .IN1(n2999), .SEL(n3000), .F(n2874) );
  MUX U812 ( .IN0(n2962), .IN1(n2960), .SEL(n2961), .F(n2835) );
  MUX U813 ( .IN0(n2944), .IN1(n2942), .SEL(n2943), .F(n516) );
  IV U814 ( .A(n516), .Z(n2814) );
  MUX U815 ( .IN0(n3043), .IN1(n3041), .SEL(n3042), .F(n2917) );
  XNOR U816 ( .A(n3334), .B(n3333), .Z(n3458) );
  MUX U817 ( .IN0(n1020), .IN1(n1018), .SEL(n1019), .F(n974) );
  MUX U818 ( .IN0(n1205), .IN1(n1203), .SEL(n1204), .F(n1144) );
  MUX U819 ( .IN0(n1376), .IN1(n1374), .SEL(n1375), .F(n1305) );
  MUX U820 ( .IN0(n517), .IN1(n1384), .SEL(n1385), .F(n1315) );
  IV U821 ( .A(n1386), .Z(n517) );
  XNOR U822 ( .A(n1505), .B(n1504), .Z(n1576) );
  MUX U823 ( .IN0(n518), .IN1(n1794), .SEL(n1795), .F(n1699) );
  IV U824 ( .A(n1796), .Z(n518) );
  XNOR U825 ( .A(n2122), .B(n2031), .Z(n2032) );
  MUX U826 ( .IN0(n2334), .IN1(n519), .SEL(n2335), .F(n2230) );
  IV U827 ( .A(n2336), .Z(n519) );
  MUX U828 ( .IN0(n2820), .IN1(n2822), .SEL(n2821), .F(n2702) );
  ANDN U829 ( .A(n1001), .B(n1005), .Z(n1004) );
  MUX U830 ( .IN0(n520), .IN1(n1235), .SEL(n1236), .F(n1176) );
  IV U831 ( .A(n1237), .Z(n520) );
  ANDN U832 ( .A(n1941), .B(n1943), .Z(n1832) );
  MUX U833 ( .IN0(n568), .IN1(n2582), .SEL(n2581), .F(n2465) );
  NANDN U834 ( .B(n987), .A(n988), .Z(n956) );
  AND U835 ( .A(n1036), .B(n1038), .Z(n995) );
  NANDN U836 ( .B(n1156), .A(n1157), .Z(n1112) );
  AND U837 ( .A(n1354), .B(n1356), .Z(n1286) );
  MUX U838 ( .IN0(n1847), .IN1(n521), .SEL(n1846), .F(n1745) );
  IV U839 ( .A(n1845), .Z(n521) );
  AND U840 ( .A(n902), .B(n903), .Z(n897) );
  MUX U841 ( .IN0(n958), .IN1(Y0[28]), .SEL(n959), .F(n929) );
  MUX U842 ( .IN0(n4135), .IN1(n4133), .SEL(n4134), .F(n4091) );
  MUX U843 ( .IN0(n4200), .IN1(n4202), .SEL(n4201), .F(n4197) );
  MUX U844 ( .IN0(n522), .IN1(n5485), .SEL(n5486), .F(n5466) );
  IV U845 ( .A(n5487), .Z(n522) );
  MUX U846 ( .IN0(n523), .IN1(n4158), .SEL(n4159), .F(n4149) );
  IV U847 ( .A(n4160), .Z(n523) );
  MUX U848 ( .IN0(n524), .IN1(n5102), .SEL(n5103), .F(n5090) );
  IV U849 ( .A(n5104), .Z(n524) );
  MUX U850 ( .IN0(n5345), .IN1(n525), .SEL(n5346), .F(n5333) );
  MUX U851 ( .IN0(n526), .IN1(n5471), .SEL(n5472), .F(n5459) );
  IV U852 ( .A(n5473), .Z(n526) );
  XNOR U853 ( .A(n4565), .B(n4564), .Z(n4584) );
  MUX U854 ( .IN0(n2155), .IN1(n2157), .SEL(n2156), .F(n2054) );
  MUX U855 ( .IN0(n2189), .IN1(n527), .SEL(n2190), .F(n2088) );
  IV U856 ( .A(n2191), .Z(n527) );
  MUX U857 ( .IN0(n2637), .IN1(n528), .SEL(n2638), .F(n2518) );
  IV U858 ( .A(n2639), .Z(n528) );
  MUX U859 ( .IN0(n2749), .IN1(n529), .SEL(n2750), .F(n2629) );
  IV U860 ( .A(n2751), .Z(n529) );
  MUX U861 ( .IN0(n2725), .IN1(n2727), .SEL(n2726), .F(n2605) );
  MUX U862 ( .IN0(n2839), .IN1(n2841), .SEL(n2840), .F(n2717) );
  MUX U863 ( .IN0(n2832), .IN1(n530), .SEL(n2833), .F(n2710) );
  IV U864 ( .A(n2834), .Z(n530) );
  MUX U865 ( .IN0(n2988), .IN1(n2990), .SEL(n2989), .F(n2863) );
  MUX U866 ( .IN0(n2922), .IN1(n531), .SEL(n2923), .F(n2800) );
  IV U867 ( .A(n2924), .Z(n531) );
  MUX U868 ( .IN0(n3236), .IN1(n3238), .SEL(n3237), .F(n3104) );
  MUX U869 ( .IN0(n3244), .IN1(n532), .SEL(n3245), .F(n3112) );
  IV U870 ( .A(n3246), .Z(n532) );
  MUX U871 ( .IN0(n3401), .IN1(n533), .SEL(n3402), .F(n3260) );
  IV U872 ( .A(n3403), .Z(n533) );
  MUX U873 ( .IN0(n3362), .IN1(n534), .SEL(n3363), .F(n3221) );
  IV U874 ( .A(n3364), .Z(n534) );
  MUX U875 ( .IN0(n3299), .IN1(n3301), .SEL(n3300), .F(n3160) );
  MUX U876 ( .IN0(n5371), .IN1(n5197), .SEL(n5199), .F(n3388) );
  MUX U877 ( .IN0(n1150), .IN1(n1152), .SEL(n1151), .F(n1108) );
  MUX U878 ( .IN0(n1954), .IN1(n1952), .SEL(n1953), .F(n1856) );
  MUX U879 ( .IN0(n1997), .IN1(n1995), .SEL(n1996), .F(n1899) );
  MUX U880 ( .IN0(n535), .IN1(n2003), .SEL(n2004), .F(n1907) );
  IV U881 ( .A(n2005), .Z(n535) );
  MUX U882 ( .IN0(n2391), .IN1(n2389), .SEL(n2390), .F(n2282) );
  MUX U883 ( .IN0(n536), .IN1(n2413), .SEL(n2414), .F(n2306) );
  IV U884 ( .A(n2415), .Z(n536) );
  MUX U885 ( .IN0(n2515), .IN1(n2513), .SEL(n2514), .F(n2405) );
  MUX U886 ( .IN0(n2476), .IN1(n2474), .SEL(n2475), .F(n2366) );
  MUX U887 ( .IN0(n2571), .IN1(n2569), .SEL(n2570), .F(n2455) );
  MUX U888 ( .IN0(n2985), .IN1(n2983), .SEL(n2984), .F(n2858) );
  MUX U889 ( .IN0(n2919), .IN1(n2917), .SEL(n2918), .F(n2795) );
  MUX U890 ( .IN0(n3133), .IN1(n3131), .SEL(n3132), .F(n2999) );
  MUX U891 ( .IN0(n537), .IN1(n3139), .SEL(n3140), .F(n3007) );
  IV U892 ( .A(n3141), .Z(n537) );
  MUX U893 ( .IN0(n3094), .IN1(n3092), .SEL(n3093), .F(n2960) );
  MUX U894 ( .IN0(n3181), .IN1(n3179), .SEL(n3180), .F(n3049) );
  XNOR U895 ( .A(n3310), .B(n3309), .Z(n3433) );
  MUX U896 ( .IN0(n1138), .IN1(n1136), .SEL(n1137), .F(n1091) );
  XNOR U897 ( .A(n1203), .B(n1202), .Z(n1260) );
  MUX U898 ( .IN0(n1444), .IN1(n1446), .SEL(n1445), .F(n1374) );
  XNOR U899 ( .A(n1394), .B(n1393), .Z(n1459) );
  XNOR U900 ( .A(n1554), .B(n1553), .Z(n1628) );
  XNOR U901 ( .A(n1583), .B(n1582), .Z(n1658) );
  MUX U902 ( .IN0(n2035), .IN1(n2037), .SEL(n2036), .F(n1934) );
  MUX U903 ( .IN0(n538), .IN1(n1773), .SEL(n1774), .F(n1682) );
  IV U904 ( .A(n1775), .Z(n538) );
  XNOR U905 ( .A(n2123), .B(n2133), .Z(n2233) );
  XOR U906 ( .A(n2551), .B(n2447), .Z(n2448) );
  MUX U907 ( .IN0(n539), .IN1(n2744), .SEL(n2745), .F(n2624) );
  IV U908 ( .A(n2746), .Z(n539) );
  MUX U909 ( .IN0(n2816), .IN1(n540), .SEL(n2815), .F(n2700) );
  IV U910 ( .A(n2814), .Z(n540) );
  MUX U911 ( .IN0(n1011), .IN1(n541), .SEL(n1010), .F(n983) );
  IV U912 ( .A(n1009), .Z(n541) );
  XNOR U913 ( .A(n1174), .B(n1173), .Z(n1227) );
  AND U914 ( .A(n1564), .B(n1566), .Z(n1486) );
  MUX U915 ( .IN0(n542), .IN1(n1672), .SEL(n1673), .F(n1592) );
  IV U916 ( .A(n1674), .Z(n542) );
  MUX U917 ( .IN0(n2826), .IN1(n2828), .SEL(n2827), .F(n2704) );
  NANDN U918 ( .B(n1028), .A(n1029), .Z(n987) );
  ANDN U919 ( .A(n1067), .B(n1038), .Z(n1027) );
  NANDN U920 ( .B(n1215), .A(n1216), .Z(n1156) );
  NAND U921 ( .A(n1832), .B(n1831), .Z(n1743) );
  MUX U922 ( .IN0(n543), .IN1(n2355), .SEL(n2356), .F(n2247) );
  IV U923 ( .A(n2357), .Z(n543) );
  ANDN U924 ( .A(n1495), .B(n1496), .Z(n1421) );
  MUX U925 ( .IN0(Y0[3]), .IN1(n3017), .SEL(n3018), .F(n2894) );
  MUX U926 ( .IN0(n894), .IN1(n896), .SEL(n895), .F(n544) );
  IV U927 ( .A(n544), .Z(n893) );
  MUX U928 ( .IN0(n989), .IN1(Y0[27]), .SEL(n990), .F(n958) );
  MUX U929 ( .IN0(n1158), .IN1(Y0[23]), .SEL(n1159), .F(n1114) );
  MUX U930 ( .IN0(n1415), .IN1(Y0[19]), .SEL(n1416), .F(n1348) );
  MUX U931 ( .IN0(n1732), .IN1(Y0[15]), .SEL(n1733), .F(n1648) );
  MUX U932 ( .IN0(n2112), .IN1(Y0[11]), .SEL(n2113), .F(n2016) );
  MUX U933 ( .IN0(n2534), .IN1(Y0[7]), .SEL(n2535), .F(n2426) );
  MUX U934 ( .IN0(n5004), .IN1(n4558), .SEL(n4559), .F(n4987) );
  MUX U935 ( .IN0(n545), .IN1(n4535), .SEL(n4100), .F(n4514) );
  IV U936 ( .A(n4098), .Z(n545) );
  MUX U937 ( .IN0(n3974), .IN1(n3972), .SEL(n3973), .F(n3928) );
  MUX U938 ( .IN0(n4695), .IN1(n4693), .SEL(n4694), .F(n4669) );
  XNOR U939 ( .A(n5270), .B(n5269), .Z(n5285) );
  MUX U940 ( .IN0(n4727), .IN1(n4729), .SEL(n4728), .F(n4724) );
  MUX U941 ( .IN0(n546), .IN1(n4163), .SEL(n4164), .F(n4142) );
  IV U942 ( .A(n4165), .Z(n546) );
  NANDN U943 ( .B(n2028), .A(n3415), .Z(n578) );
  MUX U944 ( .IN0(n547), .IN1(n5539), .SEL(n5540), .F(n3393) );
  IV U945 ( .A(n5541), .Z(n547) );
  MUX U946 ( .IN0(n5190), .IN1(n5192), .SEL(n5191), .F(n3377) );
  MUX U947 ( .IN0(n4253), .IN1(n4251), .SEL(n4252), .F(n3465) );
  MUX U948 ( .IN0(n2271), .IN1(n2273), .SEL(n2272), .F(n2163) );
  MUX U949 ( .IN0(n2394), .IN1(n2396), .SEL(n2395), .F(n2287) );
  MUX U950 ( .IN0(n2478), .IN1(n2480), .SEL(n2479), .F(n2370) );
  MUX U951 ( .IN0(n2471), .IN1(n548), .SEL(n2472), .F(n2363) );
  IV U952 ( .A(n2473), .Z(n548) );
  MUX U953 ( .IN0(n2733), .IN1(n549), .SEL(n2734), .F(n2613) );
  IV U954 ( .A(n2735), .Z(n549) );
  MUX U955 ( .IN0(n2847), .IN1(n2849), .SEL(n2848), .F(n2725) );
  MUX U956 ( .IN0(n2863), .IN1(n2865), .SEL(n2864), .F(n2741) );
  MUX U957 ( .IN0(n2996), .IN1(n550), .SEL(n2997), .F(n2871) );
  IV U958 ( .A(n2998), .Z(n550) );
  MUX U959 ( .IN0(n2957), .IN1(n551), .SEL(n2958), .F(n2832) );
  IV U960 ( .A(n2959), .Z(n551) );
  MUX U961 ( .IN0(n3046), .IN1(n552), .SEL(n3047), .F(n2922) );
  IV U962 ( .A(n3048), .Z(n552) );
  MUX U963 ( .IN0(n3136), .IN1(n553), .SEL(n3137), .F(n3004) );
  IV U964 ( .A(n3138), .Z(n553) );
  MUX U965 ( .IN0(n3096), .IN1(n3098), .SEL(n3097), .F(n2964) );
  MUX U966 ( .IN0(A[8]), .IN1(n5458), .SEL(A[31]), .F(n554) );
  IV U967 ( .A(n554), .Z(n2765) );
  MUX U968 ( .IN0(n3385), .IN1(n555), .SEL(n3386), .F(n3244) );
  IV U969 ( .A(n3387), .Z(n555) );
  MUX U970 ( .IN0(n3338), .IN1(n3340), .SEL(n3339), .F(n3199) );
  MUX U971 ( .IN0(n1259), .IN1(n1257), .SEL(n1258), .F(n1195) );
  MUX U972 ( .IN0(n2153), .IN1(n2151), .SEL(n2152), .F(n2050) );
  MUX U973 ( .IN0(n2194), .IN1(n2192), .SEL(n2193), .F(n2091) );
  MUX U974 ( .IN0(n2125), .IN1(n2123), .SEL(n2124), .F(n2031) );
  MUX U975 ( .IN0(n556), .IN1(n2306), .SEL(n2307), .F(n2200) );
  IV U976 ( .A(n2308), .Z(n556) );
  MUX U977 ( .IN0(n2499), .IN1(n2497), .SEL(n2498), .F(n2389) );
  MUX U978 ( .IN0(n2595), .IN1(n2593), .SEL(n2594), .F(n2474) );
  MUX U979 ( .IN0(n2634), .IN1(n2632), .SEL(n2633), .F(n2513) );
  MUX U980 ( .IN0(n2554), .IN1(n2552), .SEL(n2553), .F(n2447) );
  MUX U981 ( .IN0(n2685), .IN1(n2683), .SEL(n2684), .F(n2569) );
  MUX U982 ( .IN0(n557), .IN1(n2760), .SEL(n2761), .F(n2640) );
  IV U983 ( .A(n2762), .Z(n557) );
  MUX U984 ( .IN0(n3063), .IN1(n3061), .SEL(n3062), .F(n2942) );
  MUX U985 ( .IN0(n3117), .IN1(n3115), .SEL(n3116), .F(n2983) );
  MUX U986 ( .IN0(n3226), .IN1(n3224), .SEL(n3225), .F(n3092) );
  MUX U987 ( .IN0(n3265), .IN1(n3263), .SEL(n3264), .F(n3131) );
  MUX U988 ( .IN0(n558), .IN1(n3271), .SEL(n3272), .F(n3139) );
  IV U989 ( .A(n3273), .Z(n558) );
  MUX U990 ( .IN0(n3173), .IN1(n3171), .SEL(n3172), .F(n3041) );
  MUX U991 ( .IN0(n3320), .IN1(n3318), .SEL(n3319), .F(n3179) );
  MUX U992 ( .IN0(n1024), .IN1(n1026), .SEL(n1025), .F(n980) );
  MUX U993 ( .IN0(n1146), .IN1(n1144), .SEL(n1145), .F(n1102) );
  XNOR U994 ( .A(n1335), .B(n1334), .Z(n1397) );
  XNOR U995 ( .A(n1546), .B(n1545), .Z(n1618) );
  XNOR U996 ( .A(n1635), .B(n1634), .Z(n1712) );
  XNOR U997 ( .A(n1665), .B(n1664), .Z(n1749) );
  MUX U998 ( .IN0(n559), .IN1(n1891), .SEL(n1892), .F(n1794) );
  IV U999 ( .A(n1893), .Z(n559) );
  XNOR U1000 ( .A(n1883), .B(n1882), .Z(n1972) );
  MUX U1001 ( .IN0(n2438), .IN1(n560), .SEL(n2439), .F(n2334) );
  IV U1002 ( .A(n2440), .Z(n560) );
  MUX U1003 ( .IN0(n561), .IN1(n2505), .SEL(n2506), .F(n2397) );
  IV U1004 ( .A(n2507), .Z(n561) );
  MUX U1005 ( .IN0(n562), .IN1(n2728), .SEL(n2729), .F(n2608) );
  IV U1006 ( .A(n2730), .Z(n562) );
  MUX U1007 ( .IN0(n563), .IN1(n2991), .SEL(n2992), .F(n2866) );
  IV U1008 ( .A(n2993), .Z(n563) );
  MUX U1009 ( .IN0(n564), .IN1(n2909), .SEL(n2910), .F(n2785) );
  IV U1010 ( .A(n2911), .Z(n564) );
  MUX U1011 ( .IN0(n565), .IN1(n971), .SEL(n970), .F(n945) );
  IV U1012 ( .A(n969), .Z(n565) );
  AND U1013 ( .A(n1007), .B(n1008), .Z(n1003) );
  MUX U1014 ( .IN0(n1294), .IN1(n1292), .SEL(n1293), .F(n1232) );
  MUX U1015 ( .IN0(n566), .IN1(n1439), .SEL(n1440), .F(n1371) );
  IV U1016 ( .A(n1441), .Z(n566) );
  AND U1017 ( .A(n1645), .B(n1647), .Z(n1564) );
  MUX U1018 ( .IN0(n1934), .IN1(n1936), .SEL(n1935), .F(n1843) );
  MUX U1019 ( .IN0(n567), .IN1(n2158), .SEL(n2159), .F(n2057) );
  IV U1020 ( .A(n2160), .Z(n567) );
  ANDN U1021 ( .A(n2142), .B(n2144), .Z(n2041) );
  AND U1022 ( .A(n2423), .B(n2425), .Z(n2316) );
  MUX U1023 ( .IN0(n2706), .IN1(n2704), .SEL(n2705), .F(n568) );
  IV U1024 ( .A(n568), .Z(n2580) );
  NANDN U1025 ( .B(n1068), .A(n1069), .Z(n1028) );
  MUX U1026 ( .IN0(n1155), .IN1(n569), .SEL(n1154), .F(n1111) );
  IV U1027 ( .A(n1153), .Z(n569) );
  AND U1028 ( .A(n1223), .B(n1225), .Z(n1212) );
  NANDN U1029 ( .B(n1278), .A(n1279), .Z(n1215) );
  MUX U1030 ( .IN0(n570), .IN1(n1938), .SEL(n1939), .F(n1845) );
  IV U1031 ( .A(n1940), .Z(n570) );
  MUX U1032 ( .IN0(n571), .IN1(n2462), .SEL(n2463), .F(n2355) );
  IV U1033 ( .A(n2464), .Z(n571) );
  MUX U1034 ( .IN0(n2934), .IN1(n598), .SEL(n2933), .F(n572) );
  IV U1035 ( .A(n572), .Z(n2810) );
  AND U1036 ( .A(n935), .B(n937), .Z(n912) );
  ANDN U1037 ( .A(n1573), .B(n1574), .Z(n1495) );
  NAND U1038 ( .A(n883), .B(n885), .Z(n882) );
  MUX U1039 ( .IN0(n1030), .IN1(Y0[26]), .SEL(n1031), .F(n989) );
  MUX U1040 ( .IN0(n1217), .IN1(Y0[22]), .SEL(n1218), .F(n1158) );
  MUX U1041 ( .IN0(n1489), .IN1(Y0[18]), .SEL(n1490), .F(n1415) );
  MUX U1042 ( .IN0(n1823), .IN1(Y0[14]), .SEL(n1824), .F(n1732) );
  MUX U1043 ( .IN0(n2213), .IN1(Y0[10]), .SEL(n2214), .F(n2112) );
  MUX U1044 ( .IN0(n2653), .IN1(Y0[6]), .SEL(n2654), .F(n2534) );
  MUX U1045 ( .IN0(n4549), .IN1(n4547), .SEL(n4548), .F(n4526) );
  MUX U1046 ( .IN0(n4124), .IN1(n4122), .SEL(n4123), .F(n573) );
  IV U1047 ( .A(n573), .Z(n4080) );
  MUX U1048 ( .IN0(n4047), .IN1(n4045), .SEL(n4046), .F(n3999) );
  MUX U1049 ( .IN0(n4970), .IN1(n4516), .SEL(n4517), .F(n4953) );
  MUX U1050 ( .IN0(n574), .IN1(n4451), .SEL(n3918), .F(n4430) );
  IV U1051 ( .A(n3916), .Z(n574) );
  MUX U1052 ( .IN0(n5100), .IN1(n4720), .SEL(n4721), .F(n5088) );
  MUX U1053 ( .IN0(n5338), .IN1(n5336), .SEL(n5337), .F(n5316) );
  XNOR U1054 ( .A(n4669), .B(n4668), .Z(n4686) );
  MUX U1055 ( .IN0(n575), .IN1(n4367), .SEL(n3736), .F(n4346) );
  IV U1056 ( .A(n3734), .Z(n575) );
  MUX U1057 ( .IN0(n5046), .IN1(n4636), .SEL(n4638), .F(n5034) );
  MUX U1058 ( .IN0(n5608), .IN1(n5610), .SEL(n5609), .F(n5604) );
  MUX U1059 ( .IN0(n5252), .IN1(n5250), .SEL(n5251), .F(n5230) );
  MUX U1060 ( .IN0(n576), .IN1(n5564), .SEL(n5565), .F(n5539) );
  IV U1061 ( .A(n5566), .Z(n576) );
  MUX U1062 ( .IN0(n577), .IN1(n5466), .SEL(n5467), .F(n5452) );
  IV U1063 ( .A(n5468), .Z(n577) );
  MUX U1064 ( .IN0(n4218), .IN1(n578), .SEL(n4219), .F(n4104) );
  MUX U1065 ( .IN0(n579), .IN1(n4284), .SEL(n3563), .F(n4263) );
  IV U1066 ( .A(n3561), .Z(n579) );
  MUX U1067 ( .IN0(n2287), .IN1(n2289), .SEL(n2288), .F(n2181) );
  MUX U1068 ( .IN0(n3260), .IN1(n580), .SEL(n3261), .F(n3128) );
  IV U1069 ( .A(n3262), .Z(n580) );
  MUX U1070 ( .IN0(A[7]), .IN1(n5547), .SEL(A[31]), .F(n581) );
  IV U1071 ( .A(n581), .Z(n2887) );
  MUX U1072 ( .IN0(A[11]), .IN1(n5415), .SEL(A[31]), .F(n582) );
  IV U1073 ( .A(n582), .Z(n2418) );
  MUX U1074 ( .IN0(n3322), .IN1(n3324), .SEL(n3323), .F(n3183) );
  MUX U1075 ( .IN0(n3315), .IN1(n583), .SEL(n3316), .F(n3176) );
  IV U1076 ( .A(n3317), .Z(n583) );
  MUX U1077 ( .IN0(n3442), .IN1(n3440), .SEL(n3441), .F(n3310) );
  MUX U1078 ( .IN0(n1209), .IN1(n1211), .SEL(n1210), .F(n1150) );
  MUX U1079 ( .IN0(n1627), .IN1(n1625), .SEL(n1626), .F(n1546) );
  MUX U1080 ( .IN0(n1779), .IN1(n1777), .SEL(n1778), .F(n1691) );
  MUX U1081 ( .IN0(n2178), .IN1(n2176), .SEL(n2177), .F(n2075) );
  MUX U1082 ( .IN0(n2738), .IN1(n2736), .SEL(n2737), .F(n2616) );
  MUX U1083 ( .IN0(n2837), .IN1(n2835), .SEL(n2836), .F(n2713) );
  MUX U1084 ( .IN0(n3051), .IN1(n3049), .SEL(n3050), .F(n2925) );
  MUX U1085 ( .IN0(n3249), .IN1(n3247), .SEL(n3248), .F(n3115) );
  MUX U1086 ( .IN0(n584), .IN1(n3412), .SEL(n3413), .F(n3271) );
  IV U1087 ( .A(n3414), .Z(n584) );
  MUX U1088 ( .IN0(n3406), .IN1(n3404), .SEL(n3405), .F(n3263) );
  MUX U1089 ( .IN0(n3367), .IN1(n3365), .SEL(n3366), .F(n3224) );
  XNOR U1090 ( .A(n1267), .B(n1266), .Z(n1328) );
  XNOR U1091 ( .A(n1325), .B(n1324), .Z(n1387) );
  XNOR U1092 ( .A(n1476), .B(n1475), .Z(n1549) );
  MUX U1093 ( .IN0(n1605), .IN1(n585), .SEL(n1606), .F(n1526) );
  IV U1094 ( .A(n1607), .Z(n585) );
  XNOR U1095 ( .A(n1719), .B(n1718), .Z(n1805) );
  XNOR U1096 ( .A(n1754), .B(n1753), .Z(n1849) );
  XNOR U1097 ( .A(n1899), .B(n1898), .Z(n1990) );
  MUX U1098 ( .IN0(n586), .IN1(n2083), .SEL(n2084), .F(n1987) );
  IV U1099 ( .A(n2085), .Z(n586) );
  XNOR U1100 ( .A(n2003), .B(n2002), .Z(n2094) );
  XNOR U1101 ( .A(n2050), .B(n2049), .Z(n2146) );
  MUX U1102 ( .IN0(n587), .IN1(n2274), .SEL(n2275), .F(n2166) );
  IV U1103 ( .A(n2276), .Z(n587) );
  XNOR U1104 ( .A(n2298), .B(n2297), .Z(n2400) );
  XNOR U1105 ( .A(n2306), .B(n2305), .Z(n2408) );
  XNOR U1106 ( .A(n2455), .B(n2454), .Z(n2564) );
  XNOR U1107 ( .A(n2632), .B(n2631), .Z(n2747) );
  XNOR U1108 ( .A(n2640), .B(n2639), .Z(n2755) );
  XNOR U1109 ( .A(n2675), .B(n2674), .Z(n2788) );
  MUX U1110 ( .IN0(n588), .IN1(n2975), .SEL(n2976), .F(n2850) );
  IV U1111 ( .A(n2977), .Z(n588) );
  XNOR U1112 ( .A(n3061), .B(n3071), .Z(n3190) );
  MUX U1113 ( .IN0(n589), .IN1(n3163), .SEL(n3164), .F(n3033) );
  IV U1114 ( .A(n3165), .Z(n589) );
  XNOR U1115 ( .A(n974), .B(n971), .Z(n1012) );
  MUX U1116 ( .IN0(n1050), .IN1(n1048), .SEL(n1049), .F(n1001) );
  MUX U1117 ( .IN0(n590), .IN1(n1086), .SEL(n1087), .F(n1045) );
  IV U1118 ( .A(n1088), .Z(n590) );
  AND U1119 ( .A(n1305), .B(n1307), .Z(n1238) );
  MUX U1120 ( .IN0(n591), .IN1(n1514), .SEL(n1515), .F(n1439) );
  IV U1121 ( .A(n1516), .Z(n591) );
  MUX U1122 ( .IN0(n1930), .IN1(n738), .SEL(n1929), .F(n1842) );
  AND U1123 ( .A(n2013), .B(n2015), .Z(n1917) );
  ANDN U1124 ( .A(n2250), .B(n2252), .Z(n2142) );
  MUX U1125 ( .IN0(n592), .IN1(n2373), .SEL(n2374), .F(n2266) );
  IV U1126 ( .A(n2375), .Z(n592) );
  AND U1127 ( .A(n2650), .B(n2652), .Z(n2531) );
  MUX U1128 ( .IN0(n593), .IN1(n2842), .SEL(n2843), .F(n2720) );
  IV U1129 ( .A(n2844), .Z(n593) );
  MUX U1130 ( .IN0(n594), .IN1(n2953), .SEL(n2952), .F(n2826) );
  IV U1131 ( .A(n2951), .Z(n594) );
  NANDN U1132 ( .B(n956), .A(n957), .Z(n927) );
  ANDN U1133 ( .A(n1111), .B(n1078), .Z(n1067) );
  NANDN U1134 ( .B(n1112), .A(n1113), .Z(n1068) );
  MUX U1135 ( .IN0(n1234), .IN1(n1232), .SEL(n1233), .F(n595) );
  IV U1136 ( .A(n595), .Z(n1172) );
  OR U1137 ( .A(n1413), .B(n1414), .Z(n1346) );
  MUX U1138 ( .IN0(n596), .IN1(n2038), .SEL(n2039), .F(n1938) );
  IV U1139 ( .A(n2040), .Z(n596) );
  MUX U1140 ( .IN0(n597), .IN1(n2576), .SEL(n2577), .F(n2462) );
  IV U1141 ( .A(n2578), .Z(n597) );
  MUX U1142 ( .IN0(n3058), .IN1(n631), .SEL(n3057), .F(n598) );
  IV U1143 ( .A(n598), .Z(n2932) );
  AND U1144 ( .A(n1212), .B(n1214), .Z(n1120) );
  MUX U1145 ( .IN0(n599), .IN1(n1654), .SEL(n1655), .F(n1573) );
  IV U1146 ( .A(n1656), .Z(n599) );
  ANDN U1147 ( .A(n887), .B(n888), .Z(n879) );
  MUX U1148 ( .IN0(n1070), .IN1(Y0[25]), .SEL(n1071), .F(n1030) );
  MUX U1149 ( .IN0(n1280), .IN1(Y0[21]), .SEL(n1281), .F(n1217) );
  MUX U1150 ( .IN0(n1567), .IN1(Y0[17]), .SEL(n1568), .F(n1489) );
  MUX U1151 ( .IN0(n1920), .IN1(Y0[13]), .SEL(n1921), .F(n1823) );
  MUX U1152 ( .IN0(n2319), .IN1(Y0[9]), .SEL(n2320), .F(n2213) );
  MUX U1153 ( .IN0(n2773), .IN1(Y0[5]), .SEL(n2774), .F(n2653) );
  MUX U1154 ( .IN0(n906), .IN1(Y0[30]), .SEL(n907), .F(n872) );
  MUX U1155 ( .IN0(n3455), .IN1(n4136), .SEL(n3456), .F(n600) );
  IV U1156 ( .A(n600), .Z(n4094) );
  MUX U1157 ( .IN0(n601), .IN1(n4080), .SEL(n4081), .F(n4034) );
  IV U1158 ( .A(n4082), .Z(n601) );
  MUX U1159 ( .IN0(n4486), .IN1(n4484), .SEL(n4485), .F(n4463) );
  MUX U1160 ( .IN0(n4001), .IN1(n3999), .SEL(n4000), .F(n3953) );
  MUX U1161 ( .IN0(n602), .IN1(n3898), .SEL(n3899), .F(n3852) );
  IV U1162 ( .A(n3900), .Z(n602) );
  MUX U1163 ( .IN0(n4902), .IN1(n4432), .SEL(n4433), .F(n4885) );
  MUX U1164 ( .IN0(n3792), .IN1(n3790), .SEL(n3791), .F(n3746) );
  MUX U1165 ( .IN0(n4402), .IN1(n4400), .SEL(n4401), .F(n4379) );
  MUX U1166 ( .IN0(n3819), .IN1(n3817), .SEL(n3818), .F(n3771) );
  MUX U1167 ( .IN0(n5186), .IN1(n5339), .SEL(n5187), .F(n603) );
  IV U1168 ( .A(n603), .Z(n5319) );
  MUX U1169 ( .IN0(n604), .IN1(n3716), .SEL(n3717), .F(n3671) );
  IV U1170 ( .A(n3718), .Z(n604) );
  MUX U1171 ( .IN0(n4834), .IN1(n4348), .SEL(n4349), .F(n4818) );
  MUX U1172 ( .IN0(n5419), .IN1(n5277), .SEL(n5279), .F(n5407) );
  MUX U1173 ( .IN0(n3616), .IN1(n3614), .SEL(n3615), .F(n3572) );
  MUX U1174 ( .IN0(n5157), .IN1(n605), .SEL(n5158), .F(n5146) );
  IV U1175 ( .A(n5160), .Z(n605) );
  MUX U1176 ( .IN0(n4318), .IN1(n4316), .SEL(n4317), .F(n4296) );
  MUX U1177 ( .IN0(n3641), .IN1(n3639), .SEL(n3640), .F(n3596) );
  MUX U1178 ( .IN0(n5349), .IN1(n5351), .SEL(n5350), .F(n5345) );
  MUX U1179 ( .IN0(n4611), .IN1(n4609), .SEL(n4610), .F(n4589) );
  NANDN U1180 ( .B(n5628), .A(n3415), .Z(n640) );
  MUX U1181 ( .IN0(n606), .IN1(n3543), .SEL(n3544), .F(n3499) );
  IV U1182 ( .A(n3545), .Z(n606) );
  MUX U1183 ( .IN0(n2717), .IN1(n2719), .SEL(n2718), .F(n2597) );
  MUX U1184 ( .IN0(n3089), .IN1(n607), .SEL(n3090), .F(n2957) );
  IV U1185 ( .A(n3091), .Z(n607) );
  MUX U1186 ( .IN0(A[10]), .IN1(n5429), .SEL(A[31]), .F(n608) );
  IV U1187 ( .A(n608), .Z(n2526) );
  MUX U1188 ( .IN0(A[6]), .IN1(n5558), .SEL(A[31]), .F(n609) );
  IV U1189 ( .A(n609), .Z(n3012) );
  MUX U1190 ( .IN0(A[5]), .IN1(n5574), .SEL(A[31]), .F(n610) );
  IV U1191 ( .A(n610), .Z(n3144) );
  MUX U1192 ( .IN0(n4768), .IN1(n4265), .SEL(n4266), .F(n4748) );
  XNOR U1193 ( .A(n5004), .B(n5002), .Z(n5009) );
  MUX U1194 ( .IN0(n3467), .IN1(n3465), .SEL(n3466), .F(n3334) );
  MUX U1195 ( .IN0(n1141), .IN1(n611), .SEL(n1142), .F(n1099) );
  IV U1196 ( .A(n1143), .Z(n611) );
  MUX U1197 ( .IN0(n680), .IN1(n1609), .SEL(n1608), .F(n1520) );
  MUX U1198 ( .IN0(n1981), .IN1(n1979), .SEL(n1980), .F(n1883) );
  MUX U1199 ( .IN0(n612), .IN1(n2200), .SEL(n2201), .F(n2099) );
  IV U1200 ( .A(n2202), .Z(n612) );
  MUX U1201 ( .IN0(n2860), .IN1(n2858), .SEL(n2859), .F(n2736) );
  MUX U1202 ( .IN0(n2797), .IN1(n2795), .SEL(n2796), .F(n2675) );
  MUX U1203 ( .IN0(n2927), .IN1(n2925), .SEL(n2926), .F(n2803) );
  MUX U1204 ( .IN0(n3390), .IN1(n3388), .SEL(n3389), .F(n3247) );
  MUX U1205 ( .IN0(n3312), .IN1(n3310), .SEL(n3311), .F(n3171) );
  XNOR U1206 ( .A(n3404), .B(n3403), .Z(n5544) );
  XNOR U1207 ( .A(n3365), .B(n3364), .Z(n5174) );
  XNOR U1208 ( .A(n3318), .B(n3317), .Z(n3443) );
  MUX U1209 ( .IN0(n1366), .IN1(n1364), .SEL(n1365), .F(n1292) );
  MUX U1210 ( .IN0(n1197), .IN1(n1195), .SEL(n1196), .F(n1136) );
  XNOR U1211 ( .A(n1402), .B(n1401), .Z(n1469) );
  MUX U1212 ( .IN0(n1528), .IN1(n613), .SEL(n1527), .F(n1444) );
  IV U1213 ( .A(n1526), .Z(n613) );
  XNOR U1214 ( .A(n1466), .B(n1465), .Z(n1539) );
  XNOR U1215 ( .A(n1802), .B(n1801), .Z(n1894) );
  XNOR U1216 ( .A(n1810), .B(n1809), .Z(n1902) );
  XNOR U1217 ( .A(n1856), .B(n1855), .Z(n1945) );
  MUX U1218 ( .IN0(n614), .IN1(n2065), .SEL(n2066), .F(n1969) );
  IV U1219 ( .A(n2067), .Z(n614) );
  XNOR U1220 ( .A(n2091), .B(n2090), .Z(n2187) );
  MUX U1221 ( .IN0(n615), .IN1(n2290), .SEL(n2291), .F(n2184) );
  IV U1222 ( .A(n2292), .Z(n615) );
  XNOR U1223 ( .A(n2259), .B(n2258), .Z(n2361) );
  XNOR U1224 ( .A(n2348), .B(n2347), .Z(n2450) );
  XNOR U1225 ( .A(n2389), .B(n2388), .Z(n2492) );
  MUX U1226 ( .IN0(n616), .IN1(n2608), .SEL(n2609), .F(n2489) );
  IV U1227 ( .A(n2610), .Z(n616) );
  MUX U1228 ( .IN0(n617), .IN1(n2665), .SEL(n2666), .F(n2548) );
  IV U1229 ( .A(n2667), .Z(n617) );
  XNOR U1230 ( .A(n2713), .B(n2712), .Z(n2830) );
  XNOR U1231 ( .A(n2752), .B(n2751), .Z(n2869) );
  XNOR U1232 ( .A(n2760), .B(n2759), .Z(n2877) );
  XNOR U1233 ( .A(n3060), .B(n2942), .Z(n2943) );
  MUX U1234 ( .IN0(n618), .IN1(n3239), .SEL(n3240), .F(n3107) );
  IV U1235 ( .A(n3241), .Z(n618) );
  MUX U1236 ( .IN0(n3257), .IN1(n688), .SEL(n3256), .F(n619) );
  IV U1237 ( .A(n619), .Z(n3123) );
  MUX U1238 ( .IN0(n620), .IN1(n3215), .SEL(n3216), .F(n3082) );
  IV U1239 ( .A(n3217), .Z(n620) );
  MUX U1240 ( .IN0(n980), .IN1(n982), .SEL(n981), .F(n950) );
  XNOR U1241 ( .A(n1018), .B(n1017), .Z(n1051) );
  MUX U1242 ( .IN0(n621), .IN1(n1128), .SEL(n1129), .F(n1086) );
  IV U1243 ( .A(n1130), .Z(n621) );
  MUX U1244 ( .IN0(n622), .IN1(n1302), .SEL(n1303), .F(n1235) );
  IV U1245 ( .A(n1304), .Z(n622) );
  MUX U1246 ( .IN0(n623), .IN1(n1592), .SEL(n1593), .F(n1514) );
  IV U1247 ( .A(n1594), .Z(n623) );
  AND U1248 ( .A(n1820), .B(n1822), .Z(n1729) );
  MUX U1249 ( .IN0(n624), .IN1(n1959), .SEL(n1960), .F(n1863) );
  IV U1250 ( .A(n1961), .Z(n624) );
  XNOR U1251 ( .A(n1841), .B(n1842), .Z(n1838) );
  AND U1252 ( .A(n2041), .B(n2043), .Z(n1941) );
  AND U1253 ( .A(n2210), .B(n2212), .Z(n2109) );
  MUX U1254 ( .IN0(n625), .IN1(n2481), .SEL(n2482), .F(n2373) );
  IV U1255 ( .A(n2483), .Z(n625) );
  AND U1256 ( .A(n2770), .B(n2772), .Z(n2650) );
  MUX U1257 ( .IN0(n626), .IN1(n2967), .SEL(n2968), .F(n2842) );
  IV U1258 ( .A(n2969), .Z(n626) );
  MUX U1259 ( .IN0(n627), .IN1(n3079), .SEL(n3080), .F(n2951) );
  IV U1260 ( .A(n3081), .Z(n627) );
  NAND U1261 ( .A(n945), .B(n944), .Z(n939) );
  XNOR U1262 ( .A(n983), .B(n1008), .Z(n999) );
  ANDN U1263 ( .A(n1120), .B(n1121), .Z(n1076) );
  AND U1264 ( .A(n1168), .B(n1169), .Z(n1167) );
  ANDN U1265 ( .A(n1421), .B(n1422), .Z(n1354) );
  NAND U1266 ( .A(n1486), .B(n1488), .Z(n1413) );
  MUX U1267 ( .IN0(n628), .IN1(n2247), .SEL(n2248), .F(n2139) );
  IV U1268 ( .A(n2249), .Z(n628) );
  MUX U1269 ( .IN0(n629), .IN1(n2465), .SEL(n2466), .F(n2358) );
  IV U1270 ( .A(n2467), .Z(n629) );
  MUX U1271 ( .IN0(n630), .IN1(n2690), .SEL(n2691), .F(n2576) );
  IV U1272 ( .A(n2692), .Z(n630) );
  MUX U1273 ( .IN0(n3188), .IN1(n662), .SEL(n3187), .F(n631) );
  IV U1274 ( .A(n631), .Z(n3056) );
  XNOR U1275 ( .A(n956), .B(n961), .Z(n957) );
  XNOR U1276 ( .A(n1068), .B(n1073), .Z(n1069) );
  XNOR U1277 ( .A(n1215), .B(n1220), .Z(n1216) );
  XOR U1278 ( .A(n1654), .B(n1743), .Z(n1738) );
  XNOR U1279 ( .A(n3327), .B(n3326), .Z(n3156) );
  MUX U1280 ( .IN0(n1114), .IN1(Y0[24]), .SEL(n1115), .F(n1070) );
  MUX U1281 ( .IN0(n1348), .IN1(Y0[20]), .SEL(n1349), .F(n1280) );
  MUX U1282 ( .IN0(n1648), .IN1(Y0[16]), .SEL(n1649), .F(n1567) );
  MUX U1283 ( .IN0(n2016), .IN1(Y0[12]), .SEL(n2017), .F(n1920) );
  MUX U1284 ( .IN0(n2426), .IN1(Y0[8]), .SEL(n2427), .F(n2319) );
  MUX U1285 ( .IN0(Y0[4]), .IN1(n2894), .SEL(n2895), .F(n2773) );
  XNOR U1286 ( .A(n906), .B(n910), .Z(n908) );
  MUX U1287 ( .IN0(n4066), .IN1(n4064), .SEL(n4065), .F(n4018) );
  MUX U1288 ( .IN0(n4987), .IN1(n4537), .SEL(n4538), .F(n4970) );
  MUX U1289 ( .IN0(n632), .IN1(n4514), .SEL(n4054), .F(n4493) );
  IV U1290 ( .A(n4052), .Z(n632) );
  MUX U1291 ( .IN0(n4465), .IN1(n4463), .SEL(n4464), .F(n4442) );
  MUX U1292 ( .IN0(n3955), .IN1(n3953), .SEL(n3954), .F(n3909) );
  MUX U1293 ( .IN0(n633), .IN1(n3988), .SEL(n3989), .F(n3942) );
  IV U1294 ( .A(n3990), .Z(n633) );
  MUX U1295 ( .IN0(n3884), .IN1(n3882), .SEL(n3883), .F(n3836) );
  MUX U1296 ( .IN0(n4919), .IN1(n4453), .SEL(n4454), .F(n4902) );
  MUX U1297 ( .IN0(n4717), .IN1(n4715), .SEL(n4716), .F(n4693) );
  MUX U1298 ( .IN0(n634), .IN1(n4430), .SEL(n3872), .F(n4409) );
  IV U1299 ( .A(n3870), .Z(n634) );
  MUX U1300 ( .IN0(n5088), .IN1(n4700), .SEL(n4702), .F(n5076) );
  MUX U1301 ( .IN0(n4381), .IN1(n4379), .SEL(n4380), .F(n4358) );
  MUX U1302 ( .IN0(n3773), .IN1(n3771), .SEL(n3772), .F(n3727) );
  MUX U1303 ( .IN0(n635), .IN1(n3806), .SEL(n3807), .F(n3760) );
  IV U1304 ( .A(n3808), .Z(n635) );
  MUX U1305 ( .IN0(n3702), .IN1(n3700), .SEL(n3701), .F(n3657) );
  MUX U1306 ( .IN0(n4851), .IN1(n4369), .SEL(n4370), .F(n4834) );
  MUX U1307 ( .IN0(n5154), .IN1(n4740), .SEL(n4741), .F(n636) );
  IV U1308 ( .A(n636), .Z(n5140) );
  MUX U1309 ( .IN0(n5272), .IN1(n5270), .SEL(n5271), .F(n5250) );
  MUX U1310 ( .IN0(n4631), .IN1(n4629), .SEL(n4630), .F(n4609) );
  MUX U1311 ( .IN0(n637), .IN1(n4346), .SEL(n3690), .F(n4325) );
  IV U1312 ( .A(n3688), .Z(n637) );
  MUX U1313 ( .IN0(n5407), .IN1(n5257), .SEL(n5259), .F(n5395) );
  MUX U1314 ( .IN0(n4221), .IN1(n4223), .SEL(n4222), .F(n4218) );
  MUX U1315 ( .IN0(n5034), .IN1(n4616), .SEL(n4618), .F(n5024) );
  MUX U1316 ( .IN0(n4298), .IN1(n4296), .SEL(n4297), .F(n4275) );
  MUX U1317 ( .IN0(n3598), .IN1(n3596), .SEL(n3597), .F(n3554) );
  MUX U1318 ( .IN0(n638), .IN1(n3628), .SEL(n3629), .F(n3586) );
  IV U1319 ( .A(n3630), .Z(n638) );
  MUX U1320 ( .IN0(n3529), .IN1(n3527), .SEL(n3528), .F(n3487) );
  MUX U1321 ( .IN0(n639), .IN1(n4142), .SEL(n4143), .F(n4117) );
  IV U1322 ( .A(n4144), .Z(n639) );
  XNOR U1323 ( .A(n5623), .B(A[3]), .Z(n5624) );
  MUX U1324 ( .IN0(n4785), .IN1(n4286), .SEL(n4287), .F(n4768) );
  MUX U1325 ( .IN0(n5625), .IN1(n640), .SEL(n5626), .F(n3409) );
  MUX U1326 ( .IN0(n2502), .IN1(n2504), .SEL(n2503), .F(n2394) );
  MUX U1327 ( .IN0(n2757), .IN1(n641), .SEL(n2758), .F(n2637) );
  IV U1328 ( .A(n2759), .Z(n641) );
  MUX U1329 ( .IN0(n2972), .IN1(n2974), .SEL(n2973), .F(n2847) );
  MUX U1330 ( .IN0(n2929), .IN1(n2931), .SEL(n2930), .F(n2807) );
  MUX U1331 ( .IN0(n3252), .IN1(n3254), .SEL(n3253), .F(n3120) );
  XNOR U1332 ( .A(n5464), .B(n5463), .Z(n5469) );
  XNOR U1333 ( .A(n5179), .B(n5178), .Z(n5205) );
  XNOR U1334 ( .A(n4547), .B(n4545), .Z(n4560) );
  MUX U1335 ( .IN0(n642), .IN1(n4263), .SEL(n3518), .F(n4243) );
  IV U1336 ( .A(n3516), .Z(n642) );
  MUX U1337 ( .IN0(n1327), .IN1(n1325), .SEL(n1326), .F(n1257) );
  MUX U1338 ( .IN0(n1404), .IN1(n1402), .SEL(n1403), .F(n1335) );
  MUX U1339 ( .IN0(n643), .IN1(n5531), .SEL(X[31]), .F(n1523) );
  IV U1340 ( .A(X[19]), .Z(n643) );
  MUX U1341 ( .IN0(n644), .IN1(n1810), .SEL(n1811), .F(n1719) );
  IV U1342 ( .A(n1812), .Z(n644) );
  MUX U1343 ( .IN0(n645), .IN1(n4228), .SEL(X[31]), .F(n2028) );
  IV U1344 ( .A(X[13]), .Z(n645) );
  MUX U1345 ( .IN0(n2052), .IN1(n2050), .SEL(n2051), .F(n1952) );
  MUX U1346 ( .IN0(n2242), .IN1(n2240), .SEL(n2241), .F(n2123) );
  MUX U1347 ( .IN0(n646), .IN1(n2521), .SEL(n2522), .F(n2413) );
  IV U1348 ( .A(n2523), .Z(n646) );
  MUX U1349 ( .IN0(n2754), .IN1(n2752), .SEL(n2753), .F(n2632) );
  MUX U1350 ( .IN0(n3336), .IN1(n3334), .SEL(n3335), .F(n3195) );
  XNOR U1351 ( .A(n3388), .B(n3387), .Z(n5364) );
  MUX U1352 ( .IN0(n647), .IN1(n3430), .SEL(n3431), .F(n3302) );
  IV U1353 ( .A(n3432), .Z(n647) );
  XOR U1354 ( .A(n1358), .B(n1296), .Z(n1293) );
  MUX U1355 ( .IN0(n648), .IN1(n1456), .SEL(n1457), .F(n1384) );
  IV U1356 ( .A(n1458), .Z(n648) );
  ANDN U1357 ( .A(n1520), .B(n1519), .Z(n1447) );
  XNOR U1358 ( .A(n1625), .B(n1624), .Z(n1702) );
  MUX U1359 ( .IN0(n1682), .IN1(n649), .SEL(n1683), .F(n1605) );
  IV U1360 ( .A(n1684), .Z(n649) );
  XNOR U1361 ( .A(n1995), .B(n1994), .Z(n2086) );
  XNOR U1362 ( .A(n1979), .B(n1978), .Z(n2068) );
  MUX U1363 ( .IN0(n650), .IN1(n2166), .SEL(n2167), .F(n2065) );
  IV U1364 ( .A(n2168), .Z(n650) );
  MUX U1365 ( .IN0(n651), .IN1(n2184), .SEL(n2185), .F(n2083) );
  IV U1366 ( .A(n2186), .Z(n651) );
  XNOR U1367 ( .A(n2099), .B(n2098), .Z(n2195) );
  XNOR U1368 ( .A(n2282), .B(n2281), .Z(n2384) );
  MUX U1369 ( .IN0(n652), .IN1(n2624), .SEL(n2625), .F(n2505) );
  IV U1370 ( .A(n2626), .Z(n652) );
  XNOR U1371 ( .A(n2552), .B(n2562), .Z(n2668) );
  XNOR U1372 ( .A(n2569), .B(n2568), .Z(n2678) );
  XNOR U1373 ( .A(n2593), .B(n2592), .Z(n2708) );
  XNOR U1374 ( .A(n2616), .B(n2615), .Z(n2731) );
  MUX U1375 ( .IN0(n653), .IN1(n2850), .SEL(n2851), .F(n2728) );
  IV U1376 ( .A(n2852), .Z(n653) );
  XNOR U1377 ( .A(n2925), .B(n2924), .Z(n3044) );
  XNOR U1378 ( .A(n2917), .B(n2916), .Z(n3036) );
  XNOR U1379 ( .A(n2983), .B(n2982), .Z(n3110) );
  XNOR U1380 ( .A(n3092), .B(n3091), .Z(n3219) );
  XNOR U1381 ( .A(n3131), .B(n3130), .Z(n3258) );
  XNOR U1382 ( .A(n3139), .B(n3138), .Z(n3266) );
  MUX U1383 ( .IN0(n985), .IN1(n983), .SEL(n984), .F(n953) );
  NAND U1384 ( .A(n1096), .B(n1095), .Z(n1089) );
  XNOR U1385 ( .A(n1058), .B(n1057), .Z(n1097) );
  MUX U1386 ( .IN0(n654), .IN1(n1184), .SEL(n1185), .F(n1128) );
  IV U1387 ( .A(n1186), .Z(n654) );
  AND U1388 ( .A(n1729), .B(n1731), .Z(n1645) );
  MUX U1389 ( .IN0(n655), .IN1(n1763), .SEL(n1764), .F(n1672) );
  IV U1390 ( .A(n1765), .Z(n655) );
  MUX U1391 ( .IN0(n656), .IN1(n2266), .SEL(n2267), .F(n2158) );
  IV U1392 ( .A(n2268), .Z(n656) );
  AND U1393 ( .A(n2316), .B(n2318), .Z(n2210) );
  MUX U1394 ( .IN0(n657), .IN1(n2720), .SEL(n2721), .F(n2600) );
  IV U1395 ( .A(n2722), .Z(n657) );
  XNOR U1396 ( .A(n2701), .B(n2700), .Z(n2698) );
  ANDN U1397 ( .A(n2892), .B(n2893), .Z(n2770) );
  MUX U1398 ( .IN0(n3082), .IN1(n3205), .SEL(n3084), .F(n2949) );
  MUX U1399 ( .IN0(n3233), .IN1(n751), .SEL(n3232), .F(n658) );
  IV U1400 ( .A(n658), .Z(n3099) );
  MUX U1401 ( .IN0(n659), .IN1(n3202), .SEL(n3203), .F(n3079) );
  IV U1402 ( .A(n3204), .Z(n659) );
  ANDN U1403 ( .A(n1027), .B(n997), .Z(n986) );
  MUX U1404 ( .IN0(n1229), .IN1(n1231), .SEL(n1230), .F(n660) );
  IV U1405 ( .A(n660), .Z(n1174) );
  AND U1406 ( .A(n1286), .B(n1288), .Z(n1223) );
  XOR U1407 ( .A(n1238), .B(n1235), .Z(n1289) );
  NANDN U1408 ( .B(n1346), .A(n1347), .Z(n1278) );
  XNOR U1409 ( .A(n2023), .B(n2024), .Z(n2043) );
  MUX U1410 ( .IN0(n661), .IN1(n2810), .SEL(n2811), .F(n2690) );
  IV U1411 ( .A(n2812), .Z(n661) );
  MUX U1412 ( .IN0(n3327), .IN1(n3325), .SEL(n3326), .F(n662) );
  IV U1413 ( .A(n662), .Z(n3186) );
  MUX U1414 ( .IN0(n923), .IN1(n921), .SEL(n922), .F(n663) );
  IV U1415 ( .A(n663), .Z(n900) );
  NANDN U1416 ( .B(n927), .A(n928), .Z(n884) );
  XOR U1417 ( .A(n1516), .B(n1515), .Z(n1496) );
  XOR U1418 ( .A(n1745), .B(n1744), .Z(n1829) );
  XOR U1419 ( .A(n2358), .B(n2355), .Z(n2432) );
  AND U1420 ( .A(n912), .B(n914), .Z(n887) );
  MUX U1421 ( .IN0(n3281), .IN1(Y0[1]), .SEL(n3282), .F(n3149) );
  XNOR U1422 ( .A(n958), .B(n962), .Z(n960) );
  XNOR U1423 ( .A(n1070), .B(n1074), .Z(n1072) );
  XNOR U1424 ( .A(n1217), .B(n1221), .Z(n1219) );
  XNOR U1425 ( .A(n1415), .B(n1419), .Z(n1417) );
  XNOR U1426 ( .A(n1648), .B(n1652), .Z(n1650) );
  XNOR U1427 ( .A(n1920), .B(n1924), .Z(n1922) );
  XNOR U1428 ( .A(n2213), .B(n2217), .Z(n2215) );
  XNOR U1429 ( .A(n2534), .B(n2538), .Z(n2536) );
  MUX U1430 ( .IN0(n664), .IN1(n4556), .SEL(n4139), .F(n4535) );
  IV U1431 ( .A(n4138), .Z(n664) );
  MUX U1432 ( .IN0(n4020), .IN1(n4018), .SEL(n4019), .F(n3972) );
  MUX U1433 ( .IN0(n4507), .IN1(n4505), .SEL(n4506), .F(n4484) );
  MUX U1434 ( .IN0(n4953), .IN1(n4495), .SEL(n4496), .F(n4936) );
  MUX U1435 ( .IN0(n665), .IN1(n3942), .SEL(n3943), .F(n3898) );
  IV U1436 ( .A(n3944), .Z(n665) );
  MUX U1437 ( .IN0(n666), .IN1(n4472), .SEL(n3962), .F(n4451) );
  IV U1438 ( .A(n3960), .Z(n666) );
  MUX U1439 ( .IN0(n3838), .IN1(n3836), .SEL(n3837), .F(n3790) );
  MUX U1440 ( .IN0(n4423), .IN1(n4421), .SEL(n4422), .F(n4400) );
  MUX U1441 ( .IN0(n3865), .IN1(n3863), .SEL(n3864), .F(n3817) );
  MUX U1442 ( .IN0(n4885), .IN1(n4411), .SEL(n4412), .F(n4868) );
  MUX U1443 ( .IN0(n4234), .IN1(n4718), .SEL(n4235), .F(n667) );
  IV U1444 ( .A(n667), .Z(n4696) );
  MUX U1445 ( .IN0(n5076), .IN1(n4676), .SEL(n4678), .F(n5061) );
  MUX U1446 ( .IN0(n4671), .IN1(n4669), .SEL(n4670), .F(n4649) );
  MUX U1447 ( .IN0(n668), .IN1(n3760), .SEL(n3761), .F(n3716) );
  IV U1448 ( .A(n3762), .Z(n668) );
  MUX U1449 ( .IN0(n669), .IN1(n4388), .SEL(n3780), .F(n4367) );
  IV U1450 ( .A(n3778), .Z(n669) );
  MUX U1451 ( .IN0(n5294), .IN1(n5292), .SEL(n5293), .F(n5270) );
  MUX U1452 ( .IN0(n5433), .IN1(n5299), .SEL(n5301), .F(n5419) );
  MUX U1453 ( .IN0(n3659), .IN1(n3657), .SEL(n3658), .F(n3614) );
  MUX U1454 ( .IN0(n4339), .IN1(n4337), .SEL(n4338), .F(n4316) );
  MUX U1455 ( .IN0(n3683), .IN1(n3681), .SEL(n3682), .F(n3639) );
  MUX U1456 ( .IN0(n4818), .IN1(n4327), .SEL(n4328), .F(n4802) );
  MUX U1457 ( .IN0(A[1]), .IN1(n5640), .SEL(A[31]), .F(n670) );
  IV U1458 ( .A(n670), .Z(n4208) );
  MUX U1459 ( .IN0(n671), .IN1(n5559), .SEL(n5560), .F(n5548) );
  IV U1460 ( .A(n5561), .Z(n671) );
  MUX U1461 ( .IN0(n5024), .IN1(n4596), .SEL(n4598), .F(n5014) );
  MUX U1462 ( .IN0(n4591), .IN1(n4589), .SEL(n4590), .F(n4565) );
  MUX U1463 ( .IN0(n672), .IN1(n3586), .SEL(n3587), .F(n3543) );
  IV U1464 ( .A(n3588), .Z(n672) );
  MUX U1465 ( .IN0(n673), .IN1(n4305), .SEL(n3605), .F(n4284) );
  IV U1466 ( .A(n3603), .Z(n673) );
  XNOR U1467 ( .A(n5546), .B(A[7]), .Z(n5547) );
  XNOR U1468 ( .A(n5414), .B(A[11]), .Z(n5415) );
  XNOR U1469 ( .A(n5366), .B(A[15]), .Z(n5367) );
  XNOR U1470 ( .A(n4877), .B(A[23]), .Z(n4878) );
  XNOR U1471 ( .A(n4945), .B(A[19]), .Z(n4946) );
  MUX U1472 ( .IN0(A[2]), .IN1(n5633), .SEL(A[31]), .F(n674) );
  IV U1473 ( .A(n674), .Z(n4205) );
  MUX U1474 ( .IN0(n5212), .IN1(n5210), .SEL(n5211), .F(n5179) );
  MUX U1475 ( .IN0(n5383), .IN1(n5217), .SEL(n5219), .F(n5371) );
  MUX U1476 ( .IN0(n3489), .IN1(n3487), .SEL(n3488), .F(n3448) );
  MUX U1477 ( .IN0(n3511), .IN1(n3509), .SEL(n3510), .F(n3440) );
  XNOR U1478 ( .A(n4811), .B(A[27]), .Z(n4812) );
  MUX U1479 ( .IN0(n675), .IN1(n4215), .SEL(X[31]), .F(n2444) );
  IV U1480 ( .A(X[9]), .Z(n675) );
  MUX U1481 ( .IN0(n2964), .IN1(n2966), .SEL(n2965), .F(n2839) );
  MUX U1482 ( .IN0(n3183), .IN1(n3185), .SEL(n3184), .F(n3053) );
  MUX U1483 ( .IN0(A[4]), .IN1(n5592), .SEL(A[31]), .F(n3142) );
  MUX U1484 ( .IN0(n3409), .IN1(n676), .SEL(n3410), .F(n3268) );
  IV U1485 ( .A(n3411), .Z(n676) );
  MUX U1486 ( .IN0(A[9]), .IN1(n5443), .SEL(A[31]), .F(n677) );
  IV U1487 ( .A(n677), .Z(n2645) );
  MUX U1488 ( .IN0(n3377), .IN1(n3379), .SEL(n3378), .F(n3236) );
  MUX U1489 ( .IN0(X[1]), .IN1(n5172), .SEL(X[31]), .F(n678) );
  IV U1490 ( .A(n678), .Z(n4745) );
  XNOR U1491 ( .A(n4133), .B(n4131), .Z(n4147) );
  MUX U1492 ( .IN0(n1468), .IN1(n1466), .SEL(n1467), .F(n1394) );
  MUX U1493 ( .IN0(n679), .IN1(n1635), .SEL(n1636), .F(n1554) );
  IV U1494 ( .A(n1637), .Z(n679) );
  MUX U1495 ( .IN0(n1667), .IN1(n1665), .SEL(n1666), .F(n1583) );
  MUX U1496 ( .IN0(n1691), .IN1(n1693), .SEL(n1692), .F(n680) );
  MUX U1497 ( .IN0(n2093), .IN1(n2091), .SEL(n2092), .F(n1995) );
  MUX U1498 ( .IN0(n2677), .IN1(n2675), .SEL(n2676), .F(n2552) );
  MUX U1499 ( .IN0(n3197), .IN1(n3195), .SEL(n3196), .F(n3061) );
  MUX U1500 ( .IN0(n4748), .IN1(n4261), .SEL(n4262), .F(n681) );
  IV U1501 ( .A(n681), .Z(n3355) );
  XNOR U1502 ( .A(n5342), .B(n5339), .Z(n5340) );
  XNOR U1503 ( .A(n5645), .B(X[30]), .Z(n5643) );
  MUX U1504 ( .IN0(n682), .IN1(n1247), .SEL(n1248), .F(n1184) );
  IV U1505 ( .A(n1249), .Z(n682) );
  XNOR U1506 ( .A(n1709), .B(n1708), .Z(n1797) );
  MUX U1507 ( .IN0(n683), .IN1(n1873), .SEL(n1874), .F(n1773) );
  IV U1508 ( .A(n1875), .Z(n683) );
  MUX U1509 ( .IN0(n684), .IN1(n1987), .SEL(n1988), .F(n1891) );
  IV U1510 ( .A(n1989), .Z(n684) );
  XNOR U1511 ( .A(n1907), .B(n1906), .Z(n1998) );
  XNOR U1512 ( .A(n1952), .B(n1951), .Z(n2045) );
  XNOR U1513 ( .A(n2075), .B(n2074), .Z(n2169) );
  XNOR U1514 ( .A(n2240), .B(n2239), .Z(n2341) );
  XNOR U1515 ( .A(n2405), .B(n2404), .Z(n2508) );
  XNOR U1516 ( .A(n2413), .B(n2412), .Z(n2516) );
  XNOR U1517 ( .A(n2366), .B(n2365), .Z(n2469) );
  MUX U1518 ( .IN0(n685), .IN1(n2489), .SEL(n2490), .F(n2381) );
  IV U1519 ( .A(n2491), .Z(n685) );
  XNOR U1520 ( .A(n2736), .B(n2735), .Z(n2853) );
  MUX U1521 ( .IN0(n686), .IN1(n2866), .SEL(n2867), .F(n2744) );
  IV U1522 ( .A(n2868), .Z(n686) );
  XNOR U1523 ( .A(n2683), .B(n2682), .Z(n2798) );
  MUX U1524 ( .IN0(n687), .IN1(n2785), .SEL(n2786), .F(n2665) );
  IV U1525 ( .A(n2787), .Z(n687) );
  XNOR U1526 ( .A(n2999), .B(n2998), .Z(n3126) );
  XNOR U1527 ( .A(n3007), .B(n3006), .Z(n3134) );
  XNOR U1528 ( .A(n2960), .B(n2959), .Z(n3087) );
  XNOR U1529 ( .A(n3115), .B(n3114), .Z(n3242) );
  XNOR U1530 ( .A(n3049), .B(n3048), .Z(n3174) );
  XNOR U1531 ( .A(n3041), .B(n3040), .Z(n3166) );
  MUX U1532 ( .IN0(n3398), .IN1(n3396), .SEL(n3397), .F(n688) );
  IV U1533 ( .A(n688), .Z(n3255) );
  MUX U1534 ( .IN0(n689), .IN1(n3380), .SEL(n3381), .F(n3239) );
  IV U1535 ( .A(n3382), .Z(n689) );
  MUX U1536 ( .IN0(n690), .IN1(n3302), .SEL(n3303), .F(n3163) );
  IV U1537 ( .A(n3304), .Z(n690) );
  MUX U1538 ( .IN0(n3352), .IN1(n691), .SEL(n3353), .F(n3215) );
  IV U1539 ( .A(n3354), .Z(n691) );
  MUX U1540 ( .IN0(n976), .IN1(n974), .SEL(n975), .F(n941) );
  MUX U1541 ( .IN0(n692), .IN1(n1045), .SEL(n1046), .F(n1009) );
  IV U1542 ( .A(n1047), .Z(n692) );
  XNOR U1543 ( .A(n1102), .B(n1101), .Z(n1139) );
  XNOR U1544 ( .A(n1136), .B(n1134), .Z(n1187) );
  AND U1545 ( .A(n1238), .B(n1239), .Z(n1168) );
  MUX U1546 ( .IN0(n693), .IN1(n1371), .SEL(n1372), .F(n1302) );
  IV U1547 ( .A(n1373), .Z(n693) );
  XOR U1548 ( .A(n1444), .B(n1448), .Z(n1517) );
  XNOR U1549 ( .A(n1930), .B(n1929), .Z(n1928) );
  MUX U1550 ( .IN0(n694), .IN1(n2057), .SEL(n2058), .F(n1959) );
  IV U1551 ( .A(n2059), .Z(n694) );
  AND U1552 ( .A(n2109), .B(n2111), .Z(n2013) );
  MUX U1553 ( .IN0(n695), .IN1(n2121), .SEL(n2120), .F(n2024) );
  IV U1554 ( .A(n2119), .Z(n695) );
  AND U1555 ( .A(n2531), .B(n2533), .Z(n2423) );
  MUX U1556 ( .IN0(n696), .IN1(n2600), .SEL(n2601), .F(n2481) );
  IV U1557 ( .A(n2602), .Z(n696) );
  MUX U1558 ( .IN0(n697), .IN1(n3099), .SEL(n3100), .F(n2967) );
  IV U1559 ( .A(n3101), .Z(n697) );
  MUX U1560 ( .IN0(n950), .IN1(n952), .SEL(n951), .F(n918) );
  AND U1561 ( .A(n1173), .B(n1174), .Z(n1170) );
  MUX U1562 ( .IN0(n698), .IN1(n2139), .SEL(n2140), .F(n2038) );
  IV U1563 ( .A(n2141), .Z(n698) );
  XOR U1564 ( .A(n2579), .B(n2465), .Z(n2466) );
  XNOR U1565 ( .A(n2826), .B(n2824), .Z(n2935) );
  NANDN U1566 ( .B(n925), .A(n924), .Z(n896) );
  XNOR U1567 ( .A(n927), .B(n932), .Z(n928) );
  XNOR U1568 ( .A(n1028), .B(n1033), .Z(n1029) );
  XNOR U1569 ( .A(n1156), .B(n1121), .Z(n1157) );
  XNOR U1570 ( .A(n1346), .B(n1351), .Z(n1347) );
  XOR U1571 ( .A(n1594), .B(n1593), .Z(n1574) );
  MUX U1572 ( .IN0(Y0[2]), .IN1(n3149), .SEL(n3150), .F(n3017) );
  XOR U1573 ( .A(n1747), .B(n1746), .Z(n1826) );
  XOR U1574 ( .A(n2357), .B(n2356), .Z(n2429) );
  XOR U1575 ( .A(n2692), .B(n2691), .Z(n2776) );
  XNOR U1576 ( .A(n3022), .B(n2901), .Z(n2902) );
  XOR U1577 ( .A(n3188), .B(n3187), .Z(n3293) );
  XNOR U1578 ( .A(n989), .B(n993), .Z(n991) );
  XNOR U1579 ( .A(n1114), .B(n1118), .Z(n1116) );
  XNOR U1580 ( .A(n1280), .B(n1284), .Z(n1282) );
  XNOR U1581 ( .A(n1489), .B(n1493), .Z(n1491) );
  XNOR U1582 ( .A(n1732), .B(n1736), .Z(n1734) );
  XNOR U1583 ( .A(n2016), .B(n2020), .Z(n2018) );
  XNOR U1584 ( .A(n2319), .B(n2323), .Z(n2321) );
  XNOR U1585 ( .A(n2653), .B(n2657), .Z(n2655) );
  XOR U1586 ( .A(n872), .B(n873), .Z(n755) );
  MUX U1587 ( .IN0(n4110), .IN1(n4108), .SEL(n4109), .F(n4064) );
  MUX U1588 ( .IN0(n4093), .IN1(n4091), .SEL(n4092), .F(n4045) );
  MUX U1589 ( .IN0(n699), .IN1(n4034), .SEL(n4035), .F(n3988) );
  IV U1590 ( .A(n4036), .Z(n699) );
  MUX U1591 ( .IN0(n3930), .IN1(n3928), .SEL(n3929), .F(n3882) );
  MUX U1592 ( .IN0(n700), .IN1(n4493), .SEL(n4008), .F(n4472) );
  IV U1593 ( .A(n4006), .Z(n700) );
  MUX U1594 ( .IN0(n4936), .IN1(n4474), .SEL(n4475), .F(n4919) );
  MUX U1595 ( .IN0(n4444), .IN1(n4442), .SEL(n4443), .F(n4421) );
  MUX U1596 ( .IN0(n3911), .IN1(n3909), .SEL(n3910), .F(n3863) );
  MUX U1597 ( .IN0(n701), .IN1(n3852), .SEL(n3853), .F(n3806) );
  IV U1598 ( .A(n3854), .Z(n701) );
  MUX U1599 ( .IN0(n3748), .IN1(n3746), .SEL(n3747), .F(n3700) );
  MUX U1600 ( .IN0(n702), .IN1(n4409), .SEL(n3826), .F(n4388) );
  IV U1601 ( .A(n3824), .Z(n702) );
  MUX U1602 ( .IN0(n4868), .IN1(n4390), .SEL(n4391), .F(n4851) );
  MUX U1603 ( .IN0(n5318), .IN1(n5316), .SEL(n5317), .F(n5292) );
  MUX U1604 ( .IN0(n5450), .IN1(n5323), .SEL(n5325), .F(n5433) );
  MUX U1605 ( .IN0(n4360), .IN1(n4358), .SEL(n4359), .F(n4337) );
  MUX U1606 ( .IN0(n3729), .IN1(n3727), .SEL(n3728), .F(n3681) );
  MUX U1607 ( .IN0(n5061), .IN1(n4656), .SEL(n4658), .F(n5046) );
  MUX U1608 ( .IN0(n4651), .IN1(n4649), .SEL(n4650), .F(n4629) );
  MUX U1609 ( .IN0(n5518), .IN1(n5362), .SEL(n5363), .F(n703) );
  IV U1610 ( .A(n703), .Z(n5504) );
  MUX U1611 ( .IN0(n4194), .IN1(n4145), .SEL(n4146), .F(n704) );
  IV U1612 ( .A(n704), .Z(n4180) );
  MUX U1613 ( .IN0(n705), .IN1(n4177), .SEL(n4178), .F(n4163) );
  IV U1614 ( .A(n4179), .Z(n705) );
  MUX U1615 ( .IN0(n706), .IN1(n3671), .SEL(n3672), .F(n3628) );
  IV U1616 ( .A(n3673), .Z(n706) );
  MUX U1617 ( .IN0(n5601), .IN1(n5542), .SEL(n5543), .F(n707) );
  IV U1618 ( .A(n707), .Z(n5585) );
  MUX U1619 ( .IN0(n3574), .IN1(n3572), .SEL(n3573), .F(n3527) );
  MUX U1620 ( .IN0(n708), .IN1(n4325), .SEL(n3648), .F(n4305) );
  IV U1621 ( .A(n3646), .Z(n708) );
  MUX U1622 ( .IN0(n4802), .IN1(n4307), .SEL(n4308), .F(n4785) );
  MUX U1623 ( .IN0(n5629), .IN1(n5631), .SEL(n5630), .F(n5625) );
  MUX U1624 ( .IN0(n5232), .IN1(n5230), .SEL(n5231), .F(n5210) );
  MUX U1625 ( .IN0(n5395), .IN1(n5237), .SEL(n5239), .F(n5383) );
  MUX U1626 ( .IN0(n709), .IN1(n4149), .SEL(n4150), .F(n4127) );
  IV U1627 ( .A(n4151), .Z(n709) );
  MUX U1628 ( .IN0(n4277), .IN1(n4275), .SEL(n4276), .F(n4251) );
  MUX U1629 ( .IN0(n3556), .IN1(n3554), .SEL(n3555), .F(n3509) );
  XNOR U1630 ( .A(n5573), .B(A[5]), .Z(n5574) );
  XNOR U1631 ( .A(n5442), .B(A[9]), .Z(n5443) );
  MUX U1632 ( .IN0(n710), .IN1(n5356), .SEL(X[31]), .F(n5348) );
  IV U1633 ( .A(X[21]), .Z(n710) );
  XNOR U1634 ( .A(n5390), .B(A[13]), .Z(n5391) );
  XNOR U1635 ( .A(n4979), .B(A[17]), .Z(n4980) );
  XNOR U1636 ( .A(n4911), .B(A[21]), .Z(n4912) );
  AND U1637 ( .A(n5641), .B(A[0]), .Z(n3419) );
  MUX U1638 ( .IN0(n4567), .IN1(n4565), .SEL(n4566), .F(n4547) );
  MUX U1639 ( .IN0(n5014), .IN1(n4576), .SEL(n4578), .F(n5004) );
  MUX U1640 ( .IN0(n711), .IN1(n5620), .SEL(X[31]), .F(n5607) );
  IV U1641 ( .A(X[25]), .Z(n711) );
  XNOR U1642 ( .A(n4843), .B(A[25]), .Z(n4844) );
  MUX U1643 ( .IN0(n712), .IN1(n5638), .SEL(X[31]), .F(n5628) );
  IV U1644 ( .A(X[29]), .Z(n712) );
  MUX U1645 ( .IN0(A[3]), .IN1(n5624), .SEL(A[31]), .F(n3274) );
  MUX U1646 ( .IN0(n3393), .IN1(n3395), .SEL(n3394), .F(n3252) );
  MUX U1647 ( .IN0(n3369), .IN1(n3371), .SEL(n3370), .F(n3228) );
  MUX U1648 ( .IN0(X[20]), .IN1(n713), .SEL(X[31]), .F(n1426) );
  IV U1649 ( .A(n5355), .Z(n713) );
  MUX U1650 ( .IN0(X[16]), .IN1(n714), .SEL(X[31]), .F(n1788) );
  IV U1651 ( .A(n5535), .Z(n714) );
  MUX U1652 ( .IN0(X[8]), .IN1(n715), .SEL(X[31]), .F(n2563) );
  IV U1653 ( .A(n4214), .Z(n715) );
  MUX U1654 ( .IN0(X[12]), .IN1(n716), .SEL(X[31]), .F(n2134) );
  IV U1655 ( .A(n4227), .Z(n716) );
  MUX U1656 ( .IN0(X[4]), .IN1(n717), .SEL(X[31]), .F(n3072) );
  IV U1657 ( .A(n4733), .Z(n717) );
  XNOR U1658 ( .A(n4721), .B(n4718), .Z(n4719) );
  MUX U1659 ( .IN0(n718), .IN1(n3499), .SEL(n3500), .F(n3430) );
  IV U1660 ( .A(n3501), .Z(n718) );
  MUX U1661 ( .IN0(n719), .IN1(n5614), .SEL(X[31]), .F(n1041) );
  IV U1662 ( .A(X[27]), .Z(n719) );
  MUX U1663 ( .IN0(X[26]), .IN1(n720), .SEL(X[31]), .F(n1082) );
  IV U1664 ( .A(n5615), .Z(n720) );
  MUX U1665 ( .IN0(X[24]), .IN1(n721), .SEL(X[31]), .F(n1189) );
  IV U1666 ( .A(n5619), .Z(n721) );
  MUX U1667 ( .IN0(X[28]), .IN1(n722), .SEL(X[31]), .F(n1014) );
  IV U1668 ( .A(n5637), .Z(n722) );
  MUX U1669 ( .IN0(n1507), .IN1(n1505), .SEL(n1506), .F(n1432) );
  MUX U1670 ( .IN0(n723), .IN1(n1554), .SEL(n1555), .F(n1476) );
  IV U1671 ( .A(n1556), .Z(n723) );
  MUX U1672 ( .IN0(n1548), .IN1(n1546), .SEL(n1547), .F(n1466) );
  MUX U1673 ( .IN0(X[18]), .IN1(n724), .SEL(X[31]), .F(n1604) );
  IV U1674 ( .A(n5530), .Z(n724) );
  MUX U1675 ( .IN0(n725), .IN1(n5536), .SEL(X[31]), .F(n1688) );
  IV U1676 ( .A(X[17]), .Z(n725) );
  MUX U1677 ( .IN0(n1885), .IN1(n1883), .SEL(n1884), .F(n1777) );
  MUX U1678 ( .IN0(n1858), .IN1(n1856), .SEL(n1857), .F(n1754) );
  MUX U1679 ( .IN0(n1901), .IN1(n1899), .SEL(n1900), .F(n1802) );
  MUX U1680 ( .IN0(n726), .IN1(n1907), .SEL(n1908), .F(n1810) );
  IV U1681 ( .A(n1909), .Z(n726) );
  XNOR U1682 ( .A(n4777), .B(A[29]), .Z(n4778) );
  MUX U1683 ( .IN0(n727), .IN1(n4210), .SEL(X[31]), .F(n2227) );
  IV U1684 ( .A(X[11]), .Z(n727) );
  MUX U1685 ( .IN0(X[10]), .IN1(n728), .SEL(X[31]), .F(n2333) );
  IV U1686 ( .A(n4209), .Z(n728) );
  MUX U1687 ( .IN0(n2457), .IN1(n2455), .SEL(n2456), .F(n2348) );
  MUX U1688 ( .IN0(X[6]), .IN1(n729), .SEL(X[31]), .F(n2823) );
  IV U1689 ( .A(n4738), .Z(n729) );
  MUX U1690 ( .IN0(n730), .IN1(n4734), .SEL(X[31]), .F(n2939) );
  IV U1691 ( .A(X[5]), .Z(n730) );
  MUX U1692 ( .IN0(n731), .IN1(n5168), .SEL(X[31]), .F(n3212) );
  IV U1693 ( .A(X[3]), .Z(n731) );
  MUX U1694 ( .IN0(X[2]), .IN1(n732), .SEL(X[31]), .F(n3351) );
  IV U1695 ( .A(n5167), .Z(n732) );
  MUX U1696 ( .IN0(n4243), .IN1(n733), .SEL(n3480), .F(n3352) );
  IV U1697 ( .A(n3479), .Z(n733) );
  MUX U1698 ( .IN0(X[22]), .IN1(n734), .SEL(X[31]), .F(n1298) );
  IV U1699 ( .A(n5361), .Z(n734) );
  MUX U1700 ( .IN0(n735), .IN1(n5360), .SEL(X[31]), .F(n1228) );
  IV U1701 ( .A(X[23]), .Z(n735) );
  MUX U1702 ( .IN0(n736), .IN1(n1315), .SEL(n1316), .F(n1247) );
  IV U1703 ( .A(n1317), .Z(n736) );
  MUX U1704 ( .IN0(n737), .IN1(n1615), .SEL(n1616), .F(n1536) );
  IV U1705 ( .A(n1617), .Z(n737) );
  MUX U1706 ( .IN0(n2033), .IN1(n2031), .SEL(n2032), .F(n738) );
  MUX U1707 ( .IN0(X[14]), .IN1(n739), .SEL(X[31]), .F(n1937) );
  IV U1708 ( .A(n4232), .Z(n739) );
  MUX U1709 ( .IN0(n740), .IN1(n1969), .SEL(n1970), .F(n1873) );
  IV U1710 ( .A(n1971), .Z(n740) );
  XNOR U1711 ( .A(n2192), .B(n2191), .Z(n2293) );
  XNOR U1712 ( .A(n2200), .B(n2199), .Z(n2301) );
  XNOR U1713 ( .A(n2151), .B(n2150), .Z(n2254) );
  XNOR U1714 ( .A(n2176), .B(n2175), .Z(n2277) );
  MUX U1715 ( .IN0(n741), .IN1(n2381), .SEL(n2382), .F(n2274) );
  IV U1716 ( .A(n2383), .Z(n741) );
  MUX U1717 ( .IN0(n742), .IN1(n2397), .SEL(n2398), .F(n2290) );
  IV U1718 ( .A(n2399), .Z(n742) );
  MUX U1719 ( .IN0(n2337), .IN1(n2441), .SEL(n2339), .F(n2229) );
  XNOR U1720 ( .A(n2497), .B(n2496), .Z(n2611) );
  XNOR U1721 ( .A(n2474), .B(n2473), .Z(n2588) );
  XNOR U1722 ( .A(n2513), .B(n2512), .Z(n2627) );
  XNOR U1723 ( .A(n2521), .B(n2520), .Z(n2635) );
  MUX U1724 ( .IN0(n743), .IN1(n2548), .SEL(n2549), .F(n2438) );
  IV U1725 ( .A(n2550), .Z(n743) );
  MUX U1726 ( .IN0(n744), .IN1(n4739), .SEL(X[31]), .F(n2697) );
  IV U1727 ( .A(X[7]), .Z(n744) );
  XNOR U1728 ( .A(n2882), .B(n2881), .Z(n3002) );
  XNOR U1729 ( .A(n2874), .B(n2873), .Z(n2994) );
  XNOR U1730 ( .A(n2835), .B(n2834), .Z(n2955) );
  XNOR U1731 ( .A(n2858), .B(n2857), .Z(n2978) );
  XNOR U1732 ( .A(n2795), .B(n2794), .Z(n2912) );
  XNOR U1733 ( .A(n2803), .B(n2802), .Z(n2920) );
  MUX U1734 ( .IN0(n745), .IN1(n3033), .SEL(n3034), .F(n2909) );
  IV U1735 ( .A(n3035), .Z(n745) );
  MUX U1736 ( .IN0(n746), .IN1(n3123), .SEL(n3124), .F(n2991) );
  IV U1737 ( .A(n3125), .Z(n746) );
  MUX U1738 ( .IN0(n747), .IN1(n3107), .SEL(n3108), .F(n2975) );
  IV U1739 ( .A(n3109), .Z(n747) );
  XNOR U1740 ( .A(n3271), .B(n3270), .Z(n3407) );
  XNOR U1741 ( .A(n3263), .B(n3262), .Z(n3399) );
  XNOR U1742 ( .A(n3224), .B(n3223), .Z(n3360) );
  XNOR U1743 ( .A(n3247), .B(n3246), .Z(n3383) );
  XNOR U1744 ( .A(n3171), .B(n3170), .Z(n3305) );
  XNOR U1745 ( .A(n3179), .B(n3178), .Z(n3313) );
  MUX U1746 ( .IN0(n3355), .IN1(n4742), .SEL(n3357), .F(n3214) );
  XNOR U1747 ( .A(n3195), .B(n3194), .Z(n3329) );
  MUX U1748 ( .IN0(X[30]), .IN1(n748), .SEL(X[31]), .F(n948) );
  IV U1749 ( .A(n5643), .Z(n748) );
  XNOR U1750 ( .A(n1091), .B(n1095), .Z(n1131) );
  NAND U1751 ( .A(n1296), .B(n1295), .Z(n1290) );
  MUX U1752 ( .IN0(n1299), .IN1(n1301), .SEL(n1300), .F(n1229) );
  XNOR U1753 ( .A(n1144), .B(n1143), .Z(n1198) );
  NAND U1754 ( .A(n1447), .B(n1448), .Z(n1442) );
  MUX U1755 ( .IN0(n749), .IN1(n1863), .SEL(n1864), .F(n1763) );
  IV U1756 ( .A(n1865), .Z(n749) );
  MUX U1757 ( .IN0(n750), .IN1(n4233), .SEL(X[31]), .F(n1836) );
  IV U1758 ( .A(X[15]), .Z(n750) );
  AND U1759 ( .A(n1917), .B(n1919), .Z(n1820) );
  ANDN U1760 ( .A(n2358), .B(n2359), .Z(n2250) );
  MUX U1761 ( .IN0(n3374), .IN1(n3372), .SEL(n3373), .F(n751) );
  IV U1762 ( .A(n751), .Z(n3231) );
  MUX U1763 ( .IN0(n752), .IN1(n3341), .SEL(n3342), .F(n3202) );
  IV U1764 ( .A(n3343), .Z(n752) );
  MUX U1765 ( .IN0(n943), .IN1(n941), .SEL(n942), .F(n921) );
  ANDN U1766 ( .A(n953), .B(n954), .Z(n924) );
  MUX U1767 ( .IN0(n753), .IN1(n1176), .SEL(n1177), .F(n1153) );
  IV U1768 ( .A(n1178), .Z(n753) );
  XNOR U1769 ( .A(n1838), .B(n1837), .Z(n1831) );
  XNOR U1770 ( .A(n2704), .B(n2699), .Z(n2813) );
  MUX U1771 ( .IN0(n918), .IN1(n920), .SEL(n919), .F(n754) );
  IV U1772 ( .A(n754), .Z(n903) );
  XNOR U1773 ( .A(n987), .B(n992), .Z(n988) );
  XNOR U1774 ( .A(n1112), .B(n1117), .Z(n1113) );
  XNOR U1775 ( .A(n1278), .B(n1283), .Z(n1279) );
  XOR U1776 ( .A(n1441), .B(n1440), .Z(n1422) );
  XOR U1777 ( .A(n1674), .B(n1673), .Z(n1656) );
  XOR U1778 ( .A(n1940), .B(n1939), .Z(n2019) );
  XOR U1779 ( .A(n2141), .B(n2140), .Z(n2216) );
  XOR U1780 ( .A(n2249), .B(n2248), .Z(n2322) );
  XOR U1781 ( .A(n2464), .B(n2463), .Z(n2537) );
  XOR U1782 ( .A(n2578), .B(n2577), .Z(n2656) );
  XOR U1783 ( .A(n2812), .B(n2811), .Z(n2898) );
  XOR U1784 ( .A(n2934), .B(n2933), .Z(n3022) );
  XOR U1785 ( .A(n3058), .B(n3057), .Z(n3152) );
  AND U1786 ( .A(Y0[0]), .B(n3156), .Z(n3281) );
  XNOR U1787 ( .A(n929), .B(n933), .Z(n931) );
  XNOR U1788 ( .A(n1030), .B(n1034), .Z(n1032) );
  XNOR U1789 ( .A(n1158), .B(n1161), .Z(n1160) );
  XNOR U1790 ( .A(n1348), .B(n1352), .Z(n1350) );
  XNOR U1791 ( .A(n1567), .B(n1571), .Z(n1569) );
  XNOR U1792 ( .A(n1823), .B(n1827), .Z(n1825) );
  XNOR U1793 ( .A(n2112), .B(n2116), .Z(n2114) );
  XNOR U1794 ( .A(n2426), .B(n2430), .Z(n2428) );
  XNOR U1795 ( .A(n2773), .B(n2777), .Z(n2775) );
  MUX U1796 ( .IN0(n755), .IN1(n864), .SEL(n870), .F(n867) );
  ANDN U1797 ( .A(n756), .B(n[0]), .Z(n390) );
  AND U1798 ( .A(N8), .B(n756), .Z(n389) );
  AND U1799 ( .A(N9), .B(n756), .Z(n388) );
  AND U1800 ( .A(N10), .B(n756), .Z(n387) );
  AND U1801 ( .A(N11), .B(n756), .Z(n386) );
  AND U1802 ( .A(N12), .B(n756), .Z(n385) );
  AND U1803 ( .A(N13), .B(n756), .Z(n384) );
  AND U1804 ( .A(N14), .B(n756), .Z(n383) );
  AND U1805 ( .A(N15), .B(n756), .Z(n382) );
  AND U1806 ( .A(N16), .B(n756), .Z(n381) );
  AND U1807 ( .A(N17), .B(n756), .Z(n380) );
  AND U1808 ( .A(N18), .B(n756), .Z(n379) );
  AND U1809 ( .A(N19), .B(n756), .Z(n378) );
  AND U1810 ( .A(n756), .B(n757), .Z(n377) );
  XOR U1811 ( .A(n[13]), .B(\add_25/carry[13] ), .Z(n757) );
  ANDN U1812 ( .A(n758), .B(rst), .Z(n756) );
  NAND U1813 ( .A(n759), .B(n760), .Z(n758) );
  AND U1814 ( .A(n761), .B(n762), .Z(n760) );
  AND U1815 ( .A(n763), .B(n764), .Z(n762) );
  AND U1816 ( .A(n765), .B(n766), .Z(n764) );
  AND U1817 ( .A(n[13]), .B(n767), .Z(n761) );
  AND U1818 ( .A(n[10]), .B(n[0]), .Z(n767) );
  AND U1819 ( .A(n768), .B(n769), .Z(n759) );
  AND U1820 ( .A(n[3]), .B(n770), .Z(n769) );
  AND U1821 ( .A(n[1]), .B(n[2]), .Z(n770) );
  AND U1822 ( .A(n[8]), .B(n[9]), .Z(n768) );
  NAND U1823 ( .A(n771), .B(n772), .Z(n376) );
  NAND U1824 ( .A(n773), .B(n774), .Z(n772) );
  NAND U1825 ( .A(Y0[0]), .B(rst), .Z(n771) );
  NAND U1826 ( .A(n775), .B(n776), .Z(n375) );
  NAND U1827 ( .A(n777), .B(n774), .Z(n776) );
  NAND U1828 ( .A(Y0[1]), .B(rst), .Z(n775) );
  NAND U1829 ( .A(n778), .B(n779), .Z(n374) );
  NAND U1830 ( .A(n780), .B(n774), .Z(n779) );
  NAND U1831 ( .A(Y0[2]), .B(rst), .Z(n778) );
  NAND U1832 ( .A(n781), .B(n782), .Z(n373) );
  NAND U1833 ( .A(n783), .B(n774), .Z(n782) );
  NAND U1834 ( .A(Y0[3]), .B(rst), .Z(n781) );
  NAND U1835 ( .A(n784), .B(n785), .Z(n372) );
  NAND U1836 ( .A(n786), .B(n774), .Z(n785) );
  NAND U1837 ( .A(Y0[4]), .B(rst), .Z(n784) );
  NAND U1838 ( .A(n787), .B(n788), .Z(n371) );
  NAND U1839 ( .A(n789), .B(n774), .Z(n788) );
  NAND U1840 ( .A(rst), .B(Y0[5]), .Z(n787) );
  NAND U1841 ( .A(n790), .B(n791), .Z(n370) );
  NAND U1842 ( .A(n792), .B(n774), .Z(n791) );
  NAND U1843 ( .A(rst), .B(Y0[6]), .Z(n790) );
  NAND U1844 ( .A(n793), .B(n794), .Z(n369) );
  NAND U1845 ( .A(n795), .B(n774), .Z(n794) );
  NAND U1846 ( .A(rst), .B(Y0[7]), .Z(n793) );
  NAND U1847 ( .A(n796), .B(n797), .Z(n368) );
  NAND U1848 ( .A(n798), .B(n774), .Z(n797) );
  NAND U1849 ( .A(rst), .B(Y0[8]), .Z(n796) );
  NAND U1850 ( .A(n799), .B(n800), .Z(n367) );
  NAND U1851 ( .A(n801), .B(n774), .Z(n800) );
  NAND U1852 ( .A(rst), .B(Y0[9]), .Z(n799) );
  NAND U1853 ( .A(n802), .B(n803), .Z(n366) );
  NAND U1854 ( .A(n804), .B(n774), .Z(n803) );
  NAND U1855 ( .A(rst), .B(Y0[10]), .Z(n802) );
  NAND U1856 ( .A(n805), .B(n806), .Z(n365) );
  NAND U1857 ( .A(n807), .B(n774), .Z(n806) );
  NAND U1858 ( .A(rst), .B(Y0[11]), .Z(n805) );
  NAND U1859 ( .A(n808), .B(n809), .Z(n364) );
  NAND U1860 ( .A(n810), .B(n774), .Z(n809) );
  NAND U1861 ( .A(rst), .B(Y0[12]), .Z(n808) );
  NAND U1862 ( .A(n811), .B(n812), .Z(n363) );
  NAND U1863 ( .A(n813), .B(n774), .Z(n812) );
  NAND U1864 ( .A(rst), .B(Y0[13]), .Z(n811) );
  NAND U1865 ( .A(n814), .B(n815), .Z(n362) );
  NAND U1866 ( .A(n816), .B(n774), .Z(n815) );
  NAND U1867 ( .A(rst), .B(Y0[14]), .Z(n814) );
  NAND U1868 ( .A(n817), .B(n818), .Z(n361) );
  NAND U1869 ( .A(n819), .B(n774), .Z(n818) );
  NAND U1870 ( .A(rst), .B(Y0[15]), .Z(n817) );
  NAND U1871 ( .A(n820), .B(n821), .Z(n360) );
  NAND U1872 ( .A(n822), .B(n774), .Z(n821) );
  NAND U1873 ( .A(rst), .B(Y0[16]), .Z(n820) );
  NAND U1874 ( .A(n823), .B(n824), .Z(n359) );
  NAND U1875 ( .A(n825), .B(n774), .Z(n824) );
  NAND U1876 ( .A(rst), .B(Y0[17]), .Z(n823) );
  NAND U1877 ( .A(n826), .B(n827), .Z(n358) );
  NAND U1878 ( .A(n828), .B(n774), .Z(n827) );
  NAND U1879 ( .A(rst), .B(Y0[18]), .Z(n826) );
  NAND U1880 ( .A(n829), .B(n830), .Z(n357) );
  NAND U1881 ( .A(n831), .B(n774), .Z(n830) );
  NAND U1882 ( .A(rst), .B(Y0[19]), .Z(n829) );
  NAND U1883 ( .A(n832), .B(n833), .Z(n356) );
  NAND U1884 ( .A(n834), .B(n774), .Z(n833) );
  NAND U1885 ( .A(rst), .B(Y0[20]), .Z(n832) );
  NAND U1886 ( .A(n835), .B(n836), .Z(n355) );
  NAND U1887 ( .A(n837), .B(n774), .Z(n836) );
  NAND U1888 ( .A(rst), .B(Y0[21]), .Z(n835) );
  NAND U1889 ( .A(n838), .B(n839), .Z(n354) );
  NAND U1890 ( .A(n840), .B(n774), .Z(n839) );
  NAND U1891 ( .A(rst), .B(Y0[22]), .Z(n838) );
  NAND U1892 ( .A(n841), .B(n842), .Z(n353) );
  NAND U1893 ( .A(n843), .B(n774), .Z(n842) );
  NAND U1894 ( .A(rst), .B(Y0[23]), .Z(n841) );
  NAND U1895 ( .A(n844), .B(n845), .Z(n352) );
  NAND U1896 ( .A(n846), .B(n774), .Z(n845) );
  NAND U1897 ( .A(rst), .B(Y0[24]), .Z(n844) );
  NAND U1898 ( .A(n847), .B(n848), .Z(n351) );
  NAND U1899 ( .A(n849), .B(n774), .Z(n848) );
  NAND U1900 ( .A(rst), .B(Y0[25]), .Z(n847) );
  NAND U1901 ( .A(n850), .B(n851), .Z(n350) );
  NAND U1902 ( .A(n852), .B(n774), .Z(n851) );
  NAND U1903 ( .A(rst), .B(Y0[26]), .Z(n850) );
  NAND U1904 ( .A(n853), .B(n854), .Z(n349) );
  NAND U1905 ( .A(n855), .B(n774), .Z(n854) );
  NAND U1906 ( .A(rst), .B(Y0[27]), .Z(n853) );
  NAND U1907 ( .A(n856), .B(n857), .Z(n348) );
  NAND U1908 ( .A(n858), .B(n774), .Z(n857) );
  NAND U1909 ( .A(rst), .B(Y0[28]), .Z(n856) );
  NAND U1910 ( .A(n859), .B(n860), .Z(n347) );
  NAND U1911 ( .A(n861), .B(n774), .Z(n860) );
  NAND U1912 ( .A(rst), .B(Y0[29]), .Z(n859) );
  NAND U1913 ( .A(n862), .B(n863), .Z(n346) );
  NAND U1914 ( .A(n864), .B(n774), .Z(n863) );
  NAND U1915 ( .A(rst), .B(Y0[30]), .Z(n862) );
  NAND U1916 ( .A(n865), .B(n866), .Z(n345) );
  NAND U1917 ( .A(n867), .B(n774), .Z(n866) );
  NOR U1918 ( .A(rst), .B(n868), .Z(n774) );
  NAND U1919 ( .A(Y0[31]), .B(rst), .Z(n865) );
  MUX U1920 ( .IN0(Y[31]), .IN1(n867), .SEL(n869), .F(n344) );
  XNOR U1921 ( .A(Y0[31]), .B(n871), .Z(n870) );
  AND U1922 ( .A(n874), .B(n875), .Z(n873) );
  XNOR U1923 ( .A(Y0[31]), .B(n876), .Z(n875) );
  MUX U1924 ( .IN0(Y[30]), .IN1(n864), .SEL(n869), .F(n343) );
  XOR U1925 ( .A(n874), .B(Y0[31]), .Z(n864) );
  XOR U1926 ( .A(n876), .B(n871), .Z(n874) );
  XOR U1927 ( .A(n877), .B(n878), .Z(n871) );
  XOR U1928 ( .A(n879), .B(n880), .Z(n878) );
  AND U1929 ( .A(n881), .B(n882), .Z(n880) );
  XOR U1930 ( .A(n889), .B(n887), .Z(n877) );
  XOR U1931 ( .A(n890), .B(n891), .Z(n889) );
  XOR U1932 ( .A(n892), .B(n893), .Z(n891) );
  XOR U1933 ( .A(n897), .B(n898), .Z(n892) );
  ANDN U1934 ( .A(n899), .B(n900), .Z(n898) );
  XOR U1935 ( .A(n904), .B(n905), .Z(n890) );
  XOR U1936 ( .A(n894), .B(n896), .Z(n905) );
  XOR U1937 ( .A(n903), .B(n900), .Z(n904) );
  IV U1938 ( .A(n872), .Z(n876) );
  MUX U1939 ( .IN0(Y[29]), .IN1(n861), .SEL(n869), .F(n342) );
  XOR U1940 ( .A(n907), .B(Y0[30]), .Z(n861) );
  XNOR U1941 ( .A(n908), .B(n909), .Z(n907) );
  AND U1942 ( .A(n881), .B(n911), .Z(n910) );
  XNOR U1943 ( .A(n885), .B(n909), .Z(n911) );
  XOR U1944 ( .A(n883), .B(n909), .Z(n885) );
  XNOR U1945 ( .A(n888), .B(n886), .Z(n909) );
  IV U1946 ( .A(n887), .Z(n886) );
  XNOR U1947 ( .A(n894), .B(n895), .Z(n888) );
  XNOR U1948 ( .A(n896), .B(n899), .Z(n895) );
  XNOR U1949 ( .A(n900), .B(n915), .Z(n899) );
  XOR U1950 ( .A(n901), .B(n902), .Z(n915) );
  NAND U1951 ( .A(n916), .B(n917), .Z(n902) );
  IV U1952 ( .A(n903), .Z(n901) );
  IV U1953 ( .A(n884), .Z(n883) );
  MUX U1954 ( .IN0(Y[28]), .IN1(n858), .SEL(n869), .F(n341) );
  XOR U1955 ( .A(n930), .B(Y0[29]), .Z(n858) );
  XNOR U1956 ( .A(n931), .B(n932), .Z(n930) );
  AND U1957 ( .A(n881), .B(n934), .Z(n933) );
  XNOR U1958 ( .A(n928), .B(n932), .Z(n934) );
  XNOR U1959 ( .A(n914), .B(n913), .Z(n932) );
  IV U1960 ( .A(n912), .Z(n913) );
  XOR U1961 ( .A(n926), .B(n925), .Z(n914) );
  XOR U1962 ( .A(n924), .B(n938), .Z(n925) );
  XNOR U1963 ( .A(n923), .B(n922), .Z(n938) );
  XNOR U1964 ( .A(n939), .B(n940), .Z(n922) );
  IV U1965 ( .A(n921), .Z(n940) );
  XNOR U1966 ( .A(n919), .B(n920), .Z(n923) );
  NAND U1967 ( .A(n946), .B(n917), .Z(n920) );
  XNOR U1968 ( .A(n918), .B(n947), .Z(n919) );
  ANDN U1969 ( .A(n948), .B(n949), .Z(n947) );
  MUX U1970 ( .IN0(Y[27]), .IN1(n855), .SEL(n869), .F(n340) );
  XOR U1971 ( .A(n959), .B(Y0[28]), .Z(n855) );
  XNOR U1972 ( .A(n960), .B(n961), .Z(n959) );
  AND U1973 ( .A(n881), .B(n963), .Z(n962) );
  XNOR U1974 ( .A(n957), .B(n961), .Z(n963) );
  XNOR U1975 ( .A(n937), .B(n936), .Z(n961) );
  IV U1976 ( .A(n935), .Z(n936) );
  XOR U1977 ( .A(n955), .B(n954), .Z(n937) );
  XOR U1978 ( .A(n953), .B(n967), .Z(n954) );
  XNOR U1979 ( .A(n943), .B(n942), .Z(n967) );
  XOR U1980 ( .A(n972), .B(n944), .Z(n968) );
  AND U1981 ( .A(n973), .B(n916), .Z(n944) );
  IV U1982 ( .A(n941), .Z(n972) );
  XNOR U1983 ( .A(n951), .B(n952), .Z(n943) );
  NAND U1984 ( .A(n977), .B(n917), .Z(n952) );
  XNOR U1985 ( .A(n950), .B(n978), .Z(n951) );
  ANDN U1986 ( .A(n948), .B(n979), .Z(n978) );
  MUX U1987 ( .IN0(Y[26]), .IN1(n852), .SEL(n869), .F(n339) );
  XOR U1988 ( .A(n990), .B(Y0[27]), .Z(n852) );
  XNOR U1989 ( .A(n991), .B(n992), .Z(n990) );
  AND U1990 ( .A(n881), .B(n994), .Z(n993) );
  XNOR U1991 ( .A(n988), .B(n992), .Z(n994) );
  XNOR U1992 ( .A(n966), .B(n965), .Z(n992) );
  IV U1993 ( .A(n964), .Z(n965) );
  XNOR U1994 ( .A(n986), .B(n998), .Z(n966) );
  XOR U1995 ( .A(n985), .B(n984), .Z(n998) );
  XOR U1996 ( .A(n999), .B(n1000), .Z(n984) );
  XOR U1997 ( .A(n1001), .B(n1002), .Z(n1000) );
  XOR U1998 ( .A(n1003), .B(n1004), .Z(n1002) );
  XNOR U1999 ( .A(n976), .B(n975), .Z(n985) );
  XOR U2000 ( .A(n1012), .B(n970), .Z(n975) );
  XNOR U2001 ( .A(n969), .B(n1013), .Z(n970) );
  ANDN U2002 ( .A(n1014), .B(n949), .Z(n1013) );
  AND U2003 ( .A(n946), .B(n973), .Z(n971) );
  XNOR U2004 ( .A(n981), .B(n982), .Z(n976) );
  NAND U2005 ( .A(n1021), .B(n917), .Z(n982) );
  XNOR U2006 ( .A(n980), .B(n1022), .Z(n981) );
  ANDN U2007 ( .A(n948), .B(n1023), .Z(n1022) );
  MUX U2008 ( .IN0(Y[25]), .IN1(n849), .SEL(n869), .F(n338) );
  XOR U2009 ( .A(n1031), .B(Y0[26]), .Z(n849) );
  XNOR U2010 ( .A(n1032), .B(n1033), .Z(n1031) );
  AND U2011 ( .A(n881), .B(n1035), .Z(n1034) );
  XNOR U2012 ( .A(n1029), .B(n1033), .Z(n1035) );
  XNOR U2013 ( .A(n997), .B(n996), .Z(n1033) );
  IV U2014 ( .A(n995), .Z(n996) );
  XOR U2015 ( .A(n1027), .B(n1039), .Z(n997) );
  XNOR U2016 ( .A(n1011), .B(n1010), .Z(n1039) );
  XOR U2017 ( .A(n1040), .B(n1005), .Z(n1010) );
  XOR U2018 ( .A(n1006), .B(n1007), .Z(n1005) );
  NANDN U2019 ( .B(n1041), .A(n916), .Z(n1007) );
  IV U2020 ( .A(n1008), .Z(n1006) );
  XOR U2021 ( .A(n1001), .B(n1009), .Z(n1040) );
  XNOR U2022 ( .A(n1020), .B(n1019), .Z(n1011) );
  XOR U2023 ( .A(n1051), .B(n1016), .Z(n1019) );
  XNOR U2024 ( .A(n1015), .B(n1052), .Z(n1016) );
  ANDN U2025 ( .A(n1014), .B(n979), .Z(n1052) );
  XOR U2026 ( .A(n1053), .B(n1054), .Z(n1015) );
  AND U2027 ( .A(n1055), .B(n1056), .Z(n1054) );
  XNOR U2028 ( .A(n1057), .B(n1053), .Z(n1056) );
  AND U2029 ( .A(n977), .B(n973), .Z(n1017) );
  XNOR U2030 ( .A(n1025), .B(n1026), .Z(n1020) );
  NAND U2031 ( .A(n1061), .B(n917), .Z(n1026) );
  XNOR U2032 ( .A(n1024), .B(n1062), .Z(n1025) );
  ANDN U2033 ( .A(n948), .B(n1063), .Z(n1062) );
  MUX U2034 ( .IN0(Y[24]), .IN1(n846), .SEL(n869), .F(n337) );
  XOR U2035 ( .A(n1071), .B(Y0[25]), .Z(n846) );
  XNOR U2036 ( .A(n1072), .B(n1073), .Z(n1071) );
  AND U2037 ( .A(n881), .B(n1075), .Z(n1074) );
  XNOR U2038 ( .A(n1069), .B(n1073), .Z(n1075) );
  XNOR U2039 ( .A(n1038), .B(n1037), .Z(n1073) );
  IV U2040 ( .A(n1036), .Z(n1037) );
  XOR U2041 ( .A(n1067), .B(n1079), .Z(n1038) );
  XNOR U2042 ( .A(n1047), .B(n1046), .Z(n1079) );
  XOR U2043 ( .A(n1080), .B(n1050), .Z(n1046) );
  XNOR U2044 ( .A(n1043), .B(n1044), .Z(n1050) );
  NANDN U2045 ( .B(n1041), .A(n946), .Z(n1044) );
  XNOR U2046 ( .A(n1042), .B(n1081), .Z(n1043) );
  ANDN U2047 ( .A(n1082), .B(n949), .Z(n1081) );
  XNOR U2048 ( .A(n1049), .B(n1045), .Z(n1080) );
  XNOR U2049 ( .A(n1089), .B(n1090), .Z(n1049) );
  IV U2050 ( .A(n1048), .Z(n1090) );
  XNOR U2051 ( .A(n1060), .B(n1059), .Z(n1047) );
  XOR U2052 ( .A(n1097), .B(n1055), .Z(n1059) );
  XNOR U2053 ( .A(n1053), .B(n1098), .Z(n1055) );
  ANDN U2054 ( .A(n1014), .B(n1023), .Z(n1098) );
  AND U2055 ( .A(n1021), .B(n973), .Z(n1057) );
  XNOR U2056 ( .A(n1065), .B(n1066), .Z(n1060) );
  NAND U2057 ( .A(n1105), .B(n917), .Z(n1066) );
  XNOR U2058 ( .A(n1064), .B(n1106), .Z(n1065) );
  ANDN U2059 ( .A(n948), .B(n1107), .Z(n1106) );
  MUX U2060 ( .IN0(Y[23]), .IN1(n843), .SEL(n869), .F(n336) );
  XOR U2061 ( .A(n1115), .B(Y0[24]), .Z(n843) );
  XNOR U2062 ( .A(n1116), .B(n1117), .Z(n1115) );
  AND U2063 ( .A(n881), .B(n1119), .Z(n1118) );
  XNOR U2064 ( .A(n1113), .B(n1117), .Z(n1119) );
  XNOR U2065 ( .A(n1078), .B(n1077), .Z(n1117) );
  IV U2066 ( .A(n1076), .Z(n1077) );
  XOR U2067 ( .A(n1111), .B(n1122), .Z(n1078) );
  XNOR U2068 ( .A(n1088), .B(n1087), .Z(n1122) );
  XOR U2069 ( .A(n1123), .B(n1093), .Z(n1087) );
  XNOR U2070 ( .A(n1084), .B(n1085), .Z(n1093) );
  NANDN U2071 ( .B(n1041), .A(n977), .Z(n1085) );
  XNOR U2072 ( .A(n1083), .B(n1124), .Z(n1084) );
  ANDN U2073 ( .A(n1082), .B(n979), .Z(n1124) );
  XNOR U2074 ( .A(n1092), .B(n1086), .Z(n1123) );
  XNOR U2075 ( .A(n1131), .B(n1094), .Z(n1092) );
  IV U2076 ( .A(n1096), .Z(n1094) );
  AND U2077 ( .A(n1135), .B(n916), .Z(n1095) );
  XNOR U2078 ( .A(n1104), .B(n1103), .Z(n1088) );
  XOR U2079 ( .A(n1139), .B(n1100), .Z(n1103) );
  XNOR U2080 ( .A(n1099), .B(n1140), .Z(n1100) );
  ANDN U2081 ( .A(n1014), .B(n1063), .Z(n1140) );
  AND U2082 ( .A(n1061), .B(n973), .Z(n1101) );
  XNOR U2083 ( .A(n1109), .B(n1110), .Z(n1104) );
  NAND U2084 ( .A(n1147), .B(n917), .Z(n1110) );
  XNOR U2085 ( .A(n1108), .B(n1148), .Z(n1109) );
  ANDN U2086 ( .A(n948), .B(n1149), .Z(n1148) );
  MUX U2087 ( .IN0(Y[22]), .IN1(n840), .SEL(n869), .F(n335) );
  XOR U2088 ( .A(n1159), .B(Y0[23]), .Z(n840) );
  XNOR U2089 ( .A(n1160), .B(n1121), .Z(n1159) );
  AND U2090 ( .A(n881), .B(n1162), .Z(n1161) );
  XNOR U2091 ( .A(n1157), .B(n1121), .Z(n1162) );
  XOR U2092 ( .A(n1120), .B(n1163), .Z(n1121) );
  XNOR U2093 ( .A(n1155), .B(n1154), .Z(n1163) );
  XOR U2094 ( .A(n1164), .B(n1165), .Z(n1154) );
  XOR U2095 ( .A(n1166), .B(n1167), .Z(n1165) );
  XOR U2096 ( .A(n1170), .B(n1171), .Z(n1166) );
  ANDN U2097 ( .A(n1169), .B(n1172), .Z(n1171) );
  XNOR U2098 ( .A(n1175), .B(n1153), .Z(n1164) );
  XOR U2099 ( .A(n1174), .B(n1172), .Z(n1175) );
  XNOR U2100 ( .A(n1130), .B(n1129), .Z(n1155) );
  XOR U2101 ( .A(n1179), .B(n1138), .Z(n1129) );
  XNOR U2102 ( .A(n1126), .B(n1127), .Z(n1138) );
  NANDN U2103 ( .B(n1041), .A(n1021), .Z(n1127) );
  XNOR U2104 ( .A(n1125), .B(n1180), .Z(n1126) );
  ANDN U2105 ( .A(n1082), .B(n1023), .Z(n1180) );
  XNOR U2106 ( .A(n1137), .B(n1128), .Z(n1179) );
  XOR U2107 ( .A(n1187), .B(n1133), .Z(n1137) );
  XNOR U2108 ( .A(n1132), .B(n1188), .Z(n1133) );
  ANDN U2109 ( .A(n1189), .B(n949), .Z(n1188) );
  XOR U2110 ( .A(n1190), .B(n1191), .Z(n1132) );
  AND U2111 ( .A(n1192), .B(n1193), .Z(n1191) );
  XNOR U2112 ( .A(n1194), .B(n1190), .Z(n1193) );
  AND U2113 ( .A(n946), .B(n1135), .Z(n1134) );
  XNOR U2114 ( .A(n1146), .B(n1145), .Z(n1130) );
  XOR U2115 ( .A(n1198), .B(n1142), .Z(n1145) );
  XNOR U2116 ( .A(n1141), .B(n1199), .Z(n1142) );
  ANDN U2117 ( .A(n1014), .B(n1107), .Z(n1199) );
  AND U2118 ( .A(n1105), .B(n973), .Z(n1143) );
  XNOR U2119 ( .A(n1151), .B(n1152), .Z(n1146) );
  NAND U2120 ( .A(n1206), .B(n917), .Z(n1152) );
  XNOR U2121 ( .A(n1150), .B(n1207), .Z(n1151) );
  ANDN U2122 ( .A(n948), .B(n1208), .Z(n1207) );
  MUX U2123 ( .IN0(Y[21]), .IN1(n837), .SEL(n869), .F(n334) );
  XOR U2124 ( .A(n1218), .B(Y0[22]), .Z(n837) );
  XNOR U2125 ( .A(n1219), .B(n1220), .Z(n1218) );
  AND U2126 ( .A(n881), .B(n1222), .Z(n1221) );
  XNOR U2127 ( .A(n1216), .B(n1220), .Z(n1222) );
  XNOR U2128 ( .A(n1214), .B(n1213), .Z(n1220) );
  IV U2129 ( .A(n1212), .Z(n1213) );
  XNOR U2130 ( .A(n1178), .B(n1177), .Z(n1214) );
  XOR U2131 ( .A(n1226), .B(n1169), .Z(n1177) );
  XNOR U2132 ( .A(n1172), .B(n1227), .Z(n1169) );
  NANDN U2133 ( .B(n1228), .A(n916), .Z(n1173) );
  XOR U2134 ( .A(n1168), .B(n1176), .Z(n1226) );
  XNOR U2135 ( .A(n1186), .B(n1185), .Z(n1178) );
  XOR U2136 ( .A(n1240), .B(n1197), .Z(n1185) );
  XNOR U2137 ( .A(n1182), .B(n1183), .Z(n1197) );
  NANDN U2138 ( .B(n1041), .A(n1061), .Z(n1183) );
  XNOR U2139 ( .A(n1181), .B(n1241), .Z(n1182) );
  ANDN U2140 ( .A(n1082), .B(n1063), .Z(n1241) );
  XOR U2141 ( .A(n1242), .B(n1243), .Z(n1181) );
  AND U2142 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U2143 ( .A(n1246), .B(n1242), .Z(n1245) );
  XNOR U2144 ( .A(n1196), .B(n1184), .Z(n1240) );
  XOR U2145 ( .A(n1250), .B(n1192), .Z(n1196) );
  XNOR U2146 ( .A(n1190), .B(n1251), .Z(n1192) );
  ANDN U2147 ( .A(n1189), .B(n979), .Z(n1251) );
  XOR U2148 ( .A(n1252), .B(n1253), .Z(n1190) );
  AND U2149 ( .A(n1254), .B(n1255), .Z(n1253) );
  XNOR U2150 ( .A(n1256), .B(n1252), .Z(n1255) );
  AND U2151 ( .A(n977), .B(n1135), .Z(n1194) );
  XNOR U2152 ( .A(n1205), .B(n1204), .Z(n1186) );
  XOR U2153 ( .A(n1260), .B(n1201), .Z(n1204) );
  XNOR U2154 ( .A(n1200), .B(n1261), .Z(n1201) );
  ANDN U2155 ( .A(n1014), .B(n1149), .Z(n1261) );
  XOR U2156 ( .A(n1262), .B(n1263), .Z(n1200) );
  AND U2157 ( .A(n1264), .B(n1265), .Z(n1263) );
  XNOR U2158 ( .A(n1266), .B(n1262), .Z(n1265) );
  AND U2159 ( .A(n1147), .B(n973), .Z(n1202) );
  XNOR U2160 ( .A(n1210), .B(n1211), .Z(n1205) );
  NAND U2161 ( .A(n1270), .B(n917), .Z(n1211) );
  XNOR U2162 ( .A(n1209), .B(n1271), .Z(n1210) );
  ANDN U2163 ( .A(n948), .B(n1272), .Z(n1271) );
  XOR U2164 ( .A(n1273), .B(n1274), .Z(n1209) );
  AND U2165 ( .A(n1275), .B(n1276), .Z(n1274) );
  XOR U2166 ( .A(n1277), .B(n1273), .Z(n1276) );
  MUX U2167 ( .IN0(Y[20]), .IN1(n834), .SEL(n869), .F(n333) );
  XOR U2168 ( .A(n1281), .B(Y0[21]), .Z(n834) );
  XNOR U2169 ( .A(n1282), .B(n1283), .Z(n1281) );
  AND U2170 ( .A(n881), .B(n1285), .Z(n1284) );
  XNOR U2171 ( .A(n1279), .B(n1283), .Z(n1285) );
  XNOR U2172 ( .A(n1225), .B(n1224), .Z(n1283) );
  IV U2173 ( .A(n1223), .Z(n1224) );
  XNOR U2174 ( .A(n1237), .B(n1236), .Z(n1225) );
  XOR U2175 ( .A(n1289), .B(n1239), .Z(n1236) );
  XNOR U2176 ( .A(n1234), .B(n1233), .Z(n1239) );
  XNOR U2177 ( .A(n1290), .B(n1291), .Z(n1233) );
  IV U2178 ( .A(n1232), .Z(n1291) );
  XNOR U2179 ( .A(n1230), .B(n1231), .Z(n1234) );
  NANDN U2180 ( .B(n1228), .A(n946), .Z(n1231) );
  XNOR U2181 ( .A(n1229), .B(n1297), .Z(n1230) );
  ANDN U2182 ( .A(n1298), .B(n949), .Z(n1297) );
  XNOR U2183 ( .A(n1249), .B(n1248), .Z(n1237) );
  XOR U2184 ( .A(n1308), .B(n1259), .Z(n1248) );
  XNOR U2185 ( .A(n1244), .B(n1246), .Z(n1259) );
  NANDN U2186 ( .B(n1041), .A(n1105), .Z(n1246) );
  XNOR U2187 ( .A(n1242), .B(n1309), .Z(n1244) );
  ANDN U2188 ( .A(n1082), .B(n1107), .Z(n1309) );
  XOR U2189 ( .A(n1310), .B(n1311), .Z(n1242) );
  AND U2190 ( .A(n1312), .B(n1313), .Z(n1311) );
  XOR U2191 ( .A(n1314), .B(n1310), .Z(n1313) );
  XNOR U2192 ( .A(n1258), .B(n1247), .Z(n1308) );
  XOR U2193 ( .A(n1318), .B(n1254), .Z(n1258) );
  XNOR U2194 ( .A(n1252), .B(n1319), .Z(n1254) );
  ANDN U2195 ( .A(n1189), .B(n1023), .Z(n1319) );
  XOR U2196 ( .A(n1320), .B(n1321), .Z(n1252) );
  AND U2197 ( .A(n1322), .B(n1323), .Z(n1321) );
  XNOR U2198 ( .A(n1324), .B(n1320), .Z(n1323) );
  AND U2199 ( .A(n1021), .B(n1135), .Z(n1256) );
  XNOR U2200 ( .A(n1269), .B(n1268), .Z(n1249) );
  XOR U2201 ( .A(n1328), .B(n1264), .Z(n1268) );
  XNOR U2202 ( .A(n1262), .B(n1329), .Z(n1264) );
  ANDN U2203 ( .A(n1014), .B(n1208), .Z(n1329) );
  XOR U2204 ( .A(n1330), .B(n1331), .Z(n1262) );
  AND U2205 ( .A(n1332), .B(n1333), .Z(n1331) );
  XNOR U2206 ( .A(n1334), .B(n1330), .Z(n1333) );
  AND U2207 ( .A(n1206), .B(n973), .Z(n1266) );
  XNOR U2208 ( .A(n1275), .B(n1277), .Z(n1269) );
  NAND U2209 ( .A(n1338), .B(n917), .Z(n1277) );
  XNOR U2210 ( .A(n1273), .B(n1339), .Z(n1275) );
  ANDN U2211 ( .A(n948), .B(n1340), .Z(n1339) );
  XOR U2212 ( .A(n1341), .B(n1342), .Z(n1273) );
  AND U2213 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U2214 ( .A(n1345), .B(n1341), .Z(n1344) );
  MUX U2215 ( .IN0(Y[19]), .IN1(n831), .SEL(n869), .F(n332) );
  XOR U2216 ( .A(n1349), .B(Y0[20]), .Z(n831) );
  XNOR U2217 ( .A(n1350), .B(n1351), .Z(n1349) );
  AND U2218 ( .A(n881), .B(n1353), .Z(n1352) );
  XNOR U2219 ( .A(n1347), .B(n1351), .Z(n1353) );
  XNOR U2220 ( .A(n1288), .B(n1287), .Z(n1351) );
  IV U2221 ( .A(n1286), .Z(n1287) );
  XNOR U2222 ( .A(n1304), .B(n1303), .Z(n1288) );
  XOR U2223 ( .A(n1357), .B(n1307), .Z(n1303) );
  XNOR U2224 ( .A(n1294), .B(n1293), .Z(n1307) );
  XOR U2225 ( .A(n1362), .B(n1295), .Z(n1358) );
  AND U2226 ( .A(n1363), .B(n916), .Z(n1295) );
  IV U2227 ( .A(n1292), .Z(n1362) );
  XNOR U2228 ( .A(n1300), .B(n1301), .Z(n1294) );
  NANDN U2229 ( .B(n1228), .A(n977), .Z(n1301) );
  XNOR U2230 ( .A(n1299), .B(n1367), .Z(n1300) );
  ANDN U2231 ( .A(n1298), .B(n979), .Z(n1367) );
  XNOR U2232 ( .A(n1306), .B(n1302), .Z(n1357) );
  IV U2233 ( .A(n1305), .Z(n1306) );
  XNOR U2234 ( .A(n1317), .B(n1316), .Z(n1304) );
  XOR U2235 ( .A(n1377), .B(n1327), .Z(n1316) );
  XNOR U2236 ( .A(n1312), .B(n1314), .Z(n1327) );
  NANDN U2237 ( .B(n1041), .A(n1147), .Z(n1314) );
  XNOR U2238 ( .A(n1310), .B(n1378), .Z(n1312) );
  ANDN U2239 ( .A(n1082), .B(n1149), .Z(n1378) );
  XOR U2240 ( .A(n1379), .B(n1380), .Z(n1310) );
  AND U2241 ( .A(n1381), .B(n1382), .Z(n1380) );
  XOR U2242 ( .A(n1383), .B(n1379), .Z(n1382) );
  XNOR U2243 ( .A(n1326), .B(n1315), .Z(n1377) );
  XOR U2244 ( .A(n1387), .B(n1322), .Z(n1326) );
  XNOR U2245 ( .A(n1320), .B(n1388), .Z(n1322) );
  ANDN U2246 ( .A(n1189), .B(n1063), .Z(n1388) );
  XOR U2247 ( .A(n1389), .B(n1390), .Z(n1320) );
  AND U2248 ( .A(n1391), .B(n1392), .Z(n1390) );
  XNOR U2249 ( .A(n1393), .B(n1389), .Z(n1392) );
  AND U2250 ( .A(n1061), .B(n1135), .Z(n1324) );
  XNOR U2251 ( .A(n1337), .B(n1336), .Z(n1317) );
  XOR U2252 ( .A(n1397), .B(n1332), .Z(n1336) );
  XNOR U2253 ( .A(n1330), .B(n1398), .Z(n1332) );
  ANDN U2254 ( .A(n1014), .B(n1272), .Z(n1398) );
  AND U2255 ( .A(n1270), .B(n973), .Z(n1334) );
  XNOR U2256 ( .A(n1343), .B(n1345), .Z(n1337) );
  NAND U2257 ( .A(n1405), .B(n917), .Z(n1345) );
  XNOR U2258 ( .A(n1341), .B(n1406), .Z(n1343) );
  ANDN U2259 ( .A(n948), .B(n1407), .Z(n1406) );
  XOR U2260 ( .A(n1408), .B(n1409), .Z(n1341) );
  AND U2261 ( .A(n1410), .B(n1411), .Z(n1409) );
  XOR U2262 ( .A(n1412), .B(n1408), .Z(n1411) );
  MUX U2263 ( .IN0(Y[18]), .IN1(n828), .SEL(n869), .F(n331) );
  XOR U2264 ( .A(n1416), .B(Y0[19]), .Z(n828) );
  XNOR U2265 ( .A(n1417), .B(n1418), .Z(n1416) );
  AND U2266 ( .A(n881), .B(n1420), .Z(n1419) );
  XOR U2267 ( .A(n1414), .B(n1418), .Z(n1420) );
  XOR U2268 ( .A(n1413), .B(n1418), .Z(n1414) );
  XNOR U2269 ( .A(n1356), .B(n1355), .Z(n1418) );
  IV U2270 ( .A(n1354), .Z(n1355) );
  XNOR U2271 ( .A(n1373), .B(n1372), .Z(n1356) );
  XOR U2272 ( .A(n1423), .B(n1376), .Z(n1372) );
  XNOR U2273 ( .A(n1366), .B(n1365), .Z(n1376) );
  XOR U2274 ( .A(n1424), .B(n1360), .Z(n1365) );
  XNOR U2275 ( .A(n1359), .B(n1425), .Z(n1360) );
  ANDN U2276 ( .A(n1426), .B(n949), .Z(n1425) );
  XOR U2277 ( .A(n1427), .B(n1428), .Z(n1359) );
  AND U2278 ( .A(n1429), .B(n1430), .Z(n1428) );
  XNOR U2279 ( .A(n1431), .B(n1427), .Z(n1430) );
  AND U2280 ( .A(n946), .B(n1363), .Z(n1361) );
  XNOR U2281 ( .A(n1369), .B(n1370), .Z(n1366) );
  NANDN U2282 ( .B(n1228), .A(n1021), .Z(n1370) );
  XNOR U2283 ( .A(n1368), .B(n1435), .Z(n1369) );
  ANDN U2284 ( .A(n1298), .B(n1023), .Z(n1435) );
  XNOR U2285 ( .A(n1375), .B(n1371), .Z(n1423) );
  XNOR U2286 ( .A(n1442), .B(n1443), .Z(n1375) );
  IV U2287 ( .A(n1374), .Z(n1443) );
  XNOR U2288 ( .A(n1386), .B(n1385), .Z(n1373) );
  XOR U2289 ( .A(n1449), .B(n1396), .Z(n1385) );
  XNOR U2290 ( .A(n1381), .B(n1383), .Z(n1396) );
  NANDN U2291 ( .B(n1041), .A(n1206), .Z(n1383) );
  XNOR U2292 ( .A(n1379), .B(n1450), .Z(n1381) );
  ANDN U2293 ( .A(n1082), .B(n1208), .Z(n1450) );
  XOR U2294 ( .A(n1451), .B(n1452), .Z(n1379) );
  AND U2295 ( .A(n1453), .B(n1454), .Z(n1452) );
  XOR U2296 ( .A(n1455), .B(n1451), .Z(n1454) );
  XNOR U2297 ( .A(n1395), .B(n1384), .Z(n1449) );
  XOR U2298 ( .A(n1459), .B(n1391), .Z(n1395) );
  XNOR U2299 ( .A(n1389), .B(n1460), .Z(n1391) );
  ANDN U2300 ( .A(n1189), .B(n1107), .Z(n1460) );
  XOR U2301 ( .A(n1461), .B(n1462), .Z(n1389) );
  AND U2302 ( .A(n1463), .B(n1464), .Z(n1462) );
  XNOR U2303 ( .A(n1465), .B(n1461), .Z(n1464) );
  AND U2304 ( .A(n1105), .B(n1135), .Z(n1393) );
  XNOR U2305 ( .A(n1404), .B(n1403), .Z(n1386) );
  XOR U2306 ( .A(n1469), .B(n1400), .Z(n1403) );
  XNOR U2307 ( .A(n1399), .B(n1470), .Z(n1400) );
  ANDN U2308 ( .A(n1014), .B(n1340), .Z(n1470) );
  XOR U2309 ( .A(n1471), .B(n1472), .Z(n1399) );
  AND U2310 ( .A(n1473), .B(n1474), .Z(n1472) );
  XNOR U2311 ( .A(n1475), .B(n1471), .Z(n1474) );
  AND U2312 ( .A(n1338), .B(n973), .Z(n1401) );
  XNOR U2313 ( .A(n1410), .B(n1412), .Z(n1404) );
  NAND U2314 ( .A(n1479), .B(n917), .Z(n1412) );
  XNOR U2315 ( .A(n1408), .B(n1480), .Z(n1410) );
  ANDN U2316 ( .A(n948), .B(n1481), .Z(n1480) );
  NANDN U2317 ( .B(n1482), .A(n1483), .Z(n1408) );
  NAND U2318 ( .A(n1484), .B(n1485), .Z(n1483) );
  MUX U2319 ( .IN0(Y[17]), .IN1(n825), .SEL(n869), .F(n330) );
  XOR U2320 ( .A(n1490), .B(Y0[18]), .Z(n825) );
  XOR U2321 ( .A(n1491), .B(n1492), .Z(n1490) );
  AND U2322 ( .A(n881), .B(n1494), .Z(n1493) );
  XOR U2323 ( .A(n1488), .B(n1492), .Z(n1494) );
  XOR U2324 ( .A(n1487), .B(n1492), .Z(n1488) );
  XOR U2325 ( .A(n1422), .B(n1421), .Z(n1492) );
  XNOR U2326 ( .A(n1497), .B(n1446), .Z(n1440) );
  XNOR U2327 ( .A(n1434), .B(n1433), .Z(n1446) );
  XOR U2328 ( .A(n1498), .B(n1429), .Z(n1433) );
  XNOR U2329 ( .A(n1427), .B(n1499), .Z(n1429) );
  ANDN U2330 ( .A(n1426), .B(n979), .Z(n1499) );
  XOR U2331 ( .A(n1500), .B(n1501), .Z(n1427) );
  AND U2332 ( .A(n1502), .B(n1503), .Z(n1501) );
  XNOR U2333 ( .A(n1504), .B(n1500), .Z(n1503) );
  AND U2334 ( .A(n977), .B(n1363), .Z(n1431) );
  XNOR U2335 ( .A(n1437), .B(n1438), .Z(n1434) );
  NANDN U2336 ( .B(n1228), .A(n1061), .Z(n1438) );
  XNOR U2337 ( .A(n1436), .B(n1508), .Z(n1437) );
  ANDN U2338 ( .A(n1298), .B(n1063), .Z(n1508) );
  XOR U2339 ( .A(n1509), .B(n1510), .Z(n1436) );
  AND U2340 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U2341 ( .A(n1513), .B(n1509), .Z(n1512) );
  XNOR U2342 ( .A(n1445), .B(n1439), .Z(n1497) );
  XOR U2343 ( .A(n1517), .B(n1447), .Z(n1445) );
  NAND U2344 ( .A(n1521), .B(n1522), .Z(n1448) );
  NANDN U2345 ( .B(n1523), .A(n916), .Z(n1522) );
  NANDN U2346 ( .B(n1524), .A(n1525), .Z(n1521) );
  XNOR U2347 ( .A(n1458), .B(n1457), .Z(n1441) );
  XOR U2348 ( .A(n1529), .B(n1468), .Z(n1457) );
  XNOR U2349 ( .A(n1453), .B(n1455), .Z(n1468) );
  NANDN U2350 ( .B(n1041), .A(n1270), .Z(n1455) );
  XNOR U2351 ( .A(n1451), .B(n1530), .Z(n1453) );
  ANDN U2352 ( .A(n1082), .B(n1272), .Z(n1530) );
  XOR U2353 ( .A(n1531), .B(n1532), .Z(n1451) );
  AND U2354 ( .A(n1533), .B(n1534), .Z(n1532) );
  XOR U2355 ( .A(n1535), .B(n1531), .Z(n1534) );
  XNOR U2356 ( .A(n1467), .B(n1456), .Z(n1529) );
  XOR U2357 ( .A(n1539), .B(n1463), .Z(n1467) );
  XNOR U2358 ( .A(n1461), .B(n1540), .Z(n1463) );
  ANDN U2359 ( .A(n1189), .B(n1149), .Z(n1540) );
  XOR U2360 ( .A(n1541), .B(n1542), .Z(n1461) );
  AND U2361 ( .A(n1543), .B(n1544), .Z(n1542) );
  XNOR U2362 ( .A(n1545), .B(n1541), .Z(n1544) );
  AND U2363 ( .A(n1147), .B(n1135), .Z(n1465) );
  XOR U2364 ( .A(n1478), .B(n1477), .Z(n1458) );
  XOR U2365 ( .A(n1549), .B(n1473), .Z(n1477) );
  XNOR U2366 ( .A(n1471), .B(n1550), .Z(n1473) );
  ANDN U2367 ( .A(n1014), .B(n1407), .Z(n1550) );
  AND U2368 ( .A(n1405), .B(n973), .Z(n1475) );
  XOR U2369 ( .A(n1485), .B(n1484), .Z(n1478) );
  NAND U2370 ( .A(n1557), .B(n917), .Z(n1484) );
  XNOR U2371 ( .A(n1482), .B(n1558), .Z(n1485) );
  ANDN U2372 ( .A(n948), .B(n1559), .Z(n1558) );
  NANDN U2373 ( .B(n1560), .A(n1561), .Z(n1482) );
  NAND U2374 ( .A(n1562), .B(n1563), .Z(n1561) );
  IV U2375 ( .A(n1486), .Z(n1487) );
  MUX U2376 ( .IN0(Y[16]), .IN1(n822), .SEL(n869), .F(n329) );
  XOR U2377 ( .A(n1568), .B(Y0[17]), .Z(n822) );
  XOR U2378 ( .A(n1569), .B(n1570), .Z(n1568) );
  AND U2379 ( .A(n881), .B(n1572), .Z(n1571) );
  XOR U2380 ( .A(n1566), .B(n1570), .Z(n1572) );
  XOR U2381 ( .A(n1565), .B(n1570), .Z(n1566) );
  XOR U2382 ( .A(n1496), .B(n1495), .Z(n1570) );
  XNOR U2383 ( .A(n1575), .B(n1528), .Z(n1515) );
  XNOR U2384 ( .A(n1507), .B(n1506), .Z(n1528) );
  XOR U2385 ( .A(n1576), .B(n1502), .Z(n1506) );
  XNOR U2386 ( .A(n1500), .B(n1577), .Z(n1502) );
  ANDN U2387 ( .A(n1426), .B(n1023), .Z(n1577) );
  XOR U2388 ( .A(n1578), .B(n1579), .Z(n1500) );
  AND U2389 ( .A(n1580), .B(n1581), .Z(n1579) );
  XNOR U2390 ( .A(n1582), .B(n1578), .Z(n1581) );
  AND U2391 ( .A(n1021), .B(n1363), .Z(n1504) );
  XNOR U2392 ( .A(n1511), .B(n1513), .Z(n1507) );
  NANDN U2393 ( .B(n1228), .A(n1105), .Z(n1513) );
  XNOR U2394 ( .A(n1509), .B(n1586), .Z(n1511) );
  ANDN U2395 ( .A(n1298), .B(n1107), .Z(n1586) );
  XOR U2396 ( .A(n1587), .B(n1588), .Z(n1509) );
  AND U2397 ( .A(n1589), .B(n1590), .Z(n1588) );
  XOR U2398 ( .A(n1591), .B(n1587), .Z(n1590) );
  XOR U2399 ( .A(n1527), .B(n1514), .Z(n1575) );
  XNOR U2400 ( .A(n1595), .B(n1519), .Z(n1527) );
  XNOR U2401 ( .A(n1596), .B(n1525), .Z(n1519) );
  AND U2402 ( .A(n946), .B(n1597), .Z(n1525) );
  NAND U2403 ( .A(n1598), .B(n1524), .Z(n1596) );
  XOR U2404 ( .A(n1599), .B(n1600), .Z(n1524) );
  AND U2405 ( .A(n1601), .B(n1602), .Z(n1600) );
  XOR U2406 ( .A(n1603), .B(n1599), .Z(n1602) );
  NANDN U2407 ( .B(n949), .A(n1604), .Z(n1598) );
  XNOR U2408 ( .A(n1518), .B(n1526), .Z(n1595) );
  IV U2409 ( .A(n1520), .Z(n1518) );
  XNOR U2410 ( .A(n1538), .B(n1537), .Z(n1516) );
  XOR U2411 ( .A(n1610), .B(n1548), .Z(n1537) );
  XNOR U2412 ( .A(n1533), .B(n1535), .Z(n1548) );
  NANDN U2413 ( .B(n1041), .A(n1338), .Z(n1535) );
  XNOR U2414 ( .A(n1531), .B(n1611), .Z(n1533) );
  ANDN U2415 ( .A(n1082), .B(n1340), .Z(n1611) );
  XNOR U2416 ( .A(n1547), .B(n1536), .Z(n1610) );
  XOR U2417 ( .A(n1618), .B(n1543), .Z(n1547) );
  XNOR U2418 ( .A(n1541), .B(n1619), .Z(n1543) );
  ANDN U2419 ( .A(n1189), .B(n1208), .Z(n1619) );
  XOR U2420 ( .A(n1620), .B(n1621), .Z(n1541) );
  AND U2421 ( .A(n1622), .B(n1623), .Z(n1621) );
  XNOR U2422 ( .A(n1624), .B(n1620), .Z(n1623) );
  AND U2423 ( .A(n1206), .B(n1135), .Z(n1545) );
  XOR U2424 ( .A(n1556), .B(n1555), .Z(n1538) );
  XOR U2425 ( .A(n1628), .B(n1552), .Z(n1555) );
  XNOR U2426 ( .A(n1551), .B(n1629), .Z(n1552) );
  ANDN U2427 ( .A(n1014), .B(n1481), .Z(n1629) );
  XOR U2428 ( .A(n1630), .B(n1631), .Z(n1551) );
  AND U2429 ( .A(n1632), .B(n1633), .Z(n1631) );
  XNOR U2430 ( .A(n1634), .B(n1630), .Z(n1633) );
  AND U2431 ( .A(n1479), .B(n973), .Z(n1553) );
  XOR U2432 ( .A(n1563), .B(n1562), .Z(n1556) );
  NAND U2433 ( .A(n1638), .B(n917), .Z(n1562) );
  XNOR U2434 ( .A(n1560), .B(n1639), .Z(n1563) );
  ANDN U2435 ( .A(n948), .B(n1640), .Z(n1639) );
  NAND U2436 ( .A(n1641), .B(n1642), .Z(n1560) );
  NAND U2437 ( .A(n1643), .B(n1644), .Z(n1641) );
  IV U2438 ( .A(n1564), .Z(n1565) );
  MUX U2439 ( .IN0(Y[15]), .IN1(n819), .SEL(n869), .F(n328) );
  XOR U2440 ( .A(n1649), .B(Y0[16]), .Z(n819) );
  XOR U2441 ( .A(n1650), .B(n1651), .Z(n1649) );
  AND U2442 ( .A(n881), .B(n1653), .Z(n1652) );
  XOR U2443 ( .A(n1647), .B(n1651), .Z(n1653) );
  XOR U2444 ( .A(n1646), .B(n1651), .Z(n1647) );
  XOR U2445 ( .A(n1574), .B(n1573), .Z(n1651) );
  XNOR U2446 ( .A(n1657), .B(n1607), .Z(n1593) );
  XNOR U2447 ( .A(n1585), .B(n1584), .Z(n1607) );
  XOR U2448 ( .A(n1658), .B(n1580), .Z(n1584) );
  XNOR U2449 ( .A(n1578), .B(n1659), .Z(n1580) );
  ANDN U2450 ( .A(n1426), .B(n1063), .Z(n1659) );
  XOR U2451 ( .A(n1660), .B(n1661), .Z(n1578) );
  AND U2452 ( .A(n1662), .B(n1663), .Z(n1661) );
  XNOR U2453 ( .A(n1664), .B(n1660), .Z(n1663) );
  AND U2454 ( .A(n1061), .B(n1363), .Z(n1582) );
  XNOR U2455 ( .A(n1589), .B(n1591), .Z(n1585) );
  NANDN U2456 ( .B(n1228), .A(n1147), .Z(n1591) );
  XNOR U2457 ( .A(n1587), .B(n1668), .Z(n1589) );
  ANDN U2458 ( .A(n1298), .B(n1149), .Z(n1668) );
  XNOR U2459 ( .A(n1606), .B(n1592), .Z(n1657) );
  XOR U2460 ( .A(n1675), .B(n1609), .Z(n1606) );
  XNOR U2461 ( .A(n1601), .B(n1603), .Z(n1609) );
  NAND U2462 ( .A(n977), .B(n1597), .Z(n1603) );
  XNOR U2463 ( .A(n1599), .B(n1676), .Z(n1601) );
  ANDN U2464 ( .A(n1604), .B(n979), .Z(n1676) );
  XOR U2465 ( .A(n1677), .B(n1678), .Z(n1599) );
  AND U2466 ( .A(n1679), .B(n1680), .Z(n1678) );
  XOR U2467 ( .A(n1681), .B(n1677), .Z(n1680) );
  XNOR U2468 ( .A(n1608), .B(n1605), .Z(n1675) );
  AND U2469 ( .A(n1686), .B(n1687), .Z(n1685) );
  NANDN U2470 ( .B(n1688), .A(n916), .Z(n1687) );
  NANDN U2471 ( .B(n1689), .A(n1690), .Z(n1686) );
  XNOR U2472 ( .A(n1617), .B(n1616), .Z(n1594) );
  XOR U2473 ( .A(n1694), .B(n1627), .Z(n1616) );
  XNOR U2474 ( .A(n1613), .B(n1614), .Z(n1627) );
  NANDN U2475 ( .B(n1041), .A(n1405), .Z(n1614) );
  XNOR U2476 ( .A(n1612), .B(n1695), .Z(n1613) );
  ANDN U2477 ( .A(n1082), .B(n1407), .Z(n1695) );
  XNOR U2478 ( .A(n1626), .B(n1615), .Z(n1694) );
  XOR U2479 ( .A(n1702), .B(n1622), .Z(n1626) );
  XNOR U2480 ( .A(n1620), .B(n1703), .Z(n1622) );
  ANDN U2481 ( .A(n1189), .B(n1272), .Z(n1703) );
  XOR U2482 ( .A(n1704), .B(n1705), .Z(n1620) );
  AND U2483 ( .A(n1706), .B(n1707), .Z(n1705) );
  XNOR U2484 ( .A(n1708), .B(n1704), .Z(n1707) );
  AND U2485 ( .A(n1270), .B(n1135), .Z(n1624) );
  XOR U2486 ( .A(n1637), .B(n1636), .Z(n1617) );
  XOR U2487 ( .A(n1712), .B(n1632), .Z(n1636) );
  XNOR U2488 ( .A(n1630), .B(n1713), .Z(n1632) );
  ANDN U2489 ( .A(n1014), .B(n1559), .Z(n1713) );
  XOR U2490 ( .A(n1714), .B(n1715), .Z(n1630) );
  AND U2491 ( .A(n1716), .B(n1717), .Z(n1715) );
  XNOR U2492 ( .A(n1718), .B(n1714), .Z(n1717) );
  AND U2493 ( .A(n1557), .B(n973), .Z(n1634) );
  XOR U2494 ( .A(n1644), .B(n1643), .Z(n1637) );
  NAND U2495 ( .A(n1722), .B(n917), .Z(n1643) );
  XOR U2496 ( .A(n1642), .B(n1723), .Z(n1644) );
  ANDN U2497 ( .A(n948), .B(n1724), .Z(n1723) );
  ANDN U2498 ( .A(n1725), .B(n1726), .Z(n1642) );
  NAND U2499 ( .A(n1727), .B(n1728), .Z(n1725) );
  IV U2500 ( .A(n1645), .Z(n1646) );
  MUX U2501 ( .IN0(Y[14]), .IN1(n816), .SEL(n869), .F(n327) );
  XOR U2502 ( .A(n1733), .B(Y0[15]), .Z(n816) );
  XOR U2503 ( .A(n1734), .B(n1735), .Z(n1733) );
  AND U2504 ( .A(n881), .B(n1737), .Z(n1736) );
  XOR U2505 ( .A(n1731), .B(n1735), .Z(n1737) );
  XOR U2506 ( .A(n1730), .B(n1735), .Z(n1731) );
  XNOR U2507 ( .A(n1656), .B(n1655), .Z(n1735) );
  XOR U2508 ( .A(n1738), .B(n1739), .Z(n1655) );
  XOR U2509 ( .A(n1740), .B(n1741), .Z(n1739) );
  XOR U2510 ( .A(n1742), .B(n1740), .Z(n1741) );
  XNOR U2511 ( .A(n1748), .B(n1684), .Z(n1673) );
  XNOR U2512 ( .A(n1667), .B(n1666), .Z(n1684) );
  XOR U2513 ( .A(n1749), .B(n1662), .Z(n1666) );
  XNOR U2514 ( .A(n1660), .B(n1750), .Z(n1662) );
  ANDN U2515 ( .A(n1426), .B(n1107), .Z(n1750) );
  AND U2516 ( .A(n1105), .B(n1363), .Z(n1664) );
  XNOR U2517 ( .A(n1670), .B(n1671), .Z(n1667) );
  NANDN U2518 ( .B(n1228), .A(n1206), .Z(n1671) );
  XNOR U2519 ( .A(n1669), .B(n1757), .Z(n1670) );
  ANDN U2520 ( .A(n1298), .B(n1208), .Z(n1757) );
  XOR U2521 ( .A(n1758), .B(n1759), .Z(n1669) );
  AND U2522 ( .A(n1760), .B(n1761), .Z(n1759) );
  XOR U2523 ( .A(n1762), .B(n1758), .Z(n1761) );
  XNOR U2524 ( .A(n1683), .B(n1672), .Z(n1748) );
  XOR U2525 ( .A(n1766), .B(n1693), .Z(n1683) );
  XNOR U2526 ( .A(n1679), .B(n1681), .Z(n1693) );
  NAND U2527 ( .A(n1021), .B(n1597), .Z(n1681) );
  XNOR U2528 ( .A(n1677), .B(n1767), .Z(n1679) );
  ANDN U2529 ( .A(n1604), .B(n1023), .Z(n1767) );
  XOR U2530 ( .A(n1768), .B(n1769), .Z(n1677) );
  AND U2531 ( .A(n1770), .B(n1771), .Z(n1769) );
  XOR U2532 ( .A(n1772), .B(n1768), .Z(n1771) );
  XNOR U2533 ( .A(n1692), .B(n1682), .Z(n1766) );
  XOR U2534 ( .A(n1780), .B(n1690), .Z(n1776) );
  AND U2535 ( .A(n946), .B(n1781), .Z(n1690) );
  NAND U2536 ( .A(n1782), .B(n1689), .Z(n1780) );
  XOR U2537 ( .A(n1783), .B(n1784), .Z(n1689) );
  AND U2538 ( .A(n1785), .B(n1786), .Z(n1784) );
  XNOR U2539 ( .A(n1787), .B(n1783), .Z(n1786) );
  NANDN U2540 ( .B(n949), .A(n1788), .Z(n1782) );
  XNOR U2541 ( .A(n1701), .B(n1700), .Z(n1674) );
  XOR U2542 ( .A(n1789), .B(n1711), .Z(n1700) );
  XNOR U2543 ( .A(n1697), .B(n1698), .Z(n1711) );
  NANDN U2544 ( .B(n1041), .A(n1479), .Z(n1698) );
  XNOR U2545 ( .A(n1696), .B(n1790), .Z(n1697) );
  ANDN U2546 ( .A(n1082), .B(n1481), .Z(n1790) );
  XNOR U2547 ( .A(n1710), .B(n1699), .Z(n1789) );
  XOR U2548 ( .A(n1797), .B(n1706), .Z(n1710) );
  XNOR U2549 ( .A(n1704), .B(n1798), .Z(n1706) );
  ANDN U2550 ( .A(n1189), .B(n1340), .Z(n1798) );
  AND U2551 ( .A(n1338), .B(n1135), .Z(n1708) );
  XOR U2552 ( .A(n1721), .B(n1720), .Z(n1701) );
  XOR U2553 ( .A(n1805), .B(n1716), .Z(n1720) );
  XNOR U2554 ( .A(n1714), .B(n1806), .Z(n1716) );
  ANDN U2555 ( .A(n1014), .B(n1640), .Z(n1806) );
  AND U2556 ( .A(n1638), .B(n973), .Z(n1718) );
  XOR U2557 ( .A(n1728), .B(n1727), .Z(n1721) );
  NAND U2558 ( .A(n1813), .B(n917), .Z(n1727) );
  XNOR U2559 ( .A(n1726), .B(n1814), .Z(n1728) );
  ANDN U2560 ( .A(n948), .B(n1815), .Z(n1814) );
  NAND U2561 ( .A(n1816), .B(n1817), .Z(n1726) );
  NAND U2562 ( .A(n1818), .B(n1819), .Z(n1816) );
  IV U2563 ( .A(n1729), .Z(n1730) );
  MUX U2564 ( .IN0(Y[13]), .IN1(n813), .SEL(n869), .F(n326) );
  XOR U2565 ( .A(n1824), .B(Y0[14]), .Z(n813) );
  XOR U2566 ( .A(n1825), .B(n1826), .Z(n1824) );
  AND U2567 ( .A(n881), .B(n1828), .Z(n1827) );
  XOR U2568 ( .A(n1822), .B(n1826), .Z(n1828) );
  XOR U2569 ( .A(n1821), .B(n1826), .Z(n1822) );
  XOR U2570 ( .A(n1829), .B(n1743), .Z(n1746) );
  NAND U2571 ( .A(n1740), .B(n1833), .Z(n1744) );
  AND U2572 ( .A(n1834), .B(n1835), .Z(n1833) );
  NANDN U2573 ( .B(n1836), .A(n916), .Z(n1835) );
  NANDN U2574 ( .B(n1837), .A(n1838), .Z(n1834) );
  AND U2575 ( .A(n1839), .B(n1840), .Z(n1740) );
  NANDN U2576 ( .B(n1841), .A(n1842), .Z(n1840) );
  OR U2577 ( .A(n1843), .B(n1844), .Z(n1839) );
  XNOR U2578 ( .A(n1765), .B(n1764), .Z(n1747) );
  XOR U2579 ( .A(n1848), .B(n1775), .Z(n1764) );
  XNOR U2580 ( .A(n1756), .B(n1755), .Z(n1775) );
  XOR U2581 ( .A(n1849), .B(n1752), .Z(n1755) );
  XNOR U2582 ( .A(n1751), .B(n1850), .Z(n1752) );
  ANDN U2583 ( .A(n1426), .B(n1149), .Z(n1850) );
  XOR U2584 ( .A(n1851), .B(n1852), .Z(n1751) );
  AND U2585 ( .A(n1853), .B(n1854), .Z(n1852) );
  XNOR U2586 ( .A(n1855), .B(n1851), .Z(n1854) );
  AND U2587 ( .A(n1147), .B(n1363), .Z(n1753) );
  XNOR U2588 ( .A(n1760), .B(n1762), .Z(n1756) );
  NANDN U2589 ( .B(n1228), .A(n1270), .Z(n1762) );
  XNOR U2590 ( .A(n1758), .B(n1859), .Z(n1760) );
  ANDN U2591 ( .A(n1298), .B(n1272), .Z(n1859) );
  XNOR U2592 ( .A(n1774), .B(n1763), .Z(n1848) );
  XOR U2593 ( .A(n1866), .B(n1779), .Z(n1774) );
  XNOR U2594 ( .A(n1770), .B(n1772), .Z(n1779) );
  NAND U2595 ( .A(n1061), .B(n1597), .Z(n1772) );
  XNOR U2596 ( .A(n1768), .B(n1867), .Z(n1770) );
  ANDN U2597 ( .A(n1604), .B(n1063), .Z(n1867) );
  XOR U2598 ( .A(n1868), .B(n1869), .Z(n1768) );
  AND U2599 ( .A(n1870), .B(n1871), .Z(n1869) );
  XOR U2600 ( .A(n1872), .B(n1868), .Z(n1871) );
  XNOR U2601 ( .A(n1778), .B(n1773), .Z(n1866) );
  XOR U2602 ( .A(n1876), .B(n1785), .Z(n1778) );
  XNOR U2603 ( .A(n1783), .B(n1877), .Z(n1785) );
  ANDN U2604 ( .A(n1788), .B(n979), .Z(n1877) );
  XOR U2605 ( .A(n1878), .B(n1879), .Z(n1783) );
  AND U2606 ( .A(n1880), .B(n1881), .Z(n1879) );
  XNOR U2607 ( .A(n1882), .B(n1878), .Z(n1881) );
  AND U2608 ( .A(n977), .B(n1781), .Z(n1787) );
  XNOR U2609 ( .A(n1796), .B(n1795), .Z(n1765) );
  XOR U2610 ( .A(n1886), .B(n1804), .Z(n1795) );
  XNOR U2611 ( .A(n1792), .B(n1793), .Z(n1804) );
  NANDN U2612 ( .B(n1041), .A(n1557), .Z(n1793) );
  XNOR U2613 ( .A(n1791), .B(n1887), .Z(n1792) );
  ANDN U2614 ( .A(n1082), .B(n1559), .Z(n1887) );
  XNOR U2615 ( .A(n1803), .B(n1794), .Z(n1886) );
  XOR U2616 ( .A(n1894), .B(n1800), .Z(n1803) );
  XNOR U2617 ( .A(n1799), .B(n1895), .Z(n1800) );
  ANDN U2618 ( .A(n1189), .B(n1407), .Z(n1895) );
  AND U2619 ( .A(n1405), .B(n1135), .Z(n1801) );
  XOR U2620 ( .A(n1812), .B(n1811), .Z(n1796) );
  XOR U2621 ( .A(n1902), .B(n1808), .Z(n1811) );
  XNOR U2622 ( .A(n1807), .B(n1903), .Z(n1808) );
  ANDN U2623 ( .A(n1014), .B(n1724), .Z(n1903) );
  AND U2624 ( .A(n1722), .B(n973), .Z(n1809) );
  XOR U2625 ( .A(n1819), .B(n1818), .Z(n1812) );
  NAND U2626 ( .A(n1910), .B(n917), .Z(n1818) );
  XOR U2627 ( .A(n1817), .B(n1911), .Z(n1819) );
  ANDN U2628 ( .A(n948), .B(n1912), .Z(n1911) );
  ANDN U2629 ( .A(n1913), .B(n1914), .Z(n1817) );
  NAND U2630 ( .A(n1915), .B(n1916), .Z(n1913) );
  IV U2631 ( .A(n1820), .Z(n1821) );
  MUX U2632 ( .IN0(Y[12]), .IN1(n810), .SEL(n869), .F(n325) );
  XOR U2633 ( .A(n1921), .B(Y0[13]), .Z(n810) );
  XNOR U2634 ( .A(n1922), .B(n1923), .Z(n1921) );
  AND U2635 ( .A(n881), .B(n1925), .Z(n1924) );
  XNOR U2636 ( .A(n1919), .B(n1923), .Z(n1925) );
  XNOR U2637 ( .A(n1918), .B(n1923), .Z(n1919) );
  XNOR U2638 ( .A(n1847), .B(n1846), .Z(n1923) );
  XOR U2639 ( .A(n1926), .B(n1831), .Z(n1846) );
  NANDN U2640 ( .B(n1927), .A(n1928), .Z(n1837) );
  XOR U2641 ( .A(n1931), .B(n1844), .Z(n1841) );
  NAND U2642 ( .A(n1932), .B(n946), .Z(n1844) );
  NAND U2643 ( .A(n1933), .B(n1843), .Z(n1931) );
  NANDN U2644 ( .B(n949), .A(n1937), .Z(n1933) );
  XNOR U2645 ( .A(n1830), .B(n1845), .Z(n1926) );
  IV U2646 ( .A(n1832), .Z(n1830) );
  XNOR U2647 ( .A(n1865), .B(n1864), .Z(n1847) );
  XOR U2648 ( .A(n1944), .B(n1875), .Z(n1864) );
  XNOR U2649 ( .A(n1858), .B(n1857), .Z(n1875) );
  XOR U2650 ( .A(n1945), .B(n1853), .Z(n1857) );
  XNOR U2651 ( .A(n1851), .B(n1946), .Z(n1853) );
  ANDN U2652 ( .A(n1426), .B(n1208), .Z(n1946) );
  XOR U2653 ( .A(n1947), .B(n1948), .Z(n1851) );
  AND U2654 ( .A(n1949), .B(n1950), .Z(n1948) );
  XNOR U2655 ( .A(n1951), .B(n1947), .Z(n1950) );
  AND U2656 ( .A(n1206), .B(n1363), .Z(n1855) );
  XNOR U2657 ( .A(n1861), .B(n1862), .Z(n1858) );
  NANDN U2658 ( .B(n1228), .A(n1338), .Z(n1862) );
  XNOR U2659 ( .A(n1860), .B(n1955), .Z(n1861) );
  ANDN U2660 ( .A(n1298), .B(n1340), .Z(n1955) );
  XNOR U2661 ( .A(n1874), .B(n1863), .Z(n1944) );
  XOR U2662 ( .A(n1962), .B(n1885), .Z(n1874) );
  XNOR U2663 ( .A(n1870), .B(n1872), .Z(n1885) );
  NAND U2664 ( .A(n1105), .B(n1597), .Z(n1872) );
  XNOR U2665 ( .A(n1868), .B(n1963), .Z(n1870) );
  ANDN U2666 ( .A(n1604), .B(n1107), .Z(n1963) );
  XOR U2667 ( .A(n1964), .B(n1965), .Z(n1868) );
  AND U2668 ( .A(n1966), .B(n1967), .Z(n1965) );
  XOR U2669 ( .A(n1968), .B(n1964), .Z(n1967) );
  XNOR U2670 ( .A(n1884), .B(n1873), .Z(n1962) );
  XOR U2671 ( .A(n1972), .B(n1880), .Z(n1884) );
  XNOR U2672 ( .A(n1878), .B(n1973), .Z(n1880) );
  ANDN U2673 ( .A(n1788), .B(n1023), .Z(n1973) );
  XOR U2674 ( .A(n1974), .B(n1975), .Z(n1878) );
  AND U2675 ( .A(n1976), .B(n1977), .Z(n1975) );
  XNOR U2676 ( .A(n1978), .B(n1974), .Z(n1977) );
  AND U2677 ( .A(n1021), .B(n1781), .Z(n1882) );
  XNOR U2678 ( .A(n1893), .B(n1892), .Z(n1865) );
  XOR U2679 ( .A(n1982), .B(n1901), .Z(n1892) );
  XNOR U2680 ( .A(n1889), .B(n1890), .Z(n1901) );
  NANDN U2681 ( .B(n1041), .A(n1638), .Z(n1890) );
  XNOR U2682 ( .A(n1888), .B(n1983), .Z(n1889) );
  ANDN U2683 ( .A(n1082), .B(n1640), .Z(n1983) );
  XNOR U2684 ( .A(n1900), .B(n1891), .Z(n1982) );
  XOR U2685 ( .A(n1990), .B(n1897), .Z(n1900) );
  XNOR U2686 ( .A(n1896), .B(n1991), .Z(n1897) );
  ANDN U2687 ( .A(n1189), .B(n1481), .Z(n1991) );
  AND U2688 ( .A(n1479), .B(n1135), .Z(n1898) );
  XOR U2689 ( .A(n1909), .B(n1908), .Z(n1893) );
  XOR U2690 ( .A(n1998), .B(n1905), .Z(n1908) );
  XNOR U2691 ( .A(n1904), .B(n1999), .Z(n1905) );
  ANDN U2692 ( .A(n1014), .B(n1815), .Z(n1999) );
  AND U2693 ( .A(n1813), .B(n973), .Z(n1906) );
  XOR U2694 ( .A(n1916), .B(n1915), .Z(n1909) );
  NAND U2695 ( .A(n2006), .B(n917), .Z(n1915) );
  XNOR U2696 ( .A(n1914), .B(n2007), .Z(n1916) );
  ANDN U2697 ( .A(n948), .B(n2008), .Z(n2007) );
  NAND U2698 ( .A(n2009), .B(n2010), .Z(n1914) );
  NAND U2699 ( .A(n2011), .B(n2012), .Z(n2009) );
  IV U2700 ( .A(n1917), .Z(n1918) );
  MUX U2701 ( .IN0(Y[11]), .IN1(n807), .SEL(n869), .F(n324) );
  XOR U2702 ( .A(n2017), .B(Y0[12]), .Z(n807) );
  XOR U2703 ( .A(n2018), .B(n2019), .Z(n2017) );
  AND U2704 ( .A(n881), .B(n2021), .Z(n2020) );
  XOR U2705 ( .A(n2015), .B(n2019), .Z(n2021) );
  XOR U2706 ( .A(n2014), .B(n2019), .Z(n2015) );
  XNOR U2707 ( .A(n2022), .B(n1943), .Z(n1939) );
  XOR U2708 ( .A(n1928), .B(n1927), .Z(n1943) );
  NANDN U2709 ( .B(n2023), .A(n2024), .Z(n1927) );
  AND U2710 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U2711 ( .B(n2028), .A(n916), .Z(n2027) );
  NANDN U2712 ( .B(n2029), .A(n2030), .Z(n2026) );
  XNOR U2713 ( .A(n1935), .B(n1936), .Z(n1930) );
  NAND U2714 ( .A(n1932), .B(n977), .Z(n1936) );
  XNOR U2715 ( .A(n1934), .B(n2034), .Z(n1935) );
  ANDN U2716 ( .A(n1937), .B(n979), .Z(n2034) );
  XNOR U2717 ( .A(n1942), .B(n1938), .Z(n2022) );
  IV U2718 ( .A(n1941), .Z(n1942) );
  XNOR U2719 ( .A(n1961), .B(n1960), .Z(n1940) );
  XOR U2720 ( .A(n2044), .B(n1971), .Z(n1960) );
  XNOR U2721 ( .A(n1954), .B(n1953), .Z(n1971) );
  XOR U2722 ( .A(n2045), .B(n1949), .Z(n1953) );
  XNOR U2723 ( .A(n1947), .B(n2046), .Z(n1949) );
  ANDN U2724 ( .A(n1426), .B(n1272), .Z(n2046) );
  AND U2725 ( .A(n1270), .B(n1363), .Z(n1951) );
  XNOR U2726 ( .A(n1957), .B(n1958), .Z(n1954) );
  NANDN U2727 ( .B(n1228), .A(n1405), .Z(n1958) );
  XNOR U2728 ( .A(n1956), .B(n2053), .Z(n1957) );
  ANDN U2729 ( .A(n1298), .B(n1407), .Z(n2053) );
  XNOR U2730 ( .A(n1970), .B(n1959), .Z(n2044) );
  XOR U2731 ( .A(n2060), .B(n1981), .Z(n1970) );
  XNOR U2732 ( .A(n1966), .B(n1968), .Z(n1981) );
  NAND U2733 ( .A(n1147), .B(n1597), .Z(n1968) );
  XNOR U2734 ( .A(n1964), .B(n2061), .Z(n1966) );
  ANDN U2735 ( .A(n1604), .B(n1149), .Z(n2061) );
  XNOR U2736 ( .A(n1980), .B(n1969), .Z(n2060) );
  XOR U2737 ( .A(n2068), .B(n1976), .Z(n1980) );
  XNOR U2738 ( .A(n1974), .B(n2069), .Z(n1976) );
  ANDN U2739 ( .A(n1788), .B(n1063), .Z(n2069) );
  XOR U2740 ( .A(n2070), .B(n2071), .Z(n1974) );
  AND U2741 ( .A(n2072), .B(n2073), .Z(n2071) );
  XNOR U2742 ( .A(n2074), .B(n2070), .Z(n2073) );
  AND U2743 ( .A(n1061), .B(n1781), .Z(n1978) );
  XNOR U2744 ( .A(n1989), .B(n1988), .Z(n1961) );
  XOR U2745 ( .A(n2078), .B(n1997), .Z(n1988) );
  XNOR U2746 ( .A(n1985), .B(n1986), .Z(n1997) );
  NANDN U2747 ( .B(n1041), .A(n1722), .Z(n1986) );
  XNOR U2748 ( .A(n1984), .B(n2079), .Z(n1985) );
  ANDN U2749 ( .A(n1082), .B(n1724), .Z(n2079) );
  XNOR U2750 ( .A(n1996), .B(n1987), .Z(n2078) );
  XOR U2751 ( .A(n2086), .B(n1993), .Z(n1996) );
  XNOR U2752 ( .A(n1992), .B(n2087), .Z(n1993) );
  ANDN U2753 ( .A(n1189), .B(n1559), .Z(n2087) );
  AND U2754 ( .A(n1557), .B(n1135), .Z(n1994) );
  XOR U2755 ( .A(n2005), .B(n2004), .Z(n1989) );
  XOR U2756 ( .A(n2094), .B(n2001), .Z(n2004) );
  XNOR U2757 ( .A(n2000), .B(n2095), .Z(n2001) );
  ANDN U2758 ( .A(n1014), .B(n1912), .Z(n2095) );
  AND U2759 ( .A(n1910), .B(n973), .Z(n2002) );
  XOR U2760 ( .A(n2012), .B(n2011), .Z(n2005) );
  NAND U2761 ( .A(n2102), .B(n917), .Z(n2011) );
  XOR U2762 ( .A(n2010), .B(n2103), .Z(n2012) );
  ANDN U2763 ( .A(n948), .B(n2104), .Z(n2103) );
  ANDN U2764 ( .A(n2105), .B(n2106), .Z(n2010) );
  NAND U2765 ( .A(n2107), .B(n2108), .Z(n2105) );
  IV U2766 ( .A(n2013), .Z(n2014) );
  MUX U2767 ( .IN0(Y[10]), .IN1(n804), .SEL(n869), .F(n323) );
  XOR U2768 ( .A(n2113), .B(Y0[11]), .Z(n804) );
  XNOR U2769 ( .A(n2114), .B(n2115), .Z(n2113) );
  AND U2770 ( .A(n881), .B(n2117), .Z(n2116) );
  XNOR U2771 ( .A(n2111), .B(n2115), .Z(n2117) );
  XNOR U2772 ( .A(n2110), .B(n2115), .Z(n2111) );
  XNOR U2773 ( .A(n2040), .B(n2039), .Z(n2115) );
  XOR U2774 ( .A(n2118), .B(n2043), .Z(n2039) );
  XOR U2775 ( .A(n2033), .B(n2032), .Z(n2023) );
  XOR U2776 ( .A(n2126), .B(n2030), .Z(n2122) );
  AND U2777 ( .A(n2127), .B(n946), .Z(n2030) );
  NAND U2778 ( .A(n2128), .B(n2029), .Z(n2126) );
  XOR U2779 ( .A(n2129), .B(n2130), .Z(n2029) );
  AND U2780 ( .A(n2131), .B(n2132), .Z(n2130) );
  XNOR U2781 ( .A(n2133), .B(n2129), .Z(n2132) );
  NANDN U2782 ( .B(n949), .A(n2134), .Z(n2128) );
  XNOR U2783 ( .A(n2036), .B(n2037), .Z(n2033) );
  NAND U2784 ( .A(n1932), .B(n1021), .Z(n2037) );
  XNOR U2785 ( .A(n2035), .B(n2135), .Z(n2036) );
  ANDN U2786 ( .A(n1937), .B(n1023), .Z(n2135) );
  XNOR U2787 ( .A(n2042), .B(n2038), .Z(n2118) );
  IV U2788 ( .A(n2041), .Z(n2042) );
  XNOR U2789 ( .A(n2059), .B(n2058), .Z(n2040) );
  XOR U2790 ( .A(n2145), .B(n2067), .Z(n2058) );
  XNOR U2791 ( .A(n2052), .B(n2051), .Z(n2067) );
  XOR U2792 ( .A(n2146), .B(n2048), .Z(n2051) );
  XNOR U2793 ( .A(n2047), .B(n2147), .Z(n2048) );
  ANDN U2794 ( .A(n1426), .B(n1340), .Z(n2147) );
  AND U2795 ( .A(n1338), .B(n1363), .Z(n2049) );
  XNOR U2796 ( .A(n2055), .B(n2056), .Z(n2052) );
  NANDN U2797 ( .B(n1228), .A(n1479), .Z(n2056) );
  XNOR U2798 ( .A(n2054), .B(n2154), .Z(n2055) );
  ANDN U2799 ( .A(n1298), .B(n1481), .Z(n2154) );
  XNOR U2800 ( .A(n2066), .B(n2057), .Z(n2145) );
  XOR U2801 ( .A(n2161), .B(n2077), .Z(n2066) );
  XNOR U2802 ( .A(n2063), .B(n2064), .Z(n2077) );
  NAND U2803 ( .A(n1206), .B(n1597), .Z(n2064) );
  XNOR U2804 ( .A(n2062), .B(n2162), .Z(n2063) );
  ANDN U2805 ( .A(n1604), .B(n1208), .Z(n2162) );
  XNOR U2806 ( .A(n2076), .B(n2065), .Z(n2161) );
  XOR U2807 ( .A(n2169), .B(n2072), .Z(n2076) );
  XNOR U2808 ( .A(n2070), .B(n2170), .Z(n2072) );
  ANDN U2809 ( .A(n1788), .B(n1107), .Z(n2170) );
  XOR U2810 ( .A(n2171), .B(n2172), .Z(n2070) );
  AND U2811 ( .A(n2173), .B(n2174), .Z(n2172) );
  XNOR U2812 ( .A(n2175), .B(n2171), .Z(n2174) );
  AND U2813 ( .A(n1105), .B(n1781), .Z(n2074) );
  XNOR U2814 ( .A(n2085), .B(n2084), .Z(n2059) );
  XOR U2815 ( .A(n2179), .B(n2093), .Z(n2084) );
  XNOR U2816 ( .A(n2081), .B(n2082), .Z(n2093) );
  NANDN U2817 ( .B(n1041), .A(n1813), .Z(n2082) );
  XNOR U2818 ( .A(n2080), .B(n2180), .Z(n2081) );
  ANDN U2819 ( .A(n1082), .B(n1815), .Z(n2180) );
  XNOR U2820 ( .A(n2092), .B(n2083), .Z(n2179) );
  XOR U2821 ( .A(n2187), .B(n2089), .Z(n2092) );
  XNOR U2822 ( .A(n2088), .B(n2188), .Z(n2089) );
  ANDN U2823 ( .A(n1189), .B(n1640), .Z(n2188) );
  AND U2824 ( .A(n1638), .B(n1135), .Z(n2090) );
  XOR U2825 ( .A(n2101), .B(n2100), .Z(n2085) );
  XOR U2826 ( .A(n2195), .B(n2097), .Z(n2100) );
  XNOR U2827 ( .A(n2096), .B(n2196), .Z(n2097) );
  ANDN U2828 ( .A(n1014), .B(n2008), .Z(n2196) );
  AND U2829 ( .A(n2006), .B(n973), .Z(n2098) );
  XOR U2830 ( .A(n2108), .B(n2107), .Z(n2101) );
  NAND U2831 ( .A(n2203), .B(n917), .Z(n2107) );
  XNOR U2832 ( .A(n2106), .B(n2204), .Z(n2108) );
  ANDN U2833 ( .A(n948), .B(n2205), .Z(n2204) );
  NAND U2834 ( .A(n2206), .B(n2207), .Z(n2106) );
  NAND U2835 ( .A(n2208), .B(n2209), .Z(n2206) );
  IV U2836 ( .A(n2109), .Z(n2110) );
  MUX U2837 ( .IN0(Y[9]), .IN1(n801), .SEL(n869), .F(n322) );
  XOR U2838 ( .A(n2214), .B(Y0[10]), .Z(n801) );
  XOR U2839 ( .A(n2215), .B(n2216), .Z(n2214) );
  AND U2840 ( .A(n881), .B(n2218), .Z(n2217) );
  XOR U2841 ( .A(n2212), .B(n2216), .Z(n2218) );
  XOR U2842 ( .A(n2211), .B(n2216), .Z(n2212) );
  XNOR U2843 ( .A(n2219), .B(n2144), .Z(n2140) );
  XNOR U2844 ( .A(n2121), .B(n2120), .Z(n2144) );
  XOR U2845 ( .A(n2119), .B(n2220), .Z(n2120) );
  AND U2846 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2847 ( .B(n2223), .A(n2224), .Z(n2222) );
  AND U2848 ( .A(n2225), .B(n2226), .Z(n2221) );
  NANDN U2849 ( .B(n2227), .A(n916), .Z(n2226) );
  OR U2850 ( .A(n2228), .B(n2229), .Z(n2225) );
  XNOR U2851 ( .A(n2125), .B(n2124), .Z(n2121) );
  XOR U2852 ( .A(n2233), .B(n2131), .Z(n2124) );
  XNOR U2853 ( .A(n2129), .B(n2234), .Z(n2131) );
  ANDN U2854 ( .A(n2134), .B(n979), .Z(n2234) );
  XOR U2855 ( .A(n2235), .B(n2236), .Z(n2129) );
  AND U2856 ( .A(n2237), .B(n2238), .Z(n2236) );
  XNOR U2857 ( .A(n2239), .B(n2235), .Z(n2238) );
  AND U2858 ( .A(n2127), .B(n977), .Z(n2133) );
  XNOR U2859 ( .A(n2137), .B(n2138), .Z(n2125) );
  NAND U2860 ( .A(n1932), .B(n1061), .Z(n2138) );
  XNOR U2861 ( .A(n2136), .B(n2243), .Z(n2137) );
  ANDN U2862 ( .A(n1937), .B(n1063), .Z(n2243) );
  XNOR U2863 ( .A(n2143), .B(n2139), .Z(n2219) );
  IV U2864 ( .A(n2142), .Z(n2143) );
  XNOR U2865 ( .A(n2160), .B(n2159), .Z(n2141) );
  XOR U2866 ( .A(n2253), .B(n2168), .Z(n2159) );
  XNOR U2867 ( .A(n2153), .B(n2152), .Z(n2168) );
  XOR U2868 ( .A(n2254), .B(n2149), .Z(n2152) );
  XNOR U2869 ( .A(n2148), .B(n2255), .Z(n2149) );
  ANDN U2870 ( .A(n1426), .B(n1407), .Z(n2255) );
  AND U2871 ( .A(n1405), .B(n1363), .Z(n2150) );
  XNOR U2872 ( .A(n2156), .B(n2157), .Z(n2153) );
  NANDN U2873 ( .B(n1228), .A(n1557), .Z(n2157) );
  XNOR U2874 ( .A(n2155), .B(n2262), .Z(n2156) );
  ANDN U2875 ( .A(n1298), .B(n1559), .Z(n2262) );
  XNOR U2876 ( .A(n2167), .B(n2158), .Z(n2253) );
  XOR U2877 ( .A(n2269), .B(n2178), .Z(n2167) );
  XNOR U2878 ( .A(n2164), .B(n2165), .Z(n2178) );
  NAND U2879 ( .A(n1270), .B(n1597), .Z(n2165) );
  XNOR U2880 ( .A(n2163), .B(n2270), .Z(n2164) );
  ANDN U2881 ( .A(n1604), .B(n1272), .Z(n2270) );
  XNOR U2882 ( .A(n2177), .B(n2166), .Z(n2269) );
  XOR U2883 ( .A(n2277), .B(n2173), .Z(n2177) );
  XNOR U2884 ( .A(n2171), .B(n2278), .Z(n2173) );
  ANDN U2885 ( .A(n1788), .B(n1149), .Z(n2278) );
  AND U2886 ( .A(n1147), .B(n1781), .Z(n2175) );
  XNOR U2887 ( .A(n2186), .B(n2185), .Z(n2160) );
  XOR U2888 ( .A(n2285), .B(n2194), .Z(n2185) );
  XNOR U2889 ( .A(n2182), .B(n2183), .Z(n2194) );
  NANDN U2890 ( .B(n1041), .A(n1910), .Z(n2183) );
  XNOR U2891 ( .A(n2181), .B(n2286), .Z(n2182) );
  ANDN U2892 ( .A(n1082), .B(n1912), .Z(n2286) );
  XNOR U2893 ( .A(n2193), .B(n2184), .Z(n2285) );
  XOR U2894 ( .A(n2293), .B(n2190), .Z(n2193) );
  XNOR U2895 ( .A(n2189), .B(n2294), .Z(n2190) );
  ANDN U2896 ( .A(n1189), .B(n1724), .Z(n2294) );
  AND U2897 ( .A(n1722), .B(n1135), .Z(n2191) );
  XOR U2898 ( .A(n2202), .B(n2201), .Z(n2186) );
  XOR U2899 ( .A(n2301), .B(n2198), .Z(n2201) );
  XNOR U2900 ( .A(n2197), .B(n2302), .Z(n2198) );
  ANDN U2901 ( .A(n1014), .B(n2104), .Z(n2302) );
  AND U2902 ( .A(n2102), .B(n973), .Z(n2199) );
  XOR U2903 ( .A(n2209), .B(n2208), .Z(n2202) );
  NAND U2904 ( .A(n2309), .B(n917), .Z(n2208) );
  XOR U2905 ( .A(n2207), .B(n2310), .Z(n2209) );
  ANDN U2906 ( .A(n948), .B(n2311), .Z(n2310) );
  ANDN U2907 ( .A(n2312), .B(n2313), .Z(n2207) );
  NAND U2908 ( .A(n2314), .B(n2315), .Z(n2312) );
  IV U2909 ( .A(n2210), .Z(n2211) );
  MUX U2910 ( .IN0(Y[8]), .IN1(n798), .SEL(n869), .F(n321) );
  XOR U2911 ( .A(n2320), .B(Y0[9]), .Z(n798) );
  XOR U2912 ( .A(n2321), .B(n2322), .Z(n2320) );
  AND U2913 ( .A(n881), .B(n2324), .Z(n2323) );
  XOR U2914 ( .A(n2318), .B(n2322), .Z(n2324) );
  XOR U2915 ( .A(n2317), .B(n2322), .Z(n2318) );
  XNOR U2916 ( .A(n2325), .B(n2252), .Z(n2248) );
  XNOR U2917 ( .A(n2232), .B(n2231), .Z(n2252) );
  XOR U2918 ( .A(n2326), .B(n2228), .Z(n2231) );
  XNOR U2919 ( .A(n2327), .B(n2224), .Z(n2228) );
  AND U2920 ( .A(n2328), .B(n946), .Z(n2224) );
  NAND U2921 ( .A(n2329), .B(n2223), .Z(n2327) );
  NANDN U2922 ( .B(n949), .A(n2333), .Z(n2329) );
  XNOR U2923 ( .A(n2229), .B(n2230), .Z(n2326) );
  XNOR U2924 ( .A(n2337), .B(n2340), .Z(n2339) );
  XNOR U2925 ( .A(n2242), .B(n2241), .Z(n2232) );
  XOR U2926 ( .A(n2341), .B(n2237), .Z(n2241) );
  XNOR U2927 ( .A(n2235), .B(n2342), .Z(n2237) );
  ANDN U2928 ( .A(n2134), .B(n1023), .Z(n2342) );
  XOR U2929 ( .A(n2343), .B(n2344), .Z(n2235) );
  AND U2930 ( .A(n2345), .B(n2346), .Z(n2344) );
  XNOR U2931 ( .A(n2347), .B(n2343), .Z(n2346) );
  AND U2932 ( .A(n2127), .B(n1021), .Z(n2239) );
  XNOR U2933 ( .A(n2245), .B(n2246), .Z(n2242) );
  NAND U2934 ( .A(n1932), .B(n1105), .Z(n2246) );
  XNOR U2935 ( .A(n2244), .B(n2351), .Z(n2245) );
  ANDN U2936 ( .A(n1937), .B(n1107), .Z(n2351) );
  XNOR U2937 ( .A(n2251), .B(n2247), .Z(n2325) );
  IV U2938 ( .A(n2250), .Z(n2251) );
  XNOR U2939 ( .A(n2268), .B(n2267), .Z(n2249) );
  XOR U2940 ( .A(n2360), .B(n2276), .Z(n2267) );
  XNOR U2941 ( .A(n2261), .B(n2260), .Z(n2276) );
  XOR U2942 ( .A(n2361), .B(n2257), .Z(n2260) );
  XNOR U2943 ( .A(n2256), .B(n2362), .Z(n2257) );
  ANDN U2944 ( .A(n1426), .B(n1481), .Z(n2362) );
  AND U2945 ( .A(n1479), .B(n1363), .Z(n2258) );
  XNOR U2946 ( .A(n2264), .B(n2265), .Z(n2261) );
  NANDN U2947 ( .B(n1228), .A(n1638), .Z(n2265) );
  XNOR U2948 ( .A(n2263), .B(n2369), .Z(n2264) );
  ANDN U2949 ( .A(n1298), .B(n1640), .Z(n2369) );
  XNOR U2950 ( .A(n2275), .B(n2266), .Z(n2360) );
  XOR U2951 ( .A(n2376), .B(n2284), .Z(n2275) );
  XNOR U2952 ( .A(n2272), .B(n2273), .Z(n2284) );
  NAND U2953 ( .A(n1338), .B(n1597), .Z(n2273) );
  XNOR U2954 ( .A(n2271), .B(n2377), .Z(n2272) );
  ANDN U2955 ( .A(n1604), .B(n1340), .Z(n2377) );
  XNOR U2956 ( .A(n2283), .B(n2274), .Z(n2376) );
  XOR U2957 ( .A(n2384), .B(n2280), .Z(n2283) );
  XNOR U2958 ( .A(n2279), .B(n2385), .Z(n2280) );
  ANDN U2959 ( .A(n1788), .B(n1208), .Z(n2385) );
  AND U2960 ( .A(n1206), .B(n1781), .Z(n2281) );
  XNOR U2961 ( .A(n2292), .B(n2291), .Z(n2268) );
  XOR U2962 ( .A(n2392), .B(n2300), .Z(n2291) );
  XNOR U2963 ( .A(n2288), .B(n2289), .Z(n2300) );
  NANDN U2964 ( .B(n1041), .A(n2006), .Z(n2289) );
  XNOR U2965 ( .A(n2287), .B(n2393), .Z(n2288) );
  ANDN U2966 ( .A(n1082), .B(n2008), .Z(n2393) );
  XNOR U2967 ( .A(n2299), .B(n2290), .Z(n2392) );
  XOR U2968 ( .A(n2400), .B(n2296), .Z(n2299) );
  XNOR U2969 ( .A(n2295), .B(n2401), .Z(n2296) );
  ANDN U2970 ( .A(n1189), .B(n1815), .Z(n2401) );
  AND U2971 ( .A(n1813), .B(n1135), .Z(n2297) );
  XOR U2972 ( .A(n2308), .B(n2307), .Z(n2292) );
  XOR U2973 ( .A(n2408), .B(n2304), .Z(n2307) );
  XNOR U2974 ( .A(n2303), .B(n2409), .Z(n2304) );
  ANDN U2975 ( .A(n1014), .B(n2205), .Z(n2409) );
  AND U2976 ( .A(n2203), .B(n973), .Z(n2305) );
  XOR U2977 ( .A(n2315), .B(n2314), .Z(n2308) );
  NAND U2978 ( .A(n2416), .B(n917), .Z(n2314) );
  XNOR U2979 ( .A(n2313), .B(n2417), .Z(n2315) );
  ANDN U2980 ( .A(n948), .B(n2418), .Z(n2417) );
  NAND U2981 ( .A(n2419), .B(n2420), .Z(n2313) );
  NAND U2982 ( .A(n2421), .B(n2422), .Z(n2419) );
  IV U2983 ( .A(n2316), .Z(n2317) );
  MUX U2984 ( .IN0(Y[7]), .IN1(n795), .SEL(n869), .F(n320) );
  XOR U2985 ( .A(n2427), .B(Y0[8]), .Z(n795) );
  XOR U2986 ( .A(n2428), .B(n2429), .Z(n2427) );
  AND U2987 ( .A(n881), .B(n2431), .Z(n2430) );
  XOR U2988 ( .A(n2425), .B(n2429), .Z(n2431) );
  XOR U2989 ( .A(n2424), .B(n2429), .Z(n2425) );
  XNOR U2990 ( .A(n2432), .B(n2359), .Z(n2356) );
  XNOR U2991 ( .A(n2336), .B(n2335), .Z(n2359) );
  XOR U2992 ( .A(n2433), .B(n2340), .Z(n2335) );
  XNOR U2993 ( .A(n2331), .B(n2332), .Z(n2340) );
  NAND U2994 ( .A(n2328), .B(n977), .Z(n2332) );
  XNOR U2995 ( .A(n2330), .B(n2434), .Z(n2331) );
  ANDN U2996 ( .A(n2333), .B(n979), .Z(n2434) );
  XNOR U2997 ( .A(n2338), .B(n2334), .Z(n2433) );
  XOR U2998 ( .A(n2337), .B(n2441), .Z(n2338) );
  AND U2999 ( .A(n2442), .B(n2443), .Z(n2441) );
  NANDN U3000 ( .B(n2444), .A(n916), .Z(n2443) );
  NANDN U3001 ( .B(n2445), .A(n2446), .Z(n2442) );
  XNOR U3002 ( .A(n2350), .B(n2349), .Z(n2336) );
  XOR U3003 ( .A(n2450), .B(n2345), .Z(n2349) );
  XNOR U3004 ( .A(n2343), .B(n2451), .Z(n2345) );
  ANDN U3005 ( .A(n2134), .B(n1063), .Z(n2451) );
  AND U3006 ( .A(n2127), .B(n1061), .Z(n2347) );
  XNOR U3007 ( .A(n2353), .B(n2354), .Z(n2350) );
  NAND U3008 ( .A(n1932), .B(n1147), .Z(n2354) );
  XNOR U3009 ( .A(n2352), .B(n2458), .Z(n2353) );
  ANDN U3010 ( .A(n1937), .B(n1149), .Z(n2458) );
  XNOR U3011 ( .A(n2375), .B(n2374), .Z(n2357) );
  XOR U3012 ( .A(n2468), .B(n2383), .Z(n2374) );
  XNOR U3013 ( .A(n2368), .B(n2367), .Z(n2383) );
  XOR U3014 ( .A(n2469), .B(n2364), .Z(n2367) );
  XNOR U3015 ( .A(n2363), .B(n2470), .Z(n2364) );
  ANDN U3016 ( .A(n1426), .B(n1559), .Z(n2470) );
  AND U3017 ( .A(n1557), .B(n1363), .Z(n2365) );
  XNOR U3018 ( .A(n2371), .B(n2372), .Z(n2368) );
  NANDN U3019 ( .B(n1228), .A(n1722), .Z(n2372) );
  XNOR U3020 ( .A(n2370), .B(n2477), .Z(n2371) );
  ANDN U3021 ( .A(n1298), .B(n1724), .Z(n2477) );
  XNOR U3022 ( .A(n2382), .B(n2373), .Z(n2468) );
  XOR U3023 ( .A(n2484), .B(n2391), .Z(n2382) );
  XNOR U3024 ( .A(n2379), .B(n2380), .Z(n2391) );
  NAND U3025 ( .A(n1405), .B(n1597), .Z(n2380) );
  XNOR U3026 ( .A(n2378), .B(n2485), .Z(n2379) );
  ANDN U3027 ( .A(n1604), .B(n1407), .Z(n2485) );
  XNOR U3028 ( .A(n2390), .B(n2381), .Z(n2484) );
  XOR U3029 ( .A(n2492), .B(n2387), .Z(n2390) );
  XNOR U3030 ( .A(n2386), .B(n2493), .Z(n2387) );
  ANDN U3031 ( .A(n1788), .B(n1272), .Z(n2493) );
  AND U3032 ( .A(n1270), .B(n1781), .Z(n2388) );
  XNOR U3033 ( .A(n2399), .B(n2398), .Z(n2375) );
  XOR U3034 ( .A(n2500), .B(n2407), .Z(n2398) );
  XNOR U3035 ( .A(n2395), .B(n2396), .Z(n2407) );
  NANDN U3036 ( .B(n1041), .A(n2102), .Z(n2396) );
  XNOR U3037 ( .A(n2394), .B(n2501), .Z(n2395) );
  ANDN U3038 ( .A(n1082), .B(n2104), .Z(n2501) );
  XNOR U3039 ( .A(n2406), .B(n2397), .Z(n2500) );
  XOR U3040 ( .A(n2508), .B(n2403), .Z(n2406) );
  XNOR U3041 ( .A(n2402), .B(n2509), .Z(n2403) );
  ANDN U3042 ( .A(n1189), .B(n1912), .Z(n2509) );
  AND U3043 ( .A(n1910), .B(n1135), .Z(n2404) );
  XOR U3044 ( .A(n2415), .B(n2414), .Z(n2399) );
  XOR U3045 ( .A(n2516), .B(n2411), .Z(n2414) );
  XNOR U3046 ( .A(n2410), .B(n2517), .Z(n2411) );
  ANDN U3047 ( .A(n1014), .B(n2311), .Z(n2517) );
  AND U3048 ( .A(n2309), .B(n973), .Z(n2412) );
  XOR U3049 ( .A(n2422), .B(n2421), .Z(n2415) );
  NAND U3050 ( .A(n2524), .B(n917), .Z(n2421) );
  XOR U3051 ( .A(n2420), .B(n2525), .Z(n2422) );
  ANDN U3052 ( .A(n948), .B(n2526), .Z(n2525) );
  ANDN U3053 ( .A(n2527), .B(n2528), .Z(n2420) );
  NAND U3054 ( .A(n2529), .B(n2530), .Z(n2527) );
  IV U3055 ( .A(n2423), .Z(n2424) );
  MUX U3056 ( .IN0(Y[6]), .IN1(n792), .SEL(n869), .F(n319) );
  XOR U3057 ( .A(n2535), .B(Y0[7]), .Z(n792) );
  XOR U3058 ( .A(n2536), .B(n2537), .Z(n2535) );
  AND U3059 ( .A(n881), .B(n2539), .Z(n2538) );
  XOR U3060 ( .A(n2533), .B(n2537), .Z(n2539) );
  XOR U3061 ( .A(n2532), .B(n2537), .Z(n2533) );
  XNOR U3062 ( .A(n2540), .B(n2467), .Z(n2463) );
  XNOR U3063 ( .A(n2440), .B(n2439), .Z(n2467) );
  XOR U3064 ( .A(n2541), .B(n2449), .Z(n2439) );
  XNOR U3065 ( .A(n2436), .B(n2437), .Z(n2449) );
  NAND U3066 ( .A(n2328), .B(n1021), .Z(n2437) );
  XNOR U3067 ( .A(n2435), .B(n2542), .Z(n2436) );
  ANDN U3068 ( .A(n2333), .B(n1023), .Z(n2542) );
  XOR U3069 ( .A(n2543), .B(n2544), .Z(n2435) );
  AND U3070 ( .A(n2545), .B(n2546), .Z(n2544) );
  XOR U3071 ( .A(n2547), .B(n2543), .Z(n2546) );
  XNOR U3072 ( .A(n2448), .B(n2438), .Z(n2541) );
  XOR U3073 ( .A(n2555), .B(n2446), .Z(n2551) );
  AND U3074 ( .A(n2556), .B(n946), .Z(n2446) );
  NAND U3075 ( .A(n2557), .B(n2445), .Z(n2555) );
  XOR U3076 ( .A(n2558), .B(n2559), .Z(n2445) );
  AND U3077 ( .A(n2560), .B(n2561), .Z(n2559) );
  XNOR U3078 ( .A(n2562), .B(n2558), .Z(n2561) );
  NANDN U3079 ( .B(n949), .A(n2563), .Z(n2557) );
  XNOR U3080 ( .A(n2457), .B(n2456), .Z(n2440) );
  XOR U3081 ( .A(n2564), .B(n2453), .Z(n2456) );
  XNOR U3082 ( .A(n2452), .B(n2565), .Z(n2453) );
  ANDN U3083 ( .A(n2134), .B(n1107), .Z(n2565) );
  AND U3084 ( .A(n2127), .B(n1105), .Z(n2454) );
  XNOR U3085 ( .A(n2460), .B(n2461), .Z(n2457) );
  NAND U3086 ( .A(n1932), .B(n1206), .Z(n2461) );
  XNOR U3087 ( .A(n2459), .B(n2572), .Z(n2460) );
  ANDN U3088 ( .A(n1937), .B(n1208), .Z(n2572) );
  XNOR U3089 ( .A(n2466), .B(n2462), .Z(n2540) );
  XOR U3090 ( .A(n2583), .B(n2584), .Z(n2579) );
  NANDN U3091 ( .B(n2585), .A(n2586), .Z(n2583) );
  XNOR U3092 ( .A(n2483), .B(n2482), .Z(n2464) );
  XOR U3093 ( .A(n2587), .B(n2491), .Z(n2482) );
  XNOR U3094 ( .A(n2476), .B(n2475), .Z(n2491) );
  XOR U3095 ( .A(n2588), .B(n2472), .Z(n2475) );
  XNOR U3096 ( .A(n2471), .B(n2589), .Z(n2472) );
  ANDN U3097 ( .A(n1426), .B(n1640), .Z(n2589) );
  AND U3098 ( .A(n1638), .B(n1363), .Z(n2473) );
  XNOR U3099 ( .A(n2479), .B(n2480), .Z(n2476) );
  NANDN U3100 ( .B(n1228), .A(n1813), .Z(n2480) );
  XNOR U3101 ( .A(n2478), .B(n2596), .Z(n2479) );
  ANDN U3102 ( .A(n1298), .B(n1815), .Z(n2596) );
  XNOR U3103 ( .A(n2490), .B(n2481), .Z(n2587) );
  XOR U3104 ( .A(n2603), .B(n2499), .Z(n2490) );
  XNOR U3105 ( .A(n2487), .B(n2488), .Z(n2499) );
  NAND U3106 ( .A(n1479), .B(n1597), .Z(n2488) );
  XNOR U3107 ( .A(n2486), .B(n2604), .Z(n2487) );
  ANDN U3108 ( .A(n1604), .B(n1481), .Z(n2604) );
  XNOR U3109 ( .A(n2498), .B(n2489), .Z(n2603) );
  XOR U3110 ( .A(n2611), .B(n2495), .Z(n2498) );
  XNOR U3111 ( .A(n2494), .B(n2612), .Z(n2495) );
  ANDN U3112 ( .A(n1788), .B(n1340), .Z(n2612) );
  AND U3113 ( .A(n1338), .B(n1781), .Z(n2496) );
  XNOR U3114 ( .A(n2507), .B(n2506), .Z(n2483) );
  XOR U3115 ( .A(n2619), .B(n2515), .Z(n2506) );
  XNOR U3116 ( .A(n2503), .B(n2504), .Z(n2515) );
  NANDN U3117 ( .B(n1041), .A(n2203), .Z(n2504) );
  XNOR U3118 ( .A(n2502), .B(n2620), .Z(n2503) );
  ANDN U3119 ( .A(n1082), .B(n2205), .Z(n2620) );
  XNOR U3120 ( .A(n2514), .B(n2505), .Z(n2619) );
  XOR U3121 ( .A(n2627), .B(n2511), .Z(n2514) );
  XNOR U3122 ( .A(n2510), .B(n2628), .Z(n2511) );
  ANDN U3123 ( .A(n1189), .B(n2008), .Z(n2628) );
  AND U3124 ( .A(n2006), .B(n1135), .Z(n2512) );
  XOR U3125 ( .A(n2523), .B(n2522), .Z(n2507) );
  XOR U3126 ( .A(n2635), .B(n2519), .Z(n2522) );
  XNOR U3127 ( .A(n2518), .B(n2636), .Z(n2519) );
  ANDN U3128 ( .A(n1014), .B(n2418), .Z(n2636) );
  AND U3129 ( .A(n2416), .B(n973), .Z(n2520) );
  XOR U3130 ( .A(n2530), .B(n2529), .Z(n2523) );
  NAND U3131 ( .A(n2643), .B(n917), .Z(n2529) );
  XNOR U3132 ( .A(n2528), .B(n2644), .Z(n2530) );
  ANDN U3133 ( .A(n948), .B(n2645), .Z(n2644) );
  NAND U3134 ( .A(n2646), .B(n2647), .Z(n2528) );
  NAND U3135 ( .A(n2648), .B(n2649), .Z(n2646) );
  IV U3136 ( .A(n2531), .Z(n2532) );
  MUX U3137 ( .IN0(Y[5]), .IN1(n789), .SEL(n869), .F(n318) );
  XOR U3138 ( .A(n2654), .B(Y0[6]), .Z(n789) );
  XOR U3139 ( .A(n2655), .B(n2656), .Z(n2654) );
  AND U3140 ( .A(n881), .B(n2658), .Z(n2657) );
  XOR U3141 ( .A(n2652), .B(n2656), .Z(n2658) );
  XOR U3142 ( .A(n2651), .B(n2656), .Z(n2652) );
  XNOR U3143 ( .A(n2659), .B(n2582), .Z(n2577) );
  XNOR U3144 ( .A(n2550), .B(n2549), .Z(n2582) );
  XOR U3145 ( .A(n2660), .B(n2554), .Z(n2549) );
  XNOR U3146 ( .A(n2545), .B(n2547), .Z(n2554) );
  NAND U3147 ( .A(n2328), .B(n1061), .Z(n2547) );
  XNOR U3148 ( .A(n2543), .B(n2661), .Z(n2545) );
  ANDN U3149 ( .A(n2333), .B(n1063), .Z(n2661) );
  XNOR U3150 ( .A(n2553), .B(n2548), .Z(n2660) );
  XOR U3151 ( .A(n2668), .B(n2560), .Z(n2553) );
  XNOR U3152 ( .A(n2558), .B(n2669), .Z(n2560) );
  ANDN U3153 ( .A(n2563), .B(n979), .Z(n2669) );
  XOR U3154 ( .A(n2670), .B(n2671), .Z(n2558) );
  AND U3155 ( .A(n2672), .B(n2673), .Z(n2671) );
  XNOR U3156 ( .A(n2674), .B(n2670), .Z(n2673) );
  AND U3157 ( .A(n2556), .B(n977), .Z(n2562) );
  XNOR U3158 ( .A(n2571), .B(n2570), .Z(n2550) );
  XOR U3159 ( .A(n2678), .B(n2567), .Z(n2570) );
  XNOR U3160 ( .A(n2566), .B(n2679), .Z(n2567) );
  ANDN U3161 ( .A(n2134), .B(n1149), .Z(n2679) );
  AND U3162 ( .A(n2127), .B(n1147), .Z(n2568) );
  XNOR U3163 ( .A(n2574), .B(n2575), .Z(n2571) );
  NAND U3164 ( .A(n1932), .B(n1270), .Z(n2575) );
  XNOR U3165 ( .A(n2573), .B(n2686), .Z(n2574) );
  ANDN U3166 ( .A(n1937), .B(n1272), .Z(n2686) );
  XNOR U3167 ( .A(n2581), .B(n2576), .Z(n2659) );
  XOR U3168 ( .A(n2580), .B(n2693), .Z(n2581) );
  AND U3169 ( .A(n2584), .B(n2694), .Z(n2693) );
  AND U3170 ( .A(n2695), .B(n2696), .Z(n2694) );
  NANDN U3171 ( .B(n2697), .A(n916), .Z(n2696) );
  NAND U3172 ( .A(n2698), .B(n2699), .Z(n2695) );
  ANDN U3173 ( .A(n2586), .B(n2585), .Z(n2584) );
  ANDN U3174 ( .A(n2700), .B(n2701), .Z(n2585) );
  OR U3175 ( .A(n2702), .B(n2703), .Z(n2586) );
  XNOR U3176 ( .A(n2602), .B(n2601), .Z(n2578) );
  XOR U3177 ( .A(n2707), .B(n2610), .Z(n2601) );
  XNOR U3178 ( .A(n2595), .B(n2594), .Z(n2610) );
  XOR U3179 ( .A(n2708), .B(n2591), .Z(n2594) );
  XNOR U3180 ( .A(n2590), .B(n2709), .Z(n2591) );
  ANDN U3181 ( .A(n1426), .B(n1724), .Z(n2709) );
  AND U3182 ( .A(n1722), .B(n1363), .Z(n2592) );
  XNOR U3183 ( .A(n2598), .B(n2599), .Z(n2595) );
  NANDN U3184 ( .B(n1228), .A(n1910), .Z(n2599) );
  XNOR U3185 ( .A(n2597), .B(n2716), .Z(n2598) );
  ANDN U3186 ( .A(n1298), .B(n1912), .Z(n2716) );
  XNOR U3187 ( .A(n2609), .B(n2600), .Z(n2707) );
  XOR U3188 ( .A(n2723), .B(n2618), .Z(n2609) );
  XNOR U3189 ( .A(n2606), .B(n2607), .Z(n2618) );
  NAND U3190 ( .A(n1557), .B(n1597), .Z(n2607) );
  XNOR U3191 ( .A(n2605), .B(n2724), .Z(n2606) );
  ANDN U3192 ( .A(n1604), .B(n1559), .Z(n2724) );
  XNOR U3193 ( .A(n2617), .B(n2608), .Z(n2723) );
  XOR U3194 ( .A(n2731), .B(n2614), .Z(n2617) );
  XNOR U3195 ( .A(n2613), .B(n2732), .Z(n2614) );
  ANDN U3196 ( .A(n1788), .B(n1407), .Z(n2732) );
  AND U3197 ( .A(n1405), .B(n1781), .Z(n2615) );
  XNOR U3198 ( .A(n2626), .B(n2625), .Z(n2602) );
  XOR U3199 ( .A(n2739), .B(n2634), .Z(n2625) );
  XNOR U3200 ( .A(n2622), .B(n2623), .Z(n2634) );
  NANDN U3201 ( .B(n1041), .A(n2309), .Z(n2623) );
  XNOR U3202 ( .A(n2621), .B(n2740), .Z(n2622) );
  ANDN U3203 ( .A(n1082), .B(n2311), .Z(n2740) );
  XNOR U3204 ( .A(n2633), .B(n2624), .Z(n2739) );
  XOR U3205 ( .A(n2747), .B(n2630), .Z(n2633) );
  XNOR U3206 ( .A(n2629), .B(n2748), .Z(n2630) );
  ANDN U3207 ( .A(n1189), .B(n2104), .Z(n2748) );
  AND U3208 ( .A(n2102), .B(n1135), .Z(n2631) );
  XOR U3209 ( .A(n2642), .B(n2641), .Z(n2626) );
  XOR U3210 ( .A(n2755), .B(n2638), .Z(n2641) );
  XNOR U3211 ( .A(n2637), .B(n2756), .Z(n2638) );
  ANDN U3212 ( .A(n1014), .B(n2526), .Z(n2756) );
  AND U3213 ( .A(n2524), .B(n973), .Z(n2639) );
  XOR U3214 ( .A(n2649), .B(n2648), .Z(n2642) );
  NAND U3215 ( .A(n2763), .B(n917), .Z(n2648) );
  XOR U3216 ( .A(n2647), .B(n2764), .Z(n2649) );
  ANDN U3217 ( .A(n948), .B(n2765), .Z(n2764) );
  ANDN U3218 ( .A(n2766), .B(n2767), .Z(n2647) );
  NAND U3219 ( .A(n2768), .B(n2769), .Z(n2766) );
  IV U3220 ( .A(n2650), .Z(n2651) );
  MUX U3221 ( .IN0(Y[4]), .IN1(n786), .SEL(n869), .F(n317) );
  XOR U3222 ( .A(n2774), .B(Y0[5]), .Z(n786) );
  XOR U3223 ( .A(n2775), .B(n2776), .Z(n2774) );
  AND U3224 ( .A(n881), .B(n2778), .Z(n2777) );
  XOR U3225 ( .A(n2772), .B(n2776), .Z(n2778) );
  XOR U3226 ( .A(n2771), .B(n2776), .Z(n2772) );
  XNOR U3227 ( .A(n2779), .B(n2706), .Z(n2691) );
  XNOR U3228 ( .A(n2667), .B(n2666), .Z(n2706) );
  XOR U3229 ( .A(n2780), .B(n2677), .Z(n2666) );
  XNOR U3230 ( .A(n2663), .B(n2664), .Z(n2677) );
  NAND U3231 ( .A(n2328), .B(n1105), .Z(n2664) );
  XNOR U3232 ( .A(n2662), .B(n2781), .Z(n2663) );
  ANDN U3233 ( .A(n2333), .B(n1107), .Z(n2781) );
  XNOR U3234 ( .A(n2676), .B(n2665), .Z(n2780) );
  XOR U3235 ( .A(n2788), .B(n2672), .Z(n2676) );
  XNOR U3236 ( .A(n2670), .B(n2789), .Z(n2672) );
  ANDN U3237 ( .A(n2563), .B(n1023), .Z(n2789) );
  XOR U3238 ( .A(n2790), .B(n2791), .Z(n2670) );
  AND U3239 ( .A(n2792), .B(n2793), .Z(n2791) );
  XNOR U3240 ( .A(n2794), .B(n2790), .Z(n2793) );
  AND U3241 ( .A(n2556), .B(n1021), .Z(n2674) );
  XNOR U3242 ( .A(n2685), .B(n2684), .Z(n2667) );
  XOR U3243 ( .A(n2798), .B(n2681), .Z(n2684) );
  XNOR U3244 ( .A(n2680), .B(n2799), .Z(n2681) );
  ANDN U3245 ( .A(n2134), .B(n1208), .Z(n2799) );
  AND U3246 ( .A(n2127), .B(n1206), .Z(n2682) );
  XNOR U3247 ( .A(n2688), .B(n2689), .Z(n2685) );
  NAND U3248 ( .A(n1932), .B(n1338), .Z(n2689) );
  XNOR U3249 ( .A(n2687), .B(n2806), .Z(n2688) );
  ANDN U3250 ( .A(n1937), .B(n1340), .Z(n2806) );
  XOR U3251 ( .A(n2705), .B(n2690), .Z(n2779) );
  XOR U3252 ( .A(n2813), .B(n2698), .Z(n2705) );
  XOR U3253 ( .A(n2817), .B(n2703), .Z(n2701) );
  NAND U3254 ( .A(n2818), .B(n946), .Z(n2703) );
  NAND U3255 ( .A(n2819), .B(n2702), .Z(n2817) );
  NANDN U3256 ( .B(n949), .A(n2823), .Z(n2819) );
  ANDN U3257 ( .A(n2824), .B(n2825), .Z(n2699) );
  XNOR U3258 ( .A(n2722), .B(n2721), .Z(n2692) );
  XOR U3259 ( .A(n2829), .B(n2730), .Z(n2721) );
  XNOR U3260 ( .A(n2715), .B(n2714), .Z(n2730) );
  XOR U3261 ( .A(n2830), .B(n2711), .Z(n2714) );
  XNOR U3262 ( .A(n2710), .B(n2831), .Z(n2711) );
  ANDN U3263 ( .A(n1426), .B(n1815), .Z(n2831) );
  AND U3264 ( .A(n1813), .B(n1363), .Z(n2712) );
  XNOR U3265 ( .A(n2718), .B(n2719), .Z(n2715) );
  NANDN U3266 ( .B(n1228), .A(n2006), .Z(n2719) );
  XNOR U3267 ( .A(n2717), .B(n2838), .Z(n2718) );
  ANDN U3268 ( .A(n1298), .B(n2008), .Z(n2838) );
  XNOR U3269 ( .A(n2729), .B(n2720), .Z(n2829) );
  XOR U3270 ( .A(n2845), .B(n2738), .Z(n2729) );
  XNOR U3271 ( .A(n2726), .B(n2727), .Z(n2738) );
  NAND U3272 ( .A(n1638), .B(n1597), .Z(n2727) );
  XNOR U3273 ( .A(n2725), .B(n2846), .Z(n2726) );
  ANDN U3274 ( .A(n1604), .B(n1640), .Z(n2846) );
  XNOR U3275 ( .A(n2737), .B(n2728), .Z(n2845) );
  XOR U3276 ( .A(n2853), .B(n2734), .Z(n2737) );
  XNOR U3277 ( .A(n2733), .B(n2854), .Z(n2734) );
  ANDN U3278 ( .A(n1788), .B(n1481), .Z(n2854) );
  AND U3279 ( .A(n1479), .B(n1781), .Z(n2735) );
  XNOR U3280 ( .A(n2746), .B(n2745), .Z(n2722) );
  XOR U3281 ( .A(n2861), .B(n2754), .Z(n2745) );
  XNOR U3282 ( .A(n2742), .B(n2743), .Z(n2754) );
  NANDN U3283 ( .B(n1041), .A(n2416), .Z(n2743) );
  XNOR U3284 ( .A(n2741), .B(n2862), .Z(n2742) );
  ANDN U3285 ( .A(n1082), .B(n2418), .Z(n2862) );
  XNOR U3286 ( .A(n2753), .B(n2744), .Z(n2861) );
  XOR U3287 ( .A(n2869), .B(n2750), .Z(n2753) );
  XNOR U3288 ( .A(n2749), .B(n2870), .Z(n2750) );
  ANDN U3289 ( .A(n1189), .B(n2205), .Z(n2870) );
  AND U3290 ( .A(n2203), .B(n1135), .Z(n2751) );
  XOR U3291 ( .A(n2762), .B(n2761), .Z(n2746) );
  XOR U3292 ( .A(n2877), .B(n2758), .Z(n2761) );
  XNOR U3293 ( .A(n2757), .B(n2878), .Z(n2758) );
  ANDN U3294 ( .A(n1014), .B(n2645), .Z(n2878) );
  AND U3295 ( .A(n2643), .B(n973), .Z(n2759) );
  XOR U3296 ( .A(n2769), .B(n2768), .Z(n2762) );
  NAND U3297 ( .A(n2885), .B(n917), .Z(n2768) );
  XNOR U3298 ( .A(n2767), .B(n2886), .Z(n2769) );
  ANDN U3299 ( .A(n948), .B(n2887), .Z(n2886) );
  NAND U3300 ( .A(n2888), .B(n2889), .Z(n2767) );
  NAND U3301 ( .A(n2890), .B(n2891), .Z(n2888) );
  IV U3302 ( .A(n2770), .Z(n2771) );
  MUX U3303 ( .IN0(Y[3]), .IN1(n783), .SEL(n869), .F(n316) );
  XNOR U3304 ( .A(n2895), .B(Y0[4]), .Z(n783) );
  XNOR U3305 ( .A(n2897), .B(n2898), .Z(n2895) );
  XOR U3306 ( .A(n2896), .B(n2899), .Z(n2897) );
  AND U3307 ( .A(n881), .B(n2900), .Z(n2899) );
  XNOR U3308 ( .A(n2893), .B(n2898), .Z(n2900) );
  XOR U3309 ( .A(n2898), .B(n2892), .Z(n2893) );
  NOR U3310 ( .A(n2901), .B(n2902), .Z(n2892) );
  XNOR U3311 ( .A(n2903), .B(n2828), .Z(n2811) );
  XNOR U3312 ( .A(n2787), .B(n2786), .Z(n2828) );
  XOR U3313 ( .A(n2904), .B(n2797), .Z(n2786) );
  XNOR U3314 ( .A(n2783), .B(n2784), .Z(n2797) );
  NAND U3315 ( .A(n2328), .B(n1147), .Z(n2784) );
  XNOR U3316 ( .A(n2782), .B(n2905), .Z(n2783) );
  ANDN U3317 ( .A(n2333), .B(n1149), .Z(n2905) );
  XNOR U3318 ( .A(n2796), .B(n2785), .Z(n2904) );
  XOR U3319 ( .A(n2912), .B(n2792), .Z(n2796) );
  XNOR U3320 ( .A(n2790), .B(n2913), .Z(n2792) );
  ANDN U3321 ( .A(n2563), .B(n1063), .Z(n2913) );
  AND U3322 ( .A(n2556), .B(n1061), .Z(n2794) );
  XNOR U3323 ( .A(n2805), .B(n2804), .Z(n2787) );
  XOR U3324 ( .A(n2920), .B(n2801), .Z(n2804) );
  XNOR U3325 ( .A(n2800), .B(n2921), .Z(n2801) );
  ANDN U3326 ( .A(n2134), .B(n1272), .Z(n2921) );
  AND U3327 ( .A(n2127), .B(n1270), .Z(n2802) );
  XNOR U3328 ( .A(n2808), .B(n2809), .Z(n2805) );
  NAND U3329 ( .A(n1932), .B(n1405), .Z(n2809) );
  XNOR U3330 ( .A(n2807), .B(n2928), .Z(n2808) );
  ANDN U3331 ( .A(n1937), .B(n1407), .Z(n2928) );
  XNOR U3332 ( .A(n2827), .B(n2810), .Z(n2903) );
  XOR U3333 ( .A(n2935), .B(n2825), .Z(n2827) );
  XOR U3334 ( .A(n2816), .B(n2815), .Z(n2825) );
  XNOR U3335 ( .A(n2814), .B(n2936), .Z(n2815) );
  AND U3336 ( .A(n2937), .B(n2938), .Z(n2936) );
  NANDN U3337 ( .B(n2939), .A(n916), .Z(n2938) );
  NANDN U3338 ( .B(n2940), .A(n2941), .Z(n2937) );
  XNOR U3339 ( .A(n2821), .B(n2822), .Z(n2816) );
  NAND U3340 ( .A(n2818), .B(n977), .Z(n2822) );
  XNOR U3341 ( .A(n2820), .B(n2945), .Z(n2821) );
  ANDN U3342 ( .A(n2823), .B(n979), .Z(n2945) );
  NOR U3343 ( .A(n2949), .B(n2950), .Z(n2824) );
  XNOR U3344 ( .A(n2844), .B(n2843), .Z(n2812) );
  XOR U3345 ( .A(n2954), .B(n2852), .Z(n2843) );
  XNOR U3346 ( .A(n2837), .B(n2836), .Z(n2852) );
  XOR U3347 ( .A(n2955), .B(n2833), .Z(n2836) );
  XNOR U3348 ( .A(n2832), .B(n2956), .Z(n2833) );
  ANDN U3349 ( .A(n1426), .B(n1912), .Z(n2956) );
  AND U3350 ( .A(n1910), .B(n1363), .Z(n2834) );
  XNOR U3351 ( .A(n2840), .B(n2841), .Z(n2837) );
  NANDN U3352 ( .B(n1228), .A(n2102), .Z(n2841) );
  XNOR U3353 ( .A(n2839), .B(n2963), .Z(n2840) );
  ANDN U3354 ( .A(n1298), .B(n2104), .Z(n2963) );
  XNOR U3355 ( .A(n2851), .B(n2842), .Z(n2954) );
  XOR U3356 ( .A(n2970), .B(n2860), .Z(n2851) );
  XNOR U3357 ( .A(n2848), .B(n2849), .Z(n2860) );
  NAND U3358 ( .A(n1722), .B(n1597), .Z(n2849) );
  XNOR U3359 ( .A(n2847), .B(n2971), .Z(n2848) );
  ANDN U3360 ( .A(n1604), .B(n1724), .Z(n2971) );
  XNOR U3361 ( .A(n2859), .B(n2850), .Z(n2970) );
  XOR U3362 ( .A(n2978), .B(n2856), .Z(n2859) );
  XNOR U3363 ( .A(n2855), .B(n2979), .Z(n2856) );
  ANDN U3364 ( .A(n1788), .B(n1559), .Z(n2979) );
  AND U3365 ( .A(n1557), .B(n1781), .Z(n2857) );
  XNOR U3366 ( .A(n2868), .B(n2867), .Z(n2844) );
  XOR U3367 ( .A(n2986), .B(n2876), .Z(n2867) );
  XNOR U3368 ( .A(n2864), .B(n2865), .Z(n2876) );
  NANDN U3369 ( .B(n1041), .A(n2524), .Z(n2865) );
  XNOR U3370 ( .A(n2863), .B(n2987), .Z(n2864) );
  ANDN U3371 ( .A(n1082), .B(n2526), .Z(n2987) );
  XNOR U3372 ( .A(n2875), .B(n2866), .Z(n2986) );
  XOR U3373 ( .A(n2994), .B(n2872), .Z(n2875) );
  XNOR U3374 ( .A(n2871), .B(n2995), .Z(n2872) );
  ANDN U3375 ( .A(n1189), .B(n2311), .Z(n2995) );
  AND U3376 ( .A(n2309), .B(n1135), .Z(n2873) );
  XOR U3377 ( .A(n2884), .B(n2883), .Z(n2868) );
  XOR U3378 ( .A(n3002), .B(n2880), .Z(n2883) );
  XNOR U3379 ( .A(n2879), .B(n3003), .Z(n2880) );
  ANDN U3380 ( .A(n1014), .B(n2765), .Z(n3003) );
  AND U3381 ( .A(n2763), .B(n973), .Z(n2881) );
  XOR U3382 ( .A(n2891), .B(n2890), .Z(n2884) );
  NAND U3383 ( .A(n3010), .B(n917), .Z(n2890) );
  XOR U3384 ( .A(n2889), .B(n3011), .Z(n2891) );
  ANDN U3385 ( .A(n948), .B(n3012), .Z(n3011) );
  ANDN U3386 ( .A(n3013), .B(n3014), .Z(n2889) );
  NAND U3387 ( .A(n3015), .B(n3016), .Z(n3013) );
  IV U3388 ( .A(n2894), .Z(n2896) );
  MUX U3389 ( .IN0(Y[2]), .IN1(n780), .SEL(n869), .F(n315) );
  IV U3390 ( .A(n3020), .Z(n869) );
  XNOR U3391 ( .A(n3018), .B(Y0[3]), .Z(n780) );
  XNOR U3392 ( .A(n3021), .B(n3022), .Z(n3018) );
  XOR U3393 ( .A(n3019), .B(n3023), .Z(n3021) );
  AND U3394 ( .A(n881), .B(n3024), .Z(n3023) );
  XNOR U3395 ( .A(n2902), .B(n3022), .Z(n3024) );
  NANDN U3396 ( .B(n3025), .A(n3026), .Z(n2901) );
  XNOR U3397 ( .A(n3027), .B(n2953), .Z(n2933) );
  XNOR U3398 ( .A(n2911), .B(n2910), .Z(n2953) );
  XOR U3399 ( .A(n3028), .B(n2919), .Z(n2910) );
  XNOR U3400 ( .A(n2907), .B(n2908), .Z(n2919) );
  NAND U3401 ( .A(n2328), .B(n1206), .Z(n2908) );
  XNOR U3402 ( .A(n2906), .B(n3029), .Z(n2907) );
  ANDN U3403 ( .A(n2333), .B(n1208), .Z(n3029) );
  XNOR U3404 ( .A(n2918), .B(n2909), .Z(n3028) );
  XOR U3405 ( .A(n3036), .B(n2915), .Z(n2918) );
  XNOR U3406 ( .A(n2914), .B(n3037), .Z(n2915) );
  ANDN U3407 ( .A(n2563), .B(n1107), .Z(n3037) );
  AND U3408 ( .A(n2556), .B(n1105), .Z(n2916) );
  XNOR U3409 ( .A(n2927), .B(n2926), .Z(n2911) );
  XOR U3410 ( .A(n3044), .B(n2923), .Z(n2926) );
  XNOR U3411 ( .A(n2922), .B(n3045), .Z(n2923) );
  ANDN U3412 ( .A(n2134), .B(n1340), .Z(n3045) );
  AND U3413 ( .A(n2127), .B(n1338), .Z(n2924) );
  XNOR U3414 ( .A(n2930), .B(n2931), .Z(n2927) );
  NAND U3415 ( .A(n1932), .B(n1479), .Z(n2931) );
  XNOR U3416 ( .A(n2929), .B(n3052), .Z(n2930) );
  ANDN U3417 ( .A(n1937), .B(n1481), .Z(n3052) );
  XNOR U3418 ( .A(n2952), .B(n2932), .Z(n3027) );
  XOR U3419 ( .A(n3059), .B(n2950), .Z(n2952) );
  XOR U3420 ( .A(n2944), .B(n2943), .Z(n2950) );
  XOR U3421 ( .A(n3064), .B(n2941), .Z(n3060) );
  AND U3422 ( .A(n3065), .B(n946), .Z(n2941) );
  NAND U3423 ( .A(n3066), .B(n2940), .Z(n3064) );
  XOR U3424 ( .A(n3067), .B(n3068), .Z(n2940) );
  AND U3425 ( .A(n3069), .B(n3070), .Z(n3068) );
  XNOR U3426 ( .A(n3071), .B(n3067), .Z(n3070) );
  NANDN U3427 ( .B(n949), .A(n3072), .Z(n3066) );
  XNOR U3428 ( .A(n2947), .B(n2948), .Z(n2944) );
  NAND U3429 ( .A(n2818), .B(n1021), .Z(n2948) );
  XNOR U3430 ( .A(n2946), .B(n3073), .Z(n2947) );
  ANDN U3431 ( .A(n2823), .B(n1023), .Z(n3073) );
  XOR U3432 ( .A(n3074), .B(n3075), .Z(n2946) );
  AND U3433 ( .A(n3076), .B(n3077), .Z(n3075) );
  XOR U3434 ( .A(n3078), .B(n3074), .Z(n3077) );
  XNOR U3435 ( .A(n2949), .B(n2951), .Z(n3059) );
  XNOR U3436 ( .A(n3082), .B(n3085), .Z(n3084) );
  XNOR U3437 ( .A(n2969), .B(n2968), .Z(n2934) );
  XOR U3438 ( .A(n3086), .B(n2977), .Z(n2968) );
  XNOR U3439 ( .A(n2962), .B(n2961), .Z(n2977) );
  XOR U3440 ( .A(n3087), .B(n2958), .Z(n2961) );
  XNOR U3441 ( .A(n2957), .B(n3088), .Z(n2958) );
  ANDN U3442 ( .A(n1426), .B(n2008), .Z(n3088) );
  AND U3443 ( .A(n2006), .B(n1363), .Z(n2959) );
  XNOR U3444 ( .A(n2965), .B(n2966), .Z(n2962) );
  NANDN U3445 ( .B(n1228), .A(n2203), .Z(n2966) );
  XNOR U3446 ( .A(n2964), .B(n3095), .Z(n2965) );
  ANDN U3447 ( .A(n1298), .B(n2205), .Z(n3095) );
  XNOR U3448 ( .A(n2976), .B(n2967), .Z(n3086) );
  XOR U3449 ( .A(n3102), .B(n2985), .Z(n2976) );
  XNOR U3450 ( .A(n2973), .B(n2974), .Z(n2985) );
  NAND U3451 ( .A(n1813), .B(n1597), .Z(n2974) );
  XNOR U3452 ( .A(n2972), .B(n3103), .Z(n2973) );
  ANDN U3453 ( .A(n1604), .B(n1815), .Z(n3103) );
  XNOR U3454 ( .A(n2984), .B(n2975), .Z(n3102) );
  XOR U3455 ( .A(n3110), .B(n2981), .Z(n2984) );
  XNOR U3456 ( .A(n2980), .B(n3111), .Z(n2981) );
  ANDN U3457 ( .A(n1788), .B(n1640), .Z(n3111) );
  AND U3458 ( .A(n1638), .B(n1781), .Z(n2982) );
  XNOR U3459 ( .A(n2993), .B(n2992), .Z(n2969) );
  XOR U3460 ( .A(n3118), .B(n3001), .Z(n2992) );
  XNOR U3461 ( .A(n2989), .B(n2990), .Z(n3001) );
  NANDN U3462 ( .B(n1041), .A(n2643), .Z(n2990) );
  XNOR U3463 ( .A(n2988), .B(n3119), .Z(n2989) );
  ANDN U3464 ( .A(n1082), .B(n2645), .Z(n3119) );
  XNOR U3465 ( .A(n3000), .B(n2991), .Z(n3118) );
  XOR U3466 ( .A(n3126), .B(n2997), .Z(n3000) );
  XNOR U3467 ( .A(n2996), .B(n3127), .Z(n2997) );
  ANDN U3468 ( .A(n1189), .B(n2418), .Z(n3127) );
  AND U3469 ( .A(n2416), .B(n1135), .Z(n2998) );
  XOR U3470 ( .A(n3009), .B(n3008), .Z(n2993) );
  XOR U3471 ( .A(n3134), .B(n3005), .Z(n3008) );
  XNOR U3472 ( .A(n3004), .B(n3135), .Z(n3005) );
  ANDN U3473 ( .A(n1014), .B(n2887), .Z(n3135) );
  AND U3474 ( .A(n2885), .B(n973), .Z(n3006) );
  XOR U3475 ( .A(n3016), .B(n3015), .Z(n3009) );
  NAND U3476 ( .A(n3142), .B(n917), .Z(n3015) );
  XNOR U3477 ( .A(n3014), .B(n3143), .Z(n3016) );
  ANDN U3478 ( .A(n948), .B(n3144), .Z(n3143) );
  NAND U3479 ( .A(n3145), .B(n3146), .Z(n3014) );
  NAND U3480 ( .A(n3147), .B(n3148), .Z(n3145) );
  IV U3481 ( .A(n3017), .Z(n3019) );
  MUX U3482 ( .IN0(n777), .IN1(Y[1]), .SEL(n3020), .F(n314) );
  XNOR U3483 ( .A(n3150), .B(Y0[2]), .Z(n777) );
  XNOR U3484 ( .A(n3151), .B(n3152), .Z(n3150) );
  XNOR U3485 ( .A(n3149), .B(n3153), .Z(n3151) );
  AND U3486 ( .A(n881), .B(n3154), .Z(n3153) );
  XNOR U3487 ( .A(n3025), .B(n3152), .Z(n3154) );
  XOR U3488 ( .A(n3152), .B(n3026), .Z(n3025) );
  ANDN U3489 ( .A(n3155), .B(n3156), .Z(n3026) );
  XNOR U3490 ( .A(n3157), .B(n3081), .Z(n3057) );
  XNOR U3491 ( .A(n3035), .B(n3034), .Z(n3081) );
  XOR U3492 ( .A(n3158), .B(n3043), .Z(n3034) );
  XNOR U3493 ( .A(n3031), .B(n3032), .Z(n3043) );
  NAND U3494 ( .A(n2328), .B(n1270), .Z(n3032) );
  XNOR U3495 ( .A(n3030), .B(n3159), .Z(n3031) );
  ANDN U3496 ( .A(n2333), .B(n1272), .Z(n3159) );
  XNOR U3497 ( .A(n3042), .B(n3033), .Z(n3158) );
  XOR U3498 ( .A(n3166), .B(n3039), .Z(n3042) );
  XNOR U3499 ( .A(n3038), .B(n3167), .Z(n3039) );
  ANDN U3500 ( .A(n2563), .B(n1149), .Z(n3167) );
  AND U3501 ( .A(n2556), .B(n1147), .Z(n3040) );
  XNOR U3502 ( .A(n3051), .B(n3050), .Z(n3035) );
  XOR U3503 ( .A(n3174), .B(n3047), .Z(n3050) );
  XNOR U3504 ( .A(n3046), .B(n3175), .Z(n3047) );
  ANDN U3505 ( .A(n2134), .B(n1407), .Z(n3175) );
  AND U3506 ( .A(n2127), .B(n1405), .Z(n3048) );
  XNOR U3507 ( .A(n3054), .B(n3055), .Z(n3051) );
  NAND U3508 ( .A(n1932), .B(n1557), .Z(n3055) );
  XNOR U3509 ( .A(n3053), .B(n3182), .Z(n3054) );
  ANDN U3510 ( .A(n1937), .B(n1559), .Z(n3182) );
  XOR U3511 ( .A(n3080), .B(n3056), .Z(n3157) );
  XNOR U3512 ( .A(n3189), .B(n3085), .Z(n3080) );
  XNOR U3513 ( .A(n3063), .B(n3062), .Z(n3085) );
  XOR U3514 ( .A(n3190), .B(n3069), .Z(n3062) );
  XNOR U3515 ( .A(n3067), .B(n3191), .Z(n3069) );
  ANDN U3516 ( .A(n3072), .B(n979), .Z(n3191) );
  AND U3517 ( .A(n3065), .B(n977), .Z(n3071) );
  XNOR U3518 ( .A(n3076), .B(n3078), .Z(n3063) );
  NAND U3519 ( .A(n2818), .B(n1061), .Z(n3078) );
  XNOR U3520 ( .A(n3074), .B(n3198), .Z(n3076) );
  ANDN U3521 ( .A(n2823), .B(n1063), .Z(n3198) );
  XNOR U3522 ( .A(n3083), .B(n3079), .Z(n3189) );
  XOR U3523 ( .A(n3082), .B(n3205), .Z(n3083) );
  AND U3524 ( .A(n3206), .B(n3207), .Z(n3205) );
  NANDN U3525 ( .B(n3208), .A(n3209), .Z(n3207) );
  AND U3526 ( .A(n3210), .B(n3211), .Z(n3206) );
  NANDN U3527 ( .B(n3212), .A(n916), .Z(n3211) );
  OR U3528 ( .A(n3213), .B(n3214), .Z(n3210) );
  XNOR U3529 ( .A(n3101), .B(n3100), .Z(n3058) );
  XOR U3530 ( .A(n3218), .B(n3109), .Z(n3100) );
  XNOR U3531 ( .A(n3094), .B(n3093), .Z(n3109) );
  XOR U3532 ( .A(n3219), .B(n3090), .Z(n3093) );
  XNOR U3533 ( .A(n3089), .B(n3220), .Z(n3090) );
  ANDN U3534 ( .A(n1426), .B(n2104), .Z(n3220) );
  AND U3535 ( .A(n2102), .B(n1363), .Z(n3091) );
  XNOR U3536 ( .A(n3097), .B(n3098), .Z(n3094) );
  NANDN U3537 ( .B(n1228), .A(n2309), .Z(n3098) );
  XNOR U3538 ( .A(n3096), .B(n3227), .Z(n3097) );
  ANDN U3539 ( .A(n1298), .B(n2311), .Z(n3227) );
  XNOR U3540 ( .A(n3108), .B(n3099), .Z(n3218) );
  XOR U3541 ( .A(n3234), .B(n3117), .Z(n3108) );
  XNOR U3542 ( .A(n3105), .B(n3106), .Z(n3117) );
  NAND U3543 ( .A(n1910), .B(n1597), .Z(n3106) );
  XNOR U3544 ( .A(n3104), .B(n3235), .Z(n3105) );
  ANDN U3545 ( .A(n1604), .B(n1912), .Z(n3235) );
  XNOR U3546 ( .A(n3116), .B(n3107), .Z(n3234) );
  XOR U3547 ( .A(n3242), .B(n3113), .Z(n3116) );
  XNOR U3548 ( .A(n3112), .B(n3243), .Z(n3113) );
  ANDN U3549 ( .A(n1788), .B(n1724), .Z(n3243) );
  AND U3550 ( .A(n1722), .B(n1781), .Z(n3114) );
  XNOR U3551 ( .A(n3125), .B(n3124), .Z(n3101) );
  XOR U3552 ( .A(n3250), .B(n3133), .Z(n3124) );
  XNOR U3553 ( .A(n3121), .B(n3122), .Z(n3133) );
  NANDN U3554 ( .B(n1041), .A(n2763), .Z(n3122) );
  XNOR U3555 ( .A(n3120), .B(n3251), .Z(n3121) );
  ANDN U3556 ( .A(n1082), .B(n2765), .Z(n3251) );
  XNOR U3557 ( .A(n3132), .B(n3123), .Z(n3250) );
  XOR U3558 ( .A(n3258), .B(n3129), .Z(n3132) );
  XNOR U3559 ( .A(n3128), .B(n3259), .Z(n3129) );
  ANDN U3560 ( .A(n1189), .B(n2526), .Z(n3259) );
  AND U3561 ( .A(n2524), .B(n1135), .Z(n3130) );
  XOR U3562 ( .A(n3141), .B(n3140), .Z(n3125) );
  XOR U3563 ( .A(n3266), .B(n3137), .Z(n3140) );
  XNOR U3564 ( .A(n3136), .B(n3267), .Z(n3137) );
  ANDN U3565 ( .A(n1014), .B(n3012), .Z(n3267) );
  AND U3566 ( .A(n3010), .B(n973), .Z(n3138) );
  XOR U3567 ( .A(n3148), .B(n3147), .Z(n3141) );
  NAND U3568 ( .A(n3274), .B(n917), .Z(n3147) );
  XOR U3569 ( .A(n3146), .B(n3275), .Z(n3148) );
  ANDN U3570 ( .A(n948), .B(n3276), .Z(n3275) );
  ANDN U3571 ( .A(n3277), .B(n3278), .Z(n3146) );
  NAND U3572 ( .A(n3279), .B(n3280), .Z(n3277) );
  MUX U3573 ( .IN0(n773), .IN1(Y[0]), .SEL(n3020), .F(n313) );
  NANDN U3574 ( .B(rst), .A(n868), .Z(n3020) );
  AND U3575 ( .A(n3283), .B(n3284), .Z(n868) );
  AND U3576 ( .A(n3285), .B(n3286), .Z(n3284) );
  ANDN U3577 ( .A(n3287), .B(n[3]), .Z(n3286) );
  NOR U3578 ( .A(n[8]), .B(n[9]), .Z(n3287) );
  ANDN U3579 ( .A(n3288), .B(n[13]), .Z(n3285) );
  NOR U3580 ( .A(n[1]), .B(n[2]), .Z(n3288) );
  AND U3581 ( .A(n3289), .B(n3290), .Z(n3283) );
  AND U3582 ( .A(n765), .B(n3291), .Z(n3290) );
  NOR U3583 ( .A(n[0]), .B(n[10]), .Z(n3291) );
  NOR U3584 ( .A(n[6]), .B(n[7]), .Z(n765) );
  AND U3585 ( .A(n763), .B(n766), .Z(n3289) );
  NOR U3586 ( .A(n[4]), .B(n[5]), .Z(n766) );
  NOR U3587 ( .A(n[12]), .B(n[11]), .Z(n763) );
  XOR U3588 ( .A(n3282), .B(Y0[1]), .Z(n773) );
  XOR U3589 ( .A(n3292), .B(n3293), .Z(n3282) );
  XOR U3590 ( .A(n3294), .B(n3281), .Z(n3292) );
  NAND U3591 ( .A(n3295), .B(n881), .Z(n3294) );
  XOR U3592 ( .A(A[31]), .B(X[31]), .Z(n881) );
  XOR U3593 ( .A(n3155), .B(n3293), .Z(n3295) );
  XOR U3594 ( .A(n3156), .B(n3293), .Z(n3155) );
  XNOR U3595 ( .A(n3296), .B(n3204), .Z(n3187) );
  XNOR U3596 ( .A(n3165), .B(n3164), .Z(n3204) );
  XOR U3597 ( .A(n3297), .B(n3173), .Z(n3164) );
  XNOR U3598 ( .A(n3161), .B(n3162), .Z(n3173) );
  NAND U3599 ( .A(n2328), .B(n1338), .Z(n3162) );
  XNOR U3600 ( .A(n3160), .B(n3298), .Z(n3161) );
  ANDN U3601 ( .A(n2333), .B(n1340), .Z(n3298) );
  XNOR U3602 ( .A(n3172), .B(n3163), .Z(n3297) );
  XOR U3603 ( .A(n3305), .B(n3169), .Z(n3172) );
  XNOR U3604 ( .A(n3168), .B(n3306), .Z(n3169) );
  ANDN U3605 ( .A(n2563), .B(n1208), .Z(n3306) );
  AND U3606 ( .A(n2556), .B(n1206), .Z(n3170) );
  XNOR U3607 ( .A(n3181), .B(n3180), .Z(n3165) );
  XOR U3608 ( .A(n3313), .B(n3177), .Z(n3180) );
  XNOR U3609 ( .A(n3176), .B(n3314), .Z(n3177) );
  ANDN U3610 ( .A(n2134), .B(n1481), .Z(n3314) );
  AND U3611 ( .A(n2127), .B(n1479), .Z(n3178) );
  XNOR U3612 ( .A(n3184), .B(n3185), .Z(n3181) );
  NAND U3613 ( .A(n1932), .B(n1638), .Z(n3185) );
  XNOR U3614 ( .A(n3183), .B(n3321), .Z(n3184) );
  ANDN U3615 ( .A(n1937), .B(n1640), .Z(n3321) );
  XOR U3616 ( .A(n3203), .B(n3186), .Z(n3296) );
  XNOR U3617 ( .A(n3328), .B(n3217), .Z(n3203) );
  XNOR U3618 ( .A(n3197), .B(n3196), .Z(n3217) );
  XOR U3619 ( .A(n3329), .B(n3193), .Z(n3196) );
  XNOR U3620 ( .A(n3192), .B(n3330), .Z(n3193) );
  ANDN U3621 ( .A(n3072), .B(n1023), .Z(n3330) );
  AND U3622 ( .A(n3065), .B(n1021), .Z(n3194) );
  XNOR U3623 ( .A(n3200), .B(n3201), .Z(n3197) );
  NAND U3624 ( .A(n2818), .B(n1105), .Z(n3201) );
  XNOR U3625 ( .A(n3199), .B(n3337), .Z(n3200) );
  ANDN U3626 ( .A(n2823), .B(n1107), .Z(n3337) );
  XOR U3627 ( .A(n3216), .B(n3202), .Z(n3328) );
  XNOR U3628 ( .A(n3344), .B(n3213), .Z(n3216) );
  XNOR U3629 ( .A(n3345), .B(n3209), .Z(n3213) );
  AND U3630 ( .A(n3346), .B(n946), .Z(n3209) );
  NAND U3631 ( .A(n3347), .B(n3208), .Z(n3345) );
  NANDN U3632 ( .B(n949), .A(n3351), .Z(n3347) );
  XNOR U3633 ( .A(n3214), .B(n3215), .Z(n3344) );
  XNOR U3634 ( .A(n3355), .B(n3358), .Z(n3357) );
  XNOR U3635 ( .A(n3233), .B(n3232), .Z(n3188) );
  XOR U3636 ( .A(n3359), .B(n3241), .Z(n3232) );
  XNOR U3637 ( .A(n3226), .B(n3225), .Z(n3241) );
  XOR U3638 ( .A(n3360), .B(n3222), .Z(n3225) );
  XNOR U3639 ( .A(n3221), .B(n3361), .Z(n3222) );
  ANDN U3640 ( .A(n1426), .B(n2205), .Z(n3361) );
  AND U3641 ( .A(n2203), .B(n1363), .Z(n3223) );
  XNOR U3642 ( .A(n3229), .B(n3230), .Z(n3226) );
  NANDN U3643 ( .B(n1228), .A(n2416), .Z(n3230) );
  XNOR U3644 ( .A(n3228), .B(n3368), .Z(n3229) );
  ANDN U3645 ( .A(n1298), .B(n2418), .Z(n3368) );
  XNOR U3646 ( .A(n3240), .B(n3231), .Z(n3359) );
  XOR U3647 ( .A(n3375), .B(n3249), .Z(n3240) );
  XNOR U3648 ( .A(n3237), .B(n3238), .Z(n3249) );
  NAND U3649 ( .A(n2006), .B(n1597), .Z(n3238) );
  XNOR U3650 ( .A(n3236), .B(n3376), .Z(n3237) );
  ANDN U3651 ( .A(n1604), .B(n2008), .Z(n3376) );
  XNOR U3652 ( .A(n3248), .B(n3239), .Z(n3375) );
  XOR U3653 ( .A(n3383), .B(n3245), .Z(n3248) );
  XNOR U3654 ( .A(n3244), .B(n3384), .Z(n3245) );
  ANDN U3655 ( .A(n1788), .B(n1815), .Z(n3384) );
  AND U3656 ( .A(n1813), .B(n1781), .Z(n3246) );
  XNOR U3657 ( .A(n3257), .B(n3256), .Z(n3233) );
  XOR U3658 ( .A(n3391), .B(n3265), .Z(n3256) );
  XNOR U3659 ( .A(n3253), .B(n3254), .Z(n3265) );
  NANDN U3660 ( .B(n1041), .A(n2885), .Z(n3254) );
  XNOR U3661 ( .A(n3252), .B(n3392), .Z(n3253) );
  ANDN U3662 ( .A(n1082), .B(n2887), .Z(n3392) );
  XNOR U3663 ( .A(n3264), .B(n3255), .Z(n3391) );
  XOR U3664 ( .A(n3399), .B(n3261), .Z(n3264) );
  XNOR U3665 ( .A(n3260), .B(n3400), .Z(n3261) );
  ANDN U3666 ( .A(n1189), .B(n2645), .Z(n3400) );
  AND U3667 ( .A(n2643), .B(n1135), .Z(n3262) );
  XOR U3668 ( .A(n3273), .B(n3272), .Z(n3257) );
  XOR U3669 ( .A(n3407), .B(n3269), .Z(n3272) );
  XNOR U3670 ( .A(n3268), .B(n3408), .Z(n3269) );
  ANDN U3671 ( .A(n1014), .B(n3144), .Z(n3408) );
  AND U3672 ( .A(n3142), .B(n973), .Z(n3270) );
  XOR U3673 ( .A(n3280), .B(n3279), .Z(n3273) );
  NAND U3674 ( .A(n3415), .B(n917), .Z(n3279) );
  XNOR U3675 ( .A(n3278), .B(n3416), .Z(n3280) );
  ANDN U3676 ( .A(n948), .B(n3417), .Z(n3416) );
  NAND U3677 ( .A(n3418), .B(n3419), .Z(n3278) );
  NAND U3678 ( .A(n3420), .B(n3421), .Z(n3418) );
  XNOR U3679 ( .A(n3422), .B(n3343), .Z(n3326) );
  XNOR U3680 ( .A(n3304), .B(n3303), .Z(n3343) );
  XOR U3681 ( .A(n3423), .B(n3312), .Z(n3303) );
  XNOR U3682 ( .A(n3300), .B(n3301), .Z(n3312) );
  NAND U3683 ( .A(n2328), .B(n1405), .Z(n3301) );
  XNOR U3684 ( .A(n3299), .B(n3424), .Z(n3300) );
  ANDN U3685 ( .A(n2333), .B(n1407), .Z(n3424) );
  XOR U3686 ( .A(n3425), .B(n3426), .Z(n3299) );
  AND U3687 ( .A(n3427), .B(n3428), .Z(n3426) );
  XOR U3688 ( .A(n3429), .B(n3425), .Z(n3428) );
  XNOR U3689 ( .A(n3311), .B(n3302), .Z(n3423) );
  XOR U3690 ( .A(n3433), .B(n3308), .Z(n3311) );
  XNOR U3691 ( .A(n3307), .B(n3434), .Z(n3308) );
  ANDN U3692 ( .A(n2563), .B(n1272), .Z(n3434) );
  XOR U3693 ( .A(n3435), .B(n3436), .Z(n3307) );
  AND U3694 ( .A(n3437), .B(n3438), .Z(n3436) );
  XNOR U3695 ( .A(n3439), .B(n3435), .Z(n3438) );
  AND U3696 ( .A(n2556), .B(n1270), .Z(n3309) );
  XNOR U3697 ( .A(n3320), .B(n3319), .Z(n3304) );
  XOR U3698 ( .A(n3443), .B(n3316), .Z(n3319) );
  XNOR U3699 ( .A(n3315), .B(n3444), .Z(n3316) );
  ANDN U3700 ( .A(n2134), .B(n1559), .Z(n3444) );
  AND U3701 ( .A(n2127), .B(n1557), .Z(n3317) );
  XNOR U3702 ( .A(n3323), .B(n3324), .Z(n3320) );
  NAND U3703 ( .A(n1932), .B(n1722), .Z(n3324) );
  XNOR U3704 ( .A(n3322), .B(n3451), .Z(n3323) );
  ANDN U3705 ( .A(n1937), .B(n1724), .Z(n3451) );
  XNOR U3706 ( .A(n3342), .B(n3325), .Z(n3422) );
  XNOR U3707 ( .A(n3455), .B(n3456), .Z(n3325) );
  XNOR U3708 ( .A(n3457), .B(n3354), .Z(n3342) );
  XNOR U3709 ( .A(n3336), .B(n3335), .Z(n3354) );
  XOR U3710 ( .A(n3458), .B(n3332), .Z(n3335) );
  XNOR U3711 ( .A(n3331), .B(n3459), .Z(n3332) );
  ANDN U3712 ( .A(n3072), .B(n1063), .Z(n3459) );
  XOR U3713 ( .A(n3460), .B(n3461), .Z(n3331) );
  AND U3714 ( .A(n3462), .B(n3463), .Z(n3461) );
  XNOR U3715 ( .A(n3464), .B(n3460), .Z(n3463) );
  AND U3716 ( .A(n3065), .B(n1061), .Z(n3333) );
  XNOR U3717 ( .A(n3339), .B(n3340), .Z(n3336) );
  NAND U3718 ( .A(n2818), .B(n1147), .Z(n3340) );
  XNOR U3719 ( .A(n3338), .B(n3468), .Z(n3339) );
  ANDN U3720 ( .A(n2823), .B(n1149), .Z(n3468) );
  XOR U3721 ( .A(n3469), .B(n3470), .Z(n3338) );
  AND U3722 ( .A(n3471), .B(n3472), .Z(n3470) );
  XOR U3723 ( .A(n3473), .B(n3469), .Z(n3472) );
  XNOR U3724 ( .A(n3353), .B(n3341), .Z(n3457) );
  XOR U3725 ( .A(n3474), .B(n3475), .Z(n3341) );
  AND U3726 ( .A(n3476), .B(n3477), .Z(n3475) );
  XOR U3727 ( .A(n3478), .B(n3479), .Z(n3477) );
  XNOR U3728 ( .A(n3480), .B(n3474), .Z(n3478) );
  XNOR U3729 ( .A(n3431), .B(n3481), .Z(n3476) );
  XNOR U3730 ( .A(n3474), .B(n3432), .Z(n3481) );
  XNOR U3731 ( .A(n3450), .B(n3449), .Z(n3432) );
  XOR U3732 ( .A(n3482), .B(n3446), .Z(n3449) );
  XNOR U3733 ( .A(n3445), .B(n3483), .Z(n3446) );
  ANDN U3734 ( .A(n2134), .B(n1640), .Z(n3483) );
  AND U3735 ( .A(n2127), .B(n1638), .Z(n3447) );
  XNOR U3736 ( .A(n3453), .B(n3454), .Z(n3450) );
  NAND U3737 ( .A(n1813), .B(n1932), .Z(n3454) );
  XNOR U3738 ( .A(n3452), .B(n3490), .Z(n3453) );
  ANDN U3739 ( .A(n1937), .B(n1815), .Z(n3490) );
  XOR U3740 ( .A(n3494), .B(n3442), .Z(n3431) );
  XNOR U3741 ( .A(n3427), .B(n3429), .Z(n3442) );
  NAND U3742 ( .A(n2328), .B(n1479), .Z(n3429) );
  XNOR U3743 ( .A(n3425), .B(n3495), .Z(n3427) );
  ANDN U3744 ( .A(n2333), .B(n1481), .Z(n3495) );
  XNOR U3745 ( .A(n3441), .B(n3430), .Z(n3494) );
  XOR U3746 ( .A(n3502), .B(n3437), .Z(n3441) );
  XNOR U3747 ( .A(n3435), .B(n3503), .Z(n3437) );
  ANDN U3748 ( .A(n2563), .B(n1340), .Z(n3503) );
  XOR U3749 ( .A(n3504), .B(n3505), .Z(n3435) );
  AND U3750 ( .A(n3506), .B(n3507), .Z(n3505) );
  XNOR U3751 ( .A(n3508), .B(n3504), .Z(n3507) );
  AND U3752 ( .A(n2556), .B(n1338), .Z(n3439) );
  XOR U3753 ( .A(n3512), .B(n3513), .Z(n3474) );
  AND U3754 ( .A(n3514), .B(n3515), .Z(n3513) );
  XOR U3755 ( .A(n3516), .B(n3517), .Z(n3515) );
  XOR U3756 ( .A(n3512), .B(n3518), .Z(n3517) );
  XNOR U3757 ( .A(n3500), .B(n3519), .Z(n3514) );
  XNOR U3758 ( .A(n3512), .B(n3501), .Z(n3519) );
  XNOR U3759 ( .A(n3489), .B(n3488), .Z(n3501) );
  XOR U3760 ( .A(n3520), .B(n3485), .Z(n3488) );
  XNOR U3761 ( .A(n3484), .B(n3521), .Z(n3485) );
  ANDN U3762 ( .A(n2134), .B(n1724), .Z(n3521) );
  XOR U3763 ( .A(n3522), .B(n3523), .Z(n3484) );
  AND U3764 ( .A(n3524), .B(n3525), .Z(n3523) );
  XNOR U3765 ( .A(n3526), .B(n3522), .Z(n3525) );
  AND U3766 ( .A(n2127), .B(n1722), .Z(n3486) );
  XNOR U3767 ( .A(n3492), .B(n3493), .Z(n3489) );
  NAND U3768 ( .A(n1910), .B(n1932), .Z(n3493) );
  XNOR U3769 ( .A(n3491), .B(n3530), .Z(n3492) );
  ANDN U3770 ( .A(n1937), .B(n1912), .Z(n3530) );
  XOR U3771 ( .A(n3531), .B(n3532), .Z(n3491) );
  AND U3772 ( .A(n3533), .B(n3534), .Z(n3532) );
  XOR U3773 ( .A(n3535), .B(n3531), .Z(n3534) );
  XOR U3774 ( .A(n3536), .B(n3511), .Z(n3500) );
  XNOR U3775 ( .A(n3497), .B(n3498), .Z(n3511) );
  NAND U3776 ( .A(n2328), .B(n1557), .Z(n3498) );
  XNOR U3777 ( .A(n3496), .B(n3537), .Z(n3497) );
  ANDN U3778 ( .A(n2333), .B(n1559), .Z(n3537) );
  XOR U3779 ( .A(n3538), .B(n3539), .Z(n3496) );
  AND U3780 ( .A(n3540), .B(n3541), .Z(n3539) );
  XOR U3781 ( .A(n3542), .B(n3538), .Z(n3541) );
  XNOR U3782 ( .A(n3510), .B(n3499), .Z(n3536) );
  XOR U3783 ( .A(n3546), .B(n3506), .Z(n3510) );
  XNOR U3784 ( .A(n3504), .B(n3547), .Z(n3506) );
  ANDN U3785 ( .A(n2563), .B(n1407), .Z(n3547) );
  XOR U3786 ( .A(n3548), .B(n3549), .Z(n3504) );
  AND U3787 ( .A(n3550), .B(n3551), .Z(n3549) );
  XNOR U3788 ( .A(n3552), .B(n3548), .Z(n3551) );
  XOR U3789 ( .A(n3553), .B(n3508), .Z(n3546) );
  AND U3790 ( .A(n2556), .B(n1405), .Z(n3508) );
  IV U3791 ( .A(n3509), .Z(n3553) );
  XOR U3792 ( .A(n3557), .B(n3558), .Z(n3512) );
  AND U3793 ( .A(n3559), .B(n3560), .Z(n3558) );
  XOR U3794 ( .A(n3561), .B(n3562), .Z(n3560) );
  XOR U3795 ( .A(n3557), .B(n3563), .Z(n3562) );
  XNOR U3796 ( .A(n3544), .B(n3564), .Z(n3559) );
  XNOR U3797 ( .A(n3557), .B(n3545), .Z(n3564) );
  XNOR U3798 ( .A(n3529), .B(n3528), .Z(n3545) );
  XOR U3799 ( .A(n3565), .B(n3524), .Z(n3528) );
  XNOR U3800 ( .A(n3522), .B(n3566), .Z(n3524) );
  ANDN U3801 ( .A(n2134), .B(n1815), .Z(n3566) );
  XOR U3802 ( .A(n3567), .B(n3568), .Z(n3522) );
  AND U3803 ( .A(n3569), .B(n3570), .Z(n3568) );
  XNOR U3804 ( .A(n3571), .B(n3567), .Z(n3570) );
  AND U3805 ( .A(n1813), .B(n2127), .Z(n3526) );
  XNOR U3806 ( .A(n3533), .B(n3535), .Z(n3529) );
  NAND U3807 ( .A(n2006), .B(n1932), .Z(n3535) );
  XNOR U3808 ( .A(n3531), .B(n3575), .Z(n3533) );
  ANDN U3809 ( .A(n1937), .B(n2008), .Z(n3575) );
  XOR U3810 ( .A(n3579), .B(n3556), .Z(n3544) );
  XNOR U3811 ( .A(n3540), .B(n3542), .Z(n3556) );
  NAND U3812 ( .A(n2328), .B(n1638), .Z(n3542) );
  XNOR U3813 ( .A(n3538), .B(n3580), .Z(n3540) );
  ANDN U3814 ( .A(n2333), .B(n1640), .Z(n3580) );
  XOR U3815 ( .A(n3581), .B(n3582), .Z(n3538) );
  AND U3816 ( .A(n3583), .B(n3584), .Z(n3582) );
  XOR U3817 ( .A(n3585), .B(n3581), .Z(n3584) );
  XNOR U3818 ( .A(n3555), .B(n3543), .Z(n3579) );
  XOR U3819 ( .A(n3589), .B(n3550), .Z(n3555) );
  XNOR U3820 ( .A(n3548), .B(n3590), .Z(n3550) );
  ANDN U3821 ( .A(n2563), .B(n1481), .Z(n3590) );
  XOR U3822 ( .A(n3591), .B(n3592), .Z(n3548) );
  AND U3823 ( .A(n3593), .B(n3594), .Z(n3592) );
  XNOR U3824 ( .A(n3595), .B(n3591), .Z(n3594) );
  AND U3825 ( .A(n2556), .B(n1479), .Z(n3552) );
  XOR U3826 ( .A(n3599), .B(n3600), .Z(n3557) );
  AND U3827 ( .A(n3601), .B(n3602), .Z(n3600) );
  XOR U3828 ( .A(n3603), .B(n3604), .Z(n3602) );
  XOR U3829 ( .A(n3599), .B(n3605), .Z(n3604) );
  XNOR U3830 ( .A(n3587), .B(n3606), .Z(n3601) );
  XNOR U3831 ( .A(n3599), .B(n3588), .Z(n3606) );
  XNOR U3832 ( .A(n3574), .B(n3573), .Z(n3588) );
  XOR U3833 ( .A(n3607), .B(n3569), .Z(n3573) );
  XNOR U3834 ( .A(n3567), .B(n3608), .Z(n3569) );
  ANDN U3835 ( .A(n2134), .B(n1912), .Z(n3608) );
  XOR U3836 ( .A(n3609), .B(n3610), .Z(n3567) );
  AND U3837 ( .A(n3611), .B(n3612), .Z(n3610) );
  XNOR U3838 ( .A(n3613), .B(n3609), .Z(n3612) );
  AND U3839 ( .A(n1910), .B(n2127), .Z(n3571) );
  XNOR U3840 ( .A(n3577), .B(n3578), .Z(n3574) );
  NAND U3841 ( .A(n2102), .B(n1932), .Z(n3578) );
  XNOR U3842 ( .A(n3576), .B(n3617), .Z(n3577) );
  ANDN U3843 ( .A(n1937), .B(n2104), .Z(n3617) );
  XOR U3844 ( .A(n3618), .B(n3619), .Z(n3576) );
  AND U3845 ( .A(n3620), .B(n3621), .Z(n3619) );
  XOR U3846 ( .A(n3622), .B(n3618), .Z(n3621) );
  XOR U3847 ( .A(n3623), .B(n3598), .Z(n3587) );
  XNOR U3848 ( .A(n3583), .B(n3585), .Z(n3598) );
  NAND U3849 ( .A(n2328), .B(n1722), .Z(n3585) );
  XNOR U3850 ( .A(n3581), .B(n3624), .Z(n3583) );
  ANDN U3851 ( .A(n2333), .B(n1724), .Z(n3624) );
  XNOR U3852 ( .A(n3597), .B(n3586), .Z(n3623) );
  XOR U3853 ( .A(n3631), .B(n3593), .Z(n3597) );
  XNOR U3854 ( .A(n3591), .B(n3632), .Z(n3593) );
  ANDN U3855 ( .A(n2563), .B(n1559), .Z(n3632) );
  XOR U3856 ( .A(n3633), .B(n3634), .Z(n3591) );
  AND U3857 ( .A(n3635), .B(n3636), .Z(n3634) );
  XNOR U3858 ( .A(n3637), .B(n3633), .Z(n3636) );
  XOR U3859 ( .A(n3638), .B(n3595), .Z(n3631) );
  AND U3860 ( .A(n2556), .B(n1557), .Z(n3595) );
  IV U3861 ( .A(n3596), .Z(n3638) );
  XOR U3862 ( .A(n3642), .B(n3643), .Z(n3599) );
  AND U3863 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U3864 ( .A(n3646), .B(n3647), .Z(n3645) );
  XOR U3865 ( .A(n3642), .B(n3648), .Z(n3647) );
  XNOR U3866 ( .A(n3629), .B(n3649), .Z(n3644) );
  XNOR U3867 ( .A(n3642), .B(n3630), .Z(n3649) );
  XNOR U3868 ( .A(n3616), .B(n3615), .Z(n3630) );
  XOR U3869 ( .A(n3650), .B(n3611), .Z(n3615) );
  XNOR U3870 ( .A(n3609), .B(n3651), .Z(n3611) );
  ANDN U3871 ( .A(n2134), .B(n2008), .Z(n3651) );
  XOR U3872 ( .A(n3652), .B(n3653), .Z(n3609) );
  AND U3873 ( .A(n3654), .B(n3655), .Z(n3653) );
  XNOR U3874 ( .A(n3656), .B(n3652), .Z(n3655) );
  AND U3875 ( .A(n2006), .B(n2127), .Z(n3613) );
  XNOR U3876 ( .A(n3620), .B(n3622), .Z(n3616) );
  NAND U3877 ( .A(n2203), .B(n1932), .Z(n3622) );
  XNOR U3878 ( .A(n3618), .B(n3660), .Z(n3620) );
  ANDN U3879 ( .A(n1937), .B(n2205), .Z(n3660) );
  XOR U3880 ( .A(n3664), .B(n3641), .Z(n3629) );
  XNOR U3881 ( .A(n3626), .B(n3627), .Z(n3641) );
  NAND U3882 ( .A(n1813), .B(n2328), .Z(n3627) );
  XNOR U3883 ( .A(n3625), .B(n3665), .Z(n3626) );
  ANDN U3884 ( .A(n2333), .B(n1815), .Z(n3665) );
  XOR U3885 ( .A(n3666), .B(n3667), .Z(n3625) );
  AND U3886 ( .A(n3668), .B(n3669), .Z(n3667) );
  XOR U3887 ( .A(n3670), .B(n3666), .Z(n3669) );
  XNOR U3888 ( .A(n3640), .B(n3628), .Z(n3664) );
  XOR U3889 ( .A(n3674), .B(n3635), .Z(n3640) );
  XNOR U3890 ( .A(n3633), .B(n3675), .Z(n3635) );
  ANDN U3891 ( .A(n2563), .B(n1640), .Z(n3675) );
  XOR U3892 ( .A(n3676), .B(n3677), .Z(n3633) );
  AND U3893 ( .A(n3678), .B(n3679), .Z(n3677) );
  XNOR U3894 ( .A(n3680), .B(n3676), .Z(n3679) );
  AND U3895 ( .A(n2556), .B(n1638), .Z(n3637) );
  XOR U3896 ( .A(n3684), .B(n3685), .Z(n3642) );
  AND U3897 ( .A(n3686), .B(n3687), .Z(n3685) );
  XOR U3898 ( .A(n3688), .B(n3689), .Z(n3687) );
  XOR U3899 ( .A(n3684), .B(n3690), .Z(n3689) );
  XNOR U3900 ( .A(n3672), .B(n3691), .Z(n3686) );
  XNOR U3901 ( .A(n3684), .B(n3673), .Z(n3691) );
  XNOR U3902 ( .A(n3659), .B(n3658), .Z(n3673) );
  XOR U3903 ( .A(n3692), .B(n3654), .Z(n3658) );
  XNOR U3904 ( .A(n3652), .B(n3693), .Z(n3654) );
  ANDN U3905 ( .A(n2134), .B(n2104), .Z(n3693) );
  XOR U3906 ( .A(n3694), .B(n3695), .Z(n3652) );
  AND U3907 ( .A(n3696), .B(n3697), .Z(n3695) );
  XNOR U3908 ( .A(n3698), .B(n3694), .Z(n3697) );
  XOR U3909 ( .A(n3699), .B(n3656), .Z(n3692) );
  AND U3910 ( .A(n2102), .B(n2127), .Z(n3656) );
  IV U3911 ( .A(n3657), .Z(n3699) );
  XNOR U3912 ( .A(n3662), .B(n3663), .Z(n3659) );
  NAND U3913 ( .A(n2309), .B(n1932), .Z(n3663) );
  XNOR U3914 ( .A(n3661), .B(n3703), .Z(n3662) );
  ANDN U3915 ( .A(n1937), .B(n2311), .Z(n3703) );
  XOR U3916 ( .A(n3704), .B(n3705), .Z(n3661) );
  AND U3917 ( .A(n3706), .B(n3707), .Z(n3705) );
  XOR U3918 ( .A(n3708), .B(n3704), .Z(n3707) );
  XOR U3919 ( .A(n3709), .B(n3683), .Z(n3672) );
  XNOR U3920 ( .A(n3668), .B(n3670), .Z(n3683) );
  NAND U3921 ( .A(n1910), .B(n2328), .Z(n3670) );
  XNOR U3922 ( .A(n3666), .B(n3710), .Z(n3668) );
  ANDN U3923 ( .A(n2333), .B(n1912), .Z(n3710) );
  XOR U3924 ( .A(n3711), .B(n3712), .Z(n3666) );
  AND U3925 ( .A(n3713), .B(n3714), .Z(n3712) );
  XOR U3926 ( .A(n3715), .B(n3711), .Z(n3714) );
  XNOR U3927 ( .A(n3682), .B(n3671), .Z(n3709) );
  XOR U3928 ( .A(n3719), .B(n3678), .Z(n3682) );
  XNOR U3929 ( .A(n3676), .B(n3720), .Z(n3678) );
  ANDN U3930 ( .A(n2563), .B(n1724), .Z(n3720) );
  XOR U3931 ( .A(n3721), .B(n3722), .Z(n3676) );
  AND U3932 ( .A(n3723), .B(n3724), .Z(n3722) );
  XNOR U3933 ( .A(n3725), .B(n3721), .Z(n3724) );
  XOR U3934 ( .A(n3726), .B(n3680), .Z(n3719) );
  AND U3935 ( .A(n2556), .B(n1722), .Z(n3680) );
  IV U3936 ( .A(n3681), .Z(n3726) );
  XOR U3937 ( .A(n3730), .B(n3731), .Z(n3684) );
  AND U3938 ( .A(n3732), .B(n3733), .Z(n3731) );
  XOR U3939 ( .A(n3734), .B(n3735), .Z(n3733) );
  XOR U3940 ( .A(n3730), .B(n3736), .Z(n3735) );
  XNOR U3941 ( .A(n3717), .B(n3737), .Z(n3732) );
  XNOR U3942 ( .A(n3730), .B(n3718), .Z(n3737) );
  XNOR U3943 ( .A(n3702), .B(n3701), .Z(n3718) );
  XOR U3944 ( .A(n3738), .B(n3696), .Z(n3701) );
  XNOR U3945 ( .A(n3694), .B(n3739), .Z(n3696) );
  ANDN U3946 ( .A(n2134), .B(n2205), .Z(n3739) );
  XOR U3947 ( .A(n3740), .B(n3741), .Z(n3694) );
  AND U3948 ( .A(n3742), .B(n3743), .Z(n3741) );
  XNOR U3949 ( .A(n3744), .B(n3740), .Z(n3743) );
  XOR U3950 ( .A(n3745), .B(n3698), .Z(n3738) );
  AND U3951 ( .A(n2203), .B(n2127), .Z(n3698) );
  IV U3952 ( .A(n3700), .Z(n3745) );
  XNOR U3953 ( .A(n3706), .B(n3708), .Z(n3702) );
  NAND U3954 ( .A(n2416), .B(n1932), .Z(n3708) );
  XNOR U3955 ( .A(n3704), .B(n3749), .Z(n3706) );
  ANDN U3956 ( .A(n1937), .B(n2418), .Z(n3749) );
  XOR U3957 ( .A(n3750), .B(n3751), .Z(n3704) );
  AND U3958 ( .A(n3752), .B(n3753), .Z(n3751) );
  XOR U3959 ( .A(n3754), .B(n3750), .Z(n3753) );
  XOR U3960 ( .A(n3755), .B(n3729), .Z(n3717) );
  XNOR U3961 ( .A(n3713), .B(n3715), .Z(n3729) );
  NAND U3962 ( .A(n2006), .B(n2328), .Z(n3715) );
  XNOR U3963 ( .A(n3711), .B(n3756), .Z(n3713) );
  ANDN U3964 ( .A(n2333), .B(n2008), .Z(n3756) );
  XNOR U3965 ( .A(n3728), .B(n3716), .Z(n3755) );
  XOR U3966 ( .A(n3763), .B(n3723), .Z(n3728) );
  XNOR U3967 ( .A(n3721), .B(n3764), .Z(n3723) );
  ANDN U3968 ( .A(n2563), .B(n1815), .Z(n3764) );
  XOR U3969 ( .A(n3765), .B(n3766), .Z(n3721) );
  AND U3970 ( .A(n3767), .B(n3768), .Z(n3766) );
  XNOR U3971 ( .A(n3769), .B(n3765), .Z(n3768) );
  XOR U3972 ( .A(n3770), .B(n3725), .Z(n3763) );
  AND U3973 ( .A(n1813), .B(n2556), .Z(n3725) );
  IV U3974 ( .A(n3727), .Z(n3770) );
  XOR U3975 ( .A(n3774), .B(n3775), .Z(n3730) );
  AND U3976 ( .A(n3776), .B(n3777), .Z(n3775) );
  XOR U3977 ( .A(n3778), .B(n3779), .Z(n3777) );
  XOR U3978 ( .A(n3774), .B(n3780), .Z(n3779) );
  XNOR U3979 ( .A(n3761), .B(n3781), .Z(n3776) );
  XNOR U3980 ( .A(n3774), .B(n3762), .Z(n3781) );
  XNOR U3981 ( .A(n3748), .B(n3747), .Z(n3762) );
  XOR U3982 ( .A(n3782), .B(n3742), .Z(n3747) );
  XNOR U3983 ( .A(n3740), .B(n3783), .Z(n3742) );
  ANDN U3984 ( .A(n2134), .B(n2311), .Z(n3783) );
  XOR U3985 ( .A(n3784), .B(n3785), .Z(n3740) );
  AND U3986 ( .A(n3786), .B(n3787), .Z(n3785) );
  XNOR U3987 ( .A(n3788), .B(n3784), .Z(n3787) );
  XOR U3988 ( .A(n3789), .B(n3744), .Z(n3782) );
  AND U3989 ( .A(n2309), .B(n2127), .Z(n3744) );
  IV U3990 ( .A(n3746), .Z(n3789) );
  XNOR U3991 ( .A(n3752), .B(n3754), .Z(n3748) );
  NAND U3992 ( .A(n2524), .B(n1932), .Z(n3754) );
  XNOR U3993 ( .A(n3750), .B(n3793), .Z(n3752) );
  ANDN U3994 ( .A(n1937), .B(n2526), .Z(n3793) );
  XOR U3995 ( .A(n3794), .B(n3795), .Z(n3750) );
  AND U3996 ( .A(n3796), .B(n3797), .Z(n3795) );
  XOR U3997 ( .A(n3798), .B(n3794), .Z(n3797) );
  XOR U3998 ( .A(n3799), .B(n3773), .Z(n3761) );
  XNOR U3999 ( .A(n3758), .B(n3759), .Z(n3773) );
  NAND U4000 ( .A(n2102), .B(n2328), .Z(n3759) );
  XNOR U4001 ( .A(n3757), .B(n3800), .Z(n3758) );
  ANDN U4002 ( .A(n2333), .B(n2104), .Z(n3800) );
  XOR U4003 ( .A(n3801), .B(n3802), .Z(n3757) );
  AND U4004 ( .A(n3803), .B(n3804), .Z(n3802) );
  XOR U4005 ( .A(n3805), .B(n3801), .Z(n3804) );
  XNOR U4006 ( .A(n3772), .B(n3760), .Z(n3799) );
  XOR U4007 ( .A(n3809), .B(n3767), .Z(n3772) );
  XNOR U4008 ( .A(n3765), .B(n3810), .Z(n3767) );
  ANDN U4009 ( .A(n2563), .B(n1912), .Z(n3810) );
  XOR U4010 ( .A(n3811), .B(n3812), .Z(n3765) );
  AND U4011 ( .A(n3813), .B(n3814), .Z(n3812) );
  XNOR U4012 ( .A(n3815), .B(n3811), .Z(n3814) );
  XOR U4013 ( .A(n3816), .B(n3769), .Z(n3809) );
  AND U4014 ( .A(n1910), .B(n2556), .Z(n3769) );
  IV U4015 ( .A(n3771), .Z(n3816) );
  XOR U4016 ( .A(n3820), .B(n3821), .Z(n3774) );
  AND U4017 ( .A(n3822), .B(n3823), .Z(n3821) );
  XOR U4018 ( .A(n3824), .B(n3825), .Z(n3823) );
  XOR U4019 ( .A(n3820), .B(n3826), .Z(n3825) );
  XNOR U4020 ( .A(n3807), .B(n3827), .Z(n3822) );
  XNOR U4021 ( .A(n3820), .B(n3808), .Z(n3827) );
  XNOR U4022 ( .A(n3792), .B(n3791), .Z(n3808) );
  XOR U4023 ( .A(n3828), .B(n3786), .Z(n3791) );
  XNOR U4024 ( .A(n3784), .B(n3829), .Z(n3786) );
  ANDN U4025 ( .A(n2134), .B(n2418), .Z(n3829) );
  XOR U4026 ( .A(n3830), .B(n3831), .Z(n3784) );
  AND U4027 ( .A(n3832), .B(n3833), .Z(n3831) );
  XNOR U4028 ( .A(n3834), .B(n3830), .Z(n3833) );
  XOR U4029 ( .A(n3835), .B(n3788), .Z(n3828) );
  AND U4030 ( .A(n2416), .B(n2127), .Z(n3788) );
  IV U4031 ( .A(n3790), .Z(n3835) );
  XNOR U4032 ( .A(n3796), .B(n3798), .Z(n3792) );
  NAND U4033 ( .A(n2643), .B(n1932), .Z(n3798) );
  XNOR U4034 ( .A(n3794), .B(n3839), .Z(n3796) );
  ANDN U4035 ( .A(n1937), .B(n2645), .Z(n3839) );
  XOR U4036 ( .A(n3840), .B(n3841), .Z(n3794) );
  AND U4037 ( .A(n3842), .B(n3843), .Z(n3841) );
  XOR U4038 ( .A(n3844), .B(n3840), .Z(n3843) );
  XOR U4039 ( .A(n3845), .B(n3819), .Z(n3807) );
  XNOR U4040 ( .A(n3803), .B(n3805), .Z(n3819) );
  NAND U4041 ( .A(n2203), .B(n2328), .Z(n3805) );
  XNOR U4042 ( .A(n3801), .B(n3846), .Z(n3803) );
  ANDN U4043 ( .A(n2333), .B(n2205), .Z(n3846) );
  XOR U4044 ( .A(n3847), .B(n3848), .Z(n3801) );
  AND U4045 ( .A(n3849), .B(n3850), .Z(n3848) );
  XOR U4046 ( .A(n3851), .B(n3847), .Z(n3850) );
  XNOR U4047 ( .A(n3818), .B(n3806), .Z(n3845) );
  XOR U4048 ( .A(n3855), .B(n3813), .Z(n3818) );
  XNOR U4049 ( .A(n3811), .B(n3856), .Z(n3813) );
  ANDN U4050 ( .A(n2563), .B(n2008), .Z(n3856) );
  XOR U4051 ( .A(n3857), .B(n3858), .Z(n3811) );
  AND U4052 ( .A(n3859), .B(n3860), .Z(n3858) );
  XNOR U4053 ( .A(n3861), .B(n3857), .Z(n3860) );
  XOR U4054 ( .A(n3862), .B(n3815), .Z(n3855) );
  AND U4055 ( .A(n2006), .B(n2556), .Z(n3815) );
  IV U4056 ( .A(n3817), .Z(n3862) );
  XOR U4057 ( .A(n3866), .B(n3867), .Z(n3820) );
  AND U4058 ( .A(n3868), .B(n3869), .Z(n3867) );
  XOR U4059 ( .A(n3870), .B(n3871), .Z(n3869) );
  XOR U4060 ( .A(n3866), .B(n3872), .Z(n3871) );
  XNOR U4061 ( .A(n3853), .B(n3873), .Z(n3868) );
  XNOR U4062 ( .A(n3866), .B(n3854), .Z(n3873) );
  XNOR U4063 ( .A(n3838), .B(n3837), .Z(n3854) );
  XOR U4064 ( .A(n3874), .B(n3832), .Z(n3837) );
  XNOR U4065 ( .A(n3830), .B(n3875), .Z(n3832) );
  ANDN U4066 ( .A(n2134), .B(n2526), .Z(n3875) );
  XOR U4067 ( .A(n3876), .B(n3877), .Z(n3830) );
  AND U4068 ( .A(n3878), .B(n3879), .Z(n3877) );
  XNOR U4069 ( .A(n3880), .B(n3876), .Z(n3879) );
  XOR U4070 ( .A(n3881), .B(n3834), .Z(n3874) );
  AND U4071 ( .A(n2524), .B(n2127), .Z(n3834) );
  IV U4072 ( .A(n3836), .Z(n3881) );
  XNOR U4073 ( .A(n3842), .B(n3844), .Z(n3838) );
  NAND U4074 ( .A(n2763), .B(n1932), .Z(n3844) );
  XNOR U4075 ( .A(n3840), .B(n3885), .Z(n3842) );
  ANDN U4076 ( .A(n1937), .B(n2765), .Z(n3885) );
  XOR U4077 ( .A(n3886), .B(n3887), .Z(n3840) );
  AND U4078 ( .A(n3888), .B(n3889), .Z(n3887) );
  XOR U4079 ( .A(n3890), .B(n3886), .Z(n3889) );
  XOR U4080 ( .A(n3891), .B(n3865), .Z(n3853) );
  XNOR U4081 ( .A(n3849), .B(n3851), .Z(n3865) );
  NAND U4082 ( .A(n2309), .B(n2328), .Z(n3851) );
  XNOR U4083 ( .A(n3847), .B(n3892), .Z(n3849) );
  ANDN U4084 ( .A(n2333), .B(n2311), .Z(n3892) );
  XOR U4085 ( .A(n3893), .B(n3894), .Z(n3847) );
  AND U4086 ( .A(n3895), .B(n3896), .Z(n3894) );
  XOR U4087 ( .A(n3897), .B(n3893), .Z(n3896) );
  XNOR U4088 ( .A(n3864), .B(n3852), .Z(n3891) );
  XOR U4089 ( .A(n3901), .B(n3859), .Z(n3864) );
  XNOR U4090 ( .A(n3857), .B(n3902), .Z(n3859) );
  ANDN U4091 ( .A(n2563), .B(n2104), .Z(n3902) );
  XOR U4092 ( .A(n3903), .B(n3904), .Z(n3857) );
  AND U4093 ( .A(n3905), .B(n3906), .Z(n3904) );
  XNOR U4094 ( .A(n3907), .B(n3903), .Z(n3906) );
  XOR U4095 ( .A(n3908), .B(n3861), .Z(n3901) );
  AND U4096 ( .A(n2102), .B(n2556), .Z(n3861) );
  IV U4097 ( .A(n3863), .Z(n3908) );
  XOR U4098 ( .A(n3912), .B(n3913), .Z(n3866) );
  AND U4099 ( .A(n3914), .B(n3915), .Z(n3913) );
  XOR U4100 ( .A(n3916), .B(n3917), .Z(n3915) );
  XOR U4101 ( .A(n3912), .B(n3918), .Z(n3917) );
  XNOR U4102 ( .A(n3899), .B(n3919), .Z(n3914) );
  XNOR U4103 ( .A(n3912), .B(n3900), .Z(n3919) );
  XNOR U4104 ( .A(n3884), .B(n3883), .Z(n3900) );
  XOR U4105 ( .A(n3920), .B(n3878), .Z(n3883) );
  XNOR U4106 ( .A(n3876), .B(n3921), .Z(n3878) );
  ANDN U4107 ( .A(n2134), .B(n2645), .Z(n3921) );
  XOR U4108 ( .A(n3922), .B(n3923), .Z(n3876) );
  AND U4109 ( .A(n3924), .B(n3925), .Z(n3923) );
  XNOR U4110 ( .A(n3926), .B(n3922), .Z(n3925) );
  XOR U4111 ( .A(n3927), .B(n3880), .Z(n3920) );
  AND U4112 ( .A(n2643), .B(n2127), .Z(n3880) );
  IV U4113 ( .A(n3882), .Z(n3927) );
  XNOR U4114 ( .A(n3888), .B(n3890), .Z(n3884) );
  NAND U4115 ( .A(n2885), .B(n1932), .Z(n3890) );
  XNOR U4116 ( .A(n3886), .B(n3931), .Z(n3888) );
  ANDN U4117 ( .A(n1937), .B(n2887), .Z(n3931) );
  XOR U4118 ( .A(n3935), .B(n3911), .Z(n3899) );
  XNOR U4119 ( .A(n3895), .B(n3897), .Z(n3911) );
  NAND U4120 ( .A(n2416), .B(n2328), .Z(n3897) );
  XNOR U4121 ( .A(n3893), .B(n3936), .Z(n3895) );
  ANDN U4122 ( .A(n2333), .B(n2418), .Z(n3936) );
  XOR U4123 ( .A(n3937), .B(n3938), .Z(n3893) );
  AND U4124 ( .A(n3939), .B(n3940), .Z(n3938) );
  XOR U4125 ( .A(n3941), .B(n3937), .Z(n3940) );
  XNOR U4126 ( .A(n3910), .B(n3898), .Z(n3935) );
  XOR U4127 ( .A(n3945), .B(n3905), .Z(n3910) );
  XNOR U4128 ( .A(n3903), .B(n3946), .Z(n3905) );
  ANDN U4129 ( .A(n2563), .B(n2205), .Z(n3946) );
  XOR U4130 ( .A(n3947), .B(n3948), .Z(n3903) );
  AND U4131 ( .A(n3949), .B(n3950), .Z(n3948) );
  XNOR U4132 ( .A(n3951), .B(n3947), .Z(n3950) );
  XOR U4133 ( .A(n3952), .B(n3907), .Z(n3945) );
  AND U4134 ( .A(n2203), .B(n2556), .Z(n3907) );
  IV U4135 ( .A(n3909), .Z(n3952) );
  XOR U4136 ( .A(n3956), .B(n3957), .Z(n3912) );
  AND U4137 ( .A(n3958), .B(n3959), .Z(n3957) );
  XOR U4138 ( .A(n3960), .B(n3961), .Z(n3959) );
  XOR U4139 ( .A(n3956), .B(n3962), .Z(n3961) );
  XNOR U4140 ( .A(n3943), .B(n3963), .Z(n3958) );
  XNOR U4141 ( .A(n3956), .B(n3944), .Z(n3963) );
  XNOR U4142 ( .A(n3930), .B(n3929), .Z(n3944) );
  XOR U4143 ( .A(n3964), .B(n3924), .Z(n3929) );
  XNOR U4144 ( .A(n3922), .B(n3965), .Z(n3924) );
  ANDN U4145 ( .A(n2134), .B(n2765), .Z(n3965) );
  XOR U4146 ( .A(n3966), .B(n3967), .Z(n3922) );
  AND U4147 ( .A(n3968), .B(n3969), .Z(n3967) );
  XNOR U4148 ( .A(n3970), .B(n3966), .Z(n3969) );
  XOR U4149 ( .A(n3971), .B(n3926), .Z(n3964) );
  AND U4150 ( .A(n2763), .B(n2127), .Z(n3926) );
  IV U4151 ( .A(n3928), .Z(n3971) );
  XNOR U4152 ( .A(n3933), .B(n3934), .Z(n3930) );
  NAND U4153 ( .A(n3010), .B(n1932), .Z(n3934) );
  XNOR U4154 ( .A(n3932), .B(n3975), .Z(n3933) );
  ANDN U4155 ( .A(n1937), .B(n3012), .Z(n3975) );
  XOR U4156 ( .A(n3976), .B(n3977), .Z(n3932) );
  AND U4157 ( .A(n3978), .B(n3979), .Z(n3977) );
  XOR U4158 ( .A(n3980), .B(n3976), .Z(n3979) );
  XOR U4159 ( .A(n3981), .B(n3955), .Z(n3943) );
  XNOR U4160 ( .A(n3939), .B(n3941), .Z(n3955) );
  NAND U4161 ( .A(n2524), .B(n2328), .Z(n3941) );
  XNOR U4162 ( .A(n3937), .B(n3982), .Z(n3939) );
  ANDN U4163 ( .A(n2333), .B(n2526), .Z(n3982) );
  XOR U4164 ( .A(n3983), .B(n3984), .Z(n3937) );
  AND U4165 ( .A(n3985), .B(n3986), .Z(n3984) );
  XOR U4166 ( .A(n3987), .B(n3983), .Z(n3986) );
  XNOR U4167 ( .A(n3954), .B(n3942), .Z(n3981) );
  XOR U4168 ( .A(n3991), .B(n3949), .Z(n3954) );
  XNOR U4169 ( .A(n3947), .B(n3992), .Z(n3949) );
  ANDN U4170 ( .A(n2563), .B(n2311), .Z(n3992) );
  XOR U4171 ( .A(n3993), .B(n3994), .Z(n3947) );
  AND U4172 ( .A(n3995), .B(n3996), .Z(n3994) );
  XNOR U4173 ( .A(n3997), .B(n3993), .Z(n3996) );
  XOR U4174 ( .A(n3998), .B(n3951), .Z(n3991) );
  AND U4175 ( .A(n2309), .B(n2556), .Z(n3951) );
  IV U4176 ( .A(n3953), .Z(n3998) );
  XOR U4177 ( .A(n4002), .B(n4003), .Z(n3956) );
  AND U4178 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U4179 ( .A(n4006), .B(n4007), .Z(n4005) );
  XOR U4180 ( .A(n4002), .B(n4008), .Z(n4007) );
  XNOR U4181 ( .A(n3989), .B(n4009), .Z(n4004) );
  XNOR U4182 ( .A(n4002), .B(n3990), .Z(n4009) );
  XNOR U4183 ( .A(n3974), .B(n3973), .Z(n3990) );
  XOR U4184 ( .A(n4010), .B(n3968), .Z(n3973) );
  XNOR U4185 ( .A(n3966), .B(n4011), .Z(n3968) );
  ANDN U4186 ( .A(n2134), .B(n2887), .Z(n4011) );
  XOR U4187 ( .A(n4012), .B(n4013), .Z(n3966) );
  AND U4188 ( .A(n4014), .B(n4015), .Z(n4013) );
  XNOR U4189 ( .A(n4016), .B(n4012), .Z(n4015) );
  XOR U4190 ( .A(n4017), .B(n3970), .Z(n4010) );
  AND U4191 ( .A(n2885), .B(n2127), .Z(n3970) );
  IV U4192 ( .A(n3972), .Z(n4017) );
  XNOR U4193 ( .A(n3978), .B(n3980), .Z(n3974) );
  NAND U4194 ( .A(n3142), .B(n1932), .Z(n3980) );
  XNOR U4195 ( .A(n3976), .B(n4021), .Z(n3978) );
  ANDN U4196 ( .A(n1937), .B(n3144), .Z(n4021) );
  XOR U4197 ( .A(n4022), .B(n4023), .Z(n3976) );
  AND U4198 ( .A(n4024), .B(n4025), .Z(n4023) );
  XOR U4199 ( .A(n4026), .B(n4022), .Z(n4025) );
  XOR U4200 ( .A(n4027), .B(n4001), .Z(n3989) );
  XNOR U4201 ( .A(n3985), .B(n3987), .Z(n4001) );
  NAND U4202 ( .A(n2643), .B(n2328), .Z(n3987) );
  XNOR U4203 ( .A(n3983), .B(n4028), .Z(n3985) );
  ANDN U4204 ( .A(n2333), .B(n2645), .Z(n4028) );
  XOR U4205 ( .A(n4029), .B(n4030), .Z(n3983) );
  AND U4206 ( .A(n4031), .B(n4032), .Z(n4030) );
  XOR U4207 ( .A(n4033), .B(n4029), .Z(n4032) );
  XNOR U4208 ( .A(n4000), .B(n3988), .Z(n4027) );
  XOR U4209 ( .A(n4037), .B(n3995), .Z(n4000) );
  XNOR U4210 ( .A(n3993), .B(n4038), .Z(n3995) );
  ANDN U4211 ( .A(n2563), .B(n2418), .Z(n4038) );
  XOR U4212 ( .A(n4039), .B(n4040), .Z(n3993) );
  AND U4213 ( .A(n4041), .B(n4042), .Z(n4040) );
  XNOR U4214 ( .A(n4043), .B(n4039), .Z(n4042) );
  XOR U4215 ( .A(n4044), .B(n3997), .Z(n4037) );
  AND U4216 ( .A(n2416), .B(n2556), .Z(n3997) );
  IV U4217 ( .A(n3999), .Z(n4044) );
  XOR U4218 ( .A(n4048), .B(n4049), .Z(n4002) );
  AND U4219 ( .A(n4050), .B(n4051), .Z(n4049) );
  XOR U4220 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U4221 ( .A(n4048), .B(n4054), .Z(n4053) );
  XNOR U4222 ( .A(n4035), .B(n4055), .Z(n4050) );
  XNOR U4223 ( .A(n4048), .B(n4036), .Z(n4055) );
  XNOR U4224 ( .A(n4020), .B(n4019), .Z(n4036) );
  XOR U4225 ( .A(n4056), .B(n4014), .Z(n4019) );
  XNOR U4226 ( .A(n4012), .B(n4057), .Z(n4014) );
  ANDN U4227 ( .A(n2134), .B(n3012), .Z(n4057) );
  XOR U4228 ( .A(n4058), .B(n4059), .Z(n4012) );
  AND U4229 ( .A(n4060), .B(n4061), .Z(n4059) );
  XNOR U4230 ( .A(n4062), .B(n4058), .Z(n4061) );
  XOR U4231 ( .A(n4063), .B(n4016), .Z(n4056) );
  AND U4232 ( .A(n3010), .B(n2127), .Z(n4016) );
  IV U4233 ( .A(n4018), .Z(n4063) );
  XNOR U4234 ( .A(n4024), .B(n4026), .Z(n4020) );
  NAND U4235 ( .A(n3274), .B(n1932), .Z(n4026) );
  XNOR U4236 ( .A(n4022), .B(n4067), .Z(n4024) );
  ANDN U4237 ( .A(n1937), .B(n3276), .Z(n4067) );
  XOR U4238 ( .A(n4068), .B(n4069), .Z(n4022) );
  AND U4239 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR U4240 ( .A(n4072), .B(n4068), .Z(n4071) );
  XOR U4241 ( .A(n4073), .B(n4047), .Z(n4035) );
  XNOR U4242 ( .A(n4031), .B(n4033), .Z(n4047) );
  NAND U4243 ( .A(n2763), .B(n2328), .Z(n4033) );
  XNOR U4244 ( .A(n4029), .B(n4074), .Z(n4031) );
  ANDN U4245 ( .A(n2333), .B(n2765), .Z(n4074) );
  XOR U4246 ( .A(n4075), .B(n4076), .Z(n4029) );
  AND U4247 ( .A(n4077), .B(n4078), .Z(n4076) );
  XOR U4248 ( .A(n4079), .B(n4075), .Z(n4078) );
  XNOR U4249 ( .A(n4046), .B(n4034), .Z(n4073) );
  XOR U4250 ( .A(n4083), .B(n4041), .Z(n4046) );
  XNOR U4251 ( .A(n4039), .B(n4084), .Z(n4041) );
  ANDN U4252 ( .A(n2563), .B(n2526), .Z(n4084) );
  XOR U4253 ( .A(n4085), .B(n4086), .Z(n4039) );
  AND U4254 ( .A(n4087), .B(n4088), .Z(n4086) );
  XNOR U4255 ( .A(n4089), .B(n4085), .Z(n4088) );
  XOR U4256 ( .A(n4090), .B(n4043), .Z(n4083) );
  AND U4257 ( .A(n2524), .B(n2556), .Z(n4043) );
  IV U4258 ( .A(n4045), .Z(n4090) );
  XOR U4259 ( .A(n4094), .B(n4095), .Z(n4048) );
  AND U4260 ( .A(n4096), .B(n4097), .Z(n4095) );
  XOR U4261 ( .A(n4098), .B(n4099), .Z(n4097) );
  XOR U4262 ( .A(n4094), .B(n4100), .Z(n4099) );
  XNOR U4263 ( .A(n4081), .B(n4101), .Z(n4096) );
  XNOR U4264 ( .A(n4094), .B(n4082), .Z(n4101) );
  XNOR U4265 ( .A(n4066), .B(n4065), .Z(n4082) );
  XOR U4266 ( .A(n4102), .B(n4060), .Z(n4065) );
  XNOR U4267 ( .A(n4058), .B(n4103), .Z(n4060) );
  ANDN U4268 ( .A(n2134), .B(n3144), .Z(n4103) );
  XOR U4269 ( .A(n4107), .B(n4062), .Z(n4102) );
  AND U4270 ( .A(n3142), .B(n2127), .Z(n4062) );
  IV U4271 ( .A(n4064), .Z(n4107) );
  XNOR U4272 ( .A(n4070), .B(n4072), .Z(n4066) );
  NAND U4273 ( .A(n3415), .B(n1932), .Z(n4072) );
  XNOR U4274 ( .A(n4068), .B(n4111), .Z(n4070) );
  ANDN U4275 ( .A(n1937), .B(n3417), .Z(n4111) );
  XOR U4276 ( .A(n4115), .B(n4093), .Z(n4081) );
  XNOR U4277 ( .A(n4077), .B(n4079), .Z(n4093) );
  NAND U4278 ( .A(n2885), .B(n2328), .Z(n4079) );
  XNOR U4279 ( .A(n4075), .B(n4116), .Z(n4077) );
  ANDN U4280 ( .A(n2333), .B(n2887), .Z(n4116) );
  XOR U4281 ( .A(n4117), .B(n4118), .Z(n4075) );
  AND U4282 ( .A(n4119), .B(n4120), .Z(n4118) );
  XOR U4283 ( .A(n4121), .B(n4117), .Z(n4120) );
  XNOR U4284 ( .A(n4092), .B(n4080), .Z(n4115) );
  XOR U4285 ( .A(n4125), .B(n4087), .Z(n4092) );
  XNOR U4286 ( .A(n4085), .B(n4126), .Z(n4087) );
  ANDN U4287 ( .A(n2563), .B(n2645), .Z(n4126) );
  XOR U4288 ( .A(n4127), .B(n4128), .Z(n4085) );
  AND U4289 ( .A(n4129), .B(n4130), .Z(n4128) );
  XNOR U4290 ( .A(n4131), .B(n4127), .Z(n4130) );
  XOR U4291 ( .A(n4132), .B(n4089), .Z(n4125) );
  AND U4292 ( .A(n2643), .B(n2556), .Z(n4089) );
  IV U4293 ( .A(n4091), .Z(n4132) );
  XOR U4294 ( .A(n4137), .B(n4138), .Z(n3456) );
  XOR U4295 ( .A(n4139), .B(n4136), .Z(n4137) );
  XNOR U4296 ( .A(n4124), .B(n4123), .Z(n3455) );
  XOR U4297 ( .A(n4140), .B(n4135), .Z(n4123) );
  XNOR U4298 ( .A(n4119), .B(n4121), .Z(n4135) );
  NAND U4299 ( .A(n3010), .B(n2328), .Z(n4121) );
  XNOR U4300 ( .A(n4117), .B(n4141), .Z(n4119) );
  ANDN U4301 ( .A(n2333), .B(n3012), .Z(n4141) );
  XOR U4302 ( .A(n4134), .B(n4122), .Z(n4140) );
  XOR U4303 ( .A(n4145), .B(n4146), .Z(n4122) );
  XOR U4304 ( .A(n4147), .B(n4129), .Z(n4134) );
  XNOR U4305 ( .A(n4127), .B(n4148), .Z(n4129) );
  ANDN U4306 ( .A(n2563), .B(n2765), .Z(n4148) );
  AND U4307 ( .A(n2763), .B(n2556), .Z(n4131) );
  XNOR U4308 ( .A(n4152), .B(n4153), .Z(n4133) );
  AND U4309 ( .A(n4154), .B(n4155), .Z(n4153) );
  XNOR U4310 ( .A(n4150), .B(n4156), .Z(n4155) );
  XNOR U4311 ( .A(n4151), .B(n4152), .Z(n4156) );
  AND U4312 ( .A(n2885), .B(n2556), .Z(n4151) );
  XOR U4313 ( .A(n4149), .B(n4157), .Z(n4150) );
  ANDN U4314 ( .A(n2563), .B(n2887), .Z(n4157) );
  XNOR U4315 ( .A(n4143), .B(n4161), .Z(n4154) );
  XNOR U4316 ( .A(n4144), .B(n4152), .Z(n4161) );
  AND U4317 ( .A(n3142), .B(n2328), .Z(n4144) );
  XOR U4318 ( .A(n4142), .B(n4162), .Z(n4143) );
  ANDN U4319 ( .A(n2333), .B(n3144), .Z(n4162) );
  XOR U4320 ( .A(n4166), .B(n4167), .Z(n4152) );
  AND U4321 ( .A(n4168), .B(n4169), .Z(n4167) );
  XNOR U4322 ( .A(n4159), .B(n4170), .Z(n4169) );
  XNOR U4323 ( .A(n4160), .B(n4166), .Z(n4170) );
  AND U4324 ( .A(n3010), .B(n2556), .Z(n4160) );
  XOR U4325 ( .A(n4158), .B(n4171), .Z(n4159) );
  ANDN U4326 ( .A(n2563), .B(n3012), .Z(n4171) );
  XNOR U4327 ( .A(n4164), .B(n4175), .Z(n4168) );
  XNOR U4328 ( .A(n4165), .B(n4166), .Z(n4175) );
  AND U4329 ( .A(n3274), .B(n2328), .Z(n4165) );
  XOR U4330 ( .A(n4163), .B(n4176), .Z(n4164) );
  ANDN U4331 ( .A(n2333), .B(n3276), .Z(n4176) );
  XOR U4332 ( .A(n4180), .B(n4181), .Z(n4166) );
  AND U4333 ( .A(n4182), .B(n4183), .Z(n4181) );
  XNOR U4334 ( .A(n4173), .B(n4184), .Z(n4183) );
  XNOR U4335 ( .A(n4174), .B(n4180), .Z(n4184) );
  AND U4336 ( .A(n3142), .B(n2556), .Z(n4174) );
  XOR U4337 ( .A(n4172), .B(n4185), .Z(n4173) );
  ANDN U4338 ( .A(n2563), .B(n3144), .Z(n4185) );
  XNOR U4339 ( .A(n4178), .B(n4189), .Z(n4182) );
  XNOR U4340 ( .A(n4179), .B(n4180), .Z(n4189) );
  AND U4341 ( .A(n3415), .B(n2328), .Z(n4179) );
  XOR U4342 ( .A(n4177), .B(n4190), .Z(n4178) );
  ANDN U4343 ( .A(n2333), .B(n3417), .Z(n4190) );
  XNOR U4344 ( .A(n4195), .B(n4187), .Z(n4146) );
  XNOR U4345 ( .A(n4186), .B(n4196), .Z(n4187) );
  ANDN U4346 ( .A(n2563), .B(n3276), .Z(n4196) );
  XNOR U4347 ( .A(n4199), .B(n4197), .Z(n4198) );
  ANDN U4348 ( .A(n2563), .B(n3417), .Z(n4199) );
  XNOR U4349 ( .A(n4194), .B(n4188), .Z(n4195) );
  AND U4350 ( .A(n3274), .B(n2556), .Z(n4188) );
  XNOR U4351 ( .A(n4192), .B(n4193), .Z(n4145) );
  NAND U4352 ( .A(n4203), .B(n2328), .Z(n4193) );
  XNOR U4353 ( .A(n4191), .B(n4204), .Z(n4192) );
  ANDN U4354 ( .A(n2333), .B(n4205), .Z(n4204) );
  NAND U4355 ( .A(A[0]), .B(n4206), .Z(n4191) );
  NANDN U4356 ( .B(n2328), .A(n4207), .Z(n4206) );
  NANDN U4357 ( .B(n4208), .A(n2333), .Z(n4207) );
  IV U4358 ( .A(n2227), .Z(n2328) );
  XNOR U4359 ( .A(n4201), .B(n4202), .Z(n4194) );
  NAND U4360 ( .A(n4203), .B(n2556), .Z(n4202) );
  XNOR U4361 ( .A(n4200), .B(n4211), .Z(n4201) );
  ANDN U4362 ( .A(n2563), .B(n4205), .Z(n4211) );
  NAND U4363 ( .A(A[0]), .B(n4212), .Z(n4200) );
  NANDN U4364 ( .B(n2556), .A(n4213), .Z(n4212) );
  NANDN U4365 ( .B(n4208), .A(n2563), .Z(n4213) );
  IV U4366 ( .A(n2444), .Z(n2556) );
  XNOR U4367 ( .A(n4110), .B(n4109), .Z(n4124) );
  XOR U4368 ( .A(n4216), .B(n4105), .Z(n4109) );
  XNOR U4369 ( .A(n4104), .B(n4217), .Z(n4105) );
  ANDN U4370 ( .A(n2134), .B(n3276), .Z(n4217) );
  XNOR U4371 ( .A(n4220), .B(n4218), .Z(n4219) );
  ANDN U4372 ( .A(n2134), .B(n3417), .Z(n4220) );
  XNOR U4373 ( .A(n4108), .B(n4106), .Z(n4216) );
  AND U4374 ( .A(n3274), .B(n2127), .Z(n4106) );
  XNOR U4375 ( .A(n4222), .B(n4223), .Z(n4108) );
  NAND U4376 ( .A(n4203), .B(n2127), .Z(n4223) );
  XNOR U4377 ( .A(n4221), .B(n4224), .Z(n4222) );
  ANDN U4378 ( .A(n2134), .B(n4205), .Z(n4224) );
  NAND U4379 ( .A(A[0]), .B(n4225), .Z(n4221) );
  NANDN U4380 ( .B(n2127), .A(n4226), .Z(n4225) );
  NANDN U4381 ( .B(n4208), .A(n2134), .Z(n4226) );
  IV U4382 ( .A(n2028), .Z(n2127) );
  XNOR U4383 ( .A(n4113), .B(n4114), .Z(n4110) );
  NAND U4384 ( .A(n4203), .B(n1932), .Z(n4114) );
  XNOR U4385 ( .A(n4112), .B(n4229), .Z(n4113) );
  ANDN U4386 ( .A(n1937), .B(n4205), .Z(n4229) );
  NAND U4387 ( .A(A[0]), .B(n4230), .Z(n4112) );
  NANDN U4388 ( .B(n1932), .A(n4231), .Z(n4230) );
  NANDN U4389 ( .B(n4208), .A(n1937), .Z(n4231) );
  IV U4390 ( .A(n1836), .Z(n1932) );
  XNOR U4391 ( .A(n4234), .B(n4235), .Z(n4136) );
  XOR U4392 ( .A(n4236), .B(n3358), .Z(n3353) );
  XNOR U4393 ( .A(n3349), .B(n3350), .Z(n3358) );
  NAND U4394 ( .A(n3346), .B(n977), .Z(n3350) );
  XNOR U4395 ( .A(n3348), .B(n4237), .Z(n3349) );
  ANDN U4396 ( .A(n3351), .B(n979), .Z(n4237) );
  XOR U4397 ( .A(n4238), .B(n4239), .Z(n3348) );
  AND U4398 ( .A(n4240), .B(n4241), .Z(n4239) );
  XOR U4399 ( .A(n4242), .B(n4238), .Z(n4241) );
  XNOR U4400 ( .A(n3356), .B(n3352), .Z(n4236) );
  XNOR U4401 ( .A(n3467), .B(n3466), .Z(n3479) );
  XOR U4402 ( .A(n4244), .B(n3462), .Z(n3466) );
  XNOR U4403 ( .A(n3460), .B(n4245), .Z(n3462) );
  ANDN U4404 ( .A(n3072), .B(n1107), .Z(n4245) );
  XOR U4405 ( .A(n4246), .B(n4247), .Z(n3460) );
  AND U4406 ( .A(n4248), .B(n4249), .Z(n4247) );
  XNOR U4407 ( .A(n4250), .B(n4246), .Z(n4249) );
  AND U4408 ( .A(n3065), .B(n1105), .Z(n3464) );
  XNOR U4409 ( .A(n3471), .B(n3473), .Z(n3467) );
  NAND U4410 ( .A(n2818), .B(n1206), .Z(n3473) );
  XNOR U4411 ( .A(n3469), .B(n4254), .Z(n3471) );
  ANDN U4412 ( .A(n2823), .B(n1208), .Z(n4254) );
  XOR U4413 ( .A(n4255), .B(n4256), .Z(n3469) );
  AND U4414 ( .A(n4257), .B(n4258), .Z(n4256) );
  XOR U4415 ( .A(n4259), .B(n4255), .Z(n4258) );
  XOR U4416 ( .A(n4260), .B(n4261), .Z(n3480) );
  XNOR U4417 ( .A(n4262), .B(n4243), .Z(n4260) );
  XOR U4418 ( .A(n4264), .B(n4265), .Z(n3518) );
  XOR U4419 ( .A(n4266), .B(n4263), .Z(n4264) );
  XNOR U4420 ( .A(n4253), .B(n4252), .Z(n3516) );
  XOR U4421 ( .A(n4267), .B(n4248), .Z(n4252) );
  XNOR U4422 ( .A(n4246), .B(n4268), .Z(n4248) );
  ANDN U4423 ( .A(n3072), .B(n1149), .Z(n4268) );
  XOR U4424 ( .A(n4269), .B(n4270), .Z(n4246) );
  AND U4425 ( .A(n4271), .B(n4272), .Z(n4270) );
  XNOR U4426 ( .A(n4273), .B(n4269), .Z(n4272) );
  XOR U4427 ( .A(n4274), .B(n4250), .Z(n4267) );
  AND U4428 ( .A(n3065), .B(n1147), .Z(n4250) );
  IV U4429 ( .A(n4251), .Z(n4274) );
  XNOR U4430 ( .A(n4257), .B(n4259), .Z(n4253) );
  NAND U4431 ( .A(n2818), .B(n1270), .Z(n4259) );
  XNOR U4432 ( .A(n4255), .B(n4278), .Z(n4257) );
  ANDN U4433 ( .A(n2823), .B(n1272), .Z(n4278) );
  XOR U4434 ( .A(n4279), .B(n4280), .Z(n4255) );
  AND U4435 ( .A(n4281), .B(n4282), .Z(n4280) );
  XOR U4436 ( .A(n4283), .B(n4279), .Z(n4282) );
  XOR U4437 ( .A(n4285), .B(n4286), .Z(n3563) );
  XOR U4438 ( .A(n4287), .B(n4284), .Z(n4285) );
  XNOR U4439 ( .A(n4277), .B(n4276), .Z(n3561) );
  XOR U4440 ( .A(n4288), .B(n4271), .Z(n4276) );
  XNOR U4441 ( .A(n4269), .B(n4289), .Z(n4271) );
  ANDN U4442 ( .A(n3072), .B(n1208), .Z(n4289) );
  XOR U4443 ( .A(n4290), .B(n4291), .Z(n4269) );
  AND U4444 ( .A(n4292), .B(n4293), .Z(n4291) );
  XNOR U4445 ( .A(n4294), .B(n4290), .Z(n4293) );
  XOR U4446 ( .A(n4295), .B(n4273), .Z(n4288) );
  AND U4447 ( .A(n3065), .B(n1206), .Z(n4273) );
  IV U4448 ( .A(n4275), .Z(n4295) );
  XNOR U4449 ( .A(n4281), .B(n4283), .Z(n4277) );
  NAND U4450 ( .A(n2818), .B(n1338), .Z(n4283) );
  XNOR U4451 ( .A(n4279), .B(n4299), .Z(n4281) );
  ANDN U4452 ( .A(n2823), .B(n1340), .Z(n4299) );
  XOR U4453 ( .A(n4300), .B(n4301), .Z(n4279) );
  AND U4454 ( .A(n4302), .B(n4303), .Z(n4301) );
  XOR U4455 ( .A(n4304), .B(n4300), .Z(n4303) );
  XOR U4456 ( .A(n4306), .B(n4307), .Z(n3605) );
  XOR U4457 ( .A(n4308), .B(n4305), .Z(n4306) );
  XNOR U4458 ( .A(n4298), .B(n4297), .Z(n3603) );
  XOR U4459 ( .A(n4309), .B(n4292), .Z(n4297) );
  XNOR U4460 ( .A(n4290), .B(n4310), .Z(n4292) );
  ANDN U4461 ( .A(n3072), .B(n1272), .Z(n4310) );
  XOR U4462 ( .A(n4311), .B(n4312), .Z(n4290) );
  AND U4463 ( .A(n4313), .B(n4314), .Z(n4312) );
  XNOR U4464 ( .A(n4315), .B(n4311), .Z(n4314) );
  AND U4465 ( .A(n3065), .B(n1270), .Z(n4294) );
  XNOR U4466 ( .A(n4302), .B(n4304), .Z(n4298) );
  NAND U4467 ( .A(n2818), .B(n1405), .Z(n4304) );
  XNOR U4468 ( .A(n4300), .B(n4319), .Z(n4302) );
  ANDN U4469 ( .A(n2823), .B(n1407), .Z(n4319) );
  XOR U4470 ( .A(n4320), .B(n4321), .Z(n4300) );
  AND U4471 ( .A(n4322), .B(n4323), .Z(n4321) );
  XOR U4472 ( .A(n4324), .B(n4320), .Z(n4323) );
  XOR U4473 ( .A(n4326), .B(n4327), .Z(n3648) );
  XOR U4474 ( .A(n4328), .B(n4325), .Z(n4326) );
  XNOR U4475 ( .A(n4318), .B(n4317), .Z(n3646) );
  XOR U4476 ( .A(n4329), .B(n4313), .Z(n4317) );
  XNOR U4477 ( .A(n4311), .B(n4330), .Z(n4313) );
  ANDN U4478 ( .A(n3072), .B(n1340), .Z(n4330) );
  XOR U4479 ( .A(n4331), .B(n4332), .Z(n4311) );
  AND U4480 ( .A(n4333), .B(n4334), .Z(n4332) );
  XNOR U4481 ( .A(n4335), .B(n4331), .Z(n4334) );
  XOR U4482 ( .A(n4336), .B(n4315), .Z(n4329) );
  AND U4483 ( .A(n3065), .B(n1338), .Z(n4315) );
  IV U4484 ( .A(n4316), .Z(n4336) );
  XNOR U4485 ( .A(n4322), .B(n4324), .Z(n4318) );
  NAND U4486 ( .A(n2818), .B(n1479), .Z(n4324) );
  XNOR U4487 ( .A(n4320), .B(n4340), .Z(n4322) );
  ANDN U4488 ( .A(n2823), .B(n1481), .Z(n4340) );
  XOR U4489 ( .A(n4341), .B(n4342), .Z(n4320) );
  AND U4490 ( .A(n4343), .B(n4344), .Z(n4342) );
  XOR U4491 ( .A(n4345), .B(n4341), .Z(n4344) );
  XOR U4492 ( .A(n4347), .B(n4348), .Z(n3690) );
  XOR U4493 ( .A(n4349), .B(n4346), .Z(n4347) );
  XNOR U4494 ( .A(n4339), .B(n4338), .Z(n3688) );
  XOR U4495 ( .A(n4350), .B(n4333), .Z(n4338) );
  XNOR U4496 ( .A(n4331), .B(n4351), .Z(n4333) );
  ANDN U4497 ( .A(n3072), .B(n1407), .Z(n4351) );
  XOR U4498 ( .A(n4352), .B(n4353), .Z(n4331) );
  AND U4499 ( .A(n4354), .B(n4355), .Z(n4353) );
  XNOR U4500 ( .A(n4356), .B(n4352), .Z(n4355) );
  XOR U4501 ( .A(n4357), .B(n4335), .Z(n4350) );
  AND U4502 ( .A(n3065), .B(n1405), .Z(n4335) );
  IV U4503 ( .A(n4337), .Z(n4357) );
  XNOR U4504 ( .A(n4343), .B(n4345), .Z(n4339) );
  NAND U4505 ( .A(n2818), .B(n1557), .Z(n4345) );
  XNOR U4506 ( .A(n4341), .B(n4361), .Z(n4343) );
  ANDN U4507 ( .A(n2823), .B(n1559), .Z(n4361) );
  XOR U4508 ( .A(n4362), .B(n4363), .Z(n4341) );
  AND U4509 ( .A(n4364), .B(n4365), .Z(n4363) );
  XOR U4510 ( .A(n4366), .B(n4362), .Z(n4365) );
  XOR U4511 ( .A(n4368), .B(n4369), .Z(n3736) );
  XOR U4512 ( .A(n4370), .B(n4367), .Z(n4368) );
  XNOR U4513 ( .A(n4360), .B(n4359), .Z(n3734) );
  XOR U4514 ( .A(n4371), .B(n4354), .Z(n4359) );
  XNOR U4515 ( .A(n4352), .B(n4372), .Z(n4354) );
  ANDN U4516 ( .A(n3072), .B(n1481), .Z(n4372) );
  XOR U4517 ( .A(n4373), .B(n4374), .Z(n4352) );
  AND U4518 ( .A(n4375), .B(n4376), .Z(n4374) );
  XNOR U4519 ( .A(n4377), .B(n4373), .Z(n4376) );
  XOR U4520 ( .A(n4378), .B(n4356), .Z(n4371) );
  AND U4521 ( .A(n3065), .B(n1479), .Z(n4356) );
  IV U4522 ( .A(n4358), .Z(n4378) );
  XNOR U4523 ( .A(n4364), .B(n4366), .Z(n4360) );
  NAND U4524 ( .A(n2818), .B(n1638), .Z(n4366) );
  XNOR U4525 ( .A(n4362), .B(n4382), .Z(n4364) );
  ANDN U4526 ( .A(n2823), .B(n1640), .Z(n4382) );
  XOR U4527 ( .A(n4383), .B(n4384), .Z(n4362) );
  AND U4528 ( .A(n4385), .B(n4386), .Z(n4384) );
  XOR U4529 ( .A(n4387), .B(n4383), .Z(n4386) );
  XOR U4530 ( .A(n4389), .B(n4390), .Z(n3780) );
  XOR U4531 ( .A(n4391), .B(n4388), .Z(n4389) );
  XNOR U4532 ( .A(n4381), .B(n4380), .Z(n3778) );
  XOR U4533 ( .A(n4392), .B(n4375), .Z(n4380) );
  XNOR U4534 ( .A(n4373), .B(n4393), .Z(n4375) );
  ANDN U4535 ( .A(n3072), .B(n1559), .Z(n4393) );
  XOR U4536 ( .A(n4394), .B(n4395), .Z(n4373) );
  AND U4537 ( .A(n4396), .B(n4397), .Z(n4395) );
  XNOR U4538 ( .A(n4398), .B(n4394), .Z(n4397) );
  XOR U4539 ( .A(n4399), .B(n4377), .Z(n4392) );
  AND U4540 ( .A(n3065), .B(n1557), .Z(n4377) );
  IV U4541 ( .A(n4379), .Z(n4399) );
  XNOR U4542 ( .A(n4385), .B(n4387), .Z(n4381) );
  NAND U4543 ( .A(n2818), .B(n1722), .Z(n4387) );
  XNOR U4544 ( .A(n4383), .B(n4403), .Z(n4385) );
  ANDN U4545 ( .A(n2823), .B(n1724), .Z(n4403) );
  XOR U4546 ( .A(n4404), .B(n4405), .Z(n4383) );
  AND U4547 ( .A(n4406), .B(n4407), .Z(n4405) );
  XOR U4548 ( .A(n4408), .B(n4404), .Z(n4407) );
  XOR U4549 ( .A(n4410), .B(n4411), .Z(n3826) );
  XOR U4550 ( .A(n4412), .B(n4409), .Z(n4410) );
  XNOR U4551 ( .A(n4402), .B(n4401), .Z(n3824) );
  XOR U4552 ( .A(n4413), .B(n4396), .Z(n4401) );
  XNOR U4553 ( .A(n4394), .B(n4414), .Z(n4396) );
  ANDN U4554 ( .A(n3072), .B(n1640), .Z(n4414) );
  XOR U4555 ( .A(n4415), .B(n4416), .Z(n4394) );
  AND U4556 ( .A(n4417), .B(n4418), .Z(n4416) );
  XNOR U4557 ( .A(n4419), .B(n4415), .Z(n4418) );
  XOR U4558 ( .A(n4420), .B(n4398), .Z(n4413) );
  AND U4559 ( .A(n3065), .B(n1638), .Z(n4398) );
  IV U4560 ( .A(n4400), .Z(n4420) );
  XNOR U4561 ( .A(n4406), .B(n4408), .Z(n4402) );
  NAND U4562 ( .A(n2818), .B(n1813), .Z(n4408) );
  XNOR U4563 ( .A(n4404), .B(n4424), .Z(n4406) );
  ANDN U4564 ( .A(n2823), .B(n1815), .Z(n4424) );
  XOR U4565 ( .A(n4425), .B(n4426), .Z(n4404) );
  AND U4566 ( .A(n4427), .B(n4428), .Z(n4426) );
  XOR U4567 ( .A(n4429), .B(n4425), .Z(n4428) );
  XOR U4568 ( .A(n4431), .B(n4432), .Z(n3872) );
  XOR U4569 ( .A(n4433), .B(n4430), .Z(n4431) );
  XNOR U4570 ( .A(n4423), .B(n4422), .Z(n3870) );
  XOR U4571 ( .A(n4434), .B(n4417), .Z(n4422) );
  XNOR U4572 ( .A(n4415), .B(n4435), .Z(n4417) );
  ANDN U4573 ( .A(n3072), .B(n1724), .Z(n4435) );
  XOR U4574 ( .A(n4436), .B(n4437), .Z(n4415) );
  AND U4575 ( .A(n4438), .B(n4439), .Z(n4437) );
  XNOR U4576 ( .A(n4440), .B(n4436), .Z(n4439) );
  XOR U4577 ( .A(n4441), .B(n4419), .Z(n4434) );
  AND U4578 ( .A(n3065), .B(n1722), .Z(n4419) );
  IV U4579 ( .A(n4421), .Z(n4441) );
  XNOR U4580 ( .A(n4427), .B(n4429), .Z(n4423) );
  NAND U4581 ( .A(n2818), .B(n1910), .Z(n4429) );
  XNOR U4582 ( .A(n4425), .B(n4445), .Z(n4427) );
  ANDN U4583 ( .A(n2823), .B(n1912), .Z(n4445) );
  XOR U4584 ( .A(n4446), .B(n4447), .Z(n4425) );
  AND U4585 ( .A(n4448), .B(n4449), .Z(n4447) );
  XOR U4586 ( .A(n4450), .B(n4446), .Z(n4449) );
  XOR U4587 ( .A(n4452), .B(n4453), .Z(n3918) );
  XOR U4588 ( .A(n4454), .B(n4451), .Z(n4452) );
  XNOR U4589 ( .A(n4444), .B(n4443), .Z(n3916) );
  XOR U4590 ( .A(n4455), .B(n4438), .Z(n4443) );
  XNOR U4591 ( .A(n4436), .B(n4456), .Z(n4438) );
  ANDN U4592 ( .A(n3072), .B(n1815), .Z(n4456) );
  XOR U4593 ( .A(n4457), .B(n4458), .Z(n4436) );
  AND U4594 ( .A(n4459), .B(n4460), .Z(n4458) );
  XNOR U4595 ( .A(n4461), .B(n4457), .Z(n4460) );
  XOR U4596 ( .A(n4462), .B(n4440), .Z(n4455) );
  AND U4597 ( .A(n3065), .B(n1813), .Z(n4440) );
  IV U4598 ( .A(n4442), .Z(n4462) );
  XNOR U4599 ( .A(n4448), .B(n4450), .Z(n4444) );
  NAND U4600 ( .A(n2818), .B(n2006), .Z(n4450) );
  XNOR U4601 ( .A(n4446), .B(n4466), .Z(n4448) );
  ANDN U4602 ( .A(n2823), .B(n2008), .Z(n4466) );
  XOR U4603 ( .A(n4467), .B(n4468), .Z(n4446) );
  AND U4604 ( .A(n4469), .B(n4470), .Z(n4468) );
  XOR U4605 ( .A(n4471), .B(n4467), .Z(n4470) );
  XOR U4606 ( .A(n4473), .B(n4474), .Z(n3962) );
  XOR U4607 ( .A(n4475), .B(n4472), .Z(n4473) );
  XNOR U4608 ( .A(n4465), .B(n4464), .Z(n3960) );
  XOR U4609 ( .A(n4476), .B(n4459), .Z(n4464) );
  XNOR U4610 ( .A(n4457), .B(n4477), .Z(n4459) );
  ANDN U4611 ( .A(n3072), .B(n1912), .Z(n4477) );
  XOR U4612 ( .A(n4478), .B(n4479), .Z(n4457) );
  AND U4613 ( .A(n4480), .B(n4481), .Z(n4479) );
  XNOR U4614 ( .A(n4482), .B(n4478), .Z(n4481) );
  XOR U4615 ( .A(n4483), .B(n4461), .Z(n4476) );
  AND U4616 ( .A(n3065), .B(n1910), .Z(n4461) );
  IV U4617 ( .A(n4463), .Z(n4483) );
  XNOR U4618 ( .A(n4469), .B(n4471), .Z(n4465) );
  NAND U4619 ( .A(n2818), .B(n2102), .Z(n4471) );
  XNOR U4620 ( .A(n4467), .B(n4487), .Z(n4469) );
  ANDN U4621 ( .A(n2823), .B(n2104), .Z(n4487) );
  XOR U4622 ( .A(n4488), .B(n4489), .Z(n4467) );
  AND U4623 ( .A(n4490), .B(n4491), .Z(n4489) );
  XOR U4624 ( .A(n4492), .B(n4488), .Z(n4491) );
  XOR U4625 ( .A(n4494), .B(n4495), .Z(n4008) );
  XOR U4626 ( .A(n4496), .B(n4493), .Z(n4494) );
  XNOR U4627 ( .A(n4486), .B(n4485), .Z(n4006) );
  XOR U4628 ( .A(n4497), .B(n4480), .Z(n4485) );
  XNOR U4629 ( .A(n4478), .B(n4498), .Z(n4480) );
  ANDN U4630 ( .A(n3072), .B(n2008), .Z(n4498) );
  XOR U4631 ( .A(n4499), .B(n4500), .Z(n4478) );
  AND U4632 ( .A(n4501), .B(n4502), .Z(n4500) );
  XNOR U4633 ( .A(n4503), .B(n4499), .Z(n4502) );
  XOR U4634 ( .A(n4504), .B(n4482), .Z(n4497) );
  AND U4635 ( .A(n3065), .B(n2006), .Z(n4482) );
  IV U4636 ( .A(n4484), .Z(n4504) );
  XNOR U4637 ( .A(n4490), .B(n4492), .Z(n4486) );
  NAND U4638 ( .A(n2818), .B(n2203), .Z(n4492) );
  XNOR U4639 ( .A(n4488), .B(n4508), .Z(n4490) );
  ANDN U4640 ( .A(n2823), .B(n2205), .Z(n4508) );
  XOR U4641 ( .A(n4509), .B(n4510), .Z(n4488) );
  AND U4642 ( .A(n4511), .B(n4512), .Z(n4510) );
  XOR U4643 ( .A(n4513), .B(n4509), .Z(n4512) );
  XOR U4644 ( .A(n4515), .B(n4516), .Z(n4054) );
  XOR U4645 ( .A(n4517), .B(n4514), .Z(n4515) );
  XNOR U4646 ( .A(n4507), .B(n4506), .Z(n4052) );
  XOR U4647 ( .A(n4518), .B(n4501), .Z(n4506) );
  XNOR U4648 ( .A(n4499), .B(n4519), .Z(n4501) );
  ANDN U4649 ( .A(n3072), .B(n2104), .Z(n4519) );
  XOR U4650 ( .A(n4520), .B(n4521), .Z(n4499) );
  AND U4651 ( .A(n4522), .B(n4523), .Z(n4521) );
  XNOR U4652 ( .A(n4524), .B(n4520), .Z(n4523) );
  XOR U4653 ( .A(n4525), .B(n4503), .Z(n4518) );
  AND U4654 ( .A(n3065), .B(n2102), .Z(n4503) );
  IV U4655 ( .A(n4505), .Z(n4525) );
  XNOR U4656 ( .A(n4511), .B(n4513), .Z(n4507) );
  NAND U4657 ( .A(n2818), .B(n2309), .Z(n4513) );
  XNOR U4658 ( .A(n4509), .B(n4529), .Z(n4511) );
  ANDN U4659 ( .A(n2823), .B(n2311), .Z(n4529) );
  XOR U4660 ( .A(n4530), .B(n4531), .Z(n4509) );
  AND U4661 ( .A(n4532), .B(n4533), .Z(n4531) );
  XOR U4662 ( .A(n4534), .B(n4530), .Z(n4533) );
  XOR U4663 ( .A(n4536), .B(n4537), .Z(n4100) );
  XOR U4664 ( .A(n4538), .B(n4535), .Z(n4536) );
  XNOR U4665 ( .A(n4528), .B(n4527), .Z(n4098) );
  XOR U4666 ( .A(n4539), .B(n4522), .Z(n4527) );
  XNOR U4667 ( .A(n4520), .B(n4540), .Z(n4522) );
  ANDN U4668 ( .A(n3072), .B(n2205), .Z(n4540) );
  XOR U4669 ( .A(n4541), .B(n4542), .Z(n4520) );
  AND U4670 ( .A(n4543), .B(n4544), .Z(n4542) );
  XNOR U4671 ( .A(n4545), .B(n4541), .Z(n4544) );
  XOR U4672 ( .A(n4546), .B(n4524), .Z(n4539) );
  AND U4673 ( .A(n3065), .B(n2203), .Z(n4524) );
  IV U4674 ( .A(n4526), .Z(n4546) );
  XNOR U4675 ( .A(n4532), .B(n4534), .Z(n4528) );
  NAND U4676 ( .A(n2818), .B(n2416), .Z(n4534) );
  XNOR U4677 ( .A(n4530), .B(n4550), .Z(n4532) );
  ANDN U4678 ( .A(n2823), .B(n2418), .Z(n4550) );
  XOR U4679 ( .A(n4551), .B(n4552), .Z(n4530) );
  AND U4680 ( .A(n4553), .B(n4554), .Z(n4552) );
  XOR U4681 ( .A(n4555), .B(n4551), .Z(n4554) );
  XOR U4682 ( .A(n4557), .B(n4558), .Z(n4139) );
  XOR U4683 ( .A(n4559), .B(n4556), .Z(n4557) );
  XNOR U4684 ( .A(n4549), .B(n4548), .Z(n4138) );
  XOR U4685 ( .A(n4560), .B(n4543), .Z(n4548) );
  XNOR U4686 ( .A(n4541), .B(n4561), .Z(n4543) );
  ANDN U4687 ( .A(n3072), .B(n2311), .Z(n4561) );
  AND U4688 ( .A(n3065), .B(n2309), .Z(n4545) );
  XNOR U4689 ( .A(n4553), .B(n4555), .Z(n4549) );
  NAND U4690 ( .A(n2818), .B(n2524), .Z(n4555) );
  XNOR U4691 ( .A(n4551), .B(n4568), .Z(n4553) );
  ANDN U4692 ( .A(n2823), .B(n2526), .Z(n4568) );
  XOR U4693 ( .A(n4572), .B(n4573), .Z(n4556) );
  AND U4694 ( .A(n4574), .B(n4575), .Z(n4573) );
  XOR U4695 ( .A(n4576), .B(n4577), .Z(n4575) );
  XNOR U4696 ( .A(n4572), .B(n4578), .Z(n4577) );
  XNOR U4697 ( .A(n4566), .B(n4579), .Z(n4574) );
  XNOR U4698 ( .A(n4572), .B(n4567), .Z(n4579) );
  XNOR U4699 ( .A(n4570), .B(n4571), .Z(n4567) );
  NAND U4700 ( .A(n2643), .B(n2818), .Z(n4571) );
  XNOR U4701 ( .A(n4569), .B(n4580), .Z(n4570) );
  ANDN U4702 ( .A(n2823), .B(n2645), .Z(n4580) );
  XOR U4703 ( .A(n4584), .B(n4563), .Z(n4566) );
  XNOR U4704 ( .A(n4562), .B(n4585), .Z(n4563) );
  ANDN U4705 ( .A(n3072), .B(n2418), .Z(n4585) );
  AND U4706 ( .A(n3065), .B(n2416), .Z(n4564) );
  XOR U4707 ( .A(n4592), .B(n4593), .Z(n4572) );
  AND U4708 ( .A(n4594), .B(n4595), .Z(n4593) );
  XOR U4709 ( .A(n4596), .B(n4597), .Z(n4595) );
  XNOR U4710 ( .A(n4592), .B(n4598), .Z(n4597) );
  XNOR U4711 ( .A(n4590), .B(n4599), .Z(n4594) );
  XNOR U4712 ( .A(n4592), .B(n4591), .Z(n4599) );
  XNOR U4713 ( .A(n4582), .B(n4583), .Z(n4591) );
  NAND U4714 ( .A(n2763), .B(n2818), .Z(n4583) );
  XNOR U4715 ( .A(n4581), .B(n4600), .Z(n4582) );
  ANDN U4716 ( .A(n2823), .B(n2765), .Z(n4600) );
  XOR U4717 ( .A(n4604), .B(n4587), .Z(n4590) );
  XNOR U4718 ( .A(n4586), .B(n4605), .Z(n4587) );
  ANDN U4719 ( .A(n3072), .B(n2526), .Z(n4605) );
  AND U4720 ( .A(n3065), .B(n2524), .Z(n4588) );
  XOR U4721 ( .A(n4612), .B(n4613), .Z(n4592) );
  AND U4722 ( .A(n4614), .B(n4615), .Z(n4613) );
  XOR U4723 ( .A(n4616), .B(n4617), .Z(n4615) );
  XNOR U4724 ( .A(n4612), .B(n4618), .Z(n4617) );
  XNOR U4725 ( .A(n4610), .B(n4619), .Z(n4614) );
  XNOR U4726 ( .A(n4612), .B(n4611), .Z(n4619) );
  XNOR U4727 ( .A(n4602), .B(n4603), .Z(n4611) );
  NAND U4728 ( .A(n2885), .B(n2818), .Z(n4603) );
  XNOR U4729 ( .A(n4601), .B(n4620), .Z(n4602) );
  ANDN U4730 ( .A(n2823), .B(n2887), .Z(n4620) );
  XOR U4731 ( .A(n4624), .B(n4607), .Z(n4610) );
  XNOR U4732 ( .A(n4606), .B(n4625), .Z(n4607) );
  ANDN U4733 ( .A(n3072), .B(n2645), .Z(n4625) );
  AND U4734 ( .A(n2643), .B(n3065), .Z(n4608) );
  XOR U4735 ( .A(n4632), .B(n4633), .Z(n4612) );
  AND U4736 ( .A(n4634), .B(n4635), .Z(n4633) );
  XOR U4737 ( .A(n4636), .B(n4637), .Z(n4635) );
  XNOR U4738 ( .A(n4632), .B(n4638), .Z(n4637) );
  XNOR U4739 ( .A(n4630), .B(n4639), .Z(n4634) );
  XNOR U4740 ( .A(n4632), .B(n4631), .Z(n4639) );
  XNOR U4741 ( .A(n4622), .B(n4623), .Z(n4631) );
  NAND U4742 ( .A(n3010), .B(n2818), .Z(n4623) );
  XNOR U4743 ( .A(n4621), .B(n4640), .Z(n4622) );
  ANDN U4744 ( .A(n2823), .B(n3012), .Z(n4640) );
  XOR U4745 ( .A(n4644), .B(n4627), .Z(n4630) );
  XNOR U4746 ( .A(n4626), .B(n4645), .Z(n4627) );
  ANDN U4747 ( .A(n3072), .B(n2765), .Z(n4645) );
  AND U4748 ( .A(n2763), .B(n3065), .Z(n4628) );
  XOR U4749 ( .A(n4652), .B(n4653), .Z(n4632) );
  AND U4750 ( .A(n4654), .B(n4655), .Z(n4653) );
  XOR U4751 ( .A(n4656), .B(n4657), .Z(n4655) );
  XNOR U4752 ( .A(n4652), .B(n4658), .Z(n4657) );
  XNOR U4753 ( .A(n4650), .B(n4659), .Z(n4654) );
  XNOR U4754 ( .A(n4652), .B(n4651), .Z(n4659) );
  XNOR U4755 ( .A(n4642), .B(n4643), .Z(n4651) );
  NAND U4756 ( .A(n3142), .B(n2818), .Z(n4643) );
  XNOR U4757 ( .A(n4641), .B(n4660), .Z(n4642) );
  ANDN U4758 ( .A(n2823), .B(n3144), .Z(n4660) );
  XOR U4759 ( .A(n4664), .B(n4647), .Z(n4650) );
  XNOR U4760 ( .A(n4646), .B(n4665), .Z(n4647) );
  ANDN U4761 ( .A(n3072), .B(n2887), .Z(n4665) );
  AND U4762 ( .A(n2885), .B(n3065), .Z(n4648) );
  XOR U4763 ( .A(n4672), .B(n4673), .Z(n4652) );
  AND U4764 ( .A(n4674), .B(n4675), .Z(n4673) );
  XOR U4765 ( .A(n4676), .B(n4677), .Z(n4675) );
  XNOR U4766 ( .A(n4672), .B(n4678), .Z(n4677) );
  XNOR U4767 ( .A(n4670), .B(n4679), .Z(n4674) );
  XNOR U4768 ( .A(n4672), .B(n4671), .Z(n4679) );
  XNOR U4769 ( .A(n4662), .B(n4663), .Z(n4671) );
  NAND U4770 ( .A(n3274), .B(n2818), .Z(n4663) );
  XNOR U4771 ( .A(n4661), .B(n4680), .Z(n4662) );
  ANDN U4772 ( .A(n2823), .B(n3276), .Z(n4680) );
  XOR U4773 ( .A(n4681), .B(n4682), .Z(n4661) );
  AND U4774 ( .A(n4683), .B(n4684), .Z(n4682) );
  XOR U4775 ( .A(n4685), .B(n4681), .Z(n4684) );
  XOR U4776 ( .A(n4686), .B(n4667), .Z(n4670) );
  XNOR U4777 ( .A(n4666), .B(n4687), .Z(n4667) );
  ANDN U4778 ( .A(n3072), .B(n3012), .Z(n4687) );
  XOR U4779 ( .A(n4688), .B(n4689), .Z(n4666) );
  AND U4780 ( .A(n4690), .B(n4691), .Z(n4689) );
  XNOR U4781 ( .A(n4692), .B(n4688), .Z(n4691) );
  AND U4782 ( .A(n3010), .B(n3065), .Z(n4668) );
  XOR U4783 ( .A(n4696), .B(n4697), .Z(n4672) );
  AND U4784 ( .A(n4698), .B(n4699), .Z(n4697) );
  XOR U4785 ( .A(n4700), .B(n4701), .Z(n4699) );
  XNOR U4786 ( .A(n4696), .B(n4702), .Z(n4701) );
  XNOR U4787 ( .A(n4694), .B(n4703), .Z(n4698) );
  XNOR U4788 ( .A(n4696), .B(n4695), .Z(n4703) );
  XNOR U4789 ( .A(n4683), .B(n4685), .Z(n4695) );
  NAND U4790 ( .A(n3415), .B(n2818), .Z(n4685) );
  XNOR U4791 ( .A(n4681), .B(n4704), .Z(n4683) );
  ANDN U4792 ( .A(n2823), .B(n3417), .Z(n4704) );
  XOR U4793 ( .A(n4708), .B(n4690), .Z(n4694) );
  XNOR U4794 ( .A(n4688), .B(n4709), .Z(n4690) );
  ANDN U4795 ( .A(n3072), .B(n3144), .Z(n4709) );
  XOR U4796 ( .A(n4710), .B(n4711), .Z(n4688) );
  AND U4797 ( .A(n4712), .B(n4713), .Z(n4711) );
  XNOR U4798 ( .A(n4714), .B(n4710), .Z(n4713) );
  AND U4799 ( .A(n3142), .B(n3065), .Z(n4692) );
  XOR U4800 ( .A(n4719), .B(n4720), .Z(n4235) );
  XNOR U4801 ( .A(n4717), .B(n4716), .Z(n4234) );
  XOR U4802 ( .A(n4722), .B(n4712), .Z(n4716) );
  XNOR U4803 ( .A(n4710), .B(n4723), .Z(n4712) );
  ANDN U4804 ( .A(n3072), .B(n3276), .Z(n4723) );
  XNOR U4805 ( .A(n4726), .B(n4724), .Z(n4725) );
  ANDN U4806 ( .A(n3072), .B(n3417), .Z(n4726) );
  XNOR U4807 ( .A(n4715), .B(n4714), .Z(n4722) );
  AND U4808 ( .A(n3274), .B(n3065), .Z(n4714) );
  XNOR U4809 ( .A(n4728), .B(n4729), .Z(n4715) );
  NAND U4810 ( .A(n4203), .B(n3065), .Z(n4729) );
  XNOR U4811 ( .A(n4727), .B(n4730), .Z(n4728) );
  ANDN U4812 ( .A(n3072), .B(n4205), .Z(n4730) );
  NAND U4813 ( .A(A[0]), .B(n4731), .Z(n4727) );
  NANDN U4814 ( .B(n3065), .A(n4732), .Z(n4731) );
  NANDN U4815 ( .B(n4208), .A(n3072), .Z(n4732) );
  IV U4816 ( .A(n2939), .Z(n3065) );
  XNOR U4817 ( .A(n4706), .B(n4707), .Z(n4717) );
  NAND U4818 ( .A(n4203), .B(n2818), .Z(n4707) );
  XNOR U4819 ( .A(n4705), .B(n4735), .Z(n4706) );
  ANDN U4820 ( .A(n2823), .B(n4205), .Z(n4735) );
  NAND U4821 ( .A(A[0]), .B(n4736), .Z(n4705) );
  NANDN U4822 ( .B(n2818), .A(n4737), .Z(n4736) );
  NANDN U4823 ( .B(n4208), .A(n2823), .Z(n4737) );
  IV U4824 ( .A(n2697), .Z(n2818) );
  XOR U4825 ( .A(n4740), .B(n4741), .Z(n4718) );
  XOR U4826 ( .A(n3355), .B(n4742), .Z(n3356) );
  AND U4827 ( .A(n4743), .B(n4744), .Z(n4742) );
  NANDN U4828 ( .B(n4745), .A(n916), .Z(n4744) );
  NANDN U4829 ( .B(n4746), .A(n4747), .Z(n4743) );
  XNOR U4830 ( .A(n4240), .B(n4242), .Z(n4261) );
  NAND U4831 ( .A(n3346), .B(n1021), .Z(n4242) );
  XNOR U4832 ( .A(n4238), .B(n4749), .Z(n4240) );
  ANDN U4833 ( .A(n3351), .B(n1023), .Z(n4749) );
  XOR U4834 ( .A(n4750), .B(n4751), .Z(n4238) );
  AND U4835 ( .A(n4752), .B(n4753), .Z(n4751) );
  XOR U4836 ( .A(n4754), .B(n4750), .Z(n4753) );
  XNOR U4837 ( .A(n4755), .B(n4756), .Z(n4262) );
  IV U4838 ( .A(n4748), .Z(n4756) );
  XOR U4839 ( .A(n4757), .B(n4747), .Z(n4755) );
  AND U4840 ( .A(n4758), .B(n946), .Z(n4747) );
  IV U4841 ( .A(n979), .Z(n946) );
  NAND U4842 ( .A(n4759), .B(n4746), .Z(n4757) );
  XOR U4843 ( .A(n4760), .B(n4761), .Z(n4746) );
  AND U4844 ( .A(n4762), .B(n4763), .Z(n4761) );
  XNOR U4845 ( .A(n4764), .B(n4760), .Z(n4763) );
  NANDN U4846 ( .B(n949), .A(X[0]), .Z(n4759) );
  IV U4847 ( .A(n916), .Z(n949) );
  AND U4848 ( .A(n4765), .B(n4766), .Z(n916) );
  AND U4849 ( .A(A[31]), .B(n4767), .Z(n4765) );
  XNOR U4850 ( .A(n4752), .B(n4754), .Z(n4265) );
  NAND U4851 ( .A(n3346), .B(n1061), .Z(n4754) );
  XNOR U4852 ( .A(n4750), .B(n4769), .Z(n4752) );
  ANDN U4853 ( .A(n3351), .B(n1063), .Z(n4769) );
  XOR U4854 ( .A(n4770), .B(n4771), .Z(n4750) );
  AND U4855 ( .A(n4772), .B(n4773), .Z(n4771) );
  XOR U4856 ( .A(n4774), .B(n4770), .Z(n4773) );
  XNOR U4857 ( .A(n4775), .B(n4762), .Z(n4266) );
  XNOR U4858 ( .A(n4760), .B(n4776), .Z(n4762) );
  ANDN U4859 ( .A(X[0]), .B(n979), .Z(n4776) );
  XOR U4860 ( .A(n4767), .B(A[30]), .Z(n4766) );
  ANDN U4861 ( .A(n4777), .B(n4778), .Z(n4767) );
  XOR U4862 ( .A(n4779), .B(n4780), .Z(n4760) );
  AND U4863 ( .A(n4781), .B(n4782), .Z(n4780) );
  XNOR U4864 ( .A(n4783), .B(n4779), .Z(n4782) );
  XOR U4865 ( .A(n4784), .B(n4764), .Z(n4775) );
  AND U4866 ( .A(n4758), .B(n977), .Z(n4764) );
  IV U4867 ( .A(n1023), .Z(n977) );
  IV U4868 ( .A(n4768), .Z(n4784) );
  XNOR U4869 ( .A(n4772), .B(n4774), .Z(n4286) );
  NAND U4870 ( .A(n3346), .B(n1105), .Z(n4774) );
  XNOR U4871 ( .A(n4770), .B(n4786), .Z(n4772) );
  ANDN U4872 ( .A(n3351), .B(n1107), .Z(n4786) );
  XOR U4873 ( .A(n4787), .B(n4788), .Z(n4770) );
  AND U4874 ( .A(n4789), .B(n4790), .Z(n4788) );
  XOR U4875 ( .A(n4791), .B(n4787), .Z(n4790) );
  XNOR U4876 ( .A(n4792), .B(n4781), .Z(n4287) );
  XNOR U4877 ( .A(n4779), .B(n4793), .Z(n4781) );
  ANDN U4878 ( .A(X[0]), .B(n1023), .Z(n4793) );
  ANDN U4879 ( .A(n4794), .B(n4795), .Z(n4777) );
  XOR U4880 ( .A(n4796), .B(n4797), .Z(n4779) );
  AND U4881 ( .A(n4798), .B(n4799), .Z(n4797) );
  XNOR U4882 ( .A(n4800), .B(n4796), .Z(n4799) );
  XOR U4883 ( .A(n4801), .B(n4783), .Z(n4792) );
  AND U4884 ( .A(n4758), .B(n1021), .Z(n4783) );
  IV U4885 ( .A(n1063), .Z(n1021) );
  IV U4886 ( .A(n4785), .Z(n4801) );
  XNOR U4887 ( .A(n4789), .B(n4791), .Z(n4307) );
  NAND U4888 ( .A(n3346), .B(n1147), .Z(n4791) );
  XNOR U4889 ( .A(n4787), .B(n4803), .Z(n4789) );
  ANDN U4890 ( .A(n3351), .B(n1149), .Z(n4803) );
  XOR U4891 ( .A(n4804), .B(n4805), .Z(n4787) );
  AND U4892 ( .A(n4806), .B(n4807), .Z(n4805) );
  XOR U4893 ( .A(n4808), .B(n4804), .Z(n4807) );
  XNOR U4894 ( .A(n4809), .B(n4798), .Z(n4308) );
  XNOR U4895 ( .A(n4796), .B(n4810), .Z(n4798) );
  ANDN U4896 ( .A(X[0]), .B(n1063), .Z(n4810) );
  XNOR U4897 ( .A(n4794), .B(A[28]), .Z(n4795) );
  ANDN U4898 ( .A(n4811), .B(n4812), .Z(n4794) );
  XOR U4899 ( .A(n4813), .B(n4814), .Z(n4796) );
  AND U4900 ( .A(n4815), .B(n4816), .Z(n4814) );
  XNOR U4901 ( .A(n4817), .B(n4813), .Z(n4816) );
  AND U4902 ( .A(n4758), .B(n1061), .Z(n4800) );
  IV U4903 ( .A(n1107), .Z(n1061) );
  XNOR U4904 ( .A(n4806), .B(n4808), .Z(n4327) );
  NAND U4905 ( .A(n3346), .B(n1206), .Z(n4808) );
  XNOR U4906 ( .A(n4804), .B(n4819), .Z(n4806) );
  ANDN U4907 ( .A(n3351), .B(n1208), .Z(n4819) );
  XOR U4908 ( .A(n4820), .B(n4821), .Z(n4804) );
  AND U4909 ( .A(n4822), .B(n4823), .Z(n4821) );
  XOR U4910 ( .A(n4824), .B(n4820), .Z(n4823) );
  XNOR U4911 ( .A(n4825), .B(n4815), .Z(n4328) );
  XNOR U4912 ( .A(n4813), .B(n4826), .Z(n4815) );
  ANDN U4913 ( .A(X[0]), .B(n1107), .Z(n4826) );
  ANDN U4914 ( .A(n4827), .B(n4828), .Z(n4811) );
  XOR U4915 ( .A(n4829), .B(n4830), .Z(n4813) );
  AND U4916 ( .A(n4831), .B(n4832), .Z(n4830) );
  XNOR U4917 ( .A(n4833), .B(n4829), .Z(n4832) );
  AND U4918 ( .A(n4758), .B(n1105), .Z(n4817) );
  IV U4919 ( .A(n1149), .Z(n1105) );
  XNOR U4920 ( .A(n4822), .B(n4824), .Z(n4348) );
  NAND U4921 ( .A(n3346), .B(n1270), .Z(n4824) );
  XNOR U4922 ( .A(n4820), .B(n4835), .Z(n4822) );
  ANDN U4923 ( .A(n3351), .B(n1272), .Z(n4835) );
  XOR U4924 ( .A(n4836), .B(n4837), .Z(n4820) );
  AND U4925 ( .A(n4838), .B(n4839), .Z(n4837) );
  XOR U4926 ( .A(n4840), .B(n4836), .Z(n4839) );
  XNOR U4927 ( .A(n4841), .B(n4831), .Z(n4349) );
  XNOR U4928 ( .A(n4829), .B(n4842), .Z(n4831) );
  ANDN U4929 ( .A(X[0]), .B(n1149), .Z(n4842) );
  XNOR U4930 ( .A(n4827), .B(A[26]), .Z(n4828) );
  ANDN U4931 ( .A(n4843), .B(n4844), .Z(n4827) );
  XOR U4932 ( .A(n4845), .B(n4846), .Z(n4829) );
  AND U4933 ( .A(n4847), .B(n4848), .Z(n4846) );
  XNOR U4934 ( .A(n4849), .B(n4845), .Z(n4848) );
  XOR U4935 ( .A(n4850), .B(n4833), .Z(n4841) );
  AND U4936 ( .A(n4758), .B(n1147), .Z(n4833) );
  IV U4937 ( .A(n1208), .Z(n1147) );
  IV U4938 ( .A(n4834), .Z(n4850) );
  XNOR U4939 ( .A(n4838), .B(n4840), .Z(n4369) );
  NAND U4940 ( .A(n3346), .B(n1338), .Z(n4840) );
  XNOR U4941 ( .A(n4836), .B(n4852), .Z(n4838) );
  ANDN U4942 ( .A(n3351), .B(n1340), .Z(n4852) );
  XOR U4943 ( .A(n4853), .B(n4854), .Z(n4836) );
  AND U4944 ( .A(n4855), .B(n4856), .Z(n4854) );
  XOR U4945 ( .A(n4857), .B(n4853), .Z(n4856) );
  XNOR U4946 ( .A(n4858), .B(n4847), .Z(n4370) );
  XNOR U4947 ( .A(n4845), .B(n4859), .Z(n4847) );
  ANDN U4948 ( .A(X[0]), .B(n1208), .Z(n4859) );
  ANDN U4949 ( .A(n4860), .B(n4861), .Z(n4843) );
  XOR U4950 ( .A(n4862), .B(n4863), .Z(n4845) );
  AND U4951 ( .A(n4864), .B(n4865), .Z(n4863) );
  XNOR U4952 ( .A(n4866), .B(n4862), .Z(n4865) );
  XOR U4953 ( .A(n4867), .B(n4849), .Z(n4858) );
  AND U4954 ( .A(n4758), .B(n1206), .Z(n4849) );
  IV U4955 ( .A(n1272), .Z(n1206) );
  IV U4956 ( .A(n4851), .Z(n4867) );
  XNOR U4957 ( .A(n4855), .B(n4857), .Z(n4390) );
  NAND U4958 ( .A(n3346), .B(n1405), .Z(n4857) );
  XNOR U4959 ( .A(n4853), .B(n4869), .Z(n4855) );
  ANDN U4960 ( .A(n3351), .B(n1407), .Z(n4869) );
  XOR U4961 ( .A(n4870), .B(n4871), .Z(n4853) );
  AND U4962 ( .A(n4872), .B(n4873), .Z(n4871) );
  XOR U4963 ( .A(n4874), .B(n4870), .Z(n4873) );
  XNOR U4964 ( .A(n4875), .B(n4864), .Z(n4391) );
  XNOR U4965 ( .A(n4862), .B(n4876), .Z(n4864) );
  ANDN U4966 ( .A(X[0]), .B(n1272), .Z(n4876) );
  XNOR U4967 ( .A(n4860), .B(A[24]), .Z(n4861) );
  ANDN U4968 ( .A(n4877), .B(n4878), .Z(n4860) );
  XOR U4969 ( .A(n4879), .B(n4880), .Z(n4862) );
  AND U4970 ( .A(n4881), .B(n4882), .Z(n4880) );
  XNOR U4971 ( .A(n4883), .B(n4879), .Z(n4882) );
  XOR U4972 ( .A(n4884), .B(n4866), .Z(n4875) );
  AND U4973 ( .A(n4758), .B(n1270), .Z(n4866) );
  IV U4974 ( .A(n1340), .Z(n1270) );
  IV U4975 ( .A(n4868), .Z(n4884) );
  XNOR U4976 ( .A(n4872), .B(n4874), .Z(n4411) );
  NAND U4977 ( .A(n3346), .B(n1479), .Z(n4874) );
  XNOR U4978 ( .A(n4870), .B(n4886), .Z(n4872) );
  ANDN U4979 ( .A(n3351), .B(n1481), .Z(n4886) );
  XOR U4980 ( .A(n4887), .B(n4888), .Z(n4870) );
  AND U4981 ( .A(n4889), .B(n4890), .Z(n4888) );
  XOR U4982 ( .A(n4891), .B(n4887), .Z(n4890) );
  XNOR U4983 ( .A(n4892), .B(n4881), .Z(n4412) );
  XNOR U4984 ( .A(n4879), .B(n4893), .Z(n4881) );
  ANDN U4985 ( .A(X[0]), .B(n1340), .Z(n4893) );
  ANDN U4986 ( .A(n4894), .B(n4895), .Z(n4877) );
  XOR U4987 ( .A(n4896), .B(n4897), .Z(n4879) );
  AND U4988 ( .A(n4898), .B(n4899), .Z(n4897) );
  XNOR U4989 ( .A(n4900), .B(n4896), .Z(n4899) );
  XOR U4990 ( .A(n4901), .B(n4883), .Z(n4892) );
  AND U4991 ( .A(n4758), .B(n1338), .Z(n4883) );
  IV U4992 ( .A(n1407), .Z(n1338) );
  IV U4993 ( .A(n4885), .Z(n4901) );
  XNOR U4994 ( .A(n4889), .B(n4891), .Z(n4432) );
  NAND U4995 ( .A(n3346), .B(n1557), .Z(n4891) );
  XNOR U4996 ( .A(n4887), .B(n4903), .Z(n4889) );
  ANDN U4997 ( .A(n3351), .B(n1559), .Z(n4903) );
  XOR U4998 ( .A(n4904), .B(n4905), .Z(n4887) );
  AND U4999 ( .A(n4906), .B(n4907), .Z(n4905) );
  XOR U5000 ( .A(n4908), .B(n4904), .Z(n4907) );
  XNOR U5001 ( .A(n4909), .B(n4898), .Z(n4433) );
  XNOR U5002 ( .A(n4896), .B(n4910), .Z(n4898) );
  ANDN U5003 ( .A(X[0]), .B(n1407), .Z(n4910) );
  XNOR U5004 ( .A(n4894), .B(A[22]), .Z(n4895) );
  ANDN U5005 ( .A(n4911), .B(n4912), .Z(n4894) );
  XOR U5006 ( .A(n4913), .B(n4914), .Z(n4896) );
  AND U5007 ( .A(n4915), .B(n4916), .Z(n4914) );
  XNOR U5008 ( .A(n4917), .B(n4913), .Z(n4916) );
  XOR U5009 ( .A(n4918), .B(n4900), .Z(n4909) );
  AND U5010 ( .A(n4758), .B(n1405), .Z(n4900) );
  IV U5011 ( .A(n1481), .Z(n1405) );
  IV U5012 ( .A(n4902), .Z(n4918) );
  XNOR U5013 ( .A(n4906), .B(n4908), .Z(n4453) );
  NAND U5014 ( .A(n3346), .B(n1638), .Z(n4908) );
  XNOR U5015 ( .A(n4904), .B(n4920), .Z(n4906) );
  ANDN U5016 ( .A(n3351), .B(n1640), .Z(n4920) );
  XOR U5017 ( .A(n4921), .B(n4922), .Z(n4904) );
  AND U5018 ( .A(n4923), .B(n4924), .Z(n4922) );
  XOR U5019 ( .A(n4925), .B(n4921), .Z(n4924) );
  XNOR U5020 ( .A(n4926), .B(n4915), .Z(n4454) );
  XNOR U5021 ( .A(n4913), .B(n4927), .Z(n4915) );
  ANDN U5022 ( .A(X[0]), .B(n1481), .Z(n4927) );
  ANDN U5023 ( .A(n4928), .B(n4929), .Z(n4911) );
  XOR U5024 ( .A(n4930), .B(n4931), .Z(n4913) );
  AND U5025 ( .A(n4932), .B(n4933), .Z(n4931) );
  XNOR U5026 ( .A(n4934), .B(n4930), .Z(n4933) );
  XOR U5027 ( .A(n4935), .B(n4917), .Z(n4926) );
  AND U5028 ( .A(n4758), .B(n1479), .Z(n4917) );
  IV U5029 ( .A(n1559), .Z(n1479) );
  IV U5030 ( .A(n4919), .Z(n4935) );
  XNOR U5031 ( .A(n4923), .B(n4925), .Z(n4474) );
  NAND U5032 ( .A(n3346), .B(n1722), .Z(n4925) );
  XNOR U5033 ( .A(n4921), .B(n4937), .Z(n4923) );
  ANDN U5034 ( .A(n3351), .B(n1724), .Z(n4937) );
  XOR U5035 ( .A(n4938), .B(n4939), .Z(n4921) );
  AND U5036 ( .A(n4940), .B(n4941), .Z(n4939) );
  XOR U5037 ( .A(n4942), .B(n4938), .Z(n4941) );
  XNOR U5038 ( .A(n4943), .B(n4932), .Z(n4475) );
  XNOR U5039 ( .A(n4930), .B(n4944), .Z(n4932) );
  ANDN U5040 ( .A(X[0]), .B(n1559), .Z(n4944) );
  XNOR U5041 ( .A(n4928), .B(A[20]), .Z(n4929) );
  ANDN U5042 ( .A(n4945), .B(n4946), .Z(n4928) );
  XOR U5043 ( .A(n4947), .B(n4948), .Z(n4930) );
  AND U5044 ( .A(n4949), .B(n4950), .Z(n4948) );
  XNOR U5045 ( .A(n4951), .B(n4947), .Z(n4950) );
  XOR U5046 ( .A(n4952), .B(n4934), .Z(n4943) );
  AND U5047 ( .A(n4758), .B(n1557), .Z(n4934) );
  IV U5048 ( .A(n1640), .Z(n1557) );
  IV U5049 ( .A(n4936), .Z(n4952) );
  XNOR U5050 ( .A(n4940), .B(n4942), .Z(n4495) );
  NAND U5051 ( .A(n3346), .B(n1813), .Z(n4942) );
  XNOR U5052 ( .A(n4938), .B(n4954), .Z(n4940) );
  ANDN U5053 ( .A(n3351), .B(n1815), .Z(n4954) );
  XOR U5054 ( .A(n4955), .B(n4956), .Z(n4938) );
  AND U5055 ( .A(n4957), .B(n4958), .Z(n4956) );
  XOR U5056 ( .A(n4959), .B(n4955), .Z(n4958) );
  XNOR U5057 ( .A(n4960), .B(n4949), .Z(n4496) );
  XNOR U5058 ( .A(n4947), .B(n4961), .Z(n4949) );
  ANDN U5059 ( .A(X[0]), .B(n1640), .Z(n4961) );
  ANDN U5060 ( .A(n4962), .B(n4963), .Z(n4945) );
  XOR U5061 ( .A(n4964), .B(n4965), .Z(n4947) );
  AND U5062 ( .A(n4966), .B(n4967), .Z(n4965) );
  XNOR U5063 ( .A(n4968), .B(n4964), .Z(n4967) );
  XOR U5064 ( .A(n4969), .B(n4951), .Z(n4960) );
  AND U5065 ( .A(n4758), .B(n1638), .Z(n4951) );
  IV U5066 ( .A(n1724), .Z(n1638) );
  IV U5067 ( .A(n4953), .Z(n4969) );
  XNOR U5068 ( .A(n4957), .B(n4959), .Z(n4516) );
  NAND U5069 ( .A(n3346), .B(n1910), .Z(n4959) );
  XNOR U5070 ( .A(n4955), .B(n4971), .Z(n4957) );
  ANDN U5071 ( .A(n3351), .B(n1912), .Z(n4971) );
  XOR U5072 ( .A(n4972), .B(n4973), .Z(n4955) );
  AND U5073 ( .A(n4974), .B(n4975), .Z(n4973) );
  XOR U5074 ( .A(n4976), .B(n4972), .Z(n4975) );
  XNOR U5075 ( .A(n4977), .B(n4966), .Z(n4517) );
  XNOR U5076 ( .A(n4964), .B(n4978), .Z(n4966) );
  ANDN U5077 ( .A(X[0]), .B(n1724), .Z(n4978) );
  XNOR U5078 ( .A(n4962), .B(A[18]), .Z(n4963) );
  ANDN U5079 ( .A(n4979), .B(n4980), .Z(n4962) );
  XOR U5080 ( .A(n4981), .B(n4982), .Z(n4964) );
  AND U5081 ( .A(n4983), .B(n4984), .Z(n4982) );
  XNOR U5082 ( .A(n4985), .B(n4981), .Z(n4984) );
  XOR U5083 ( .A(n4986), .B(n4968), .Z(n4977) );
  AND U5084 ( .A(n4758), .B(n1722), .Z(n4968) );
  IV U5085 ( .A(n1815), .Z(n1722) );
  IV U5086 ( .A(n4970), .Z(n4986) );
  XNOR U5087 ( .A(n4974), .B(n4976), .Z(n4537) );
  NAND U5088 ( .A(n3346), .B(n2006), .Z(n4976) );
  XNOR U5089 ( .A(n4972), .B(n4988), .Z(n4974) );
  ANDN U5090 ( .A(n3351), .B(n2008), .Z(n4988) );
  XOR U5091 ( .A(n4989), .B(n4990), .Z(n4972) );
  AND U5092 ( .A(n4991), .B(n4992), .Z(n4990) );
  XOR U5093 ( .A(n4993), .B(n4989), .Z(n4992) );
  XNOR U5094 ( .A(n4994), .B(n4983), .Z(n4538) );
  XNOR U5095 ( .A(n4981), .B(n4995), .Z(n4983) );
  ANDN U5096 ( .A(X[0]), .B(n1815), .Z(n4995) );
  ANDN U5097 ( .A(n4996), .B(n4997), .Z(n4979) );
  XOR U5098 ( .A(n4998), .B(n4999), .Z(n4981) );
  AND U5099 ( .A(n5000), .B(n5001), .Z(n4999) );
  XNOR U5100 ( .A(n5002), .B(n4998), .Z(n5001) );
  XOR U5101 ( .A(n5003), .B(n4985), .Z(n4994) );
  AND U5102 ( .A(n4758), .B(n1813), .Z(n4985) );
  IV U5103 ( .A(n1912), .Z(n1813) );
  IV U5104 ( .A(n4987), .Z(n5003) );
  XNOR U5105 ( .A(n4991), .B(n4993), .Z(n4558) );
  NAND U5106 ( .A(n3346), .B(n2102), .Z(n4993) );
  XNOR U5107 ( .A(n4989), .B(n5005), .Z(n4991) );
  ANDN U5108 ( .A(n3351), .B(n2104), .Z(n5005) );
  XNOR U5109 ( .A(n5009), .B(n5000), .Z(n4559) );
  XNOR U5110 ( .A(n4998), .B(n5010), .Z(n5000) );
  ANDN U5111 ( .A(X[0]), .B(n1912), .Z(n5010) );
  AND U5112 ( .A(n4758), .B(n1910), .Z(n5002) );
  XNOR U5113 ( .A(n5007), .B(n5008), .Z(n4576) );
  NAND U5114 ( .A(n3346), .B(n2203), .Z(n5008) );
  XNOR U5115 ( .A(n5006), .B(n5015), .Z(n5007) );
  ANDN U5116 ( .A(n3351), .B(n2205), .Z(n5015) );
  XNOR U5117 ( .A(n5019), .B(n5012), .Z(n4578) );
  XNOR U5118 ( .A(n5011), .B(n5020), .Z(n5012) );
  ANDN U5119 ( .A(X[0]), .B(n2008), .Z(n5020) );
  AND U5120 ( .A(n4758), .B(n2006), .Z(n5013) );
  XNOR U5121 ( .A(n5017), .B(n5018), .Z(n4596) );
  NAND U5122 ( .A(n3346), .B(n2309), .Z(n5018) );
  XNOR U5123 ( .A(n5016), .B(n5025), .Z(n5017) );
  ANDN U5124 ( .A(n3351), .B(n2311), .Z(n5025) );
  XNOR U5125 ( .A(n5029), .B(n5022), .Z(n4598) );
  XNOR U5126 ( .A(n5021), .B(n5030), .Z(n5022) );
  ANDN U5127 ( .A(X[0]), .B(n2104), .Z(n5030) );
  AND U5128 ( .A(n4758), .B(n2102), .Z(n5023) );
  XNOR U5129 ( .A(n5027), .B(n5028), .Z(n4616) );
  NAND U5130 ( .A(n3346), .B(n2416), .Z(n5028) );
  XNOR U5131 ( .A(n5026), .B(n5035), .Z(n5027) );
  ANDN U5132 ( .A(n3351), .B(n2418), .Z(n5035) );
  XNOR U5133 ( .A(n5039), .B(n5032), .Z(n4618) );
  XNOR U5134 ( .A(n5031), .B(n5040), .Z(n5032) );
  ANDN U5135 ( .A(X[0]), .B(n2205), .Z(n5040) );
  XOR U5136 ( .A(n5041), .B(n5042), .Z(n5031) );
  AND U5137 ( .A(n5043), .B(n5044), .Z(n5042) );
  XNOR U5138 ( .A(n5045), .B(n5041), .Z(n5044) );
  AND U5139 ( .A(n4758), .B(n2203), .Z(n5033) );
  XNOR U5140 ( .A(n5037), .B(n5038), .Z(n4636) );
  NAND U5141 ( .A(n3346), .B(n2524), .Z(n5038) );
  XNOR U5142 ( .A(n5036), .B(n5047), .Z(n5037) );
  ANDN U5143 ( .A(n3351), .B(n2526), .Z(n5047) );
  XOR U5144 ( .A(n5048), .B(n5049), .Z(n5036) );
  AND U5145 ( .A(n5050), .B(n5051), .Z(n5049) );
  XOR U5146 ( .A(n5052), .B(n5048), .Z(n5051) );
  XNOR U5147 ( .A(n5053), .B(n5043), .Z(n4638) );
  XNOR U5148 ( .A(n5041), .B(n5054), .Z(n5043) );
  ANDN U5149 ( .A(X[0]), .B(n2311), .Z(n5054) );
  XOR U5150 ( .A(n5055), .B(n5056), .Z(n5041) );
  AND U5151 ( .A(n5057), .B(n5058), .Z(n5056) );
  XNOR U5152 ( .A(n5059), .B(n5055), .Z(n5058) );
  XOR U5153 ( .A(n5060), .B(n5045), .Z(n5053) );
  AND U5154 ( .A(n4758), .B(n2309), .Z(n5045) );
  IV U5155 ( .A(n5046), .Z(n5060) );
  XNOR U5156 ( .A(n5050), .B(n5052), .Z(n4656) );
  NAND U5157 ( .A(n3346), .B(n2643), .Z(n5052) );
  XNOR U5158 ( .A(n5048), .B(n5062), .Z(n5050) );
  ANDN U5159 ( .A(n3351), .B(n2645), .Z(n5062) );
  XOR U5160 ( .A(n5063), .B(n5064), .Z(n5048) );
  AND U5161 ( .A(n5065), .B(n5066), .Z(n5064) );
  XOR U5162 ( .A(n5067), .B(n5063), .Z(n5066) );
  XNOR U5163 ( .A(n5068), .B(n5057), .Z(n4658) );
  XNOR U5164 ( .A(n5055), .B(n5069), .Z(n5057) );
  ANDN U5165 ( .A(X[0]), .B(n2418), .Z(n5069) );
  XOR U5166 ( .A(n5070), .B(n5071), .Z(n5055) );
  AND U5167 ( .A(n5072), .B(n5073), .Z(n5071) );
  XNOR U5168 ( .A(n5074), .B(n5070), .Z(n5073) );
  XOR U5169 ( .A(n5075), .B(n5059), .Z(n5068) );
  AND U5170 ( .A(n4758), .B(n2416), .Z(n5059) );
  IV U5171 ( .A(n5061), .Z(n5075) );
  XNOR U5172 ( .A(n5065), .B(n5067), .Z(n4676) );
  NAND U5173 ( .A(n3346), .B(n2763), .Z(n5067) );
  XNOR U5174 ( .A(n5063), .B(n5077), .Z(n5065) );
  ANDN U5175 ( .A(n3351), .B(n2765), .Z(n5077) );
  XNOR U5176 ( .A(n5081), .B(n5072), .Z(n4678) );
  XNOR U5177 ( .A(n5070), .B(n5082), .Z(n5072) );
  ANDN U5178 ( .A(X[0]), .B(n2526), .Z(n5082) );
  XOR U5179 ( .A(n5083), .B(n5084), .Z(n5070) );
  AND U5180 ( .A(n5085), .B(n5086), .Z(n5084) );
  XNOR U5181 ( .A(n5087), .B(n5083), .Z(n5086) );
  AND U5182 ( .A(n4758), .B(n2524), .Z(n5074) );
  XNOR U5183 ( .A(n5079), .B(n5080), .Z(n4700) );
  NAND U5184 ( .A(n3346), .B(n2885), .Z(n5080) );
  XNOR U5185 ( .A(n5078), .B(n5089), .Z(n5079) );
  ANDN U5186 ( .A(n3351), .B(n2887), .Z(n5089) );
  XNOR U5187 ( .A(n5093), .B(n5085), .Z(n4702) );
  XNOR U5188 ( .A(n5083), .B(n5094), .Z(n5085) );
  ANDN U5189 ( .A(X[0]), .B(n2645), .Z(n5094) );
  XOR U5190 ( .A(n5095), .B(n5096), .Z(n5083) );
  AND U5191 ( .A(n5097), .B(n5098), .Z(n5096) );
  XNOR U5192 ( .A(n5099), .B(n5095), .Z(n5098) );
  AND U5193 ( .A(n4758), .B(n2643), .Z(n5087) );
  XNOR U5194 ( .A(n5091), .B(n5092), .Z(n4720) );
  NAND U5195 ( .A(n3346), .B(n3010), .Z(n5092) );
  XNOR U5196 ( .A(n5090), .B(n5101), .Z(n5091) );
  ANDN U5197 ( .A(n3351), .B(n3012), .Z(n5101) );
  XNOR U5198 ( .A(n5105), .B(n5097), .Z(n4721) );
  XNOR U5199 ( .A(n5095), .B(n5106), .Z(n5097) );
  ANDN U5200 ( .A(X[0]), .B(n2765), .Z(n5106) );
  AND U5201 ( .A(n4758), .B(n2763), .Z(n5099) );
  XNOR U5202 ( .A(n5110), .B(n5111), .Z(n5100) );
  AND U5203 ( .A(n5112), .B(n5113), .Z(n5111) );
  XNOR U5204 ( .A(n5108), .B(n5114), .Z(n5113) );
  XNOR U5205 ( .A(n5109), .B(n5110), .Z(n5114) );
  AND U5206 ( .A(n4758), .B(n2885), .Z(n5109) );
  XOR U5207 ( .A(n5107), .B(n5115), .Z(n5108) );
  ANDN U5208 ( .A(X[0]), .B(n2887), .Z(n5115) );
  XNOR U5209 ( .A(n5103), .B(n5119), .Z(n5112) );
  XNOR U5210 ( .A(n5104), .B(n5110), .Z(n5119) );
  AND U5211 ( .A(n3142), .B(n3346), .Z(n5104) );
  XOR U5212 ( .A(n5102), .B(n5120), .Z(n5103) );
  ANDN U5213 ( .A(n3351), .B(n3144), .Z(n5120) );
  XOR U5214 ( .A(n5124), .B(n5125), .Z(n5110) );
  AND U5215 ( .A(n5126), .B(n5127), .Z(n5125) );
  XNOR U5216 ( .A(n5117), .B(n5128), .Z(n5127) );
  XNOR U5217 ( .A(n5118), .B(n5124), .Z(n5128) );
  AND U5218 ( .A(n4758), .B(n3010), .Z(n5118) );
  XOR U5219 ( .A(n5116), .B(n5129), .Z(n5117) );
  ANDN U5220 ( .A(X[0]), .B(n3012), .Z(n5129) );
  XNOR U5221 ( .A(n5122), .B(n5133), .Z(n5126) );
  XNOR U5222 ( .A(n5123), .B(n5124), .Z(n5133) );
  AND U5223 ( .A(n3274), .B(n3346), .Z(n5123) );
  XOR U5224 ( .A(n5121), .B(n5134), .Z(n5122) );
  ANDN U5225 ( .A(n3351), .B(n3276), .Z(n5134) );
  XOR U5226 ( .A(n5135), .B(n5136), .Z(n5121) );
  ANDN U5227 ( .A(n5137), .B(n5138), .Z(n5136) );
  XNOR U5228 ( .A(n5139), .B(n5135), .Z(n5137) );
  XOR U5229 ( .A(n5140), .B(n5141), .Z(n5124) );
  AND U5230 ( .A(n5142), .B(n5143), .Z(n5141) );
  XNOR U5231 ( .A(n5131), .B(n5144), .Z(n5143) );
  XNOR U5232 ( .A(n5132), .B(n5140), .Z(n5144) );
  AND U5233 ( .A(n4758), .B(n3142), .Z(n5132) );
  XOR U5234 ( .A(n5130), .B(n5145), .Z(n5131) );
  ANDN U5235 ( .A(X[0]), .B(n3144), .Z(n5145) );
  XNOR U5236 ( .A(n5138), .B(n5149), .Z(n5142) );
  XNOR U5237 ( .A(n5139), .B(n5140), .Z(n5149) );
  AND U5238 ( .A(n3415), .B(n3346), .Z(n5139) );
  XOR U5239 ( .A(n5135), .B(n5150), .Z(n5138) );
  ANDN U5240 ( .A(n3351), .B(n3417), .Z(n5150) );
  XNOR U5241 ( .A(n5155), .B(n5147), .Z(n4741) );
  XNOR U5242 ( .A(n5146), .B(n5156), .Z(n5147) );
  ANDN U5243 ( .A(X[0]), .B(n3276), .Z(n5156) );
  XNOR U5244 ( .A(n5159), .B(n5157), .Z(n5158) );
  ANDN U5245 ( .A(X[0]), .B(n3417), .Z(n5159) );
  ANDN U5246 ( .A(n4758), .B(n4205), .Z(n5160) );
  XNOR U5247 ( .A(n5154), .B(n5148), .Z(n5155) );
  AND U5248 ( .A(n4758), .B(n3274), .Z(n5148) );
  XNOR U5249 ( .A(n5152), .B(n5153), .Z(n4740) );
  NAND U5250 ( .A(n4203), .B(n3346), .Z(n5153) );
  XNOR U5251 ( .A(n5151), .B(n5164), .Z(n5152) );
  ANDN U5252 ( .A(n3351), .B(n4205), .Z(n5164) );
  NAND U5253 ( .A(A[0]), .B(n5165), .Z(n5151) );
  NANDN U5254 ( .B(n3346), .A(n5166), .Z(n5165) );
  NANDN U5255 ( .B(n4208), .A(n3351), .Z(n5166) );
  IV U5256 ( .A(n3212), .Z(n3346) );
  XNOR U5257 ( .A(n5162), .B(n5163), .Z(n5154) );
  NAND U5258 ( .A(n4203), .B(n4758), .Z(n5163) );
  XNOR U5259 ( .A(n5161), .B(n5169), .Z(n5162) );
  ANDN U5260 ( .A(X[0]), .B(n4205), .Z(n5169) );
  NAND U5261 ( .A(A[0]), .B(n5170), .Z(n5161) );
  NANDN U5262 ( .B(n4758), .A(n5171), .Z(n5170) );
  NANDN U5263 ( .B(n4208), .A(X[0]), .Z(n5171) );
  IV U5264 ( .A(n4745), .Z(n4758) );
  XNOR U5265 ( .A(n3374), .B(n3373), .Z(n3327) );
  XOR U5266 ( .A(n5173), .B(n3382), .Z(n3373) );
  XNOR U5267 ( .A(n3367), .B(n3366), .Z(n3382) );
  XOR U5268 ( .A(n5174), .B(n3363), .Z(n3366) );
  XNOR U5269 ( .A(n3362), .B(n5175), .Z(n3363) );
  ANDN U5270 ( .A(n1426), .B(n2311), .Z(n5175) );
  AND U5271 ( .A(n2309), .B(n1363), .Z(n3364) );
  XNOR U5272 ( .A(n3370), .B(n3371), .Z(n3367) );
  NANDN U5273 ( .B(n1228), .A(n2524), .Z(n3371) );
  XNOR U5274 ( .A(n3369), .B(n5182), .Z(n3370) );
  ANDN U5275 ( .A(n1298), .B(n2526), .Z(n5182) );
  XOR U5276 ( .A(n3381), .B(n3372), .Z(n5173) );
  XNOR U5277 ( .A(n5186), .B(n5187), .Z(n3372) );
  XOR U5278 ( .A(n5188), .B(n3390), .Z(n3381) );
  XNOR U5279 ( .A(n3378), .B(n3379), .Z(n3390) );
  NAND U5280 ( .A(n2102), .B(n1597), .Z(n3379) );
  XNOR U5281 ( .A(n3377), .B(n5189), .Z(n3378) );
  ANDN U5282 ( .A(n1604), .B(n2104), .Z(n5189) );
  XNOR U5283 ( .A(n3389), .B(n3380), .Z(n5188) );
  XOR U5284 ( .A(n5193), .B(n5194), .Z(n3380) );
  AND U5285 ( .A(n5195), .B(n5196), .Z(n5194) );
  XOR U5286 ( .A(n5197), .B(n5198), .Z(n5196) );
  XNOR U5287 ( .A(n5193), .B(n5199), .Z(n5198) );
  XNOR U5288 ( .A(n5180), .B(n5200), .Z(n5195) );
  XNOR U5289 ( .A(n5193), .B(n5181), .Z(n5200) );
  XNOR U5290 ( .A(n5184), .B(n5185), .Z(n5181) );
  NANDN U5291 ( .B(n1228), .A(n2643), .Z(n5185) );
  XNOR U5292 ( .A(n5183), .B(n5201), .Z(n5184) );
  ANDN U5293 ( .A(n1298), .B(n2645), .Z(n5201) );
  XOR U5294 ( .A(n5205), .B(n5177), .Z(n5180) );
  XNOR U5295 ( .A(n5176), .B(n5206), .Z(n5177) );
  ANDN U5296 ( .A(n1426), .B(n2418), .Z(n5206) );
  AND U5297 ( .A(n2416), .B(n1363), .Z(n5178) );
  XOR U5298 ( .A(n5213), .B(n5214), .Z(n5193) );
  AND U5299 ( .A(n5215), .B(n5216), .Z(n5214) );
  XOR U5300 ( .A(n5217), .B(n5218), .Z(n5216) );
  XNOR U5301 ( .A(n5213), .B(n5219), .Z(n5218) );
  XNOR U5302 ( .A(n5211), .B(n5220), .Z(n5215) );
  XNOR U5303 ( .A(n5213), .B(n5212), .Z(n5220) );
  XNOR U5304 ( .A(n5203), .B(n5204), .Z(n5212) );
  NANDN U5305 ( .B(n1228), .A(n2763), .Z(n5204) );
  XNOR U5306 ( .A(n5202), .B(n5221), .Z(n5203) );
  ANDN U5307 ( .A(n1298), .B(n2765), .Z(n5221) );
  XOR U5308 ( .A(n5225), .B(n5208), .Z(n5211) );
  XNOR U5309 ( .A(n5207), .B(n5226), .Z(n5208) );
  ANDN U5310 ( .A(n1426), .B(n2526), .Z(n5226) );
  AND U5311 ( .A(n2524), .B(n1363), .Z(n5209) );
  XOR U5312 ( .A(n5233), .B(n5234), .Z(n5213) );
  AND U5313 ( .A(n5235), .B(n5236), .Z(n5234) );
  XOR U5314 ( .A(n5237), .B(n5238), .Z(n5236) );
  XNOR U5315 ( .A(n5233), .B(n5239), .Z(n5238) );
  XNOR U5316 ( .A(n5231), .B(n5240), .Z(n5235) );
  XNOR U5317 ( .A(n5233), .B(n5232), .Z(n5240) );
  XNOR U5318 ( .A(n5223), .B(n5224), .Z(n5232) );
  NANDN U5319 ( .B(n1228), .A(n2885), .Z(n5224) );
  XNOR U5320 ( .A(n5222), .B(n5241), .Z(n5223) );
  ANDN U5321 ( .A(n1298), .B(n2887), .Z(n5241) );
  XOR U5322 ( .A(n5245), .B(n5228), .Z(n5231) );
  XNOR U5323 ( .A(n5227), .B(n5246), .Z(n5228) );
  ANDN U5324 ( .A(n1426), .B(n2645), .Z(n5246) );
  AND U5325 ( .A(n2643), .B(n1363), .Z(n5229) );
  XOR U5326 ( .A(n5253), .B(n5254), .Z(n5233) );
  AND U5327 ( .A(n5255), .B(n5256), .Z(n5254) );
  XOR U5328 ( .A(n5257), .B(n5258), .Z(n5256) );
  XNOR U5329 ( .A(n5253), .B(n5259), .Z(n5258) );
  XNOR U5330 ( .A(n5251), .B(n5260), .Z(n5255) );
  XNOR U5331 ( .A(n5253), .B(n5252), .Z(n5260) );
  XNOR U5332 ( .A(n5243), .B(n5244), .Z(n5252) );
  NANDN U5333 ( .B(n1228), .A(n3010), .Z(n5244) );
  XNOR U5334 ( .A(n5242), .B(n5261), .Z(n5243) );
  ANDN U5335 ( .A(n1298), .B(n3012), .Z(n5261) );
  XOR U5336 ( .A(n5265), .B(n5248), .Z(n5251) );
  XNOR U5337 ( .A(n5247), .B(n5266), .Z(n5248) );
  ANDN U5338 ( .A(n1426), .B(n2765), .Z(n5266) );
  AND U5339 ( .A(n2763), .B(n1363), .Z(n5249) );
  XOR U5340 ( .A(n5273), .B(n5274), .Z(n5253) );
  AND U5341 ( .A(n5275), .B(n5276), .Z(n5274) );
  XOR U5342 ( .A(n5277), .B(n5278), .Z(n5276) );
  XNOR U5343 ( .A(n5273), .B(n5279), .Z(n5278) );
  XNOR U5344 ( .A(n5271), .B(n5280), .Z(n5275) );
  XNOR U5345 ( .A(n5273), .B(n5272), .Z(n5280) );
  XNOR U5346 ( .A(n5263), .B(n5264), .Z(n5272) );
  NANDN U5347 ( .B(n1228), .A(n3142), .Z(n5264) );
  XNOR U5348 ( .A(n5262), .B(n5281), .Z(n5263) );
  ANDN U5349 ( .A(n1298), .B(n3144), .Z(n5281) );
  XOR U5350 ( .A(n5285), .B(n5268), .Z(n5271) );
  XNOR U5351 ( .A(n5267), .B(n5286), .Z(n5268) );
  ANDN U5352 ( .A(n1426), .B(n2887), .Z(n5286) );
  XOR U5353 ( .A(n5287), .B(n5288), .Z(n5267) );
  AND U5354 ( .A(n5289), .B(n5290), .Z(n5288) );
  XNOR U5355 ( .A(n5291), .B(n5287), .Z(n5290) );
  AND U5356 ( .A(n2885), .B(n1363), .Z(n5269) );
  XOR U5357 ( .A(n5295), .B(n5296), .Z(n5273) );
  AND U5358 ( .A(n5297), .B(n5298), .Z(n5296) );
  XOR U5359 ( .A(n5299), .B(n5300), .Z(n5298) );
  XNOR U5360 ( .A(n5295), .B(n5301), .Z(n5300) );
  XNOR U5361 ( .A(n5293), .B(n5302), .Z(n5297) );
  XNOR U5362 ( .A(n5295), .B(n5294), .Z(n5302) );
  XNOR U5363 ( .A(n5283), .B(n5284), .Z(n5294) );
  NANDN U5364 ( .B(n1228), .A(n3274), .Z(n5284) );
  XNOR U5365 ( .A(n5282), .B(n5303), .Z(n5283) );
  ANDN U5366 ( .A(n1298), .B(n3276), .Z(n5303) );
  XOR U5367 ( .A(n5304), .B(n5305), .Z(n5282) );
  AND U5368 ( .A(n5306), .B(n5307), .Z(n5305) );
  XOR U5369 ( .A(n5308), .B(n5304), .Z(n5307) );
  XOR U5370 ( .A(n5309), .B(n5289), .Z(n5293) );
  XNOR U5371 ( .A(n5287), .B(n5310), .Z(n5289) );
  ANDN U5372 ( .A(n1426), .B(n3012), .Z(n5310) );
  XOR U5373 ( .A(n5311), .B(n5312), .Z(n5287) );
  AND U5374 ( .A(n5313), .B(n5314), .Z(n5312) );
  XNOR U5375 ( .A(n5315), .B(n5311), .Z(n5314) );
  AND U5376 ( .A(n3010), .B(n1363), .Z(n5291) );
  XOR U5377 ( .A(n5319), .B(n5320), .Z(n5295) );
  AND U5378 ( .A(n5321), .B(n5322), .Z(n5320) );
  XOR U5379 ( .A(n5323), .B(n5324), .Z(n5322) );
  XNOR U5380 ( .A(n5319), .B(n5325), .Z(n5324) );
  XNOR U5381 ( .A(n5317), .B(n5326), .Z(n5321) );
  XNOR U5382 ( .A(n5319), .B(n5318), .Z(n5326) );
  XNOR U5383 ( .A(n5306), .B(n5308), .Z(n5318) );
  NANDN U5384 ( .B(n1228), .A(n3415), .Z(n5308) );
  XNOR U5385 ( .A(n5304), .B(n5327), .Z(n5306) );
  ANDN U5386 ( .A(n1298), .B(n3417), .Z(n5327) );
  XOR U5387 ( .A(n5331), .B(n5313), .Z(n5317) );
  XNOR U5388 ( .A(n5311), .B(n5332), .Z(n5313) );
  ANDN U5389 ( .A(n1426), .B(n3144), .Z(n5332) );
  AND U5390 ( .A(n3142), .B(n1363), .Z(n5315) );
  XOR U5391 ( .A(n5340), .B(n5341), .Z(n5187) );
  XNOR U5392 ( .A(n5338), .B(n5337), .Z(n5186) );
  XOR U5393 ( .A(n5343), .B(n5334), .Z(n5337) );
  XNOR U5394 ( .A(n5333), .B(n5344), .Z(n5334) );
  ANDN U5395 ( .A(n1426), .B(n3276), .Z(n5344) );
  XNOR U5396 ( .A(n5347), .B(n5345), .Z(n5346) );
  ANDN U5397 ( .A(n1426), .B(n3417), .Z(n5347) );
  XNOR U5398 ( .A(n5336), .B(n5335), .Z(n5343) );
  AND U5399 ( .A(n3274), .B(n1363), .Z(n5335) );
  XNOR U5400 ( .A(n5350), .B(n5351), .Z(n5336) );
  NAND U5401 ( .A(n4203), .B(n1363), .Z(n5351) );
  XNOR U5402 ( .A(n5349), .B(n5352), .Z(n5350) );
  ANDN U5403 ( .A(n1426), .B(n4205), .Z(n5352) );
  NAND U5404 ( .A(A[0]), .B(n5353), .Z(n5349) );
  NANDN U5405 ( .B(n1363), .A(n5354), .Z(n5353) );
  NANDN U5406 ( .B(n4208), .A(n1426), .Z(n5354) );
  IV U5407 ( .A(n5348), .Z(n1363) );
  XNOR U5408 ( .A(n5329), .B(n5330), .Z(n5338) );
  NANDN U5409 ( .B(n1228), .A(n4203), .Z(n5330) );
  XNOR U5410 ( .A(n5328), .B(n5357), .Z(n5329) );
  ANDN U5411 ( .A(n1298), .B(n4205), .Z(n5357) );
  NAND U5412 ( .A(A[0]), .B(n5358), .Z(n5328) );
  NAND U5413 ( .A(n5359), .B(n1228), .Z(n5358) );
  NANDN U5414 ( .B(n4208), .A(n1298), .Z(n5359) );
  XOR U5415 ( .A(n5362), .B(n5363), .Z(n5339) );
  XOR U5416 ( .A(n5364), .B(n3386), .Z(n3389) );
  XNOR U5417 ( .A(n3385), .B(n5365), .Z(n3386) );
  ANDN U5418 ( .A(n1788), .B(n1912), .Z(n5365) );
  XNOR U5419 ( .A(n4996), .B(A[16]), .Z(n4997) );
  ANDN U5420 ( .A(n5366), .B(n5367), .Z(n4996) );
  AND U5421 ( .A(n1910), .B(n1781), .Z(n3387) );
  IV U5422 ( .A(n2008), .Z(n1910) );
  XNOR U5423 ( .A(n5191), .B(n5192), .Z(n5197) );
  NAND U5424 ( .A(n2203), .B(n1597), .Z(n5192) );
  XNOR U5425 ( .A(n5190), .B(n5372), .Z(n5191) );
  ANDN U5426 ( .A(n1604), .B(n2205), .Z(n5372) );
  XNOR U5427 ( .A(n5376), .B(n5369), .Z(n5199) );
  XNOR U5428 ( .A(n5368), .B(n5377), .Z(n5369) );
  ANDN U5429 ( .A(n1788), .B(n2008), .Z(n5377) );
  ANDN U5430 ( .A(n5378), .B(n5379), .Z(n5366) );
  AND U5431 ( .A(n2006), .B(n1781), .Z(n5370) );
  IV U5432 ( .A(n2104), .Z(n2006) );
  XNOR U5433 ( .A(n5374), .B(n5375), .Z(n5217) );
  NAND U5434 ( .A(n2309), .B(n1597), .Z(n5375) );
  XNOR U5435 ( .A(n5373), .B(n5384), .Z(n5374) );
  ANDN U5436 ( .A(n1604), .B(n2311), .Z(n5384) );
  XNOR U5437 ( .A(n5388), .B(n5381), .Z(n5219) );
  XNOR U5438 ( .A(n5380), .B(n5389), .Z(n5381) );
  ANDN U5439 ( .A(n1788), .B(n2104), .Z(n5389) );
  XNOR U5440 ( .A(n5378), .B(A[14]), .Z(n5379) );
  ANDN U5441 ( .A(n5390), .B(n5391), .Z(n5378) );
  AND U5442 ( .A(n2102), .B(n1781), .Z(n5382) );
  IV U5443 ( .A(n2205), .Z(n2102) );
  XNOR U5444 ( .A(n5386), .B(n5387), .Z(n5237) );
  NAND U5445 ( .A(n2416), .B(n1597), .Z(n5387) );
  XNOR U5446 ( .A(n5385), .B(n5396), .Z(n5386) );
  ANDN U5447 ( .A(n1604), .B(n2418), .Z(n5396) );
  XNOR U5448 ( .A(n5400), .B(n5393), .Z(n5239) );
  XNOR U5449 ( .A(n5392), .B(n5401), .Z(n5393) );
  ANDN U5450 ( .A(n1788), .B(n2205), .Z(n5401) );
  ANDN U5451 ( .A(n5402), .B(n5403), .Z(n5390) );
  AND U5452 ( .A(n2203), .B(n1781), .Z(n5394) );
  IV U5453 ( .A(n2311), .Z(n2203) );
  XNOR U5454 ( .A(n5398), .B(n5399), .Z(n5257) );
  NAND U5455 ( .A(n2524), .B(n1597), .Z(n5399) );
  XNOR U5456 ( .A(n5397), .B(n5408), .Z(n5398) );
  ANDN U5457 ( .A(n1604), .B(n2526), .Z(n5408) );
  XNOR U5458 ( .A(n5412), .B(n5405), .Z(n5259) );
  XNOR U5459 ( .A(n5404), .B(n5413), .Z(n5405) );
  ANDN U5460 ( .A(n1788), .B(n2311), .Z(n5413) );
  XNOR U5461 ( .A(n5402), .B(A[12]), .Z(n5403) );
  ANDN U5462 ( .A(n5414), .B(n5415), .Z(n5402) );
  AND U5463 ( .A(n2309), .B(n1781), .Z(n5406) );
  IV U5464 ( .A(n2418), .Z(n2309) );
  XNOR U5465 ( .A(n5410), .B(n5411), .Z(n5277) );
  NAND U5466 ( .A(n2643), .B(n1597), .Z(n5411) );
  XNOR U5467 ( .A(n5409), .B(n5420), .Z(n5410) );
  ANDN U5468 ( .A(n1604), .B(n2645), .Z(n5420) );
  XOR U5469 ( .A(n5421), .B(n5422), .Z(n5409) );
  AND U5470 ( .A(n5423), .B(n5424), .Z(n5422) );
  XOR U5471 ( .A(n5425), .B(n5421), .Z(n5424) );
  XNOR U5472 ( .A(n5426), .B(n5417), .Z(n5279) );
  XNOR U5473 ( .A(n5416), .B(n5427), .Z(n5417) );
  ANDN U5474 ( .A(n1788), .B(n2418), .Z(n5427) );
  ANDN U5475 ( .A(n5428), .B(n5429), .Z(n5414) );
  AND U5476 ( .A(n2416), .B(n1781), .Z(n5418) );
  IV U5477 ( .A(n2526), .Z(n2416) );
  XNOR U5478 ( .A(n5423), .B(n5425), .Z(n5299) );
  NAND U5479 ( .A(n2763), .B(n1597), .Z(n5425) );
  XNOR U5480 ( .A(n5421), .B(n5434), .Z(n5423) );
  ANDN U5481 ( .A(n1604), .B(n2765), .Z(n5434) );
  XOR U5482 ( .A(n5435), .B(n5436), .Z(n5421) );
  AND U5483 ( .A(n5437), .B(n5438), .Z(n5436) );
  XOR U5484 ( .A(n5439), .B(n5435), .Z(n5438) );
  XNOR U5485 ( .A(n5440), .B(n5431), .Z(n5301) );
  XNOR U5486 ( .A(n5430), .B(n5441), .Z(n5431) );
  ANDN U5487 ( .A(n1788), .B(n2526), .Z(n5441) );
  XNOR U5488 ( .A(n5428), .B(A[10]), .Z(n5429) );
  ANDN U5489 ( .A(n5442), .B(n5443), .Z(n5428) );
  XOR U5490 ( .A(n5444), .B(n5445), .Z(n5430) );
  AND U5491 ( .A(n5446), .B(n5447), .Z(n5445) );
  XNOR U5492 ( .A(n5448), .B(n5444), .Z(n5447) );
  XOR U5493 ( .A(n5449), .B(n5432), .Z(n5440) );
  AND U5494 ( .A(n2524), .B(n1781), .Z(n5432) );
  IV U5495 ( .A(n2645), .Z(n2524) );
  IV U5496 ( .A(n5433), .Z(n5449) );
  XNOR U5497 ( .A(n5437), .B(n5439), .Z(n5323) );
  NAND U5498 ( .A(n2885), .B(n1597), .Z(n5439) );
  XNOR U5499 ( .A(n5435), .B(n5451), .Z(n5437) );
  ANDN U5500 ( .A(n1604), .B(n2887), .Z(n5451) );
  XNOR U5501 ( .A(n5455), .B(n5446), .Z(n5325) );
  XNOR U5502 ( .A(n5444), .B(n5456), .Z(n5446) );
  ANDN U5503 ( .A(n1788), .B(n2645), .Z(n5456) );
  ANDN U5504 ( .A(n5457), .B(n5458), .Z(n5442) );
  XOR U5505 ( .A(n5459), .B(n5460), .Z(n5444) );
  AND U5506 ( .A(n5461), .B(n5462), .Z(n5460) );
  XNOR U5507 ( .A(n5463), .B(n5459), .Z(n5462) );
  AND U5508 ( .A(n2643), .B(n1781), .Z(n5448) );
  IV U5509 ( .A(n2765), .Z(n2643) );
  XNOR U5510 ( .A(n5453), .B(n5454), .Z(n5341) );
  NAND U5511 ( .A(n3010), .B(n1597), .Z(n5454) );
  XNOR U5512 ( .A(n5452), .B(n5465), .Z(n5453) );
  ANDN U5513 ( .A(n1604), .B(n3012), .Z(n5465) );
  XNOR U5514 ( .A(n5469), .B(n5461), .Z(n5342) );
  XNOR U5515 ( .A(n5459), .B(n5470), .Z(n5461) );
  ANDN U5516 ( .A(n1788), .B(n2765), .Z(n5470) );
  AND U5517 ( .A(n2763), .B(n1781), .Z(n5463) );
  XNOR U5518 ( .A(n5474), .B(n5475), .Z(n5464) );
  AND U5519 ( .A(n5476), .B(n5477), .Z(n5475) );
  XNOR U5520 ( .A(n5472), .B(n5478), .Z(n5477) );
  XNOR U5521 ( .A(n5473), .B(n5474), .Z(n5478) );
  AND U5522 ( .A(n2885), .B(n1781), .Z(n5473) );
  XOR U5523 ( .A(n5471), .B(n5479), .Z(n5472) );
  ANDN U5524 ( .A(n1788), .B(n2887), .Z(n5479) );
  XNOR U5525 ( .A(n5467), .B(n5483), .Z(n5476) );
  XNOR U5526 ( .A(n5468), .B(n5474), .Z(n5483) );
  AND U5527 ( .A(n3142), .B(n1597), .Z(n5468) );
  XOR U5528 ( .A(n5466), .B(n5484), .Z(n5467) );
  ANDN U5529 ( .A(n1604), .B(n3144), .Z(n5484) );
  XOR U5530 ( .A(n5488), .B(n5489), .Z(n5474) );
  AND U5531 ( .A(n5490), .B(n5491), .Z(n5489) );
  XNOR U5532 ( .A(n5481), .B(n5492), .Z(n5491) );
  XNOR U5533 ( .A(n5482), .B(n5488), .Z(n5492) );
  AND U5534 ( .A(n3010), .B(n1781), .Z(n5482) );
  XOR U5535 ( .A(n5480), .B(n5493), .Z(n5481) );
  ANDN U5536 ( .A(n1788), .B(n3012), .Z(n5493) );
  XNOR U5537 ( .A(n5486), .B(n5497), .Z(n5490) );
  XNOR U5538 ( .A(n5487), .B(n5488), .Z(n5497) );
  AND U5539 ( .A(n3274), .B(n1597), .Z(n5487) );
  XOR U5540 ( .A(n5485), .B(n5498), .Z(n5486) );
  ANDN U5541 ( .A(n1604), .B(n3276), .Z(n5498) );
  XOR U5542 ( .A(n5499), .B(n5500), .Z(n5485) );
  ANDN U5543 ( .A(n5501), .B(n5502), .Z(n5500) );
  XNOR U5544 ( .A(n5503), .B(n5499), .Z(n5501) );
  XOR U5545 ( .A(n5504), .B(n5505), .Z(n5488) );
  AND U5546 ( .A(n5506), .B(n5507), .Z(n5505) );
  XNOR U5547 ( .A(n5495), .B(n5508), .Z(n5507) );
  XNOR U5548 ( .A(n5496), .B(n5504), .Z(n5508) );
  AND U5549 ( .A(n3142), .B(n1781), .Z(n5496) );
  XOR U5550 ( .A(n5494), .B(n5509), .Z(n5495) );
  ANDN U5551 ( .A(n1788), .B(n3144), .Z(n5509) );
  XNOR U5552 ( .A(n5502), .B(n5513), .Z(n5506) );
  XNOR U5553 ( .A(n5503), .B(n5504), .Z(n5513) );
  AND U5554 ( .A(n3415), .B(n1597), .Z(n5503) );
  XOR U5555 ( .A(n5499), .B(n5514), .Z(n5502) );
  ANDN U5556 ( .A(n1604), .B(n3417), .Z(n5514) );
  XNOR U5557 ( .A(n5519), .B(n5511), .Z(n5363) );
  XNOR U5558 ( .A(n5510), .B(n5520), .Z(n5511) );
  ANDN U5559 ( .A(n1788), .B(n3276), .Z(n5520) );
  XNOR U5560 ( .A(n5523), .B(n5521), .Z(n5522) );
  ANDN U5561 ( .A(n1788), .B(n3417), .Z(n5523) );
  XNOR U5562 ( .A(n5518), .B(n5512), .Z(n5519) );
  AND U5563 ( .A(n3274), .B(n1781), .Z(n5512) );
  XNOR U5564 ( .A(n5516), .B(n5517), .Z(n5362) );
  NAND U5565 ( .A(n4203), .B(n1597), .Z(n5517) );
  XNOR U5566 ( .A(n5515), .B(n5527), .Z(n5516) );
  ANDN U5567 ( .A(n1604), .B(n4205), .Z(n5527) );
  NAND U5568 ( .A(A[0]), .B(n5528), .Z(n5515) );
  NANDN U5569 ( .B(n1597), .A(n5529), .Z(n5528) );
  NANDN U5570 ( .B(n4208), .A(n1604), .Z(n5529) );
  IV U5571 ( .A(n1523), .Z(n1597) );
  XNOR U5572 ( .A(n5525), .B(n5526), .Z(n5518) );
  NAND U5573 ( .A(n4203), .B(n1781), .Z(n5526) );
  XNOR U5574 ( .A(n5524), .B(n5532), .Z(n5525) );
  ANDN U5575 ( .A(n1788), .B(n4205), .Z(n5532) );
  NAND U5576 ( .A(A[0]), .B(n5533), .Z(n5524) );
  NANDN U5577 ( .B(n1781), .A(n5534), .Z(n5533) );
  NANDN U5578 ( .B(n4208), .A(n1788), .Z(n5534) );
  IV U5579 ( .A(n1688), .Z(n1781) );
  XNOR U5580 ( .A(n3398), .B(n3397), .Z(n3374) );
  XOR U5581 ( .A(n5537), .B(n3406), .Z(n3397) );
  XNOR U5582 ( .A(n3394), .B(n3395), .Z(n3406) );
  NANDN U5583 ( .B(n1041), .A(n3010), .Z(n3395) );
  XNOR U5584 ( .A(n3393), .B(n5538), .Z(n3394) );
  ANDN U5585 ( .A(n1082), .B(n3012), .Z(n5538) );
  XOR U5586 ( .A(n3405), .B(n3396), .Z(n5537) );
  XOR U5587 ( .A(n5542), .B(n5543), .Z(n3396) );
  XOR U5588 ( .A(n5544), .B(n3402), .Z(n3405) );
  XNOR U5589 ( .A(n3401), .B(n5545), .Z(n3402) );
  ANDN U5590 ( .A(n1189), .B(n2765), .Z(n5545) );
  XNOR U5591 ( .A(n5457), .B(A[8]), .Z(n5458) );
  ANDN U5592 ( .A(n5546), .B(n5547), .Z(n5457) );
  AND U5593 ( .A(n2763), .B(n1135), .Z(n3403) );
  IV U5594 ( .A(n2887), .Z(n2763) );
  XNOR U5595 ( .A(n5551), .B(n5552), .Z(n3404) );
  AND U5596 ( .A(n5553), .B(n5554), .Z(n5552) );
  XNOR U5597 ( .A(n5549), .B(n5555), .Z(n5554) );
  XNOR U5598 ( .A(n5550), .B(n5551), .Z(n5555) );
  AND U5599 ( .A(n2885), .B(n1135), .Z(n5550) );
  IV U5600 ( .A(n3012), .Z(n2885) );
  XOR U5601 ( .A(n5548), .B(n5556), .Z(n5549) );
  ANDN U5602 ( .A(n1189), .B(n2887), .Z(n5556) );
  ANDN U5603 ( .A(n5557), .B(n5558), .Z(n5546) );
  XNOR U5604 ( .A(n5540), .B(n5562), .Z(n5553) );
  XNOR U5605 ( .A(n5541), .B(n5551), .Z(n5562) );
  ANDN U5606 ( .A(n3142), .B(n1041), .Z(n5541) );
  XOR U5607 ( .A(n5539), .B(n5563), .Z(n5540) );
  ANDN U5608 ( .A(n1082), .B(n3144), .Z(n5563) );
  XOR U5609 ( .A(n5567), .B(n5568), .Z(n5551) );
  AND U5610 ( .A(n5569), .B(n5570), .Z(n5568) );
  XNOR U5611 ( .A(n5560), .B(n5571), .Z(n5570) );
  XNOR U5612 ( .A(n5561), .B(n5567), .Z(n5571) );
  AND U5613 ( .A(n3010), .B(n1135), .Z(n5561) );
  IV U5614 ( .A(n3144), .Z(n3010) );
  XOR U5615 ( .A(n5559), .B(n5572), .Z(n5560) );
  ANDN U5616 ( .A(n1189), .B(n3012), .Z(n5572) );
  XNOR U5617 ( .A(n5557), .B(A[6]), .Z(n5558) );
  ANDN U5618 ( .A(n5573), .B(n5574), .Z(n5557) );
  XNOR U5619 ( .A(n5565), .B(n5578), .Z(n5569) );
  XNOR U5620 ( .A(n5566), .B(n5567), .Z(n5578) );
  ANDN U5621 ( .A(n3274), .B(n1041), .Z(n5566) );
  XOR U5622 ( .A(n5564), .B(n5579), .Z(n5565) );
  ANDN U5623 ( .A(n1082), .B(n3276), .Z(n5579) );
  XOR U5624 ( .A(n5580), .B(n5581), .Z(n5564) );
  ANDN U5625 ( .A(n5582), .B(n5583), .Z(n5581) );
  XNOR U5626 ( .A(n5584), .B(n5580), .Z(n5582) );
  XOR U5627 ( .A(n5585), .B(n5586), .Z(n5567) );
  AND U5628 ( .A(n5587), .B(n5588), .Z(n5586) );
  XNOR U5629 ( .A(n5576), .B(n5589), .Z(n5588) );
  XNOR U5630 ( .A(n5577), .B(n5585), .Z(n5589) );
  AND U5631 ( .A(n3142), .B(n1135), .Z(n5577) );
  XOR U5632 ( .A(n5575), .B(n5590), .Z(n5576) );
  ANDN U5633 ( .A(n1189), .B(n3144), .Z(n5590) );
  ANDN U5634 ( .A(n5591), .B(n5592), .Z(n5573) );
  XNOR U5635 ( .A(n5583), .B(n5596), .Z(n5587) );
  XNOR U5636 ( .A(n5584), .B(n5585), .Z(n5596) );
  ANDN U5637 ( .A(n3415), .B(n1041), .Z(n5584) );
  XOR U5638 ( .A(n5580), .B(n5597), .Z(n5583) );
  ANDN U5639 ( .A(n1082), .B(n3417), .Z(n5597) );
  XNOR U5640 ( .A(n5602), .B(n5594), .Z(n5543) );
  XNOR U5641 ( .A(n5593), .B(n5603), .Z(n5594) );
  ANDN U5642 ( .A(n1189), .B(n3276), .Z(n5603) );
  XNOR U5643 ( .A(n5606), .B(n5604), .Z(n5605) );
  ANDN U5644 ( .A(n1189), .B(n3417), .Z(n5606) );
  XNOR U5645 ( .A(n5601), .B(n5595), .Z(n5602) );
  AND U5646 ( .A(n3274), .B(n1135), .Z(n5595) );
  XNOR U5647 ( .A(n5599), .B(n5600), .Z(n5542) );
  NANDN U5648 ( .B(n1041), .A(n4203), .Z(n5600) );
  XNOR U5649 ( .A(n5598), .B(n5611), .Z(n5599) );
  ANDN U5650 ( .A(n1082), .B(n4205), .Z(n5611) );
  NAND U5651 ( .A(A[0]), .B(n5612), .Z(n5598) );
  NAND U5652 ( .A(n5613), .B(n1041), .Z(n5612) );
  NANDN U5653 ( .B(n4208), .A(n1082), .Z(n5613) );
  XNOR U5654 ( .A(n5609), .B(n5610), .Z(n5601) );
  NAND U5655 ( .A(n4203), .B(n1135), .Z(n5610) );
  XNOR U5656 ( .A(n5608), .B(n5616), .Z(n5609) );
  ANDN U5657 ( .A(n1189), .B(n4205), .Z(n5616) );
  NAND U5658 ( .A(A[0]), .B(n5617), .Z(n5608) );
  NANDN U5659 ( .B(n1135), .A(n5618), .Z(n5617) );
  NANDN U5660 ( .B(n4208), .A(n1189), .Z(n5618) );
  IV U5661 ( .A(n5607), .Z(n1135) );
  XOR U5662 ( .A(n3414), .B(n3413), .Z(n3398) );
  XOR U5663 ( .A(n5621), .B(n3410), .Z(n3413) );
  XNOR U5664 ( .A(n3409), .B(n5622), .Z(n3410) );
  ANDN U5665 ( .A(n1014), .B(n3276), .Z(n5622) );
  IV U5666 ( .A(n3142), .Z(n3276) );
  XNOR U5667 ( .A(n5591), .B(A[4]), .Z(n5592) );
  ANDN U5668 ( .A(n5623), .B(n5624), .Z(n5591) );
  XNOR U5669 ( .A(n5627), .B(n5625), .Z(n5626) );
  ANDN U5670 ( .A(n1014), .B(n3417), .Z(n5627) );
  IV U5671 ( .A(n3274), .Z(n3417) );
  IV U5672 ( .A(n4205), .Z(n3415) );
  XNOR U5673 ( .A(n3412), .B(n3411), .Z(n5621) );
  AND U5674 ( .A(n3274), .B(n973), .Z(n3411) );
  ANDN U5675 ( .A(n5632), .B(n5633), .Z(n5623) );
  XNOR U5676 ( .A(n5630), .B(n5631), .Z(n3412) );
  NAND U5677 ( .A(n4203), .B(n973), .Z(n5631) );
  XNOR U5678 ( .A(n5629), .B(n5634), .Z(n5630) );
  ANDN U5679 ( .A(n1014), .B(n4205), .Z(n5634) );
  NAND U5680 ( .A(A[0]), .B(n5635), .Z(n5629) );
  NANDN U5681 ( .B(n973), .A(n5636), .Z(n5635) );
  NANDN U5682 ( .B(n4208), .A(n1014), .Z(n5636) );
  IV U5683 ( .A(n5628), .Z(n973) );
  XOR U5684 ( .A(n3421), .B(n3420), .Z(n3414) );
  NAND U5685 ( .A(n4203), .B(n917), .Z(n3420) );
  IV U5686 ( .A(n4208), .Z(n4203) );
  XOR U5687 ( .A(n3419), .B(n5639), .Z(n3421) );
  ANDN U5688 ( .A(n948), .B(n4205), .Z(n5639) );
  XNOR U5689 ( .A(n5632), .B(A[2]), .Z(n5633) );
  NOR U5690 ( .A(A[0]), .B(n5640), .Z(n5632) );
  NANDN U5691 ( .B(n917), .A(n5642), .Z(n5641) );
  NANDN U5692 ( .B(n4208), .A(n948), .Z(n5642) );
  XOR U5693 ( .A(A[0]), .B(A[1]), .Z(n5640) );
  AND U5694 ( .A(n5644), .B(n5643), .Z(n917) );
  ANDN U5695 ( .A(X[31]), .B(n5645), .Z(n5644) );
  NANDN U5696 ( .B(n5646), .A(n5638), .Z(n5645) );
  XNOR U5697 ( .A(n5646), .B(X[29]), .Z(n5638) );
  NAND U5698 ( .A(n5637), .B(n5647), .Z(n5646) );
  XOR U5699 ( .A(n5647), .B(X[28]), .Z(n5637) );
  ANDN U5700 ( .A(n5614), .B(n5648), .Z(n5647) );
  XNOR U5701 ( .A(n5648), .B(X[27]), .Z(n5614) );
  NAND U5702 ( .A(n5615), .B(n5649), .Z(n5648) );
  XOR U5703 ( .A(n5649), .B(X[26]), .Z(n5615) );
  ANDN U5704 ( .A(n5620), .B(n5650), .Z(n5649) );
  XNOR U5705 ( .A(n5650), .B(X[25]), .Z(n5620) );
  NAND U5706 ( .A(n5619), .B(n5651), .Z(n5650) );
  XOR U5707 ( .A(n5651), .B(X[24]), .Z(n5619) );
  ANDN U5708 ( .A(n5360), .B(n5652), .Z(n5651) );
  XNOR U5709 ( .A(n5652), .B(X[23]), .Z(n5360) );
  NAND U5710 ( .A(n5361), .B(n5653), .Z(n5652) );
  XOR U5711 ( .A(n5653), .B(X[22]), .Z(n5361) );
  ANDN U5712 ( .A(n5356), .B(n5654), .Z(n5653) );
  XNOR U5713 ( .A(n5654), .B(X[21]), .Z(n5356) );
  NAND U5714 ( .A(n5355), .B(n5655), .Z(n5654) );
  XOR U5715 ( .A(n5655), .B(X[20]), .Z(n5355) );
  ANDN U5716 ( .A(n5531), .B(n5656), .Z(n5655) );
  XNOR U5717 ( .A(n5656), .B(X[19]), .Z(n5531) );
  NAND U5718 ( .A(n5530), .B(n5657), .Z(n5656) );
  XOR U5719 ( .A(n5657), .B(X[18]), .Z(n5530) );
  ANDN U5720 ( .A(n5536), .B(n5658), .Z(n5657) );
  XNOR U5721 ( .A(n5658), .B(X[17]), .Z(n5536) );
  NAND U5722 ( .A(n5535), .B(n5659), .Z(n5658) );
  XOR U5723 ( .A(n5659), .B(X[16]), .Z(n5535) );
  ANDN U5724 ( .A(n4233), .B(n5660), .Z(n5659) );
  XNOR U5725 ( .A(n5660), .B(X[15]), .Z(n4233) );
  NAND U5726 ( .A(n4232), .B(n5661), .Z(n5660) );
  XOR U5727 ( .A(n5661), .B(X[14]), .Z(n4232) );
  ANDN U5728 ( .A(n4228), .B(n5662), .Z(n5661) );
  XNOR U5729 ( .A(n5662), .B(X[13]), .Z(n4228) );
  NAND U5730 ( .A(n4227), .B(n5663), .Z(n5662) );
  XOR U5731 ( .A(n5663), .B(X[12]), .Z(n4227) );
  ANDN U5732 ( .A(n4210), .B(n5664), .Z(n5663) );
  XNOR U5733 ( .A(n5664), .B(X[11]), .Z(n4210) );
  NAND U5734 ( .A(n4209), .B(n5665), .Z(n5664) );
  XOR U5735 ( .A(n5665), .B(X[10]), .Z(n4209) );
  ANDN U5736 ( .A(n4215), .B(n5666), .Z(n5665) );
  XNOR U5737 ( .A(n5666), .B(X[9]), .Z(n4215) );
  NAND U5738 ( .A(n4214), .B(n5667), .Z(n5666) );
  XOR U5739 ( .A(n5667), .B(X[8]), .Z(n4214) );
  ANDN U5740 ( .A(n4739), .B(n5668), .Z(n5667) );
  XNOR U5741 ( .A(n5668), .B(X[7]), .Z(n4739) );
  NAND U5742 ( .A(n4738), .B(n5669), .Z(n5668) );
  XOR U5743 ( .A(n5669), .B(X[6]), .Z(n4738) );
  ANDN U5744 ( .A(n4734), .B(n5670), .Z(n5669) );
  XNOR U5745 ( .A(n5670), .B(X[5]), .Z(n4734) );
  NAND U5746 ( .A(n4733), .B(n5671), .Z(n5670) );
  XOR U5747 ( .A(n5671), .B(X[4]), .Z(n4733) );
  ANDN U5748 ( .A(n5168), .B(n5672), .Z(n5671) );
  XNOR U5749 ( .A(n5672), .B(X[3]), .Z(n5168) );
  NAND U5750 ( .A(n5167), .B(n5673), .Z(n5672) );
  XOR U5751 ( .A(n5673), .B(X[2]), .Z(n5167) );
  NOR U5752 ( .A(n5172), .B(X[0]), .Z(n5673) );
  XOR U5753 ( .A(X[0]), .B(X[1]), .Z(n5172) );
endmodule

