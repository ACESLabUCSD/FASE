
module MxM_W32_N100 ( clk, rst, A, X, Y );
  input [31:0] A;
  input [31:0] X;
  output [31:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, \add_25/carry[6] ,
         \add_25/carry[5] , \add_25/carry[4] , \add_25/carry[3] ,
         \add_25/carry[2] , n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628;
  wire   [31:0] Y0;
  wire   [6:0] n;

  DFF \n_reg[0]  ( .D(n357), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n356), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n355), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n354), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n353), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n352), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n351), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \Y0_reg[0]  ( .D(n350), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n349), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n348), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n347), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n346), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n345), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n344), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n343), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y0_reg[8]  ( .D(n342), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[8]) );
  DFF \Y0_reg[9]  ( .D(n341), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[9]) );
  DFF \Y0_reg[10]  ( .D(n340), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[10]) );
  DFF \Y0_reg[11]  ( .D(n339), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[11]) );
  DFF \Y0_reg[12]  ( .D(n338), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[12]) );
  DFF \Y0_reg[13]  ( .D(n337), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[13]) );
  DFF \Y0_reg[14]  ( .D(n336), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[14]) );
  DFF \Y0_reg[15]  ( .D(n335), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[15]) );
  DFF \Y0_reg[16]  ( .D(n334), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[16]) );
  DFF \Y0_reg[17]  ( .D(n333), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[17]) );
  DFF \Y0_reg[18]  ( .D(n332), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[18]) );
  DFF \Y0_reg[19]  ( .D(n331), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[19]) );
  DFF \Y0_reg[20]  ( .D(n330), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[20]) );
  DFF \Y0_reg[21]  ( .D(n329), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[21]) );
  DFF \Y0_reg[22]  ( .D(n328), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[22]) );
  DFF \Y0_reg[23]  ( .D(n327), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[23]) );
  DFF \Y0_reg[24]  ( .D(n326), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[24]) );
  DFF \Y0_reg[25]  ( .D(n325), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[25]) );
  DFF \Y0_reg[26]  ( .D(n324), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[26]) );
  DFF \Y0_reg[27]  ( .D(n323), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[27]) );
  DFF \Y0_reg[28]  ( .D(n322), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[28]) );
  DFF \Y0_reg[29]  ( .D(n321), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[29]) );
  DFF \Y0_reg[30]  ( .D(n320), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[30]) );
  DFF \Y0_reg[31]  ( .D(n319), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[31]) );
  DFF \Y_reg[31]  ( .D(n318), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[31]) );
  DFF \Y_reg[30]  ( .D(n317), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[30]) );
  DFF \Y_reg[29]  ( .D(n316), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[29]) );
  DFF \Y_reg[28]  ( .D(n315), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[28]) );
  DFF \Y_reg[27]  ( .D(n314), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[27]) );
  DFF \Y_reg[26]  ( .D(n313), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[26]) );
  DFF \Y_reg[25]  ( .D(n312), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[25]) );
  DFF \Y_reg[24]  ( .D(n311), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[24]) );
  DFF \Y_reg[23]  ( .D(n310), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[23]) );
  DFF \Y_reg[22]  ( .D(n309), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[22]) );
  DFF \Y_reg[21]  ( .D(n308), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[21]) );
  DFF \Y_reg[20]  ( .D(n307), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[20]) );
  DFF \Y_reg[19]  ( .D(n306), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[19]) );
  DFF \Y_reg[18]  ( .D(n305), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[18]) );
  DFF \Y_reg[17]  ( .D(n304), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[17]) );
  DFF \Y_reg[16]  ( .D(n303), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[16]) );
  DFF \Y_reg[15]  ( .D(n302), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[15]) );
  DFF \Y_reg[14]  ( .D(n301), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[14]) );
  DFF \Y_reg[13]  ( .D(n300), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[13]) );
  DFF \Y_reg[12]  ( .D(n299), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[12]) );
  DFF \Y_reg[11]  ( .D(n298), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[11]) );
  DFF \Y_reg[10]  ( .D(n297), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[10]) );
  DFF \Y_reg[9]  ( .D(n296), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[9]) );
  DFF \Y_reg[8]  ( .D(n295), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[8]) );
  DFF \Y_reg[7]  ( .D(n294), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n293), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n292), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n291), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n290), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n289), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n288), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n287), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  MUX U360 ( .IN0(n4059), .IN1(n358), .SEL(n4060), .F(n4013) );
  IV U361 ( .A(n4061), .Z(n358) );
  MUX U362 ( .IN0(n3887), .IN1(n3889), .SEL(n3888), .F(n3841) );
  MUX U363 ( .IN0(n4660), .IN1(n4662), .SEL(n4661), .F(n4636) );
  MUX U364 ( .IN0(n3712), .IN1(n3714), .SEL(n3713), .F(n3666) );
  XNOR U365 ( .A(n4648), .B(n4647), .Z(n4663) );
  XNOR U366 ( .A(n5031), .B(n5029), .Z(n5036) );
  MUX U367 ( .IN0(n3616), .IN1(n3618), .SEL(n3617), .F(n3573) );
  MUX U368 ( .IN0(n5364), .IN1(n5366), .SEL(n5365), .F(n5352) );
  MUX U369 ( .IN0(n5222), .IN1(n359), .SEL(n5223), .F(n5202) );
  IV U370 ( .A(n5224), .Z(n359) );
  MUX U371 ( .IN0(n5371), .IN1(n360), .SEL(n5372), .F(n5359) );
  IV U372 ( .A(n5373), .Z(n360) );
  MUX U373 ( .IN0(n4581), .IN1(n361), .SEL(n4582), .F(n4561) );
  IV U374 ( .A(n4583), .Z(n361) );
  XNOR U375 ( .A(n3569), .B(n3568), .Z(n3605) );
  MUX U376 ( .IN0(n4986), .IN1(n362), .SEL(n4987), .F(n4976) );
  IV U377 ( .A(n4988), .Z(n362) );
  XNOR U378 ( .A(n3594), .B(n3592), .Z(n3629) );
  XNOR U379 ( .A(n4757), .B(n4755), .Z(n4764) );
  NANDN U380 ( .B(n1648), .A(n3370), .Z(n375) );
  MUX U381 ( .IN0(n3446), .IN1(n3448), .SEL(n3447), .F(n3407) );
  MUX U382 ( .IN0(n3439), .IN1(n363), .SEL(n3440), .F(n3400) );
  IV U383 ( .A(n3441), .Z(n363) );
  MUX U384 ( .IN0(n3451), .IN1(n3453), .SEL(n3452), .F(n3380) );
  MUX U385 ( .IN0(n1359), .IN1(n364), .SEL(n1360), .F(n1290) );
  IV U386 ( .A(n1361), .Z(n364) );
  MUX U387 ( .IN0(n1656), .IN1(n1658), .SEL(n1657), .F(n1572) );
  MUX U388 ( .IN0(n1711), .IN1(n365), .SEL(n1712), .F(n1620) );
  IV U389 ( .A(n1713), .Z(n365) );
  MUX U390 ( .IN0(n1759), .IN1(n366), .SEL(n1760), .F(n1664) );
  IV U391 ( .A(n1761), .Z(n366) );
  MUX U392 ( .IN0(n1864), .IN1(n367), .SEL(n1865), .F(n1767) );
  IV U393 ( .A(n1866), .Z(n367) );
  MUX U394 ( .IN0(n2123), .IN1(n2125), .SEL(n2124), .F(n2022) );
  MUX U395 ( .IN0(n2239), .IN1(n368), .SEL(n2240), .F(n2131) );
  IV U396 ( .A(n2241), .Z(n368) );
  MUX U397 ( .IN0(n2412), .IN1(n369), .SEL(n2413), .F(n2303) );
  IV U398 ( .A(n2414), .Z(n369) );
  MUX U399 ( .IN0(A[29]), .IN1(n4733), .SEL(A[31]), .F(n370) );
  IV U400 ( .A(n370), .Z(n983) );
  MUX U401 ( .IN0(n371), .IN1(n4721), .SEL(A[31]), .F(n939) );
  IV U402 ( .A(A[30]), .Z(n371) );
  MUX U403 ( .IN0(n5283), .IN1(n5285), .SEL(n5284), .F(n5259) );
  MUX U404 ( .IN0(n5033), .IN1(n5035), .SEL(n5034), .F(n5018) );
  XNOR U405 ( .A(n5405), .B(n5403), .Z(n5410) );
  MUX U406 ( .IN0(n4616), .IN1(n4618), .SEL(n4617), .F(n4596) );
  MUX U407 ( .IN0(n4621), .IN1(n372), .SEL(n4622), .F(n4601) );
  IV U408 ( .A(n4623), .Z(n372) );
  XNOR U409 ( .A(n5271), .B(n5270), .Z(n5286) );
  MUX U410 ( .IN0(n5352), .IN1(n5354), .SEL(n5353), .F(n5340) );
  MUX U411 ( .IN0(n5202), .IN1(n373), .SEL(n5203), .F(n5182) );
  IV U412 ( .A(n5204), .Z(n373) );
  MUX U413 ( .IN0(n5359), .IN1(n374), .SEL(n5360), .F(n5347) );
  IV U414 ( .A(n5361), .Z(n374) );
  MUX U415 ( .IN0(n3531), .IN1(n3533), .SEL(n3532), .F(n3486) );
  XNOR U416 ( .A(n4989), .B(n4988), .Z(n4994) );
  MUX U417 ( .IN0(n4981), .IN1(n4983), .SEL(n4982), .F(n4971) );
  MUX U418 ( .IN0(n5476), .IN1(n375), .SEL(n5477), .F(n5465) );
  XNOR U419 ( .A(n3482), .B(n3481), .Z(n3520) );
  MUX U420 ( .IN0(n4966), .IN1(n376), .SEL(n4967), .F(n4953) );
  IV U421 ( .A(n4968), .Z(n376) );
  MUX U422 ( .IN0(n3400), .IN1(n377), .SEL(n3401), .F(n3270) );
  IV U423 ( .A(n3402), .Z(n377) );
  MUX U424 ( .IN0(n1511), .IN1(n378), .SEL(n1512), .F(n1431) );
  IV U425 ( .A(n1513), .Z(n378) );
  MUX U426 ( .IN0(n1572), .IN1(n1574), .SEL(n1573), .F(n1491) );
  MUX U427 ( .IN0(n1629), .IN1(n1631), .SEL(n1630), .F(n1547) );
  MUX U428 ( .IN0(n1944), .IN1(n1946), .SEL(n1945), .F(n1848) );
  MUX U429 ( .IN0(n1952), .IN1(n379), .SEL(n1953), .F(n1856) );
  IV U430 ( .A(n1954), .Z(n379) );
  MUX U431 ( .IN0(n1960), .IN1(n380), .SEL(n1961), .F(n1864) );
  IV U432 ( .A(n1962), .Z(n380) );
  MUX U433 ( .IN0(n2007), .IN1(n381), .SEL(n2008), .F(n1907) );
  IV U434 ( .A(n2009), .Z(n381) );
  MUX U435 ( .IN0(n2204), .IN1(n2206), .SEL(n2205), .F(n2096) );
  MUX U436 ( .IN0(n2346), .IN1(n382), .SEL(n2347), .F(n2239) );
  IV U437 ( .A(n2348), .Z(n382) );
  MUX U438 ( .IN0(n2526), .IN1(n383), .SEL(n2527), .F(n2412) );
  IV U439 ( .A(n2528), .Z(n383) );
  MUX U440 ( .IN0(n3152), .IN1(n384), .SEL(n3153), .F(n3027) );
  IV U441 ( .A(n3154), .Z(n384) );
  MUX U442 ( .IN0(n1059), .IN1(n385), .SEL(n1060), .F(n1013) );
  IV U443 ( .A(n1061), .Z(n385) );
  MUX U444 ( .IN0(n3303), .IN1(n3305), .SEL(n3304), .F(n3168) );
  MUX U445 ( .IN0(n386), .IN1(n1094), .SEL(n1093), .F(n1056) );
  IV U446 ( .A(n1092), .Z(n386) );
  MUX U447 ( .IN0(n4067), .IN1(n4069), .SEL(n4068), .F(n4023) );
  MUX U448 ( .IN0(n5045), .IN1(n5047), .SEL(n5046), .F(n5033) );
  XNOR U449 ( .A(n5043), .B(n5042), .Z(n5048) );
  MUX U450 ( .IN0(n5237), .IN1(n5239), .SEL(n5238), .F(n5217) );
  MUX U451 ( .IN0(n5385), .IN1(n387), .SEL(n5386), .F(n5371) );
  IV U452 ( .A(n5387), .Z(n387) );
  MUX U453 ( .IN0(n4596), .IN1(n4598), .SEL(n4597), .F(n4576) );
  MUX U454 ( .IN0(n4601), .IN1(n388), .SEL(n4602), .F(n4581) );
  IV U455 ( .A(n4603), .Z(n388) );
  MUX U456 ( .IN0(n3580), .IN1(n3582), .SEL(n3581), .F(n3536) );
  XNOR U457 ( .A(n5205), .B(n5204), .Z(n5220) );
  MUX U458 ( .IN0(n5340), .IN1(n5342), .SEL(n5341), .F(n5328) );
  XNOR U459 ( .A(n5350), .B(n5349), .Z(n5355) );
  NANDN U460 ( .B(n2404), .A(n3370), .Z(n401) );
  MUX U461 ( .IN0(n4976), .IN1(n389), .SEL(n4977), .F(n4966) );
  IV U462 ( .A(n4978), .Z(n389) );
  MUX U463 ( .IN0(n4971), .IN1(n4973), .SEL(n4972), .F(n4961) );
  XNOR U464 ( .A(n3442), .B(n3441), .Z(n3475) );
  MUX U465 ( .IN0(n1751), .IN1(n1753), .SEL(n1752), .F(n1656) );
  MUX U466 ( .IN0(n2048), .IN1(n390), .SEL(n2049), .F(n1952) );
  IV U467 ( .A(n2050), .Z(n390) );
  MUX U468 ( .IN0(n2056), .IN1(n391), .SEL(n2057), .F(n1960) );
  IV U469 ( .A(n2058), .Z(n391) );
  MUX U470 ( .IN0(n2014), .IN1(n2016), .SEL(n2015), .F(n1916) );
  MUX U471 ( .IN0(n2022), .IN1(n2024), .SEL(n2023), .F(n1924) );
  MUX U472 ( .IN0(n2108), .IN1(n392), .SEL(n2109), .F(n2007) );
  IV U473 ( .A(n2110), .Z(n392) );
  MUX U474 ( .IN0(n2141), .IN1(n2143), .SEL(n2142), .F(n2040) );
  MUX U475 ( .IN0(n2312), .IN1(n2314), .SEL(n2313), .F(n2204) );
  MUX U476 ( .IN0(n2454), .IN1(n393), .SEL(n2455), .F(n2346) );
  IV U477 ( .A(n2456), .Z(n393) );
  MUX U478 ( .IN0(n2622), .IN1(n2624), .SEL(n2623), .F(n2503) );
  MUX U479 ( .IN0(n2760), .IN1(n394), .SEL(n2761), .F(n2640) );
  IV U480 ( .A(n2762), .Z(n394) );
  MUX U481 ( .IN0(n3286), .IN1(n395), .SEL(n3287), .F(n3152) );
  IV U482 ( .A(n3288), .Z(n395) );
  MUX U483 ( .IN0(n1085), .IN1(n1087), .SEL(n1086), .F(n1043) );
  MUX U484 ( .IN0(n975), .IN1(n396), .SEL(n976), .F(n929) );
  IV U485 ( .A(n977), .Z(n396) );
  MUX U486 ( .IN0(n397), .IN1(n1321), .SEL(n1320), .F(n1256) );
  IV U487 ( .A(n1319), .Z(n397) );
  MUX U488 ( .IN0(n5407), .IN1(n5409), .SEL(n5408), .F(n5390) );
  MUX U489 ( .IN0(n5288), .IN1(n398), .SEL(n5289), .F(n5266) );
  IV U490 ( .A(n5290), .Z(n398) );
  MUX U491 ( .IN0(n5106), .IN1(n5108), .SEL(n5107), .F(n5090) );
  MUX U492 ( .IN0(n5217), .IN1(n5219), .SEL(n5218), .F(n5197) );
  MUX U493 ( .IN0(n4991), .IN1(n4993), .SEL(n4992), .F(n4981) );
  XNOR U494 ( .A(n4773), .B(n4772), .Z(n4780) );
  MUX U495 ( .IN0(n4556), .IN1(n4558), .SEL(n4557), .F(n4536) );
  XNOR U496 ( .A(n4584), .B(n4583), .Z(n4599) );
  MUX U497 ( .IN0(n5182), .IN1(n399), .SEL(n5183), .F(n5162) );
  IV U498 ( .A(n5184), .Z(n399) );
  MUX U499 ( .IN0(n5347), .IN1(n400), .SEL(n5348), .F(n5335) );
  IV U500 ( .A(n5349), .Z(n400) );
  MUX U501 ( .IN0(n4152), .IN1(n401), .SEL(n4153), .F(n4141) );
  MUX U502 ( .IN0(n5328), .IN1(n5330), .SEL(n5329), .F(n5145) );
  MUX U503 ( .IN0(n4517), .IN1(n402), .SEL(n4518), .F(n4496) );
  IV U504 ( .A(n4519), .Z(n402) );
  XNOR U505 ( .A(n4969), .B(n4968), .Z(n4974) );
  MUX U506 ( .IN0(n3407), .IN1(n3409), .SEL(n3408), .F(n3277) );
  MUX U507 ( .IN0(n1820), .IN1(n1822), .SEL(n1821), .F(n1718) );
  MUX U508 ( .IN0(n1856), .IN1(n403), .SEL(n1857), .F(n1759) );
  IV U509 ( .A(n1858), .Z(n403) );
  MUX U510 ( .IN0(n1848), .IN1(n1850), .SEL(n1849), .F(n1751) );
  MUX U511 ( .IN0(n2157), .IN1(n404), .SEL(n2158), .F(n2056) );
  IV U512 ( .A(n2159), .Z(n404) );
  MUX U513 ( .IN0(n2330), .IN1(n2332), .SEL(n2331), .F(n2223) );
  MUX U514 ( .IN0(n2323), .IN1(n405), .SEL(n2324), .F(n2216) );
  IV U515 ( .A(n2325), .Z(n405) );
  MUX U516 ( .IN0(n2362), .IN1(n406), .SEL(n2363), .F(n2255) );
  IV U517 ( .A(n2364), .Z(n406) );
  MUX U518 ( .IN0(n2419), .IN1(n2421), .SEL(n2420), .F(n2312) );
  MUX U519 ( .IN0(n2573), .IN1(n407), .SEL(n2574), .F(n2454) );
  IV U520 ( .A(n2575), .Z(n407) );
  MUX U521 ( .IN0(n2990), .IN1(n2992), .SEL(n2991), .F(n2866) );
  MUX U522 ( .IN0(n2998), .IN1(n408), .SEL(n2999), .F(n2874) );
  IV U523 ( .A(n3000), .Z(n408) );
  MUX U524 ( .IN0(A[28]), .IN1(n4750), .SEL(A[31]), .F(n409) );
  IV U525 ( .A(n409), .Z(n1023) );
  MUX U526 ( .IN0(n1043), .IN1(n1045), .SEL(n1044), .F(n1002) );
  XNOR U527 ( .A(n1324), .B(n1321), .Z(n1384) );
  MUX U528 ( .IN0(n5470), .IN1(n5472), .SEL(n5471), .F(n5454) );
  MUX U529 ( .IN0(n410), .IN1(n5085), .SEL(n5086), .F(n5071) );
  IV U530 ( .A(n5087), .Z(n410) );
  XNOR U531 ( .A(n4604), .B(n4603), .Z(n4619) );
  MUX U532 ( .IN0(n5548), .IN1(n411), .SEL(n5549), .F(n5530) );
  IV U533 ( .A(n5550), .Z(n411) );
  MUX U534 ( .IN0(n5197), .IN1(n5199), .SEL(n5198), .F(n5177) );
  MUX U535 ( .IN0(n4536), .IN1(n4538), .SEL(n4537), .F(n4524) );
  NANDN U536 ( .B(n2899), .A(n3370), .Z(n424) );
  MUX U537 ( .IN0(n4541), .IN1(n412), .SEL(n4542), .F(n4517) );
  IV U538 ( .A(n4543), .Z(n412) );
  XNOR U539 ( .A(n4251), .B(n4249), .Z(n4264) );
  XNOR U540 ( .A(n5185), .B(n5184), .Z(n5200) );
  MUX U541 ( .IN0(n5335), .IN1(n413), .SEL(n5336), .F(n5323) );
  IV U542 ( .A(n5337), .Z(n413) );
  MUX U543 ( .IN0(n4961), .IN1(n4963), .SEL(n4962), .F(n4944) );
  MUX U544 ( .IN0(n5131), .IN1(n414), .SEL(n5132), .F(n3317) );
  IV U545 ( .A(n5133), .Z(n414) );
  MUX U546 ( .IN0(n1767), .IN1(n415), .SEL(n1768), .F(n1674) );
  IV U547 ( .A(n1769), .Z(n415) );
  MUX U548 ( .IN0(n1916), .IN1(n1918), .SEL(n1917), .F(n1820) );
  MUX U549 ( .IN0(n2040), .IN1(n2042), .SEL(n2041), .F(n1944) );
  MUX U550 ( .IN0(n2216), .IN1(n416), .SEL(n2217), .F(n2108) );
  IV U551 ( .A(n2218), .Z(n416) );
  MUX U552 ( .IN0(n2370), .IN1(n417), .SEL(n2371), .F(n2263) );
  IV U553 ( .A(n2372), .Z(n417) );
  MUX U554 ( .IN0(n2470), .IN1(n418), .SEL(n2471), .F(n2362) );
  IV U555 ( .A(n2472), .Z(n418) );
  MUX U556 ( .IN0(n2565), .IN1(n2567), .SEL(n2566), .F(n2446) );
  MUX U557 ( .IN0(n2557), .IN1(n2559), .SEL(n2558), .F(n2438) );
  MUX U558 ( .IN0(n2647), .IN1(n2649), .SEL(n2648), .F(n2533) );
  MUX U559 ( .IN0(n2940), .IN1(n419), .SEL(n2941), .F(n2815) );
  IV U560 ( .A(n2942), .Z(n419) );
  MUX U561 ( .IN0(n1024), .IN1(n1026), .SEL(n1025), .F(n984) );
  MUX U562 ( .IN0(n1396), .IN1(n1398), .SEL(n1397), .F(n1328) );
  MUX U563 ( .IN0(A[25]), .IN1(n4799), .SEL(A[31]), .F(n420) );
  IV U564 ( .A(n420), .Z(n1168) );
  MUX U565 ( .IN0(n2395), .IN1(n2397), .SEL(n2396), .F(n2290) );
  XNOR U566 ( .A(n1155), .B(n1154), .Z(n1210) );
  XNOR U567 ( .A(n647), .B(n1645), .Z(n1568) );
  AND U568 ( .A(n924), .B(n926), .Z(n895) );
  MUX U569 ( .IN0(n5101), .IN1(n421), .SEL(n5102), .F(n5085) );
  IV U570 ( .A(n5103), .Z(n421) );
  XNOR U571 ( .A(n5247), .B(n5246), .Z(n5264) );
  MUX U572 ( .IN0(n4146), .IN1(n4148), .SEL(n4147), .F(n4132) );
  MUX U573 ( .IN0(n4561), .IN1(n422), .SEL(n4562), .F(n4541) );
  IV U574 ( .A(n4563), .Z(n422) );
  XNOR U575 ( .A(n3527), .B(n3526), .Z(n3562) );
  MUX U576 ( .IN0(n423), .IN1(n5530), .SEL(n5531), .F(n5514) );
  IV U577 ( .A(n5532), .Z(n423) );
  MUX U578 ( .IN0(n5177), .IN1(n5179), .SEL(n5178), .F(n5157) );
  MUX U579 ( .IN0(n4679), .IN1(n424), .SEL(n4680), .F(n4665) );
  XNOR U580 ( .A(n4979), .B(n4978), .Z(n4984) );
  MUX U581 ( .IN0(n5162), .IN1(n425), .SEL(n5163), .F(n5131) );
  IV U582 ( .A(n5164), .Z(n425) );
  XNOR U583 ( .A(n3509), .B(n3507), .Z(n3544) );
  MUX U584 ( .IN0(n5323), .IN1(n426), .SEL(n5324), .F(n3340) );
  IV U585 ( .A(n5325), .Z(n426) );
  MUX U586 ( .IN0(n2263), .IN1(n427), .SEL(n2264), .F(n2157) );
  IV U587 ( .A(n2265), .Z(n427) );
  MUX U588 ( .IN0(n2701), .IN1(n2703), .SEL(n2702), .F(n2581) );
  MUX U589 ( .IN0(n2831), .IN1(n428), .SEL(n2832), .F(n2709) );
  IV U590 ( .A(n2833), .Z(n428) );
  MUX U591 ( .IN0(n2839), .IN1(n429), .SEL(n2840), .F(n2717) );
  IV U592 ( .A(n2841), .Z(n429) );
  MUX U593 ( .IN0(A[22]), .IN1(n4850), .SEL(A[31]), .F(n430) );
  IV U594 ( .A(n430), .Z(n1367) );
  MUX U595 ( .IN0(A[24]), .IN1(n4816), .SEL(A[31]), .F(n431) );
  IV U596 ( .A(n431), .Z(n1232) );
  MUX U597 ( .IN0(A[17]), .IN1(n4935), .SEL(A[31]), .F(n432) );
  IV U598 ( .A(n432), .Z(n1775) );
  MUX U599 ( .IN0(A[19]), .IN1(n4901), .SEL(A[31]), .F(n433) );
  IV U600 ( .A(n433), .Z(n1600) );
  MUX U601 ( .IN0(A[26]), .IN1(n4783), .SEL(A[31]), .F(n434) );
  IV U602 ( .A(n434), .Z(n1109) );
  MUX U603 ( .IN0(A[27]), .IN1(n4767), .SEL(A[31]), .F(n435) );
  IV U604 ( .A(n435), .Z(n1067) );
  MUX U605 ( .IN0(n1229), .IN1(n1227), .SEL(n1228), .F(n1163) );
  MUX U606 ( .IN0(n2906), .IN1(n2908), .SEL(n2907), .F(n2780) );
  XNOR U607 ( .A(n1392), .B(n1391), .Z(n1458) );
  XOR U608 ( .A(n1736), .B(n1651), .Z(n1652) );
  ANDN U609 ( .A(n946), .B(n926), .Z(n915) );
  XNOR U610 ( .A(n5374), .B(n5373), .Z(n5381) );
  MUX U611 ( .IN0(n4141), .IN1(n436), .SEL(n4142), .F(n4127) );
  IV U612 ( .A(n4143), .Z(n436) );
  MUX U613 ( .IN0(n5116), .IN1(n5118), .SEL(n5117), .F(n5112) );
  MUX U614 ( .IN0(n437), .IN1(n5449), .SEL(n5450), .F(n5435) );
  IV U615 ( .A(n5451), .Z(n437) );
  MUX U616 ( .IN0(n438), .IN1(n5071), .SEL(n5072), .F(n5062) );
  IV U617 ( .A(n5073), .Z(n438) );
  XNOR U618 ( .A(n4564), .B(n4563), .Z(n4579) );
  NANDN U619 ( .B(n5562), .A(n3370), .Z(n454) );
  MUX U620 ( .IN0(n5157), .IN1(n5159), .SEL(n5158), .F(n5138) );
  XNOR U621 ( .A(n5338), .B(n5337), .Z(n5343) );
  XNOR U622 ( .A(n5165), .B(n5164), .Z(n5180) );
  XNOR U623 ( .A(n3403), .B(n3402), .Z(n3437) );
  MUX U624 ( .IN0(n2255), .IN1(n439), .SEL(n2256), .F(n2149) );
  IV U625 ( .A(n2257), .Z(n439) );
  MUX U626 ( .IN0(n2550), .IN1(n440), .SEL(n2551), .F(n2431) );
  IV U627 ( .A(n2552), .Z(n440) );
  MUX U628 ( .IN0(n2742), .IN1(n2744), .SEL(n2743), .F(n2622) );
  MUX U629 ( .IN0(n2964), .IN1(n441), .SEL(n2965), .F(n2839) );
  IV U630 ( .A(n2966), .Z(n441) );
  MUX U631 ( .IN0(A[12]), .IN1(n5358), .SEL(A[31]), .F(n442) );
  IV U632 ( .A(n442), .Z(n2271) );
  MUX U633 ( .IN0(n3159), .IN1(n3161), .SEL(n3160), .F(n3034) );
  MUX U634 ( .IN0(A[20]), .IN1(n4884), .SEL(A[31]), .F(n443) );
  IV U635 ( .A(n443), .Z(n1519) );
  MUX U636 ( .IN0(n3128), .IN1(n444), .SEL(n3129), .F(n2998) );
  IV U637 ( .A(n3130), .Z(n444) );
  MUX U638 ( .IN0(A[15]), .IN1(n5322), .SEL(A[31]), .F(n445) );
  IV U639 ( .A(n445), .Z(n1968) );
  MUX U640 ( .IN0(A[23]), .IN1(n4833), .SEL(A[31]), .F(n446) );
  IV U641 ( .A(n446), .Z(n1300) );
  MUX U642 ( .IN0(A[21]), .IN1(n4867), .SEL(A[31]), .F(n447) );
  IV U643 ( .A(n447), .Z(n1441) );
  MUX U644 ( .IN0(n1141), .IN1(n1143), .SEL(n1142), .F(n1085) );
  MUX U645 ( .IN0(n1297), .IN1(n1295), .SEL(n1296), .F(n1227) );
  MUX U646 ( .IN0(n1356), .IN1(n1354), .SEL(n1355), .F(n1285) );
  MUX U647 ( .IN0(n1545), .IN1(n1543), .SEL(n1544), .F(n1465) );
  MUX U648 ( .IN0(n448), .IN1(n1679), .SEL(n1680), .F(n1595) );
  IV U649 ( .A(n1681), .Z(n448) );
  MUX U650 ( .IN0(n2310), .IN1(n2308), .SEL(n2309), .F(n2200) );
  MUX U651 ( .IN0(n449), .IN1(n2600), .SEL(n2601), .F(n2481) );
  IV U652 ( .A(n2602), .Z(n449) );
  MUX U653 ( .IN0(n1020), .IN1(n1018), .SEL(n1019), .F(n978) );
  MUX U654 ( .IN0(n1328), .IN1(n1330), .SEL(n1329), .F(n1259) );
  MUX U655 ( .IN0(n450), .IN1(n1496), .SEL(n1497), .F(n1416) );
  IV U656 ( .A(n1498), .Z(n450) );
  XOR U657 ( .A(n705), .B(n1985), .Z(n1889) );
  MUX U658 ( .IN0(n2290), .IN1(n2292), .SEL(n2291), .F(n2183) );
  ANDN U659 ( .A(n915), .B(n897), .Z(n886) );
  AND U660 ( .A(n955), .B(n957), .Z(n924) );
  MUX U661 ( .IN0(n1707), .IN1(n1705), .SEL(n1706), .F(n1614) );
  MUX U662 ( .IN0(n5465), .IN1(n451), .SEL(n5466), .F(n5449) );
  IV U663 ( .A(n5467), .Z(n451) );
  MUX U664 ( .IN0(n4576), .IN1(n4578), .SEL(n4577), .F(n4556) );
  MUX U665 ( .IN0(n5553), .IN1(n5555), .SEL(n5554), .F(n5535) );
  XNOR U666 ( .A(n5362), .B(n5361), .Z(n5367) );
  MUX U667 ( .IN0(n452), .IN1(n4127), .SEL(n4128), .F(n4113) );
  IV U668 ( .A(n4129), .Z(n452) );
  MUX U669 ( .IN0(n453), .IN1(n5062), .SEL(n5063), .F(n5050) );
  IV U670 ( .A(n5064), .Z(n453) );
  MUX U671 ( .IN0(n5559), .IN1(n454), .SEL(n5560), .F(n5548) );
  MUX U672 ( .IN0(n5138), .IN1(n5140), .SEL(n5139), .F(n3324) );
  MUX U673 ( .IN0(n2478), .IN1(n455), .SEL(n2479), .F(n2370) );
  IV U674 ( .A(n2480), .Z(n455) );
  MUX U675 ( .IN0(n2446), .IN1(n2448), .SEL(n2447), .F(n2338) );
  MUX U676 ( .IN0(n2640), .IN1(n456), .SEL(n2641), .F(n2526) );
  IV U677 ( .A(n2642), .Z(n456) );
  MUX U678 ( .IN0(n2815), .IN1(n457), .SEL(n2816), .F(n2693) );
  IV U679 ( .A(n2817), .Z(n457) );
  MUX U680 ( .IN0(n2767), .IN1(n2769), .SEL(n2768), .F(n2647) );
  MUX U681 ( .IN0(n3080), .IN1(n3082), .SEL(n3081), .F(n2948) );
  MUX U682 ( .IN0(n3088), .IN1(n458), .SEL(n3089), .F(n2956) );
  IV U683 ( .A(n3090), .Z(n458) );
  MUX U684 ( .IN0(A[16]), .IN1(n4952), .SEL(A[31]), .F(n459) );
  IV U685 ( .A(n459), .Z(n1872) );
  MUX U686 ( .IN0(A[18]), .IN1(n4918), .SEL(A[31]), .F(n460) );
  IV U687 ( .A(n460), .Z(n1684) );
  MUX U688 ( .IN0(A[14]), .IN1(n5334), .SEL(A[31]), .F(n461) );
  IV U689 ( .A(n461), .Z(n2064) );
  MUX U690 ( .IN0(n3120), .IN1(n3122), .SEL(n3121), .F(n2990) );
  MUX U691 ( .IN0(A[13]), .IN1(n5346), .SEL(A[31]), .F(n462) );
  IV U692 ( .A(n462), .Z(n2165) );
  MUX U693 ( .IN0(n3262), .IN1(n463), .SEL(n3263), .F(n3128) );
  IV U694 ( .A(n3264), .Z(n463) );
  XNOR U695 ( .A(n3420), .B(n3419), .Z(n4199) );
  MUX U696 ( .IN0(n1160), .IN1(n464), .SEL(n1161), .F(n1101) );
  IV U697 ( .A(n1162), .Z(n464) );
  MUX U698 ( .IN0(n1394), .IN1(n1392), .SEL(n1393), .F(n1324) );
  MUX U699 ( .IN0(n465), .IN1(n1436), .SEL(n1437), .F(n1362) );
  IV U700 ( .A(n1438), .Z(n465) );
  MUX U701 ( .IN0(n2096), .IN1(n2098), .SEL(n2097), .F(n1995) );
  MUX U702 ( .IN0(n1716), .IN1(n1714), .SEL(n1715), .F(n1625) );
  MUX U703 ( .IN0(n1764), .IN1(n1762), .SEL(n1763), .F(n1669) );
  MUX U704 ( .IN0(n2260), .IN1(n2258), .SEL(n2259), .F(n2152) );
  MUX U705 ( .IN0(n2221), .IN1(n2219), .SEL(n2220), .F(n2111) );
  MUX U706 ( .IN0(n2244), .IN1(n2242), .SEL(n2243), .F(n2136) );
  MUX U707 ( .IN0(n2675), .IN1(n2673), .SEL(n2674), .F(n2553) );
  MUX U708 ( .IN0(n2836), .IN1(n2834), .SEL(n2835), .F(n2712) );
  MUX U709 ( .IN0(n466), .IN1(n2842), .SEL(n2843), .F(n2720) );
  IV U710 ( .A(n2844), .Z(n466) );
  MUX U711 ( .IN0(n1053), .IN1(n1051), .SEL(n1052), .F(n1008) );
  MUX U712 ( .IN0(n1064), .IN1(n1062), .SEL(n1063), .F(n1018) );
  XNOR U713 ( .A(n1217), .B(n1216), .Z(n1278) );
  MUX U714 ( .IN0(n467), .IN1(n1659), .SEL(n1660), .F(n1575) );
  IV U715 ( .A(n1661), .Z(n467) );
  XNOR U716 ( .A(n1737), .B(n1747), .Z(n1836) );
  MUX U717 ( .IN0(n2190), .IN1(n468), .SEL(n2191), .F(n2079) );
  IV U718 ( .A(n2192), .Z(n468) );
  XOR U719 ( .A(n928), .B(n905), .Z(n902) );
  MUX U720 ( .IN0(n1002), .IN1(n1004), .SEL(n1003), .F(n469) );
  IV U721 ( .A(n469), .Z(n968) );
  AND U722 ( .A(n1036), .B(n1038), .Z(n996) );
  NOR U723 ( .A(n1703), .B(n1704), .Z(n1702) );
  NANDN U724 ( .B(n874), .A(n886), .Z(n854) );
  MUX U725 ( .IN0(n889), .IN1(Y0[29]), .SEL(n890), .F(n866) );
  MUX U726 ( .IN0(n4483), .IN1(n4481), .SEL(n4482), .F(n4460) );
  MUX U727 ( .IN0(n5419), .IN1(n5296), .SEL(n5297), .F(n5405) );
  MUX U728 ( .IN0(n5479), .IN1(n5481), .SEL(n5480), .F(n5476) );
  MUX U729 ( .IN0(n470), .IN1(n5076), .SEL(n5077), .F(n5057) );
  IV U730 ( .A(n5078), .Z(n470) );
  MUX U731 ( .IN0(n471), .IN1(n5435), .SEL(n5436), .F(n5426) );
  IV U732 ( .A(n5437), .Z(n471) );
  NANDN U733 ( .B(n5303), .A(n3370), .Z(n492) );
  MUX U734 ( .IN0(n4524), .IN1(n4526), .SEL(n4525), .F(n4506) );
  XNOR U735 ( .A(n4544), .B(n4543), .Z(n4559) );
  MUX U736 ( .IN0(n472), .IN1(n5503), .SEL(n5504), .F(n3356) );
  IV U737 ( .A(n5505), .Z(n472) );
  XNOR U738 ( .A(n5326), .B(n5325), .Z(n5331) );
  XNOR U739 ( .A(n5055), .B(n5054), .Z(n5060) );
  MUX U740 ( .IN0(n2223), .IN1(n2225), .SEL(n2224), .F(n2115) );
  MUX U741 ( .IN0(n2338), .IN1(n2340), .SEL(n2339), .F(n2231) );
  MUX U742 ( .IN0(n2581), .IN1(n2583), .SEL(n2582), .F(n2462) );
  MUX U743 ( .IN0(n2589), .IN1(n473), .SEL(n2590), .F(n2470) );
  IV U744 ( .A(n2591), .Z(n473) );
  MUX U745 ( .IN0(n2533), .IN1(n2535), .SEL(n2534), .F(n2419) );
  MUX U746 ( .IN0(n2670), .IN1(n474), .SEL(n2671), .F(n2550) );
  IV U747 ( .A(n2672), .Z(n474) );
  MUX U748 ( .IN0(n2866), .IN1(n2868), .SEL(n2867), .F(n2742) );
  MUX U749 ( .IN0(n2874), .IN1(n475), .SEL(n2875), .F(n2750) );
  IV U750 ( .A(n2876), .Z(n475) );
  MUX U751 ( .IN0(n3013), .IN1(n3015), .SEL(n3014), .F(n2889) );
  MUX U752 ( .IN0(n3064), .IN1(n3066), .SEL(n3065), .F(n2932) );
  MUX U753 ( .IN0(n3072), .IN1(n476), .SEL(n3073), .F(n2940) );
  IV U754 ( .A(n3074), .Z(n476) );
  MUX U755 ( .IN0(n3188), .IN1(n3190), .SEL(n3189), .F(n3056) );
  MUX U756 ( .IN0(n3181), .IN1(n477), .SEL(n3182), .F(n3049) );
  IV U757 ( .A(n3183), .Z(n477) );
  MUX U758 ( .IN0(n3228), .IN1(n478), .SEL(n3229), .F(n3096) );
  IV U759 ( .A(n3230), .Z(n478) );
  MUX U760 ( .IN0(n3136), .IN1(n479), .SEL(n3137), .F(n3006) );
  IV U761 ( .A(n3138), .Z(n479) );
  MUX U762 ( .IN0(n5136), .IN1(n5134), .SEL(n5135), .F(n3320) );
  MUX U763 ( .IN0(n3405), .IN1(n3403), .SEL(n3404), .F(n3273) );
  XNOR U764 ( .A(n3395), .B(n3394), .Z(n3457) );
  MUX U765 ( .IN0(n1068), .IN1(n1070), .SEL(n1069), .F(n1024) );
  MUX U766 ( .IN0(n1671), .IN1(n1669), .SEL(n1670), .F(n1585) );
  MUX U767 ( .IN0(n480), .IN1(n2059), .SEL(n2060), .F(n1963) );
  IV U768 ( .A(n2061), .Z(n480) );
  MUX U769 ( .IN0(n2037), .IN1(n2035), .SEL(n2036), .F(n1939) );
  MUX U770 ( .IN0(n2328), .IN1(n2326), .SEL(n2327), .F(n2219) );
  MUX U771 ( .IN0(n2367), .IN1(n2365), .SEL(n2366), .F(n2258) );
  MUX U772 ( .IN0(n2407), .IN1(n2409), .SEL(n2408), .F(n481) );
  IV U773 ( .A(n481), .Z(n2297) );
  MUX U774 ( .IN0(n2578), .IN1(n2576), .SEL(n2577), .F(n2457) );
  MUX U775 ( .IN0(n2765), .IN1(n2763), .SEL(n2764), .F(n2643) );
  MUX U776 ( .IN0(n482), .IN1(n2967), .SEL(n2968), .F(n2842) );
  IV U777 ( .A(n2969), .Z(n482) );
  MUX U778 ( .IN0(n2961), .IN1(n2959), .SEL(n2960), .F(n2834) );
  MUX U779 ( .IN0(n2922), .IN1(n2920), .SEL(n2921), .F(n2795) );
  MUX U780 ( .IN0(n2904), .IN1(n2902), .SEL(n2903), .F(n483) );
  IV U781 ( .A(n483), .Z(n2774) );
  MUX U782 ( .IN0(n3003), .IN1(n3001), .SEL(n3002), .F(n2877) );
  XNOR U783 ( .A(n3289), .B(n3288), .Z(n3413) );
  MUX U784 ( .IN0(n980), .IN1(n978), .SEL(n979), .F(n934) );
  MUX U785 ( .IN0(n1165), .IN1(n1163), .SEL(n1164), .F(n1104) );
  MUX U786 ( .IN0(n1336), .IN1(n1334), .SEL(n1335), .F(n1265) );
  MUX U787 ( .IN0(n484), .IN1(n1344), .SEL(n1345), .F(n1275) );
  IV U788 ( .A(n1346), .Z(n484) );
  XNOR U789 ( .A(n1465), .B(n1464), .Z(n1536) );
  MUX U790 ( .IN0(n485), .IN1(n1754), .SEL(n1755), .F(n1659) );
  IV U791 ( .A(n1756), .Z(n485) );
  XNOR U792 ( .A(n2082), .B(n1991), .Z(n1992) );
  MUX U793 ( .IN0(n2294), .IN1(n486), .SEL(n2295), .F(n2190) );
  IV U794 ( .A(n2296), .Z(n486) );
  MUX U795 ( .IN0(n2780), .IN1(n2782), .SEL(n2781), .F(n2662) );
  ANDN U796 ( .A(n961), .B(n965), .Z(n964) );
  MUX U797 ( .IN0(n487), .IN1(n1195), .SEL(n1196), .F(n1136) );
  IV U798 ( .A(n1197), .Z(n487) );
  ANDN U799 ( .A(n1901), .B(n1903), .Z(n1792) );
  MUX U800 ( .IN0(n535), .IN1(n2542), .SEL(n2541), .F(n2425) );
  NANDN U801 ( .B(n947), .A(n948), .Z(n916) );
  AND U802 ( .A(n996), .B(n998), .Z(n955) );
  NANDN U803 ( .B(n1116), .A(n1117), .Z(n1072) );
  AND U804 ( .A(n1314), .B(n1316), .Z(n1246) );
  MUX U805 ( .IN0(n1807), .IN1(n488), .SEL(n1806), .F(n1705) );
  IV U806 ( .A(n1805), .Z(n488) );
  AND U807 ( .A(n862), .B(n863), .Z(n857) );
  MUX U808 ( .IN0(n918), .IN1(Y0[28]), .SEL(n919), .F(n889) );
  MUX U809 ( .IN0(n4090), .IN1(n4088), .SEL(n4089), .F(n4046) );
  MUX U810 ( .IN0(n4155), .IN1(n4157), .SEL(n4156), .F(n4152) );
  MUX U811 ( .IN0(n489), .IN1(n5440), .SEL(n5441), .F(n5421) );
  IV U812 ( .A(n5442), .Z(n489) );
  MUX U813 ( .IN0(n490), .IN1(n4113), .SEL(n4114), .F(n4104) );
  IV U814 ( .A(n4115), .Z(n490) );
  MUX U815 ( .IN0(n491), .IN1(n5057), .SEL(n5058), .F(n5045) );
  IV U816 ( .A(n5059), .Z(n491) );
  MUX U817 ( .IN0(n5300), .IN1(n492), .SEL(n5301), .F(n5288) );
  MUX U818 ( .IN0(n493), .IN1(n5426), .SEL(n5427), .F(n5414) );
  IV U819 ( .A(n5428), .Z(n493) );
  XNOR U820 ( .A(n4520), .B(n4519), .Z(n4539) );
  MUX U821 ( .IN0(n2115), .IN1(n2117), .SEL(n2116), .F(n2014) );
  MUX U822 ( .IN0(n2149), .IN1(n494), .SEL(n2150), .F(n2048) );
  IV U823 ( .A(n2151), .Z(n494) );
  MUX U824 ( .IN0(n2597), .IN1(n495), .SEL(n2598), .F(n2478) );
  IV U825 ( .A(n2599), .Z(n495) );
  MUX U826 ( .IN0(n2709), .IN1(n496), .SEL(n2710), .F(n2589) );
  IV U827 ( .A(n2711), .Z(n496) );
  MUX U828 ( .IN0(n2685), .IN1(n2687), .SEL(n2686), .F(n2565) );
  MUX U829 ( .IN0(n2799), .IN1(n2801), .SEL(n2800), .F(n2677) );
  MUX U830 ( .IN0(n2792), .IN1(n497), .SEL(n2793), .F(n2670) );
  IV U831 ( .A(n2794), .Z(n497) );
  MUX U832 ( .IN0(n2948), .IN1(n2950), .SEL(n2949), .F(n2823) );
  MUX U833 ( .IN0(n2882), .IN1(n498), .SEL(n2883), .F(n2760) );
  IV U834 ( .A(n2884), .Z(n498) );
  MUX U835 ( .IN0(n3196), .IN1(n3198), .SEL(n3197), .F(n3064) );
  MUX U836 ( .IN0(n3204), .IN1(n499), .SEL(n3205), .F(n3072) );
  IV U837 ( .A(n3206), .Z(n499) );
  MUX U838 ( .IN0(n3356), .IN1(n500), .SEL(n3357), .F(n3220) );
  IV U839 ( .A(n3358), .Z(n500) );
  MUX U840 ( .IN0(n3317), .IN1(n501), .SEL(n3318), .F(n3181) );
  IV U841 ( .A(n3319), .Z(n501) );
  MUX U842 ( .IN0(n3254), .IN1(n3256), .SEL(n3255), .F(n3120) );
  MUX U843 ( .IN0(n5326), .IN1(n5152), .SEL(n5154), .F(n3343) );
  MUX U844 ( .IN0(n1110), .IN1(n1112), .SEL(n1111), .F(n1068) );
  MUX U845 ( .IN0(n1914), .IN1(n1912), .SEL(n1913), .F(n1816) );
  MUX U846 ( .IN0(n1957), .IN1(n1955), .SEL(n1956), .F(n1859) );
  MUX U847 ( .IN0(n502), .IN1(n1963), .SEL(n1964), .F(n1867) );
  IV U848 ( .A(n1965), .Z(n502) );
  MUX U849 ( .IN0(n2351), .IN1(n2349), .SEL(n2350), .F(n2242) );
  MUX U850 ( .IN0(n503), .IN1(n2373), .SEL(n2374), .F(n2266) );
  IV U851 ( .A(n2375), .Z(n503) );
  MUX U852 ( .IN0(n2475), .IN1(n2473), .SEL(n2474), .F(n2365) );
  MUX U853 ( .IN0(n2436), .IN1(n2434), .SEL(n2435), .F(n2326) );
  MUX U854 ( .IN0(n2531), .IN1(n2529), .SEL(n2530), .F(n2415) );
  MUX U855 ( .IN0(n2945), .IN1(n2943), .SEL(n2944), .F(n2818) );
  MUX U856 ( .IN0(n2879), .IN1(n2877), .SEL(n2878), .F(n2755) );
  MUX U857 ( .IN0(n3093), .IN1(n3091), .SEL(n3092), .F(n2959) );
  MUX U858 ( .IN0(n504), .IN1(n3099), .SEL(n3100), .F(n2967) );
  IV U859 ( .A(n3101), .Z(n504) );
  MUX U860 ( .IN0(n3054), .IN1(n3052), .SEL(n3053), .F(n2920) );
  MUX U861 ( .IN0(n3141), .IN1(n3139), .SEL(n3140), .F(n3009) );
  XNOR U862 ( .A(n3265), .B(n3264), .Z(n3388) );
  MUX U863 ( .IN0(n1098), .IN1(n1096), .SEL(n1097), .F(n1051) );
  XNOR U864 ( .A(n1163), .B(n1162), .Z(n1220) );
  MUX U865 ( .IN0(n1404), .IN1(n1406), .SEL(n1405), .F(n1334) );
  XNOR U866 ( .A(n1354), .B(n1353), .Z(n1419) );
  XNOR U867 ( .A(n1514), .B(n1513), .Z(n1588) );
  XNOR U868 ( .A(n1543), .B(n1542), .Z(n1618) );
  MUX U869 ( .IN0(n1995), .IN1(n1997), .SEL(n1996), .F(n1894) );
  MUX U870 ( .IN0(n505), .IN1(n1733), .SEL(n1734), .F(n1642) );
  IV U871 ( .A(n1735), .Z(n505) );
  XNOR U872 ( .A(n2083), .B(n2093), .Z(n2193) );
  XOR U873 ( .A(n2511), .B(n2407), .Z(n2408) );
  MUX U874 ( .IN0(n506), .IN1(n2704), .SEL(n2705), .F(n2584) );
  IV U875 ( .A(n2706), .Z(n506) );
  MUX U876 ( .IN0(n2776), .IN1(n507), .SEL(n2775), .F(n2660) );
  IV U877 ( .A(n2774), .Z(n507) );
  MUX U878 ( .IN0(n971), .IN1(n508), .SEL(n970), .F(n943) );
  IV U879 ( .A(n969), .Z(n508) );
  XNOR U880 ( .A(n1134), .B(n1133), .Z(n1187) );
  AND U881 ( .A(n1524), .B(n1526), .Z(n1446) );
  MUX U882 ( .IN0(n509), .IN1(n1632), .SEL(n1633), .F(n1552) );
  IV U883 ( .A(n1634), .Z(n509) );
  MUX U884 ( .IN0(n2786), .IN1(n2788), .SEL(n2787), .F(n2664) );
  NANDN U885 ( .B(n988), .A(n989), .Z(n947) );
  ANDN U886 ( .A(n1027), .B(n998), .Z(n987) );
  NANDN U887 ( .B(n1175), .A(n1176), .Z(n1116) );
  NAND U888 ( .A(n1792), .B(n1791), .Z(n1703) );
  MUX U889 ( .IN0(n510), .IN1(n2315), .SEL(n2316), .F(n2207) );
  IV U890 ( .A(n2317), .Z(n510) );
  ANDN U891 ( .A(n1455), .B(n1456), .Z(n1381) );
  MUX U892 ( .IN0(Y0[3]), .IN1(n2977), .SEL(n2978), .F(n2854) );
  MUX U893 ( .IN0(n854), .IN1(n856), .SEL(n855), .F(n511) );
  IV U894 ( .A(n511), .Z(n853) );
  MUX U895 ( .IN0(n949), .IN1(Y0[27]), .SEL(n950), .F(n918) );
  MUX U896 ( .IN0(n1118), .IN1(Y0[23]), .SEL(n1119), .F(n1074) );
  MUX U897 ( .IN0(n1375), .IN1(Y0[19]), .SEL(n1376), .F(n1308) );
  MUX U898 ( .IN0(n1692), .IN1(Y0[15]), .SEL(n1693), .F(n1608) );
  MUX U899 ( .IN0(n2072), .IN1(Y0[11]), .SEL(n2073), .F(n1976) );
  MUX U900 ( .IN0(n2494), .IN1(Y0[7]), .SEL(n2495), .F(n2386) );
  MUX U901 ( .IN0(n4959), .IN1(n4513), .SEL(n4514), .F(n4942) );
  MUX U902 ( .IN0(n512), .IN1(n4490), .SEL(n4055), .F(n4469) );
  IV U903 ( .A(n4053), .Z(n512) );
  MUX U904 ( .IN0(n3929), .IN1(n3927), .SEL(n3928), .F(n3883) );
  MUX U905 ( .IN0(n4650), .IN1(n4648), .SEL(n4649), .F(n4624) );
  XNOR U906 ( .A(n5225), .B(n5224), .Z(n5240) );
  MUX U907 ( .IN0(n4682), .IN1(n4684), .SEL(n4683), .F(n4679) );
  MUX U908 ( .IN0(n513), .IN1(n4118), .SEL(n4119), .F(n4097) );
  IV U909 ( .A(n4120), .Z(n513) );
  NANDN U910 ( .B(n1988), .A(n3370), .Z(n545) );
  MUX U911 ( .IN0(n514), .IN1(n5494), .SEL(n5495), .F(n3348) );
  IV U912 ( .A(n5496), .Z(n514) );
  MUX U913 ( .IN0(n5145), .IN1(n5147), .SEL(n5146), .F(n3332) );
  MUX U914 ( .IN0(n4208), .IN1(n4206), .SEL(n4207), .F(n3420) );
  MUX U915 ( .IN0(n2231), .IN1(n2233), .SEL(n2232), .F(n2123) );
  MUX U916 ( .IN0(n2354), .IN1(n2356), .SEL(n2355), .F(n2247) );
  MUX U917 ( .IN0(n2438), .IN1(n2440), .SEL(n2439), .F(n2330) );
  MUX U918 ( .IN0(n2431), .IN1(n515), .SEL(n2432), .F(n2323) );
  IV U919 ( .A(n2433), .Z(n515) );
  MUX U920 ( .IN0(n2693), .IN1(n516), .SEL(n2694), .F(n2573) );
  IV U921 ( .A(n2695), .Z(n516) );
  MUX U922 ( .IN0(n2807), .IN1(n2809), .SEL(n2808), .F(n2685) );
  MUX U923 ( .IN0(n2823), .IN1(n2825), .SEL(n2824), .F(n2701) );
  MUX U924 ( .IN0(n2956), .IN1(n517), .SEL(n2957), .F(n2831) );
  IV U925 ( .A(n2958), .Z(n517) );
  MUX U926 ( .IN0(n2917), .IN1(n518), .SEL(n2918), .F(n2792) );
  IV U927 ( .A(n2919), .Z(n518) );
  MUX U928 ( .IN0(n3006), .IN1(n519), .SEL(n3007), .F(n2882) );
  IV U929 ( .A(n3008), .Z(n519) );
  MUX U930 ( .IN0(n3096), .IN1(n520), .SEL(n3097), .F(n2964) );
  IV U931 ( .A(n3098), .Z(n520) );
  MUX U932 ( .IN0(n3056), .IN1(n3058), .SEL(n3057), .F(n2924) );
  MUX U933 ( .IN0(A[8]), .IN1(n5413), .SEL(A[31]), .F(n521) );
  IV U934 ( .A(n521), .Z(n2725) );
  MUX U935 ( .IN0(n3340), .IN1(n522), .SEL(n3341), .F(n3204) );
  IV U936 ( .A(n3342), .Z(n522) );
  MUX U937 ( .IN0(n3293), .IN1(n3295), .SEL(n3294), .F(n3159) );
  MUX U938 ( .IN0(n1219), .IN1(n1217), .SEL(n1218), .F(n1155) );
  MUX U939 ( .IN0(n2113), .IN1(n2111), .SEL(n2112), .F(n2010) );
  MUX U940 ( .IN0(n2154), .IN1(n2152), .SEL(n2153), .F(n2051) );
  MUX U941 ( .IN0(n2085), .IN1(n2083), .SEL(n2084), .F(n1991) );
  MUX U942 ( .IN0(n523), .IN1(n2266), .SEL(n2267), .F(n2160) );
  IV U943 ( .A(n2268), .Z(n523) );
  MUX U944 ( .IN0(n2459), .IN1(n2457), .SEL(n2458), .F(n2349) );
  MUX U945 ( .IN0(n2555), .IN1(n2553), .SEL(n2554), .F(n2434) );
  MUX U946 ( .IN0(n2594), .IN1(n2592), .SEL(n2593), .F(n2473) );
  MUX U947 ( .IN0(n2514), .IN1(n2512), .SEL(n2513), .F(n2407) );
  MUX U948 ( .IN0(n2645), .IN1(n2643), .SEL(n2644), .F(n2529) );
  MUX U949 ( .IN0(n524), .IN1(n2720), .SEL(n2721), .F(n2600) );
  IV U950 ( .A(n2722), .Z(n524) );
  MUX U951 ( .IN0(n3023), .IN1(n3021), .SEL(n3022), .F(n2902) );
  MUX U952 ( .IN0(n3077), .IN1(n3075), .SEL(n3076), .F(n2943) );
  MUX U953 ( .IN0(n3186), .IN1(n3184), .SEL(n3185), .F(n3052) );
  MUX U954 ( .IN0(n3225), .IN1(n3223), .SEL(n3224), .F(n3091) );
  MUX U955 ( .IN0(n525), .IN1(n3231), .SEL(n3232), .F(n3099) );
  IV U956 ( .A(n3233), .Z(n525) );
  MUX U957 ( .IN0(n3133), .IN1(n3131), .SEL(n3132), .F(n3001) );
  MUX U958 ( .IN0(n3275), .IN1(n3273), .SEL(n3274), .F(n3139) );
  MUX U959 ( .IN0(n984), .IN1(n986), .SEL(n985), .F(n940) );
  MUX U960 ( .IN0(n1106), .IN1(n1104), .SEL(n1105), .F(n1062) );
  XNOR U961 ( .A(n1295), .B(n1294), .Z(n1357) );
  XNOR U962 ( .A(n1506), .B(n1505), .Z(n1578) );
  XNOR U963 ( .A(n1595), .B(n1594), .Z(n1672) );
  XNOR U964 ( .A(n1625), .B(n1624), .Z(n1709) );
  MUX U965 ( .IN0(n526), .IN1(n1851), .SEL(n1852), .F(n1754) );
  IV U966 ( .A(n1853), .Z(n526) );
  XNOR U967 ( .A(n1843), .B(n1842), .Z(n1932) );
  MUX U968 ( .IN0(n2398), .IN1(n527), .SEL(n2399), .F(n2294) );
  IV U969 ( .A(n2400), .Z(n527) );
  MUX U970 ( .IN0(n528), .IN1(n2465), .SEL(n2466), .F(n2357) );
  IV U971 ( .A(n2467), .Z(n528) );
  MUX U972 ( .IN0(n529), .IN1(n2688), .SEL(n2689), .F(n2568) );
  IV U973 ( .A(n2690), .Z(n529) );
  MUX U974 ( .IN0(n530), .IN1(n2951), .SEL(n2952), .F(n2826) );
  IV U975 ( .A(n2953), .Z(n530) );
  MUX U976 ( .IN0(n531), .IN1(n2869), .SEL(n2870), .F(n2745) );
  IV U977 ( .A(n2871), .Z(n531) );
  MUX U978 ( .IN0(n532), .IN1(n931), .SEL(n930), .F(n905) );
  IV U979 ( .A(n929), .Z(n532) );
  AND U980 ( .A(n967), .B(n968), .Z(n963) );
  MUX U981 ( .IN0(n1254), .IN1(n1252), .SEL(n1253), .F(n1192) );
  MUX U982 ( .IN0(n533), .IN1(n1399), .SEL(n1400), .F(n1331) );
  IV U983 ( .A(n1401), .Z(n533) );
  AND U984 ( .A(n1605), .B(n1607), .Z(n1524) );
  MUX U985 ( .IN0(n1894), .IN1(n1896), .SEL(n1895), .F(n1803) );
  MUX U986 ( .IN0(n534), .IN1(n2118), .SEL(n2119), .F(n2017) );
  IV U987 ( .A(n2120), .Z(n534) );
  ANDN U988 ( .A(n2102), .B(n2104), .Z(n2001) );
  AND U989 ( .A(n2383), .B(n2385), .Z(n2276) );
  MUX U990 ( .IN0(n2666), .IN1(n2664), .SEL(n2665), .F(n535) );
  IV U991 ( .A(n535), .Z(n2540) );
  NANDN U992 ( .B(n1028), .A(n1029), .Z(n988) );
  MUX U993 ( .IN0(n1115), .IN1(n536), .SEL(n1114), .F(n1071) );
  IV U994 ( .A(n1113), .Z(n536) );
  AND U995 ( .A(n1183), .B(n1185), .Z(n1172) );
  NANDN U996 ( .B(n1238), .A(n1239), .Z(n1175) );
  MUX U997 ( .IN0(n537), .IN1(n1898), .SEL(n1899), .F(n1805) );
  IV U998 ( .A(n1900), .Z(n537) );
  MUX U999 ( .IN0(n538), .IN1(n2422), .SEL(n2423), .F(n2315) );
  IV U1000 ( .A(n2424), .Z(n538) );
  MUX U1001 ( .IN0(n2894), .IN1(n565), .SEL(n2893), .F(n539) );
  IV U1002 ( .A(n539), .Z(n2770) );
  AND U1003 ( .A(n895), .B(n897), .Z(n872) );
  ANDN U1004 ( .A(n1533), .B(n1534), .Z(n1455) );
  NAND U1005 ( .A(n843), .B(n845), .Z(n842) );
  MUX U1006 ( .IN0(n990), .IN1(Y0[26]), .SEL(n991), .F(n949) );
  MUX U1007 ( .IN0(n1177), .IN1(Y0[22]), .SEL(n1178), .F(n1118) );
  MUX U1008 ( .IN0(n1449), .IN1(Y0[18]), .SEL(n1450), .F(n1375) );
  MUX U1009 ( .IN0(n1783), .IN1(Y0[14]), .SEL(n1784), .F(n1692) );
  MUX U1010 ( .IN0(n2173), .IN1(Y0[10]), .SEL(n2174), .F(n2072) );
  MUX U1011 ( .IN0(n2613), .IN1(Y0[6]), .SEL(n2614), .F(n2494) );
  MUX U1012 ( .IN0(n4504), .IN1(n4502), .SEL(n4503), .F(n4481) );
  MUX U1013 ( .IN0(n4079), .IN1(n4077), .SEL(n4078), .F(n540) );
  IV U1014 ( .A(n540), .Z(n4035) );
  MUX U1015 ( .IN0(n4002), .IN1(n4000), .SEL(n4001), .F(n3954) );
  MUX U1016 ( .IN0(n4925), .IN1(n4471), .SEL(n4472), .F(n4908) );
  MUX U1017 ( .IN0(n541), .IN1(n4406), .SEL(n3873), .F(n4385) );
  IV U1018 ( .A(n3871), .Z(n541) );
  MUX U1019 ( .IN0(n5055), .IN1(n4675), .SEL(n4676), .F(n5043) );
  MUX U1020 ( .IN0(n5293), .IN1(n5291), .SEL(n5292), .F(n5271) );
  XNOR U1021 ( .A(n4624), .B(n4623), .Z(n4641) );
  MUX U1022 ( .IN0(n542), .IN1(n4322), .SEL(n3691), .F(n4301) );
  IV U1023 ( .A(n3689), .Z(n542) );
  MUX U1024 ( .IN0(n5001), .IN1(n4591), .SEL(n4593), .F(n4989) );
  MUX U1025 ( .IN0(n5563), .IN1(n5565), .SEL(n5564), .F(n5559) );
  MUX U1026 ( .IN0(n5207), .IN1(n5205), .SEL(n5206), .F(n5185) );
  MUX U1027 ( .IN0(n543), .IN1(n5519), .SEL(n5520), .F(n5494) );
  IV U1028 ( .A(n5521), .Z(n543) );
  MUX U1029 ( .IN0(n544), .IN1(n5421), .SEL(n5422), .F(n5407) );
  IV U1030 ( .A(n5423), .Z(n544) );
  MUX U1031 ( .IN0(n4173), .IN1(n545), .SEL(n4174), .F(n4059) );
  MUX U1032 ( .IN0(n546), .IN1(n4239), .SEL(n3518), .F(n4218) );
  IV U1033 ( .A(n3516), .Z(n546) );
  MUX U1034 ( .IN0(n2247), .IN1(n2249), .SEL(n2248), .F(n2141) );
  MUX U1035 ( .IN0(n3220), .IN1(n547), .SEL(n3221), .F(n3088) );
  IV U1036 ( .A(n3222), .Z(n547) );
  MUX U1037 ( .IN0(A[7]), .IN1(n5502), .SEL(A[31]), .F(n548) );
  IV U1038 ( .A(n548), .Z(n2847) );
  MUX U1039 ( .IN0(A[11]), .IN1(n5370), .SEL(A[31]), .F(n549) );
  IV U1040 ( .A(n549), .Z(n2378) );
  MUX U1041 ( .IN0(n3277), .IN1(n3279), .SEL(n3278), .F(n3143) );
  MUX U1042 ( .IN0(n3270), .IN1(n550), .SEL(n3271), .F(n3136) );
  IV U1043 ( .A(n3272), .Z(n550) );
  MUX U1044 ( .IN0(n3397), .IN1(n3395), .SEL(n3396), .F(n3265) );
  MUX U1045 ( .IN0(n1169), .IN1(n1171), .SEL(n1170), .F(n1110) );
  MUX U1046 ( .IN0(n1587), .IN1(n1585), .SEL(n1586), .F(n1506) );
  MUX U1047 ( .IN0(n1739), .IN1(n1737), .SEL(n1738), .F(n1651) );
  MUX U1048 ( .IN0(n2138), .IN1(n2136), .SEL(n2137), .F(n2035) );
  MUX U1049 ( .IN0(n2698), .IN1(n2696), .SEL(n2697), .F(n2576) );
  MUX U1050 ( .IN0(n2797), .IN1(n2795), .SEL(n2796), .F(n2673) );
  MUX U1051 ( .IN0(n3011), .IN1(n3009), .SEL(n3010), .F(n2885) );
  MUX U1052 ( .IN0(n3209), .IN1(n3207), .SEL(n3208), .F(n3075) );
  MUX U1053 ( .IN0(n551), .IN1(n3367), .SEL(n3368), .F(n3231) );
  IV U1054 ( .A(n3369), .Z(n551) );
  MUX U1055 ( .IN0(n3361), .IN1(n3359), .SEL(n3360), .F(n3223) );
  MUX U1056 ( .IN0(n3322), .IN1(n3320), .SEL(n3321), .F(n3184) );
  XNOR U1057 ( .A(n1227), .B(n1226), .Z(n1288) );
  XNOR U1058 ( .A(n1285), .B(n1284), .Z(n1347) );
  XNOR U1059 ( .A(n1436), .B(n1435), .Z(n1509) );
  MUX U1060 ( .IN0(n1565), .IN1(n552), .SEL(n1566), .F(n1486) );
  IV U1061 ( .A(n1567), .Z(n552) );
  XNOR U1062 ( .A(n1679), .B(n1678), .Z(n1765) );
  XNOR U1063 ( .A(n1714), .B(n1713), .Z(n1809) );
  XNOR U1064 ( .A(n1859), .B(n1858), .Z(n1950) );
  MUX U1065 ( .IN0(n553), .IN1(n2043), .SEL(n2044), .F(n1947) );
  IV U1066 ( .A(n2045), .Z(n553) );
  XNOR U1067 ( .A(n1963), .B(n1962), .Z(n2054) );
  XNOR U1068 ( .A(n2010), .B(n2009), .Z(n2106) );
  MUX U1069 ( .IN0(n554), .IN1(n2234), .SEL(n2235), .F(n2126) );
  IV U1070 ( .A(n2236), .Z(n554) );
  XNOR U1071 ( .A(n2258), .B(n2257), .Z(n2360) );
  XNOR U1072 ( .A(n2266), .B(n2265), .Z(n2368) );
  XNOR U1073 ( .A(n2415), .B(n2414), .Z(n2524) );
  XNOR U1074 ( .A(n2592), .B(n2591), .Z(n2707) );
  XNOR U1075 ( .A(n2600), .B(n2599), .Z(n2715) );
  XNOR U1076 ( .A(n2635), .B(n2634), .Z(n2748) );
  MUX U1077 ( .IN0(n555), .IN1(n2935), .SEL(n2936), .F(n2810) );
  IV U1078 ( .A(n2937), .Z(n555) );
  XNOR U1079 ( .A(n3021), .B(n3031), .Z(n3150) );
  MUX U1080 ( .IN0(n556), .IN1(n3123), .SEL(n3124), .F(n2993) );
  IV U1081 ( .A(n3125), .Z(n556) );
  XNOR U1082 ( .A(n934), .B(n931), .Z(n972) );
  MUX U1083 ( .IN0(n1010), .IN1(n1008), .SEL(n1009), .F(n961) );
  MUX U1084 ( .IN0(n557), .IN1(n1046), .SEL(n1047), .F(n1005) );
  IV U1085 ( .A(n1048), .Z(n557) );
  AND U1086 ( .A(n1265), .B(n1267), .Z(n1198) );
  MUX U1087 ( .IN0(n558), .IN1(n1474), .SEL(n1475), .F(n1399) );
  IV U1088 ( .A(n1476), .Z(n558) );
  MUX U1089 ( .IN0(n1890), .IN1(n705), .SEL(n1889), .F(n1802) );
  AND U1090 ( .A(n1973), .B(n1975), .Z(n1877) );
  ANDN U1091 ( .A(n2210), .B(n2212), .Z(n2102) );
  MUX U1092 ( .IN0(n559), .IN1(n2333), .SEL(n2334), .F(n2226) );
  IV U1093 ( .A(n2335), .Z(n559) );
  AND U1094 ( .A(n2610), .B(n2612), .Z(n2491) );
  MUX U1095 ( .IN0(n560), .IN1(n2802), .SEL(n2803), .F(n2680) );
  IV U1096 ( .A(n2804), .Z(n560) );
  MUX U1097 ( .IN0(n561), .IN1(n2913), .SEL(n2912), .F(n2786) );
  IV U1098 ( .A(n2911), .Z(n561) );
  NANDN U1099 ( .B(n916), .A(n917), .Z(n887) );
  ANDN U1100 ( .A(n1071), .B(n1038), .Z(n1027) );
  NANDN U1101 ( .B(n1072), .A(n1073), .Z(n1028) );
  MUX U1102 ( .IN0(n1194), .IN1(n1192), .SEL(n1193), .F(n562) );
  IV U1103 ( .A(n562), .Z(n1132) );
  OR U1104 ( .A(n1373), .B(n1374), .Z(n1306) );
  MUX U1105 ( .IN0(n563), .IN1(n1998), .SEL(n1999), .F(n1898) );
  IV U1106 ( .A(n2000), .Z(n563) );
  MUX U1107 ( .IN0(n564), .IN1(n2536), .SEL(n2537), .F(n2422) );
  IV U1108 ( .A(n2538), .Z(n564) );
  MUX U1109 ( .IN0(n3018), .IN1(n598), .SEL(n3017), .F(n565) );
  IV U1110 ( .A(n565), .Z(n2892) );
  AND U1111 ( .A(n1172), .B(n1174), .Z(n1080) );
  MUX U1112 ( .IN0(n566), .IN1(n1614), .SEL(n1615), .F(n1533) );
  IV U1113 ( .A(n1616), .Z(n566) );
  ANDN U1114 ( .A(n847), .B(n848), .Z(n839) );
  MUX U1115 ( .IN0(n1030), .IN1(Y0[25]), .SEL(n1031), .F(n990) );
  MUX U1116 ( .IN0(n1240), .IN1(Y0[21]), .SEL(n1241), .F(n1177) );
  MUX U1117 ( .IN0(n1527), .IN1(Y0[17]), .SEL(n1528), .F(n1449) );
  MUX U1118 ( .IN0(n1880), .IN1(Y0[13]), .SEL(n1881), .F(n1783) );
  MUX U1119 ( .IN0(n2279), .IN1(Y0[9]), .SEL(n2280), .F(n2173) );
  MUX U1120 ( .IN0(n2733), .IN1(Y0[5]), .SEL(n2734), .F(n2613) );
  MUX U1121 ( .IN0(n866), .IN1(Y0[30]), .SEL(n867), .F(n832) );
  MUX U1122 ( .IN0(n3410), .IN1(n4091), .SEL(n3411), .F(n567) );
  IV U1123 ( .A(n567), .Z(n4049) );
  MUX U1124 ( .IN0(n568), .IN1(n4035), .SEL(n4036), .F(n3989) );
  IV U1125 ( .A(n4037), .Z(n568) );
  MUX U1126 ( .IN0(n4441), .IN1(n4439), .SEL(n4440), .F(n4418) );
  MUX U1127 ( .IN0(n3956), .IN1(n3954), .SEL(n3955), .F(n3908) );
  MUX U1128 ( .IN0(n569), .IN1(n3853), .SEL(n3854), .F(n3807) );
  IV U1129 ( .A(n3855), .Z(n569) );
  MUX U1130 ( .IN0(n4857), .IN1(n4387), .SEL(n4388), .F(n4840) );
  MUX U1131 ( .IN0(n3747), .IN1(n3745), .SEL(n3746), .F(n3701) );
  MUX U1132 ( .IN0(n4357), .IN1(n4355), .SEL(n4356), .F(n4334) );
  MUX U1133 ( .IN0(n3774), .IN1(n3772), .SEL(n3773), .F(n3726) );
  MUX U1134 ( .IN0(n5141), .IN1(n5294), .SEL(n5142), .F(n570) );
  IV U1135 ( .A(n570), .Z(n5274) );
  MUX U1136 ( .IN0(n571), .IN1(n3671), .SEL(n3672), .F(n3626) );
  IV U1137 ( .A(n3673), .Z(n571) );
  MUX U1138 ( .IN0(n4789), .IN1(n4303), .SEL(n4304), .F(n4773) );
  MUX U1139 ( .IN0(n5374), .IN1(n5232), .SEL(n5234), .F(n5362) );
  MUX U1140 ( .IN0(n3571), .IN1(n3569), .SEL(n3570), .F(n3527) );
  MUX U1141 ( .IN0(n5112), .IN1(n572), .SEL(n5113), .F(n5101) );
  IV U1142 ( .A(n5115), .Z(n572) );
  MUX U1143 ( .IN0(n4273), .IN1(n4271), .SEL(n4272), .F(n4251) );
  MUX U1144 ( .IN0(n3596), .IN1(n3594), .SEL(n3595), .F(n3551) );
  MUX U1145 ( .IN0(n5304), .IN1(n5306), .SEL(n5305), .F(n5300) );
  MUX U1146 ( .IN0(n4566), .IN1(n4564), .SEL(n4565), .F(n4544) );
  NANDN U1147 ( .B(n5583), .A(n3370), .Z(n607) );
  MUX U1148 ( .IN0(n573), .IN1(n3498), .SEL(n3499), .F(n3454) );
  IV U1149 ( .A(n3500), .Z(n573) );
  MUX U1150 ( .IN0(n2677), .IN1(n2679), .SEL(n2678), .F(n2557) );
  MUX U1151 ( .IN0(n3049), .IN1(n574), .SEL(n3050), .F(n2917) );
  IV U1152 ( .A(n3051), .Z(n574) );
  MUX U1153 ( .IN0(A[10]), .IN1(n5384), .SEL(A[31]), .F(n575) );
  IV U1154 ( .A(n575), .Z(n2486) );
  MUX U1155 ( .IN0(A[6]), .IN1(n5513), .SEL(A[31]), .F(n576) );
  IV U1156 ( .A(n576), .Z(n2972) );
  MUX U1157 ( .IN0(A[5]), .IN1(n5529), .SEL(A[31]), .F(n577) );
  IV U1158 ( .A(n577), .Z(n3104) );
  MUX U1159 ( .IN0(n4723), .IN1(n4220), .SEL(n4221), .F(n4703) );
  XNOR U1160 ( .A(n4959), .B(n4957), .Z(n4964) );
  MUX U1161 ( .IN0(n3422), .IN1(n3420), .SEL(n3421), .F(n3289) );
  MUX U1162 ( .IN0(n1101), .IN1(n578), .SEL(n1102), .F(n1059) );
  IV U1163 ( .A(n1103), .Z(n578) );
  MUX U1164 ( .IN0(n647), .IN1(n1569), .SEL(n1568), .F(n1480) );
  MUX U1165 ( .IN0(n1941), .IN1(n1939), .SEL(n1940), .F(n1843) );
  MUX U1166 ( .IN0(n579), .IN1(n2160), .SEL(n2161), .F(n2059) );
  IV U1167 ( .A(n2162), .Z(n579) );
  MUX U1168 ( .IN0(n2820), .IN1(n2818), .SEL(n2819), .F(n2696) );
  MUX U1169 ( .IN0(n2757), .IN1(n2755), .SEL(n2756), .F(n2635) );
  MUX U1170 ( .IN0(n2887), .IN1(n2885), .SEL(n2886), .F(n2763) );
  MUX U1171 ( .IN0(n3345), .IN1(n3343), .SEL(n3344), .F(n3207) );
  MUX U1172 ( .IN0(n3267), .IN1(n3265), .SEL(n3266), .F(n3131) );
  XNOR U1173 ( .A(n3359), .B(n3358), .Z(n5499) );
  XNOR U1174 ( .A(n3320), .B(n3319), .Z(n5129) );
  XNOR U1175 ( .A(n3273), .B(n3272), .Z(n3398) );
  MUX U1176 ( .IN0(n1326), .IN1(n1324), .SEL(n1325), .F(n1252) );
  MUX U1177 ( .IN0(n1157), .IN1(n1155), .SEL(n1156), .F(n1096) );
  XNOR U1178 ( .A(n1362), .B(n1361), .Z(n1429) );
  MUX U1179 ( .IN0(n1488), .IN1(n580), .SEL(n1487), .F(n1404) );
  IV U1180 ( .A(n1486), .Z(n580) );
  XNOR U1181 ( .A(n1426), .B(n1425), .Z(n1499) );
  XNOR U1182 ( .A(n1762), .B(n1761), .Z(n1854) );
  XNOR U1183 ( .A(n1770), .B(n1769), .Z(n1862) );
  XNOR U1184 ( .A(n1816), .B(n1815), .Z(n1905) );
  MUX U1185 ( .IN0(n581), .IN1(n2025), .SEL(n2026), .F(n1929) );
  IV U1186 ( .A(n2027), .Z(n581) );
  XNOR U1187 ( .A(n2051), .B(n2050), .Z(n2147) );
  MUX U1188 ( .IN0(n582), .IN1(n2250), .SEL(n2251), .F(n2144) );
  IV U1189 ( .A(n2252), .Z(n582) );
  XNOR U1190 ( .A(n2219), .B(n2218), .Z(n2321) );
  XNOR U1191 ( .A(n2308), .B(n2307), .Z(n2410) );
  XNOR U1192 ( .A(n2349), .B(n2348), .Z(n2452) );
  MUX U1193 ( .IN0(n583), .IN1(n2568), .SEL(n2569), .F(n2449) );
  IV U1194 ( .A(n2570), .Z(n583) );
  MUX U1195 ( .IN0(n584), .IN1(n2625), .SEL(n2626), .F(n2508) );
  IV U1196 ( .A(n2627), .Z(n584) );
  XNOR U1197 ( .A(n2673), .B(n2672), .Z(n2790) );
  XNOR U1198 ( .A(n2712), .B(n2711), .Z(n2829) );
  XNOR U1199 ( .A(n2720), .B(n2719), .Z(n2837) );
  XNOR U1200 ( .A(n3020), .B(n2902), .Z(n2903) );
  MUX U1201 ( .IN0(n585), .IN1(n3199), .SEL(n3200), .F(n3067) );
  IV U1202 ( .A(n3201), .Z(n585) );
  MUX U1203 ( .IN0(n3217), .IN1(n655), .SEL(n3216), .F(n586) );
  IV U1204 ( .A(n586), .Z(n3083) );
  MUX U1205 ( .IN0(n587), .IN1(n3175), .SEL(n3176), .F(n3042) );
  IV U1206 ( .A(n3177), .Z(n587) );
  MUX U1207 ( .IN0(n940), .IN1(n942), .SEL(n941), .F(n910) );
  XNOR U1208 ( .A(n978), .B(n977), .Z(n1011) );
  MUX U1209 ( .IN0(n588), .IN1(n1088), .SEL(n1089), .F(n1046) );
  IV U1210 ( .A(n1090), .Z(n588) );
  MUX U1211 ( .IN0(n589), .IN1(n1262), .SEL(n1263), .F(n1195) );
  IV U1212 ( .A(n1264), .Z(n589) );
  MUX U1213 ( .IN0(n590), .IN1(n1552), .SEL(n1553), .F(n1474) );
  IV U1214 ( .A(n1554), .Z(n590) );
  AND U1215 ( .A(n1780), .B(n1782), .Z(n1689) );
  MUX U1216 ( .IN0(n591), .IN1(n1919), .SEL(n1920), .F(n1823) );
  IV U1217 ( .A(n1921), .Z(n591) );
  XNOR U1218 ( .A(n1801), .B(n1802), .Z(n1798) );
  AND U1219 ( .A(n2001), .B(n2003), .Z(n1901) );
  AND U1220 ( .A(n2170), .B(n2172), .Z(n2069) );
  MUX U1221 ( .IN0(n592), .IN1(n2441), .SEL(n2442), .F(n2333) );
  IV U1222 ( .A(n2443), .Z(n592) );
  AND U1223 ( .A(n2730), .B(n2732), .Z(n2610) );
  MUX U1224 ( .IN0(n593), .IN1(n2927), .SEL(n2928), .F(n2802) );
  IV U1225 ( .A(n2929), .Z(n593) );
  MUX U1226 ( .IN0(n594), .IN1(n3039), .SEL(n3040), .F(n2911) );
  IV U1227 ( .A(n3041), .Z(n594) );
  NAND U1228 ( .A(n905), .B(n904), .Z(n899) );
  XNOR U1229 ( .A(n943), .B(n968), .Z(n959) );
  ANDN U1230 ( .A(n1080), .B(n1081), .Z(n1036) );
  AND U1231 ( .A(n1128), .B(n1129), .Z(n1127) );
  ANDN U1232 ( .A(n1381), .B(n1382), .Z(n1314) );
  NAND U1233 ( .A(n1446), .B(n1448), .Z(n1373) );
  MUX U1234 ( .IN0(n595), .IN1(n2207), .SEL(n2208), .F(n2099) );
  IV U1235 ( .A(n2209), .Z(n595) );
  MUX U1236 ( .IN0(n596), .IN1(n2425), .SEL(n2426), .F(n2318) );
  IV U1237 ( .A(n2427), .Z(n596) );
  MUX U1238 ( .IN0(n597), .IN1(n2650), .SEL(n2651), .F(n2536) );
  IV U1239 ( .A(n2652), .Z(n597) );
  MUX U1240 ( .IN0(n3148), .IN1(n629), .SEL(n3147), .F(n598) );
  IV U1241 ( .A(n598), .Z(n3016) );
  XNOR U1242 ( .A(n916), .B(n921), .Z(n917) );
  XNOR U1243 ( .A(n1028), .B(n1033), .Z(n1029) );
  XNOR U1244 ( .A(n1175), .B(n1180), .Z(n1176) );
  XOR U1245 ( .A(n1614), .B(n1703), .Z(n1698) );
  XNOR U1246 ( .A(n3282), .B(n3281), .Z(n3116) );
  MUX U1247 ( .IN0(n1074), .IN1(Y0[24]), .SEL(n1075), .F(n1030) );
  MUX U1248 ( .IN0(n1308), .IN1(Y0[20]), .SEL(n1309), .F(n1240) );
  MUX U1249 ( .IN0(n1608), .IN1(Y0[16]), .SEL(n1609), .F(n1527) );
  MUX U1250 ( .IN0(n1976), .IN1(Y0[12]), .SEL(n1977), .F(n1880) );
  MUX U1251 ( .IN0(n2386), .IN1(Y0[8]), .SEL(n2387), .F(n2279) );
  MUX U1252 ( .IN0(Y0[4]), .IN1(n2854), .SEL(n2855), .F(n2733) );
  XNOR U1253 ( .A(n866), .B(n870), .Z(n868) );
  MUX U1254 ( .IN0(n4021), .IN1(n4019), .SEL(n4020), .F(n3973) );
  MUX U1255 ( .IN0(n4942), .IN1(n4492), .SEL(n4493), .F(n4925) );
  MUX U1256 ( .IN0(n599), .IN1(n4469), .SEL(n4009), .F(n4448) );
  IV U1257 ( .A(n4007), .Z(n599) );
  MUX U1258 ( .IN0(n4420), .IN1(n4418), .SEL(n4419), .F(n4397) );
  MUX U1259 ( .IN0(n3910), .IN1(n3908), .SEL(n3909), .F(n3864) );
  MUX U1260 ( .IN0(n600), .IN1(n3943), .SEL(n3944), .F(n3897) );
  IV U1261 ( .A(n3945), .Z(n600) );
  MUX U1262 ( .IN0(n3839), .IN1(n3837), .SEL(n3838), .F(n3791) );
  MUX U1263 ( .IN0(n4874), .IN1(n4408), .SEL(n4409), .F(n4857) );
  MUX U1264 ( .IN0(n4672), .IN1(n4670), .SEL(n4671), .F(n4648) );
  MUX U1265 ( .IN0(n601), .IN1(n4385), .SEL(n3827), .F(n4364) );
  IV U1266 ( .A(n3825), .Z(n601) );
  MUX U1267 ( .IN0(n5043), .IN1(n4655), .SEL(n4657), .F(n5031) );
  MUX U1268 ( .IN0(n4336), .IN1(n4334), .SEL(n4335), .F(n4313) );
  MUX U1269 ( .IN0(n3728), .IN1(n3726), .SEL(n3727), .F(n3682) );
  MUX U1270 ( .IN0(n602), .IN1(n3761), .SEL(n3762), .F(n3715) );
  IV U1271 ( .A(n3763), .Z(n602) );
  MUX U1272 ( .IN0(n3657), .IN1(n3655), .SEL(n3656), .F(n3612) );
  MUX U1273 ( .IN0(n4806), .IN1(n4324), .SEL(n4325), .F(n4789) );
  MUX U1274 ( .IN0(n5109), .IN1(n4695), .SEL(n4696), .F(n603) );
  IV U1275 ( .A(n603), .Z(n5095) );
  MUX U1276 ( .IN0(n5227), .IN1(n5225), .SEL(n5226), .F(n5205) );
  MUX U1277 ( .IN0(n4586), .IN1(n4584), .SEL(n4585), .F(n4564) );
  MUX U1278 ( .IN0(n604), .IN1(n4301), .SEL(n3645), .F(n4280) );
  IV U1279 ( .A(n3643), .Z(n604) );
  MUX U1280 ( .IN0(n5362), .IN1(n5212), .SEL(n5214), .F(n5350) );
  MUX U1281 ( .IN0(n4176), .IN1(n4178), .SEL(n4177), .F(n4173) );
  MUX U1282 ( .IN0(n4989), .IN1(n4571), .SEL(n4573), .F(n4979) );
  MUX U1283 ( .IN0(n4253), .IN1(n4251), .SEL(n4252), .F(n4230) );
  MUX U1284 ( .IN0(n3553), .IN1(n3551), .SEL(n3552), .F(n3509) );
  MUX U1285 ( .IN0(n605), .IN1(n3583), .SEL(n3584), .F(n3541) );
  IV U1286 ( .A(n3585), .Z(n605) );
  MUX U1287 ( .IN0(n3484), .IN1(n3482), .SEL(n3483), .F(n3442) );
  MUX U1288 ( .IN0(n606), .IN1(n4097), .SEL(n4098), .F(n4072) );
  IV U1289 ( .A(n4099), .Z(n606) );
  XNOR U1290 ( .A(n5578), .B(A[3]), .Z(n5579) );
  MUX U1291 ( .IN0(n4740), .IN1(n4241), .SEL(n4242), .F(n4723) );
  MUX U1292 ( .IN0(n5580), .IN1(n607), .SEL(n5581), .F(n3364) );
  MUX U1293 ( .IN0(n2462), .IN1(n2464), .SEL(n2463), .F(n2354) );
  MUX U1294 ( .IN0(n2717), .IN1(n608), .SEL(n2718), .F(n2597) );
  IV U1295 ( .A(n2719), .Z(n608) );
  MUX U1296 ( .IN0(n2932), .IN1(n2934), .SEL(n2933), .F(n2807) );
  MUX U1297 ( .IN0(n2889), .IN1(n2891), .SEL(n2890), .F(n2767) );
  MUX U1298 ( .IN0(n3212), .IN1(n3214), .SEL(n3213), .F(n3080) );
  XNOR U1299 ( .A(n5419), .B(n5418), .Z(n5424) );
  XNOR U1300 ( .A(n5134), .B(n5133), .Z(n5160) );
  XNOR U1301 ( .A(n4502), .B(n4500), .Z(n4515) );
  MUX U1302 ( .IN0(n609), .IN1(n4218), .SEL(n3473), .F(n4198) );
  IV U1303 ( .A(n3471), .Z(n609) );
  MUX U1304 ( .IN0(n1287), .IN1(n1285), .SEL(n1286), .F(n1217) );
  MUX U1305 ( .IN0(n1364), .IN1(n1362), .SEL(n1363), .F(n1295) );
  MUX U1306 ( .IN0(n610), .IN1(n5486), .SEL(X[31]), .F(n1483) );
  IV U1307 ( .A(X[19]), .Z(n610) );
  MUX U1308 ( .IN0(n611), .IN1(n1770), .SEL(n1771), .F(n1679) );
  IV U1309 ( .A(n1772), .Z(n611) );
  MUX U1310 ( .IN0(n612), .IN1(n4183), .SEL(X[31]), .F(n1988) );
  IV U1311 ( .A(X[13]), .Z(n612) );
  MUX U1312 ( .IN0(n2012), .IN1(n2010), .SEL(n2011), .F(n1912) );
  MUX U1313 ( .IN0(n2202), .IN1(n2200), .SEL(n2201), .F(n2083) );
  MUX U1314 ( .IN0(n613), .IN1(n2481), .SEL(n2482), .F(n2373) );
  IV U1315 ( .A(n2483), .Z(n613) );
  MUX U1316 ( .IN0(n2714), .IN1(n2712), .SEL(n2713), .F(n2592) );
  MUX U1317 ( .IN0(n3291), .IN1(n3289), .SEL(n3290), .F(n3155) );
  XNOR U1318 ( .A(n3343), .B(n3342), .Z(n5319) );
  MUX U1319 ( .IN0(n614), .IN1(n3385), .SEL(n3386), .F(n3257) );
  IV U1320 ( .A(n3387), .Z(n614) );
  XOR U1321 ( .A(n1318), .B(n1256), .Z(n1253) );
  MUX U1322 ( .IN0(n615), .IN1(n1416), .SEL(n1417), .F(n1344) );
  IV U1323 ( .A(n1418), .Z(n615) );
  ANDN U1324 ( .A(n1480), .B(n1479), .Z(n1407) );
  XNOR U1325 ( .A(n1585), .B(n1584), .Z(n1662) );
  MUX U1326 ( .IN0(n1642), .IN1(n616), .SEL(n1643), .F(n1565) );
  IV U1327 ( .A(n1644), .Z(n616) );
  XNOR U1328 ( .A(n1955), .B(n1954), .Z(n2046) );
  XNOR U1329 ( .A(n1939), .B(n1938), .Z(n2028) );
  MUX U1330 ( .IN0(n617), .IN1(n2126), .SEL(n2127), .F(n2025) );
  IV U1331 ( .A(n2128), .Z(n617) );
  MUX U1332 ( .IN0(n618), .IN1(n2144), .SEL(n2145), .F(n2043) );
  IV U1333 ( .A(n2146), .Z(n618) );
  XNOR U1334 ( .A(n2059), .B(n2058), .Z(n2155) );
  XNOR U1335 ( .A(n2242), .B(n2241), .Z(n2344) );
  MUX U1336 ( .IN0(n619), .IN1(n2584), .SEL(n2585), .F(n2465) );
  IV U1337 ( .A(n2586), .Z(n619) );
  XNOR U1338 ( .A(n2512), .B(n2522), .Z(n2628) );
  XNOR U1339 ( .A(n2529), .B(n2528), .Z(n2638) );
  XNOR U1340 ( .A(n2553), .B(n2552), .Z(n2668) );
  XNOR U1341 ( .A(n2576), .B(n2575), .Z(n2691) );
  MUX U1342 ( .IN0(n620), .IN1(n2810), .SEL(n2811), .F(n2688) );
  IV U1343 ( .A(n2812), .Z(n620) );
  XNOR U1344 ( .A(n2885), .B(n2884), .Z(n3004) );
  XNOR U1345 ( .A(n2877), .B(n2876), .Z(n2996) );
  XNOR U1346 ( .A(n2943), .B(n2942), .Z(n3070) );
  XNOR U1347 ( .A(n3052), .B(n3051), .Z(n3179) );
  XNOR U1348 ( .A(n3091), .B(n3090), .Z(n3218) );
  XNOR U1349 ( .A(n3099), .B(n3098), .Z(n3226) );
  MUX U1350 ( .IN0(n945), .IN1(n943), .SEL(n944), .F(n913) );
  NAND U1351 ( .A(n1056), .B(n1055), .Z(n1049) );
  XNOR U1352 ( .A(n1018), .B(n1017), .Z(n1057) );
  MUX U1353 ( .IN0(n621), .IN1(n1144), .SEL(n1145), .F(n1088) );
  IV U1354 ( .A(n1146), .Z(n621) );
  AND U1355 ( .A(n1689), .B(n1691), .Z(n1605) );
  MUX U1356 ( .IN0(n622), .IN1(n1723), .SEL(n1724), .F(n1632) );
  IV U1357 ( .A(n1725), .Z(n622) );
  MUX U1358 ( .IN0(n623), .IN1(n2226), .SEL(n2227), .F(n2118) );
  IV U1359 ( .A(n2228), .Z(n623) );
  AND U1360 ( .A(n2276), .B(n2278), .Z(n2170) );
  MUX U1361 ( .IN0(n624), .IN1(n2680), .SEL(n2681), .F(n2560) );
  IV U1362 ( .A(n2682), .Z(n624) );
  XNOR U1363 ( .A(n2661), .B(n2660), .Z(n2658) );
  ANDN U1364 ( .A(n2852), .B(n2853), .Z(n2730) );
  MUX U1365 ( .IN0(n3042), .IN1(n3165), .SEL(n3044), .F(n2909) );
  MUX U1366 ( .IN0(n3193), .IN1(n718), .SEL(n3192), .F(n625) );
  IV U1367 ( .A(n625), .Z(n3059) );
  MUX U1368 ( .IN0(n626), .IN1(n3162), .SEL(n3163), .F(n3039) );
  IV U1369 ( .A(n3164), .Z(n626) );
  ANDN U1370 ( .A(n987), .B(n957), .Z(n946) );
  MUX U1371 ( .IN0(n1189), .IN1(n1191), .SEL(n1190), .F(n627) );
  IV U1372 ( .A(n627), .Z(n1134) );
  AND U1373 ( .A(n1246), .B(n1248), .Z(n1183) );
  XOR U1374 ( .A(n1198), .B(n1195), .Z(n1249) );
  NANDN U1375 ( .B(n1306), .A(n1307), .Z(n1238) );
  XNOR U1376 ( .A(n1983), .B(n1984), .Z(n2003) );
  MUX U1377 ( .IN0(n628), .IN1(n2770), .SEL(n2771), .F(n2650) );
  IV U1378 ( .A(n2772), .Z(n628) );
  MUX U1379 ( .IN0(n3282), .IN1(n3280), .SEL(n3281), .F(n629) );
  IV U1380 ( .A(n629), .Z(n3146) );
  MUX U1381 ( .IN0(n883), .IN1(n881), .SEL(n882), .F(n630) );
  IV U1382 ( .A(n630), .Z(n860) );
  NANDN U1383 ( .B(n887), .A(n888), .Z(n844) );
  XOR U1384 ( .A(n1476), .B(n1475), .Z(n1456) );
  XOR U1385 ( .A(n1705), .B(n1704), .Z(n1789) );
  XOR U1386 ( .A(n2318), .B(n2315), .Z(n2392) );
  AND U1387 ( .A(n872), .B(n874), .Z(n847) );
  MUX U1388 ( .IN0(n3241), .IN1(Y0[1]), .SEL(n3242), .F(n3109) );
  XNOR U1389 ( .A(n918), .B(n922), .Z(n920) );
  XNOR U1390 ( .A(n1030), .B(n1034), .Z(n1032) );
  XNOR U1391 ( .A(n1177), .B(n1181), .Z(n1179) );
  XNOR U1392 ( .A(n1375), .B(n1379), .Z(n1377) );
  XNOR U1393 ( .A(n1608), .B(n1612), .Z(n1610) );
  XNOR U1394 ( .A(n1880), .B(n1884), .Z(n1882) );
  XNOR U1395 ( .A(n2173), .B(n2177), .Z(n2175) );
  XNOR U1396 ( .A(n2494), .B(n2498), .Z(n2496) );
  MUX U1397 ( .IN0(n631), .IN1(n4511), .SEL(n4094), .F(n4490) );
  IV U1398 ( .A(n4093), .Z(n631) );
  MUX U1399 ( .IN0(n3975), .IN1(n3973), .SEL(n3974), .F(n3927) );
  MUX U1400 ( .IN0(n4462), .IN1(n4460), .SEL(n4461), .F(n4439) );
  MUX U1401 ( .IN0(n4908), .IN1(n4450), .SEL(n4451), .F(n4891) );
  MUX U1402 ( .IN0(n632), .IN1(n3897), .SEL(n3898), .F(n3853) );
  IV U1403 ( .A(n3899), .Z(n632) );
  MUX U1404 ( .IN0(n633), .IN1(n4427), .SEL(n3917), .F(n4406) );
  IV U1405 ( .A(n3915), .Z(n633) );
  MUX U1406 ( .IN0(n3793), .IN1(n3791), .SEL(n3792), .F(n3745) );
  MUX U1407 ( .IN0(n4378), .IN1(n4376), .SEL(n4377), .F(n4355) );
  MUX U1408 ( .IN0(n3820), .IN1(n3818), .SEL(n3819), .F(n3772) );
  MUX U1409 ( .IN0(n4840), .IN1(n4366), .SEL(n4367), .F(n4823) );
  MUX U1410 ( .IN0(n4189), .IN1(n4673), .SEL(n4190), .F(n634) );
  IV U1411 ( .A(n634), .Z(n4651) );
  MUX U1412 ( .IN0(n5031), .IN1(n4631), .SEL(n4633), .F(n5016) );
  MUX U1413 ( .IN0(n4626), .IN1(n4624), .SEL(n4625), .F(n4604) );
  MUX U1414 ( .IN0(n635), .IN1(n3715), .SEL(n3716), .F(n3671) );
  IV U1415 ( .A(n3717), .Z(n635) );
  MUX U1416 ( .IN0(n636), .IN1(n4343), .SEL(n3735), .F(n4322) );
  IV U1417 ( .A(n3733), .Z(n636) );
  MUX U1418 ( .IN0(n5249), .IN1(n5247), .SEL(n5248), .F(n5225) );
  MUX U1419 ( .IN0(n5388), .IN1(n5254), .SEL(n5256), .F(n5374) );
  MUX U1420 ( .IN0(n3614), .IN1(n3612), .SEL(n3613), .F(n3569) );
  MUX U1421 ( .IN0(n4294), .IN1(n4292), .SEL(n4293), .F(n4271) );
  MUX U1422 ( .IN0(n3638), .IN1(n3636), .SEL(n3637), .F(n3594) );
  MUX U1423 ( .IN0(n4773), .IN1(n4282), .SEL(n4283), .F(n4757) );
  MUX U1424 ( .IN0(A[1]), .IN1(n5595), .SEL(A[31]), .F(n637) );
  IV U1425 ( .A(n637), .Z(n4163) );
  MUX U1426 ( .IN0(n638), .IN1(n5514), .SEL(n5515), .F(n5503) );
  IV U1427 ( .A(n5516), .Z(n638) );
  MUX U1428 ( .IN0(n4979), .IN1(n4551), .SEL(n4553), .F(n4969) );
  MUX U1429 ( .IN0(n4546), .IN1(n4544), .SEL(n4545), .F(n4520) );
  MUX U1430 ( .IN0(n639), .IN1(n3541), .SEL(n3542), .F(n3498) );
  IV U1431 ( .A(n3543), .Z(n639) );
  MUX U1432 ( .IN0(n640), .IN1(n4260), .SEL(n3560), .F(n4239) );
  IV U1433 ( .A(n3558), .Z(n640) );
  XNOR U1434 ( .A(n5501), .B(A[7]), .Z(n5502) );
  XNOR U1435 ( .A(n5369), .B(A[11]), .Z(n5370) );
  XNOR U1436 ( .A(n5321), .B(A[15]), .Z(n5322) );
  XNOR U1437 ( .A(n4832), .B(A[23]), .Z(n4833) );
  XNOR U1438 ( .A(n4900), .B(A[19]), .Z(n4901) );
  MUX U1439 ( .IN0(A[2]), .IN1(n5588), .SEL(A[31]), .F(n641) );
  IV U1440 ( .A(n641), .Z(n4160) );
  MUX U1441 ( .IN0(n5167), .IN1(n5165), .SEL(n5166), .F(n5134) );
  MUX U1442 ( .IN0(n5338), .IN1(n5172), .SEL(n5174), .F(n5326) );
  MUX U1443 ( .IN0(n3444), .IN1(n3442), .SEL(n3443), .F(n3403) );
  MUX U1444 ( .IN0(n3466), .IN1(n3464), .SEL(n3465), .F(n3395) );
  XNOR U1445 ( .A(n4766), .B(A[27]), .Z(n4767) );
  MUX U1446 ( .IN0(n642), .IN1(n4170), .SEL(X[31]), .F(n2404) );
  IV U1447 ( .A(X[9]), .Z(n642) );
  MUX U1448 ( .IN0(n2924), .IN1(n2926), .SEL(n2925), .F(n2799) );
  MUX U1449 ( .IN0(n3143), .IN1(n3145), .SEL(n3144), .F(n3013) );
  MUX U1450 ( .IN0(A[4]), .IN1(n5547), .SEL(A[31]), .F(n3102) );
  MUX U1451 ( .IN0(n3364), .IN1(n643), .SEL(n3365), .F(n3228) );
  IV U1452 ( .A(n3366), .Z(n643) );
  MUX U1453 ( .IN0(A[9]), .IN1(n5398), .SEL(A[31]), .F(n644) );
  IV U1454 ( .A(n644), .Z(n2605) );
  MUX U1455 ( .IN0(n3332), .IN1(n3334), .SEL(n3333), .F(n3196) );
  MUX U1456 ( .IN0(X[1]), .IN1(n5127), .SEL(X[31]), .F(n645) );
  IV U1457 ( .A(n645), .Z(n4700) );
  XNOR U1458 ( .A(n4088), .B(n4086), .Z(n4102) );
  MUX U1459 ( .IN0(n1428), .IN1(n1426), .SEL(n1427), .F(n1354) );
  MUX U1460 ( .IN0(n646), .IN1(n1595), .SEL(n1596), .F(n1514) );
  IV U1461 ( .A(n1597), .Z(n646) );
  MUX U1462 ( .IN0(n1627), .IN1(n1625), .SEL(n1626), .F(n1543) );
  MUX U1463 ( .IN0(n1651), .IN1(n1653), .SEL(n1652), .F(n647) );
  MUX U1464 ( .IN0(n2053), .IN1(n2051), .SEL(n2052), .F(n1955) );
  MUX U1465 ( .IN0(n2637), .IN1(n2635), .SEL(n2636), .F(n2512) );
  MUX U1466 ( .IN0(n3157), .IN1(n3155), .SEL(n3156), .F(n3021) );
  MUX U1467 ( .IN0(n4703), .IN1(n4216), .SEL(n4217), .F(n648) );
  IV U1468 ( .A(n648), .Z(n3310) );
  XNOR U1469 ( .A(n5297), .B(n5294), .Z(n5295) );
  XNOR U1470 ( .A(n5600), .B(X[30]), .Z(n5598) );
  MUX U1471 ( .IN0(n649), .IN1(n1207), .SEL(n1208), .F(n1144) );
  IV U1472 ( .A(n1209), .Z(n649) );
  XNOR U1473 ( .A(n1669), .B(n1668), .Z(n1757) );
  MUX U1474 ( .IN0(n650), .IN1(n1833), .SEL(n1834), .F(n1733) );
  IV U1475 ( .A(n1835), .Z(n650) );
  MUX U1476 ( .IN0(n651), .IN1(n1947), .SEL(n1948), .F(n1851) );
  IV U1477 ( .A(n1949), .Z(n651) );
  XNOR U1478 ( .A(n1867), .B(n1866), .Z(n1958) );
  XNOR U1479 ( .A(n1912), .B(n1911), .Z(n2005) );
  XNOR U1480 ( .A(n2035), .B(n2034), .Z(n2129) );
  XNOR U1481 ( .A(n2200), .B(n2199), .Z(n2301) );
  XNOR U1482 ( .A(n2365), .B(n2364), .Z(n2468) );
  XNOR U1483 ( .A(n2373), .B(n2372), .Z(n2476) );
  XNOR U1484 ( .A(n2326), .B(n2325), .Z(n2429) );
  MUX U1485 ( .IN0(n652), .IN1(n2449), .SEL(n2450), .F(n2341) );
  IV U1486 ( .A(n2451), .Z(n652) );
  XNOR U1487 ( .A(n2696), .B(n2695), .Z(n2813) );
  MUX U1488 ( .IN0(n653), .IN1(n2826), .SEL(n2827), .F(n2704) );
  IV U1489 ( .A(n2828), .Z(n653) );
  XNOR U1490 ( .A(n2643), .B(n2642), .Z(n2758) );
  MUX U1491 ( .IN0(n654), .IN1(n2745), .SEL(n2746), .F(n2625) );
  IV U1492 ( .A(n2747), .Z(n654) );
  XNOR U1493 ( .A(n2959), .B(n2958), .Z(n3086) );
  XNOR U1494 ( .A(n2967), .B(n2966), .Z(n3094) );
  XNOR U1495 ( .A(n2920), .B(n2919), .Z(n3047) );
  XNOR U1496 ( .A(n3075), .B(n3074), .Z(n3202) );
  XNOR U1497 ( .A(n3009), .B(n3008), .Z(n3134) );
  XNOR U1498 ( .A(n3001), .B(n3000), .Z(n3126) );
  MUX U1499 ( .IN0(n3353), .IN1(n3351), .SEL(n3352), .F(n655) );
  IV U1500 ( .A(n655), .Z(n3215) );
  MUX U1501 ( .IN0(n656), .IN1(n3335), .SEL(n3336), .F(n3199) );
  IV U1502 ( .A(n3337), .Z(n656) );
  MUX U1503 ( .IN0(n657), .IN1(n3257), .SEL(n3258), .F(n3123) );
  IV U1504 ( .A(n3259), .Z(n657) );
  MUX U1505 ( .IN0(n3307), .IN1(n658), .SEL(n3308), .F(n3175) );
  IV U1506 ( .A(n3309), .Z(n658) );
  MUX U1507 ( .IN0(n936), .IN1(n934), .SEL(n935), .F(n901) );
  MUX U1508 ( .IN0(n659), .IN1(n1005), .SEL(n1006), .F(n969) );
  IV U1509 ( .A(n1007), .Z(n659) );
  XNOR U1510 ( .A(n1062), .B(n1061), .Z(n1099) );
  XNOR U1511 ( .A(n1096), .B(n1094), .Z(n1147) );
  AND U1512 ( .A(n1198), .B(n1199), .Z(n1128) );
  MUX U1513 ( .IN0(n660), .IN1(n1331), .SEL(n1332), .F(n1262) );
  IV U1514 ( .A(n1333), .Z(n660) );
  XOR U1515 ( .A(n1404), .B(n1408), .Z(n1477) );
  XNOR U1516 ( .A(n1890), .B(n1889), .Z(n1888) );
  MUX U1517 ( .IN0(n661), .IN1(n2017), .SEL(n2018), .F(n1919) );
  IV U1518 ( .A(n2019), .Z(n661) );
  AND U1519 ( .A(n2069), .B(n2071), .Z(n1973) );
  MUX U1520 ( .IN0(n662), .IN1(n2081), .SEL(n2080), .F(n1984) );
  IV U1521 ( .A(n2079), .Z(n662) );
  AND U1522 ( .A(n2491), .B(n2493), .Z(n2383) );
  MUX U1523 ( .IN0(n663), .IN1(n2560), .SEL(n2561), .F(n2441) );
  IV U1524 ( .A(n2562), .Z(n663) );
  MUX U1525 ( .IN0(n664), .IN1(n3059), .SEL(n3060), .F(n2927) );
  IV U1526 ( .A(n3061), .Z(n664) );
  MUX U1527 ( .IN0(n910), .IN1(n912), .SEL(n911), .F(n878) );
  AND U1528 ( .A(n1133), .B(n1134), .Z(n1130) );
  MUX U1529 ( .IN0(n665), .IN1(n2099), .SEL(n2100), .F(n1998) );
  IV U1530 ( .A(n2101), .Z(n665) );
  XOR U1531 ( .A(n2539), .B(n2425), .Z(n2426) );
  XNOR U1532 ( .A(n2786), .B(n2784), .Z(n2895) );
  NANDN U1533 ( .B(n885), .A(n884), .Z(n856) );
  XNOR U1534 ( .A(n887), .B(n892), .Z(n888) );
  XNOR U1535 ( .A(n988), .B(n993), .Z(n989) );
  XNOR U1536 ( .A(n1116), .B(n1081), .Z(n1117) );
  XNOR U1537 ( .A(n1306), .B(n1311), .Z(n1307) );
  XOR U1538 ( .A(n1554), .B(n1553), .Z(n1534) );
  MUX U1539 ( .IN0(Y0[2]), .IN1(n3109), .SEL(n3110), .F(n2977) );
  XOR U1540 ( .A(n1707), .B(n1706), .Z(n1786) );
  XOR U1541 ( .A(n2317), .B(n2316), .Z(n2389) );
  XOR U1542 ( .A(n2652), .B(n2651), .Z(n2736) );
  XNOR U1543 ( .A(n2982), .B(n2861), .Z(n2862) );
  XOR U1544 ( .A(n3148), .B(n3147), .Z(n3248) );
  XNOR U1545 ( .A(n949), .B(n953), .Z(n951) );
  XNOR U1546 ( .A(n1074), .B(n1078), .Z(n1076) );
  XNOR U1547 ( .A(n1240), .B(n1244), .Z(n1242) );
  XNOR U1548 ( .A(n1449), .B(n1453), .Z(n1451) );
  XNOR U1549 ( .A(n1692), .B(n1696), .Z(n1694) );
  XNOR U1550 ( .A(n1976), .B(n1980), .Z(n1978) );
  XNOR U1551 ( .A(n2279), .B(n2283), .Z(n2281) );
  XNOR U1552 ( .A(n2613), .B(n2617), .Z(n2615) );
  XOR U1553 ( .A(n832), .B(n833), .Z(n722) );
  MUX U1554 ( .IN0(n4065), .IN1(n4063), .SEL(n4064), .F(n4019) );
  MUX U1555 ( .IN0(n4048), .IN1(n4046), .SEL(n4047), .F(n4000) );
  MUX U1556 ( .IN0(n666), .IN1(n3989), .SEL(n3990), .F(n3943) );
  IV U1557 ( .A(n3991), .Z(n666) );
  MUX U1558 ( .IN0(n3885), .IN1(n3883), .SEL(n3884), .F(n3837) );
  MUX U1559 ( .IN0(n667), .IN1(n4448), .SEL(n3963), .F(n4427) );
  IV U1560 ( .A(n3961), .Z(n667) );
  MUX U1561 ( .IN0(n4891), .IN1(n4429), .SEL(n4430), .F(n4874) );
  MUX U1562 ( .IN0(n4399), .IN1(n4397), .SEL(n4398), .F(n4376) );
  MUX U1563 ( .IN0(n3866), .IN1(n3864), .SEL(n3865), .F(n3818) );
  MUX U1564 ( .IN0(n668), .IN1(n3807), .SEL(n3808), .F(n3761) );
  IV U1565 ( .A(n3809), .Z(n668) );
  MUX U1566 ( .IN0(n3703), .IN1(n3701), .SEL(n3702), .F(n3655) );
  MUX U1567 ( .IN0(n669), .IN1(n4364), .SEL(n3781), .F(n4343) );
  IV U1568 ( .A(n3779), .Z(n669) );
  MUX U1569 ( .IN0(n4823), .IN1(n4345), .SEL(n4346), .F(n4806) );
  MUX U1570 ( .IN0(n5273), .IN1(n5271), .SEL(n5272), .F(n5247) );
  MUX U1571 ( .IN0(n5405), .IN1(n5278), .SEL(n5280), .F(n5388) );
  MUX U1572 ( .IN0(n4315), .IN1(n4313), .SEL(n4314), .F(n4292) );
  MUX U1573 ( .IN0(n3684), .IN1(n3682), .SEL(n3683), .F(n3636) );
  MUX U1574 ( .IN0(n5016), .IN1(n4611), .SEL(n4613), .F(n5001) );
  MUX U1575 ( .IN0(n4606), .IN1(n4604), .SEL(n4605), .F(n4584) );
  MUX U1576 ( .IN0(n5473), .IN1(n5317), .SEL(n5318), .F(n670) );
  IV U1577 ( .A(n670), .Z(n5459) );
  MUX U1578 ( .IN0(n4149), .IN1(n4100), .SEL(n4101), .F(n671) );
  IV U1579 ( .A(n671), .Z(n4135) );
  MUX U1580 ( .IN0(n672), .IN1(n4132), .SEL(n4133), .F(n4118) );
  IV U1581 ( .A(n4134), .Z(n672) );
  MUX U1582 ( .IN0(n673), .IN1(n3626), .SEL(n3627), .F(n3583) );
  IV U1583 ( .A(n3628), .Z(n673) );
  MUX U1584 ( .IN0(n5556), .IN1(n5497), .SEL(n5498), .F(n674) );
  IV U1585 ( .A(n674), .Z(n5540) );
  MUX U1586 ( .IN0(n3529), .IN1(n3527), .SEL(n3528), .F(n3482) );
  MUX U1587 ( .IN0(n675), .IN1(n4280), .SEL(n3603), .F(n4260) );
  IV U1588 ( .A(n3601), .Z(n675) );
  MUX U1589 ( .IN0(n4757), .IN1(n4262), .SEL(n4263), .F(n4740) );
  MUX U1590 ( .IN0(n5584), .IN1(n5586), .SEL(n5585), .F(n5580) );
  MUX U1591 ( .IN0(n5187), .IN1(n5185), .SEL(n5186), .F(n5165) );
  MUX U1592 ( .IN0(n5350), .IN1(n5192), .SEL(n5194), .F(n5338) );
  MUX U1593 ( .IN0(n676), .IN1(n4104), .SEL(n4105), .F(n4082) );
  IV U1594 ( .A(n4106), .Z(n676) );
  MUX U1595 ( .IN0(n4232), .IN1(n4230), .SEL(n4231), .F(n4206) );
  MUX U1596 ( .IN0(n3511), .IN1(n3509), .SEL(n3510), .F(n3464) );
  XNOR U1597 ( .A(n5528), .B(A[5]), .Z(n5529) );
  XNOR U1598 ( .A(n5397), .B(A[9]), .Z(n5398) );
  MUX U1599 ( .IN0(n677), .IN1(n5311), .SEL(X[31]), .F(n5303) );
  IV U1600 ( .A(X[21]), .Z(n677) );
  XNOR U1601 ( .A(n5345), .B(A[13]), .Z(n5346) );
  XNOR U1602 ( .A(n4934), .B(A[17]), .Z(n4935) );
  XNOR U1603 ( .A(n4866), .B(A[21]), .Z(n4867) );
  AND U1604 ( .A(n5596), .B(A[0]), .Z(n3374) );
  MUX U1605 ( .IN0(n4522), .IN1(n4520), .SEL(n4521), .F(n4502) );
  MUX U1606 ( .IN0(n4969), .IN1(n4531), .SEL(n4533), .F(n4959) );
  MUX U1607 ( .IN0(n678), .IN1(n5575), .SEL(X[31]), .F(n5562) );
  IV U1608 ( .A(X[25]), .Z(n678) );
  XNOR U1609 ( .A(n4798), .B(A[25]), .Z(n4799) );
  MUX U1610 ( .IN0(n679), .IN1(n5593), .SEL(X[31]), .F(n5583) );
  IV U1611 ( .A(X[29]), .Z(n679) );
  MUX U1612 ( .IN0(A[3]), .IN1(n5579), .SEL(A[31]), .F(n3234) );
  MUX U1613 ( .IN0(n3348), .IN1(n3350), .SEL(n3349), .F(n3212) );
  MUX U1614 ( .IN0(n3324), .IN1(n3326), .SEL(n3325), .F(n3188) );
  MUX U1615 ( .IN0(X[20]), .IN1(n680), .SEL(X[31]), .F(n1386) );
  IV U1616 ( .A(n5310), .Z(n680) );
  MUX U1617 ( .IN0(X[16]), .IN1(n681), .SEL(X[31]), .F(n1748) );
  IV U1618 ( .A(n5490), .Z(n681) );
  MUX U1619 ( .IN0(X[8]), .IN1(n682), .SEL(X[31]), .F(n2523) );
  IV U1620 ( .A(n4169), .Z(n682) );
  MUX U1621 ( .IN0(X[12]), .IN1(n683), .SEL(X[31]), .F(n2094) );
  IV U1622 ( .A(n4182), .Z(n683) );
  MUX U1623 ( .IN0(X[4]), .IN1(n684), .SEL(X[31]), .F(n3032) );
  IV U1624 ( .A(n4688), .Z(n684) );
  XNOR U1625 ( .A(n4676), .B(n4673), .Z(n4674) );
  MUX U1626 ( .IN0(n685), .IN1(n3454), .SEL(n3455), .F(n3385) );
  IV U1627 ( .A(n3456), .Z(n685) );
  MUX U1628 ( .IN0(n686), .IN1(n5569), .SEL(X[31]), .F(n1001) );
  IV U1629 ( .A(X[27]), .Z(n686) );
  MUX U1630 ( .IN0(X[26]), .IN1(n687), .SEL(X[31]), .F(n1042) );
  IV U1631 ( .A(n5570), .Z(n687) );
  MUX U1632 ( .IN0(X[24]), .IN1(n688), .SEL(X[31]), .F(n1149) );
  IV U1633 ( .A(n5574), .Z(n688) );
  MUX U1634 ( .IN0(X[28]), .IN1(n689), .SEL(X[31]), .F(n974) );
  IV U1635 ( .A(n5592), .Z(n689) );
  MUX U1636 ( .IN0(n1467), .IN1(n1465), .SEL(n1466), .F(n1392) );
  MUX U1637 ( .IN0(n690), .IN1(n1514), .SEL(n1515), .F(n1436) );
  IV U1638 ( .A(n1516), .Z(n690) );
  MUX U1639 ( .IN0(n1508), .IN1(n1506), .SEL(n1507), .F(n1426) );
  MUX U1640 ( .IN0(X[18]), .IN1(n691), .SEL(X[31]), .F(n1564) );
  IV U1641 ( .A(n5485), .Z(n691) );
  MUX U1642 ( .IN0(n692), .IN1(n5491), .SEL(X[31]), .F(n1648) );
  IV U1643 ( .A(X[17]), .Z(n692) );
  MUX U1644 ( .IN0(n1845), .IN1(n1843), .SEL(n1844), .F(n1737) );
  MUX U1645 ( .IN0(n1818), .IN1(n1816), .SEL(n1817), .F(n1714) );
  MUX U1646 ( .IN0(n1861), .IN1(n1859), .SEL(n1860), .F(n1762) );
  MUX U1647 ( .IN0(n693), .IN1(n1867), .SEL(n1868), .F(n1770) );
  IV U1648 ( .A(n1869), .Z(n693) );
  XNOR U1649 ( .A(n4732), .B(A[29]), .Z(n4733) );
  MUX U1650 ( .IN0(n694), .IN1(n4165), .SEL(X[31]), .F(n2187) );
  IV U1651 ( .A(X[11]), .Z(n694) );
  MUX U1652 ( .IN0(X[10]), .IN1(n695), .SEL(X[31]), .F(n2293) );
  IV U1653 ( .A(n4164), .Z(n695) );
  MUX U1654 ( .IN0(n2417), .IN1(n2415), .SEL(n2416), .F(n2308) );
  MUX U1655 ( .IN0(X[6]), .IN1(n696), .SEL(X[31]), .F(n2783) );
  IV U1656 ( .A(n4693), .Z(n696) );
  MUX U1657 ( .IN0(n697), .IN1(n4689), .SEL(X[31]), .F(n2899) );
  IV U1658 ( .A(X[5]), .Z(n697) );
  MUX U1659 ( .IN0(n698), .IN1(n5123), .SEL(X[31]), .F(n3172) );
  IV U1660 ( .A(X[3]), .Z(n698) );
  MUX U1661 ( .IN0(X[2]), .IN1(n699), .SEL(X[31]), .F(n3306) );
  IV U1662 ( .A(n5122), .Z(n699) );
  MUX U1663 ( .IN0(n4198), .IN1(n700), .SEL(n3435), .F(n3307) );
  IV U1664 ( .A(n3434), .Z(n700) );
  MUX U1665 ( .IN0(X[22]), .IN1(n701), .SEL(X[31]), .F(n1258) );
  IV U1666 ( .A(n5316), .Z(n701) );
  MUX U1667 ( .IN0(n702), .IN1(n5315), .SEL(X[31]), .F(n1188) );
  IV U1668 ( .A(X[23]), .Z(n702) );
  MUX U1669 ( .IN0(n703), .IN1(n1275), .SEL(n1276), .F(n1207) );
  IV U1670 ( .A(n1277), .Z(n703) );
  MUX U1671 ( .IN0(n704), .IN1(n1575), .SEL(n1576), .F(n1496) );
  IV U1672 ( .A(n1577), .Z(n704) );
  MUX U1673 ( .IN0(n1993), .IN1(n1991), .SEL(n1992), .F(n705) );
  MUX U1674 ( .IN0(X[14]), .IN1(n706), .SEL(X[31]), .F(n1897) );
  IV U1675 ( .A(n4187), .Z(n706) );
  MUX U1676 ( .IN0(n707), .IN1(n1929), .SEL(n1930), .F(n1833) );
  IV U1677 ( .A(n1931), .Z(n707) );
  XNOR U1678 ( .A(n2152), .B(n2151), .Z(n2253) );
  XNOR U1679 ( .A(n2160), .B(n2159), .Z(n2261) );
  XNOR U1680 ( .A(n2111), .B(n2110), .Z(n2214) );
  XNOR U1681 ( .A(n2136), .B(n2135), .Z(n2237) );
  MUX U1682 ( .IN0(n708), .IN1(n2341), .SEL(n2342), .F(n2234) );
  IV U1683 ( .A(n2343), .Z(n708) );
  MUX U1684 ( .IN0(n709), .IN1(n2357), .SEL(n2358), .F(n2250) );
  IV U1685 ( .A(n2359), .Z(n709) );
  MUX U1686 ( .IN0(n2297), .IN1(n2401), .SEL(n2299), .F(n2189) );
  XNOR U1687 ( .A(n2457), .B(n2456), .Z(n2571) );
  XNOR U1688 ( .A(n2434), .B(n2433), .Z(n2548) );
  XNOR U1689 ( .A(n2473), .B(n2472), .Z(n2587) );
  XNOR U1690 ( .A(n2481), .B(n2480), .Z(n2595) );
  MUX U1691 ( .IN0(n710), .IN1(n2508), .SEL(n2509), .F(n2398) );
  IV U1692 ( .A(n2510), .Z(n710) );
  MUX U1693 ( .IN0(n711), .IN1(n4694), .SEL(X[31]), .F(n2657) );
  IV U1694 ( .A(X[7]), .Z(n711) );
  XNOR U1695 ( .A(n2842), .B(n2841), .Z(n2962) );
  XNOR U1696 ( .A(n2834), .B(n2833), .Z(n2954) );
  XNOR U1697 ( .A(n2795), .B(n2794), .Z(n2915) );
  XNOR U1698 ( .A(n2818), .B(n2817), .Z(n2938) );
  XNOR U1699 ( .A(n2755), .B(n2754), .Z(n2872) );
  XNOR U1700 ( .A(n2763), .B(n2762), .Z(n2880) );
  MUX U1701 ( .IN0(n712), .IN1(n2993), .SEL(n2994), .F(n2869) );
  IV U1702 ( .A(n2995), .Z(n712) );
  MUX U1703 ( .IN0(n713), .IN1(n3083), .SEL(n3084), .F(n2951) );
  IV U1704 ( .A(n3085), .Z(n713) );
  MUX U1705 ( .IN0(n714), .IN1(n3067), .SEL(n3068), .F(n2935) );
  IV U1706 ( .A(n3069), .Z(n714) );
  XNOR U1707 ( .A(n3231), .B(n3230), .Z(n3362) );
  XNOR U1708 ( .A(n3223), .B(n3222), .Z(n3354) );
  XNOR U1709 ( .A(n3184), .B(n3183), .Z(n3315) );
  XNOR U1710 ( .A(n3207), .B(n3206), .Z(n3338) );
  XNOR U1711 ( .A(n3131), .B(n3130), .Z(n3260) );
  XNOR U1712 ( .A(n3139), .B(n3138), .Z(n3268) );
  MUX U1713 ( .IN0(n3310), .IN1(n4697), .SEL(n3312), .F(n3174) );
  XNOR U1714 ( .A(n3155), .B(n3154), .Z(n3284) );
  MUX U1715 ( .IN0(X[30]), .IN1(n715), .SEL(X[31]), .F(n908) );
  IV U1716 ( .A(n5598), .Z(n715) );
  XNOR U1717 ( .A(n1051), .B(n1055), .Z(n1091) );
  NAND U1718 ( .A(n1256), .B(n1255), .Z(n1250) );
  MUX U1719 ( .IN0(n1259), .IN1(n1261), .SEL(n1260), .F(n1189) );
  XNOR U1720 ( .A(n1104), .B(n1103), .Z(n1158) );
  NAND U1721 ( .A(n1407), .B(n1408), .Z(n1402) );
  MUX U1722 ( .IN0(n716), .IN1(n1823), .SEL(n1824), .F(n1723) );
  IV U1723 ( .A(n1825), .Z(n716) );
  MUX U1724 ( .IN0(n717), .IN1(n4188), .SEL(X[31]), .F(n1796) );
  IV U1725 ( .A(X[15]), .Z(n717) );
  AND U1726 ( .A(n1877), .B(n1879), .Z(n1780) );
  ANDN U1727 ( .A(n2318), .B(n2319), .Z(n2210) );
  MUX U1728 ( .IN0(n3329), .IN1(n3327), .SEL(n3328), .F(n718) );
  IV U1729 ( .A(n718), .Z(n3191) );
  MUX U1730 ( .IN0(n719), .IN1(n3296), .SEL(n3297), .F(n3162) );
  IV U1731 ( .A(n3298), .Z(n719) );
  MUX U1732 ( .IN0(n903), .IN1(n901), .SEL(n902), .F(n881) );
  ANDN U1733 ( .A(n913), .B(n914), .Z(n884) );
  MUX U1734 ( .IN0(n720), .IN1(n1136), .SEL(n1137), .F(n1113) );
  IV U1735 ( .A(n1138), .Z(n720) );
  XNOR U1736 ( .A(n1798), .B(n1797), .Z(n1791) );
  XNOR U1737 ( .A(n2664), .B(n2659), .Z(n2773) );
  MUX U1738 ( .IN0(n878), .IN1(n880), .SEL(n879), .F(n721) );
  IV U1739 ( .A(n721), .Z(n863) );
  XNOR U1740 ( .A(n947), .B(n952), .Z(n948) );
  XNOR U1741 ( .A(n1072), .B(n1077), .Z(n1073) );
  XNOR U1742 ( .A(n1238), .B(n1243), .Z(n1239) );
  XOR U1743 ( .A(n1401), .B(n1400), .Z(n1382) );
  XOR U1744 ( .A(n1634), .B(n1633), .Z(n1616) );
  XOR U1745 ( .A(n1900), .B(n1899), .Z(n1979) );
  XOR U1746 ( .A(n2101), .B(n2100), .Z(n2176) );
  XOR U1747 ( .A(n2209), .B(n2208), .Z(n2282) );
  XOR U1748 ( .A(n2424), .B(n2423), .Z(n2497) );
  XOR U1749 ( .A(n2538), .B(n2537), .Z(n2616) );
  XOR U1750 ( .A(n2772), .B(n2771), .Z(n2858) );
  XOR U1751 ( .A(n2894), .B(n2893), .Z(n2982) );
  XOR U1752 ( .A(n3018), .B(n3017), .Z(n3112) );
  AND U1753 ( .A(Y0[0]), .B(n3116), .Z(n3241) );
  XNOR U1754 ( .A(n889), .B(n893), .Z(n891) );
  XNOR U1755 ( .A(n990), .B(n994), .Z(n992) );
  XNOR U1756 ( .A(n1118), .B(n1121), .Z(n1120) );
  XNOR U1757 ( .A(n1308), .B(n1312), .Z(n1310) );
  XNOR U1758 ( .A(n1527), .B(n1531), .Z(n1529) );
  XNOR U1759 ( .A(n1783), .B(n1787), .Z(n1785) );
  XNOR U1760 ( .A(n2072), .B(n2076), .Z(n2074) );
  XNOR U1761 ( .A(n2386), .B(n2390), .Z(n2388) );
  XNOR U1762 ( .A(n2733), .B(n2737), .Z(n2735) );
  MUX U1763 ( .IN0(n722), .IN1(n824), .SEL(n830), .F(n827) );
  ANDN U1764 ( .A(n723), .B(n[0]), .Z(n357) );
  AND U1765 ( .A(N8), .B(n723), .Z(n356) );
  AND U1766 ( .A(N9), .B(n723), .Z(n355) );
  AND U1767 ( .A(N10), .B(n723), .Z(n354) );
  AND U1768 ( .A(N11), .B(n723), .Z(n353) );
  AND U1769 ( .A(N12), .B(n723), .Z(n352) );
  AND U1770 ( .A(n723), .B(n724), .Z(n351) );
  XOR U1771 ( .A(n[6]), .B(\add_25/carry[6] ), .Z(n724) );
  ANDN U1772 ( .A(n725), .B(rst), .Z(n723) );
  NAND U1773 ( .A(n726), .B(n727), .Z(n725) );
  AND U1774 ( .A(n728), .B(n[0]), .Z(n727) );
  ANDN U1775 ( .A(n729), .B(n[2]), .Z(n728) );
  AND U1776 ( .A(n[6]), .B(n730), .Z(n726) );
  AND U1777 ( .A(n[5]), .B(n[1]), .Z(n730) );
  NAND U1778 ( .A(n731), .B(n732), .Z(n350) );
  NAND U1779 ( .A(n733), .B(n734), .Z(n732) );
  NAND U1780 ( .A(Y0[0]), .B(rst), .Z(n731) );
  NAND U1781 ( .A(n735), .B(n736), .Z(n349) );
  NAND U1782 ( .A(n737), .B(n734), .Z(n736) );
  NAND U1783 ( .A(Y0[1]), .B(rst), .Z(n735) );
  NAND U1784 ( .A(n738), .B(n739), .Z(n348) );
  NAND U1785 ( .A(n740), .B(n734), .Z(n739) );
  NAND U1786 ( .A(Y0[2]), .B(rst), .Z(n738) );
  NAND U1787 ( .A(n741), .B(n742), .Z(n347) );
  NAND U1788 ( .A(n743), .B(n734), .Z(n742) );
  NAND U1789 ( .A(Y0[3]), .B(rst), .Z(n741) );
  NAND U1790 ( .A(n744), .B(n745), .Z(n346) );
  NAND U1791 ( .A(n746), .B(n734), .Z(n745) );
  NAND U1792 ( .A(Y0[4]), .B(rst), .Z(n744) );
  NAND U1793 ( .A(n747), .B(n748), .Z(n345) );
  NAND U1794 ( .A(n749), .B(n734), .Z(n748) );
  NAND U1795 ( .A(rst), .B(Y0[5]), .Z(n747) );
  NAND U1796 ( .A(n750), .B(n751), .Z(n344) );
  NAND U1797 ( .A(n752), .B(n734), .Z(n751) );
  NAND U1798 ( .A(rst), .B(Y0[6]), .Z(n750) );
  NAND U1799 ( .A(n753), .B(n754), .Z(n343) );
  NAND U1800 ( .A(n755), .B(n734), .Z(n754) );
  NAND U1801 ( .A(rst), .B(Y0[7]), .Z(n753) );
  NAND U1802 ( .A(n756), .B(n757), .Z(n342) );
  NAND U1803 ( .A(n758), .B(n734), .Z(n757) );
  NAND U1804 ( .A(rst), .B(Y0[8]), .Z(n756) );
  NAND U1805 ( .A(n759), .B(n760), .Z(n341) );
  NAND U1806 ( .A(n761), .B(n734), .Z(n760) );
  NAND U1807 ( .A(rst), .B(Y0[9]), .Z(n759) );
  NAND U1808 ( .A(n762), .B(n763), .Z(n340) );
  NAND U1809 ( .A(n764), .B(n734), .Z(n763) );
  NAND U1810 ( .A(rst), .B(Y0[10]), .Z(n762) );
  NAND U1811 ( .A(n765), .B(n766), .Z(n339) );
  NAND U1812 ( .A(n767), .B(n734), .Z(n766) );
  NAND U1813 ( .A(rst), .B(Y0[11]), .Z(n765) );
  NAND U1814 ( .A(n768), .B(n769), .Z(n338) );
  NAND U1815 ( .A(n770), .B(n734), .Z(n769) );
  NAND U1816 ( .A(rst), .B(Y0[12]), .Z(n768) );
  NAND U1817 ( .A(n771), .B(n772), .Z(n337) );
  NAND U1818 ( .A(n773), .B(n734), .Z(n772) );
  NAND U1819 ( .A(rst), .B(Y0[13]), .Z(n771) );
  NAND U1820 ( .A(n774), .B(n775), .Z(n336) );
  NAND U1821 ( .A(n776), .B(n734), .Z(n775) );
  NAND U1822 ( .A(rst), .B(Y0[14]), .Z(n774) );
  NAND U1823 ( .A(n777), .B(n778), .Z(n335) );
  NAND U1824 ( .A(n779), .B(n734), .Z(n778) );
  NAND U1825 ( .A(rst), .B(Y0[15]), .Z(n777) );
  NAND U1826 ( .A(n780), .B(n781), .Z(n334) );
  NAND U1827 ( .A(n782), .B(n734), .Z(n781) );
  NAND U1828 ( .A(rst), .B(Y0[16]), .Z(n780) );
  NAND U1829 ( .A(n783), .B(n784), .Z(n333) );
  NAND U1830 ( .A(n785), .B(n734), .Z(n784) );
  NAND U1831 ( .A(rst), .B(Y0[17]), .Z(n783) );
  NAND U1832 ( .A(n786), .B(n787), .Z(n332) );
  NAND U1833 ( .A(n788), .B(n734), .Z(n787) );
  NAND U1834 ( .A(rst), .B(Y0[18]), .Z(n786) );
  NAND U1835 ( .A(n789), .B(n790), .Z(n331) );
  NAND U1836 ( .A(n791), .B(n734), .Z(n790) );
  NAND U1837 ( .A(rst), .B(Y0[19]), .Z(n789) );
  NAND U1838 ( .A(n792), .B(n793), .Z(n330) );
  NAND U1839 ( .A(n794), .B(n734), .Z(n793) );
  NAND U1840 ( .A(rst), .B(Y0[20]), .Z(n792) );
  NAND U1841 ( .A(n795), .B(n796), .Z(n329) );
  NAND U1842 ( .A(n797), .B(n734), .Z(n796) );
  NAND U1843 ( .A(rst), .B(Y0[21]), .Z(n795) );
  NAND U1844 ( .A(n798), .B(n799), .Z(n328) );
  NAND U1845 ( .A(n800), .B(n734), .Z(n799) );
  NAND U1846 ( .A(rst), .B(Y0[22]), .Z(n798) );
  NAND U1847 ( .A(n801), .B(n802), .Z(n327) );
  NAND U1848 ( .A(n803), .B(n734), .Z(n802) );
  NAND U1849 ( .A(rst), .B(Y0[23]), .Z(n801) );
  NAND U1850 ( .A(n804), .B(n805), .Z(n326) );
  NAND U1851 ( .A(n806), .B(n734), .Z(n805) );
  NAND U1852 ( .A(rst), .B(Y0[24]), .Z(n804) );
  NAND U1853 ( .A(n807), .B(n808), .Z(n325) );
  NAND U1854 ( .A(n809), .B(n734), .Z(n808) );
  NAND U1855 ( .A(rst), .B(Y0[25]), .Z(n807) );
  NAND U1856 ( .A(n810), .B(n811), .Z(n324) );
  NAND U1857 ( .A(n812), .B(n734), .Z(n811) );
  NAND U1858 ( .A(rst), .B(Y0[26]), .Z(n810) );
  NAND U1859 ( .A(n813), .B(n814), .Z(n323) );
  NAND U1860 ( .A(n815), .B(n734), .Z(n814) );
  NAND U1861 ( .A(rst), .B(Y0[27]), .Z(n813) );
  NAND U1862 ( .A(n816), .B(n817), .Z(n322) );
  NAND U1863 ( .A(n818), .B(n734), .Z(n817) );
  NAND U1864 ( .A(rst), .B(Y0[28]), .Z(n816) );
  NAND U1865 ( .A(n819), .B(n820), .Z(n321) );
  NAND U1866 ( .A(n821), .B(n734), .Z(n820) );
  NAND U1867 ( .A(rst), .B(Y0[29]), .Z(n819) );
  NAND U1868 ( .A(n822), .B(n823), .Z(n320) );
  NAND U1869 ( .A(n824), .B(n734), .Z(n823) );
  NAND U1870 ( .A(rst), .B(Y0[30]), .Z(n822) );
  NAND U1871 ( .A(n825), .B(n826), .Z(n319) );
  NAND U1872 ( .A(n827), .B(n734), .Z(n826) );
  NOR U1873 ( .A(rst), .B(n828), .Z(n734) );
  NAND U1874 ( .A(Y0[31]), .B(rst), .Z(n825) );
  MUX U1875 ( .IN0(Y[31]), .IN1(n827), .SEL(n829), .F(n318) );
  XNOR U1876 ( .A(Y0[31]), .B(n831), .Z(n830) );
  AND U1877 ( .A(n834), .B(n835), .Z(n833) );
  XNOR U1878 ( .A(Y0[31]), .B(n836), .Z(n835) );
  MUX U1879 ( .IN0(Y[30]), .IN1(n824), .SEL(n829), .F(n317) );
  XOR U1880 ( .A(n834), .B(Y0[31]), .Z(n824) );
  XOR U1881 ( .A(n836), .B(n831), .Z(n834) );
  XOR U1882 ( .A(n837), .B(n838), .Z(n831) );
  XOR U1883 ( .A(n839), .B(n840), .Z(n838) );
  AND U1884 ( .A(n841), .B(n842), .Z(n840) );
  XOR U1885 ( .A(n849), .B(n847), .Z(n837) );
  XOR U1886 ( .A(n850), .B(n851), .Z(n849) );
  XOR U1887 ( .A(n852), .B(n853), .Z(n851) );
  XOR U1888 ( .A(n857), .B(n858), .Z(n852) );
  ANDN U1889 ( .A(n859), .B(n860), .Z(n858) );
  XOR U1890 ( .A(n864), .B(n865), .Z(n850) );
  XOR U1891 ( .A(n854), .B(n856), .Z(n865) );
  XOR U1892 ( .A(n863), .B(n860), .Z(n864) );
  IV U1893 ( .A(n832), .Z(n836) );
  MUX U1894 ( .IN0(Y[29]), .IN1(n821), .SEL(n829), .F(n316) );
  XOR U1895 ( .A(n867), .B(Y0[30]), .Z(n821) );
  XNOR U1896 ( .A(n868), .B(n869), .Z(n867) );
  AND U1897 ( .A(n841), .B(n871), .Z(n870) );
  XNOR U1898 ( .A(n845), .B(n869), .Z(n871) );
  XOR U1899 ( .A(n843), .B(n869), .Z(n845) );
  XNOR U1900 ( .A(n848), .B(n846), .Z(n869) );
  IV U1901 ( .A(n847), .Z(n846) );
  XNOR U1902 ( .A(n854), .B(n855), .Z(n848) );
  XNOR U1903 ( .A(n856), .B(n859), .Z(n855) );
  XNOR U1904 ( .A(n860), .B(n875), .Z(n859) );
  XOR U1905 ( .A(n861), .B(n862), .Z(n875) );
  NAND U1906 ( .A(n876), .B(n877), .Z(n862) );
  IV U1907 ( .A(n863), .Z(n861) );
  IV U1908 ( .A(n844), .Z(n843) );
  MUX U1909 ( .IN0(Y[28]), .IN1(n818), .SEL(n829), .F(n315) );
  XOR U1910 ( .A(n890), .B(Y0[29]), .Z(n818) );
  XNOR U1911 ( .A(n891), .B(n892), .Z(n890) );
  AND U1912 ( .A(n841), .B(n894), .Z(n893) );
  XNOR U1913 ( .A(n888), .B(n892), .Z(n894) );
  XNOR U1914 ( .A(n874), .B(n873), .Z(n892) );
  IV U1915 ( .A(n872), .Z(n873) );
  XOR U1916 ( .A(n886), .B(n885), .Z(n874) );
  XOR U1917 ( .A(n884), .B(n898), .Z(n885) );
  XNOR U1918 ( .A(n883), .B(n882), .Z(n898) );
  XNOR U1919 ( .A(n899), .B(n900), .Z(n882) );
  IV U1920 ( .A(n881), .Z(n900) );
  XNOR U1921 ( .A(n879), .B(n880), .Z(n883) );
  NAND U1922 ( .A(n906), .B(n877), .Z(n880) );
  XNOR U1923 ( .A(n878), .B(n907), .Z(n879) );
  ANDN U1924 ( .A(n908), .B(n909), .Z(n907) );
  MUX U1925 ( .IN0(Y[27]), .IN1(n815), .SEL(n829), .F(n314) );
  XOR U1926 ( .A(n919), .B(Y0[28]), .Z(n815) );
  XNOR U1927 ( .A(n920), .B(n921), .Z(n919) );
  AND U1928 ( .A(n841), .B(n923), .Z(n922) );
  XNOR U1929 ( .A(n917), .B(n921), .Z(n923) );
  XNOR U1930 ( .A(n897), .B(n896), .Z(n921) );
  IV U1931 ( .A(n895), .Z(n896) );
  XOR U1932 ( .A(n915), .B(n914), .Z(n897) );
  XOR U1933 ( .A(n913), .B(n927), .Z(n914) );
  XNOR U1934 ( .A(n903), .B(n902), .Z(n927) );
  XOR U1935 ( .A(n932), .B(n904), .Z(n928) );
  AND U1936 ( .A(n933), .B(n876), .Z(n904) );
  IV U1937 ( .A(n901), .Z(n932) );
  XNOR U1938 ( .A(n911), .B(n912), .Z(n903) );
  NAND U1939 ( .A(n937), .B(n877), .Z(n912) );
  XNOR U1940 ( .A(n910), .B(n938), .Z(n911) );
  ANDN U1941 ( .A(n908), .B(n939), .Z(n938) );
  MUX U1942 ( .IN0(Y[26]), .IN1(n812), .SEL(n829), .F(n313) );
  XOR U1943 ( .A(n950), .B(Y0[27]), .Z(n812) );
  XNOR U1944 ( .A(n951), .B(n952), .Z(n950) );
  AND U1945 ( .A(n841), .B(n954), .Z(n953) );
  XNOR U1946 ( .A(n948), .B(n952), .Z(n954) );
  XNOR U1947 ( .A(n926), .B(n925), .Z(n952) );
  IV U1948 ( .A(n924), .Z(n925) );
  XNOR U1949 ( .A(n946), .B(n958), .Z(n926) );
  XOR U1950 ( .A(n945), .B(n944), .Z(n958) );
  XOR U1951 ( .A(n959), .B(n960), .Z(n944) );
  XOR U1952 ( .A(n961), .B(n962), .Z(n960) );
  XOR U1953 ( .A(n963), .B(n964), .Z(n962) );
  XNOR U1954 ( .A(n936), .B(n935), .Z(n945) );
  XOR U1955 ( .A(n972), .B(n930), .Z(n935) );
  XNOR U1956 ( .A(n929), .B(n973), .Z(n930) );
  ANDN U1957 ( .A(n974), .B(n909), .Z(n973) );
  AND U1958 ( .A(n906), .B(n933), .Z(n931) );
  XNOR U1959 ( .A(n941), .B(n942), .Z(n936) );
  NAND U1960 ( .A(n981), .B(n877), .Z(n942) );
  XNOR U1961 ( .A(n940), .B(n982), .Z(n941) );
  ANDN U1962 ( .A(n908), .B(n983), .Z(n982) );
  MUX U1963 ( .IN0(Y[25]), .IN1(n809), .SEL(n829), .F(n312) );
  XOR U1964 ( .A(n991), .B(Y0[26]), .Z(n809) );
  XNOR U1965 ( .A(n992), .B(n993), .Z(n991) );
  AND U1966 ( .A(n841), .B(n995), .Z(n994) );
  XNOR U1967 ( .A(n989), .B(n993), .Z(n995) );
  XNOR U1968 ( .A(n957), .B(n956), .Z(n993) );
  IV U1969 ( .A(n955), .Z(n956) );
  XOR U1970 ( .A(n987), .B(n999), .Z(n957) );
  XNOR U1971 ( .A(n971), .B(n970), .Z(n999) );
  XOR U1972 ( .A(n1000), .B(n965), .Z(n970) );
  XOR U1973 ( .A(n966), .B(n967), .Z(n965) );
  NANDN U1974 ( .B(n1001), .A(n876), .Z(n967) );
  IV U1975 ( .A(n968), .Z(n966) );
  XOR U1976 ( .A(n961), .B(n969), .Z(n1000) );
  XNOR U1977 ( .A(n980), .B(n979), .Z(n971) );
  XOR U1978 ( .A(n1011), .B(n976), .Z(n979) );
  XNOR U1979 ( .A(n975), .B(n1012), .Z(n976) );
  ANDN U1980 ( .A(n974), .B(n939), .Z(n1012) );
  XOR U1981 ( .A(n1013), .B(n1014), .Z(n975) );
  AND U1982 ( .A(n1015), .B(n1016), .Z(n1014) );
  XNOR U1983 ( .A(n1017), .B(n1013), .Z(n1016) );
  AND U1984 ( .A(n937), .B(n933), .Z(n977) );
  XNOR U1985 ( .A(n985), .B(n986), .Z(n980) );
  NAND U1986 ( .A(n1021), .B(n877), .Z(n986) );
  XNOR U1987 ( .A(n984), .B(n1022), .Z(n985) );
  ANDN U1988 ( .A(n908), .B(n1023), .Z(n1022) );
  MUX U1989 ( .IN0(Y[24]), .IN1(n806), .SEL(n829), .F(n311) );
  XOR U1990 ( .A(n1031), .B(Y0[25]), .Z(n806) );
  XNOR U1991 ( .A(n1032), .B(n1033), .Z(n1031) );
  AND U1992 ( .A(n841), .B(n1035), .Z(n1034) );
  XNOR U1993 ( .A(n1029), .B(n1033), .Z(n1035) );
  XNOR U1994 ( .A(n998), .B(n997), .Z(n1033) );
  IV U1995 ( .A(n996), .Z(n997) );
  XOR U1996 ( .A(n1027), .B(n1039), .Z(n998) );
  XNOR U1997 ( .A(n1007), .B(n1006), .Z(n1039) );
  XOR U1998 ( .A(n1040), .B(n1010), .Z(n1006) );
  XNOR U1999 ( .A(n1003), .B(n1004), .Z(n1010) );
  NANDN U2000 ( .B(n1001), .A(n906), .Z(n1004) );
  XNOR U2001 ( .A(n1002), .B(n1041), .Z(n1003) );
  ANDN U2002 ( .A(n1042), .B(n909), .Z(n1041) );
  XNOR U2003 ( .A(n1009), .B(n1005), .Z(n1040) );
  XNOR U2004 ( .A(n1049), .B(n1050), .Z(n1009) );
  IV U2005 ( .A(n1008), .Z(n1050) );
  XNOR U2006 ( .A(n1020), .B(n1019), .Z(n1007) );
  XOR U2007 ( .A(n1057), .B(n1015), .Z(n1019) );
  XNOR U2008 ( .A(n1013), .B(n1058), .Z(n1015) );
  ANDN U2009 ( .A(n974), .B(n983), .Z(n1058) );
  AND U2010 ( .A(n981), .B(n933), .Z(n1017) );
  XNOR U2011 ( .A(n1025), .B(n1026), .Z(n1020) );
  NAND U2012 ( .A(n1065), .B(n877), .Z(n1026) );
  XNOR U2013 ( .A(n1024), .B(n1066), .Z(n1025) );
  ANDN U2014 ( .A(n908), .B(n1067), .Z(n1066) );
  MUX U2015 ( .IN0(Y[23]), .IN1(n803), .SEL(n829), .F(n310) );
  XOR U2016 ( .A(n1075), .B(Y0[24]), .Z(n803) );
  XNOR U2017 ( .A(n1076), .B(n1077), .Z(n1075) );
  AND U2018 ( .A(n841), .B(n1079), .Z(n1078) );
  XNOR U2019 ( .A(n1073), .B(n1077), .Z(n1079) );
  XNOR U2020 ( .A(n1038), .B(n1037), .Z(n1077) );
  IV U2021 ( .A(n1036), .Z(n1037) );
  XOR U2022 ( .A(n1071), .B(n1082), .Z(n1038) );
  XNOR U2023 ( .A(n1048), .B(n1047), .Z(n1082) );
  XOR U2024 ( .A(n1083), .B(n1053), .Z(n1047) );
  XNOR U2025 ( .A(n1044), .B(n1045), .Z(n1053) );
  NANDN U2026 ( .B(n1001), .A(n937), .Z(n1045) );
  XNOR U2027 ( .A(n1043), .B(n1084), .Z(n1044) );
  ANDN U2028 ( .A(n1042), .B(n939), .Z(n1084) );
  XNOR U2029 ( .A(n1052), .B(n1046), .Z(n1083) );
  XNOR U2030 ( .A(n1091), .B(n1054), .Z(n1052) );
  IV U2031 ( .A(n1056), .Z(n1054) );
  AND U2032 ( .A(n1095), .B(n876), .Z(n1055) );
  XNOR U2033 ( .A(n1064), .B(n1063), .Z(n1048) );
  XOR U2034 ( .A(n1099), .B(n1060), .Z(n1063) );
  XNOR U2035 ( .A(n1059), .B(n1100), .Z(n1060) );
  ANDN U2036 ( .A(n974), .B(n1023), .Z(n1100) );
  AND U2037 ( .A(n1021), .B(n933), .Z(n1061) );
  XNOR U2038 ( .A(n1069), .B(n1070), .Z(n1064) );
  NAND U2039 ( .A(n1107), .B(n877), .Z(n1070) );
  XNOR U2040 ( .A(n1068), .B(n1108), .Z(n1069) );
  ANDN U2041 ( .A(n908), .B(n1109), .Z(n1108) );
  MUX U2042 ( .IN0(Y[22]), .IN1(n800), .SEL(n829), .F(n309) );
  XOR U2043 ( .A(n1119), .B(Y0[23]), .Z(n800) );
  XNOR U2044 ( .A(n1120), .B(n1081), .Z(n1119) );
  AND U2045 ( .A(n841), .B(n1122), .Z(n1121) );
  XNOR U2046 ( .A(n1117), .B(n1081), .Z(n1122) );
  XOR U2047 ( .A(n1080), .B(n1123), .Z(n1081) );
  XNOR U2048 ( .A(n1115), .B(n1114), .Z(n1123) );
  XOR U2049 ( .A(n1124), .B(n1125), .Z(n1114) );
  XOR U2050 ( .A(n1126), .B(n1127), .Z(n1125) );
  XOR U2051 ( .A(n1130), .B(n1131), .Z(n1126) );
  ANDN U2052 ( .A(n1129), .B(n1132), .Z(n1131) );
  XNOR U2053 ( .A(n1135), .B(n1113), .Z(n1124) );
  XOR U2054 ( .A(n1134), .B(n1132), .Z(n1135) );
  XNOR U2055 ( .A(n1090), .B(n1089), .Z(n1115) );
  XOR U2056 ( .A(n1139), .B(n1098), .Z(n1089) );
  XNOR U2057 ( .A(n1086), .B(n1087), .Z(n1098) );
  NANDN U2058 ( .B(n1001), .A(n981), .Z(n1087) );
  XNOR U2059 ( .A(n1085), .B(n1140), .Z(n1086) );
  ANDN U2060 ( .A(n1042), .B(n983), .Z(n1140) );
  XNOR U2061 ( .A(n1097), .B(n1088), .Z(n1139) );
  XOR U2062 ( .A(n1147), .B(n1093), .Z(n1097) );
  XNOR U2063 ( .A(n1092), .B(n1148), .Z(n1093) );
  ANDN U2064 ( .A(n1149), .B(n909), .Z(n1148) );
  XOR U2065 ( .A(n1150), .B(n1151), .Z(n1092) );
  AND U2066 ( .A(n1152), .B(n1153), .Z(n1151) );
  XNOR U2067 ( .A(n1154), .B(n1150), .Z(n1153) );
  AND U2068 ( .A(n906), .B(n1095), .Z(n1094) );
  XNOR U2069 ( .A(n1106), .B(n1105), .Z(n1090) );
  XOR U2070 ( .A(n1158), .B(n1102), .Z(n1105) );
  XNOR U2071 ( .A(n1101), .B(n1159), .Z(n1102) );
  ANDN U2072 ( .A(n974), .B(n1067), .Z(n1159) );
  AND U2073 ( .A(n1065), .B(n933), .Z(n1103) );
  XNOR U2074 ( .A(n1111), .B(n1112), .Z(n1106) );
  NAND U2075 ( .A(n1166), .B(n877), .Z(n1112) );
  XNOR U2076 ( .A(n1110), .B(n1167), .Z(n1111) );
  ANDN U2077 ( .A(n908), .B(n1168), .Z(n1167) );
  MUX U2078 ( .IN0(Y[21]), .IN1(n797), .SEL(n829), .F(n308) );
  XOR U2079 ( .A(n1178), .B(Y0[22]), .Z(n797) );
  XNOR U2080 ( .A(n1179), .B(n1180), .Z(n1178) );
  AND U2081 ( .A(n841), .B(n1182), .Z(n1181) );
  XNOR U2082 ( .A(n1176), .B(n1180), .Z(n1182) );
  XNOR U2083 ( .A(n1174), .B(n1173), .Z(n1180) );
  IV U2084 ( .A(n1172), .Z(n1173) );
  XNOR U2085 ( .A(n1138), .B(n1137), .Z(n1174) );
  XOR U2086 ( .A(n1186), .B(n1129), .Z(n1137) );
  XNOR U2087 ( .A(n1132), .B(n1187), .Z(n1129) );
  NANDN U2088 ( .B(n1188), .A(n876), .Z(n1133) );
  XOR U2089 ( .A(n1128), .B(n1136), .Z(n1186) );
  XNOR U2090 ( .A(n1146), .B(n1145), .Z(n1138) );
  XOR U2091 ( .A(n1200), .B(n1157), .Z(n1145) );
  XNOR U2092 ( .A(n1142), .B(n1143), .Z(n1157) );
  NANDN U2093 ( .B(n1001), .A(n1021), .Z(n1143) );
  XNOR U2094 ( .A(n1141), .B(n1201), .Z(n1142) );
  ANDN U2095 ( .A(n1042), .B(n1023), .Z(n1201) );
  XOR U2096 ( .A(n1202), .B(n1203), .Z(n1141) );
  AND U2097 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U2098 ( .A(n1206), .B(n1202), .Z(n1205) );
  XNOR U2099 ( .A(n1156), .B(n1144), .Z(n1200) );
  XOR U2100 ( .A(n1210), .B(n1152), .Z(n1156) );
  XNOR U2101 ( .A(n1150), .B(n1211), .Z(n1152) );
  ANDN U2102 ( .A(n1149), .B(n939), .Z(n1211) );
  XOR U2103 ( .A(n1212), .B(n1213), .Z(n1150) );
  AND U2104 ( .A(n1214), .B(n1215), .Z(n1213) );
  XNOR U2105 ( .A(n1216), .B(n1212), .Z(n1215) );
  AND U2106 ( .A(n937), .B(n1095), .Z(n1154) );
  XNOR U2107 ( .A(n1165), .B(n1164), .Z(n1146) );
  XOR U2108 ( .A(n1220), .B(n1161), .Z(n1164) );
  XNOR U2109 ( .A(n1160), .B(n1221), .Z(n1161) );
  ANDN U2110 ( .A(n974), .B(n1109), .Z(n1221) );
  XOR U2111 ( .A(n1222), .B(n1223), .Z(n1160) );
  AND U2112 ( .A(n1224), .B(n1225), .Z(n1223) );
  XNOR U2113 ( .A(n1226), .B(n1222), .Z(n1225) );
  AND U2114 ( .A(n1107), .B(n933), .Z(n1162) );
  XNOR U2115 ( .A(n1170), .B(n1171), .Z(n1165) );
  NAND U2116 ( .A(n1230), .B(n877), .Z(n1171) );
  XNOR U2117 ( .A(n1169), .B(n1231), .Z(n1170) );
  ANDN U2118 ( .A(n908), .B(n1232), .Z(n1231) );
  XOR U2119 ( .A(n1233), .B(n1234), .Z(n1169) );
  AND U2120 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U2121 ( .A(n1237), .B(n1233), .Z(n1236) );
  MUX U2122 ( .IN0(Y[20]), .IN1(n794), .SEL(n829), .F(n307) );
  XOR U2123 ( .A(n1241), .B(Y0[21]), .Z(n794) );
  XNOR U2124 ( .A(n1242), .B(n1243), .Z(n1241) );
  AND U2125 ( .A(n841), .B(n1245), .Z(n1244) );
  XNOR U2126 ( .A(n1239), .B(n1243), .Z(n1245) );
  XNOR U2127 ( .A(n1185), .B(n1184), .Z(n1243) );
  IV U2128 ( .A(n1183), .Z(n1184) );
  XNOR U2129 ( .A(n1197), .B(n1196), .Z(n1185) );
  XOR U2130 ( .A(n1249), .B(n1199), .Z(n1196) );
  XNOR U2131 ( .A(n1194), .B(n1193), .Z(n1199) );
  XNOR U2132 ( .A(n1250), .B(n1251), .Z(n1193) );
  IV U2133 ( .A(n1192), .Z(n1251) );
  XNOR U2134 ( .A(n1190), .B(n1191), .Z(n1194) );
  NANDN U2135 ( .B(n1188), .A(n906), .Z(n1191) );
  XNOR U2136 ( .A(n1189), .B(n1257), .Z(n1190) );
  ANDN U2137 ( .A(n1258), .B(n909), .Z(n1257) );
  XNOR U2138 ( .A(n1209), .B(n1208), .Z(n1197) );
  XOR U2139 ( .A(n1268), .B(n1219), .Z(n1208) );
  XNOR U2140 ( .A(n1204), .B(n1206), .Z(n1219) );
  NANDN U2141 ( .B(n1001), .A(n1065), .Z(n1206) );
  XNOR U2142 ( .A(n1202), .B(n1269), .Z(n1204) );
  ANDN U2143 ( .A(n1042), .B(n1067), .Z(n1269) );
  XOR U2144 ( .A(n1270), .B(n1271), .Z(n1202) );
  AND U2145 ( .A(n1272), .B(n1273), .Z(n1271) );
  XOR U2146 ( .A(n1274), .B(n1270), .Z(n1273) );
  XNOR U2147 ( .A(n1218), .B(n1207), .Z(n1268) );
  XOR U2148 ( .A(n1278), .B(n1214), .Z(n1218) );
  XNOR U2149 ( .A(n1212), .B(n1279), .Z(n1214) );
  ANDN U2150 ( .A(n1149), .B(n983), .Z(n1279) );
  XOR U2151 ( .A(n1280), .B(n1281), .Z(n1212) );
  AND U2152 ( .A(n1282), .B(n1283), .Z(n1281) );
  XNOR U2153 ( .A(n1284), .B(n1280), .Z(n1283) );
  AND U2154 ( .A(n981), .B(n1095), .Z(n1216) );
  XNOR U2155 ( .A(n1229), .B(n1228), .Z(n1209) );
  XOR U2156 ( .A(n1288), .B(n1224), .Z(n1228) );
  XNOR U2157 ( .A(n1222), .B(n1289), .Z(n1224) );
  ANDN U2158 ( .A(n974), .B(n1168), .Z(n1289) );
  XOR U2159 ( .A(n1290), .B(n1291), .Z(n1222) );
  AND U2160 ( .A(n1292), .B(n1293), .Z(n1291) );
  XNOR U2161 ( .A(n1294), .B(n1290), .Z(n1293) );
  AND U2162 ( .A(n1166), .B(n933), .Z(n1226) );
  XNOR U2163 ( .A(n1235), .B(n1237), .Z(n1229) );
  NAND U2164 ( .A(n1298), .B(n877), .Z(n1237) );
  XNOR U2165 ( .A(n1233), .B(n1299), .Z(n1235) );
  ANDN U2166 ( .A(n908), .B(n1300), .Z(n1299) );
  XOR U2167 ( .A(n1301), .B(n1302), .Z(n1233) );
  AND U2168 ( .A(n1303), .B(n1304), .Z(n1302) );
  XOR U2169 ( .A(n1305), .B(n1301), .Z(n1304) );
  MUX U2170 ( .IN0(Y[19]), .IN1(n791), .SEL(n829), .F(n306) );
  XOR U2171 ( .A(n1309), .B(Y0[20]), .Z(n791) );
  XNOR U2172 ( .A(n1310), .B(n1311), .Z(n1309) );
  AND U2173 ( .A(n841), .B(n1313), .Z(n1312) );
  XNOR U2174 ( .A(n1307), .B(n1311), .Z(n1313) );
  XNOR U2175 ( .A(n1248), .B(n1247), .Z(n1311) );
  IV U2176 ( .A(n1246), .Z(n1247) );
  XNOR U2177 ( .A(n1264), .B(n1263), .Z(n1248) );
  XOR U2178 ( .A(n1317), .B(n1267), .Z(n1263) );
  XNOR U2179 ( .A(n1254), .B(n1253), .Z(n1267) );
  XOR U2180 ( .A(n1322), .B(n1255), .Z(n1318) );
  AND U2181 ( .A(n1323), .B(n876), .Z(n1255) );
  IV U2182 ( .A(n1252), .Z(n1322) );
  XNOR U2183 ( .A(n1260), .B(n1261), .Z(n1254) );
  NANDN U2184 ( .B(n1188), .A(n937), .Z(n1261) );
  XNOR U2185 ( .A(n1259), .B(n1327), .Z(n1260) );
  ANDN U2186 ( .A(n1258), .B(n939), .Z(n1327) );
  XNOR U2187 ( .A(n1266), .B(n1262), .Z(n1317) );
  IV U2188 ( .A(n1265), .Z(n1266) );
  XNOR U2189 ( .A(n1277), .B(n1276), .Z(n1264) );
  XOR U2190 ( .A(n1337), .B(n1287), .Z(n1276) );
  XNOR U2191 ( .A(n1272), .B(n1274), .Z(n1287) );
  NANDN U2192 ( .B(n1001), .A(n1107), .Z(n1274) );
  XNOR U2193 ( .A(n1270), .B(n1338), .Z(n1272) );
  ANDN U2194 ( .A(n1042), .B(n1109), .Z(n1338) );
  XOR U2195 ( .A(n1339), .B(n1340), .Z(n1270) );
  AND U2196 ( .A(n1341), .B(n1342), .Z(n1340) );
  XOR U2197 ( .A(n1343), .B(n1339), .Z(n1342) );
  XNOR U2198 ( .A(n1286), .B(n1275), .Z(n1337) );
  XOR U2199 ( .A(n1347), .B(n1282), .Z(n1286) );
  XNOR U2200 ( .A(n1280), .B(n1348), .Z(n1282) );
  ANDN U2201 ( .A(n1149), .B(n1023), .Z(n1348) );
  XOR U2202 ( .A(n1349), .B(n1350), .Z(n1280) );
  AND U2203 ( .A(n1351), .B(n1352), .Z(n1350) );
  XNOR U2204 ( .A(n1353), .B(n1349), .Z(n1352) );
  AND U2205 ( .A(n1021), .B(n1095), .Z(n1284) );
  XNOR U2206 ( .A(n1297), .B(n1296), .Z(n1277) );
  XOR U2207 ( .A(n1357), .B(n1292), .Z(n1296) );
  XNOR U2208 ( .A(n1290), .B(n1358), .Z(n1292) );
  ANDN U2209 ( .A(n974), .B(n1232), .Z(n1358) );
  AND U2210 ( .A(n1230), .B(n933), .Z(n1294) );
  XNOR U2211 ( .A(n1303), .B(n1305), .Z(n1297) );
  NAND U2212 ( .A(n1365), .B(n877), .Z(n1305) );
  XNOR U2213 ( .A(n1301), .B(n1366), .Z(n1303) );
  ANDN U2214 ( .A(n908), .B(n1367), .Z(n1366) );
  XOR U2215 ( .A(n1368), .B(n1369), .Z(n1301) );
  AND U2216 ( .A(n1370), .B(n1371), .Z(n1369) );
  XOR U2217 ( .A(n1372), .B(n1368), .Z(n1371) );
  MUX U2218 ( .IN0(Y[18]), .IN1(n788), .SEL(n829), .F(n305) );
  XOR U2219 ( .A(n1376), .B(Y0[19]), .Z(n788) );
  XNOR U2220 ( .A(n1377), .B(n1378), .Z(n1376) );
  AND U2221 ( .A(n841), .B(n1380), .Z(n1379) );
  XOR U2222 ( .A(n1374), .B(n1378), .Z(n1380) );
  XOR U2223 ( .A(n1373), .B(n1378), .Z(n1374) );
  XNOR U2224 ( .A(n1316), .B(n1315), .Z(n1378) );
  IV U2225 ( .A(n1314), .Z(n1315) );
  XNOR U2226 ( .A(n1333), .B(n1332), .Z(n1316) );
  XOR U2227 ( .A(n1383), .B(n1336), .Z(n1332) );
  XNOR U2228 ( .A(n1326), .B(n1325), .Z(n1336) );
  XOR U2229 ( .A(n1384), .B(n1320), .Z(n1325) );
  XNOR U2230 ( .A(n1319), .B(n1385), .Z(n1320) );
  ANDN U2231 ( .A(n1386), .B(n909), .Z(n1385) );
  XOR U2232 ( .A(n1387), .B(n1388), .Z(n1319) );
  AND U2233 ( .A(n1389), .B(n1390), .Z(n1388) );
  XNOR U2234 ( .A(n1391), .B(n1387), .Z(n1390) );
  AND U2235 ( .A(n906), .B(n1323), .Z(n1321) );
  XNOR U2236 ( .A(n1329), .B(n1330), .Z(n1326) );
  NANDN U2237 ( .B(n1188), .A(n981), .Z(n1330) );
  XNOR U2238 ( .A(n1328), .B(n1395), .Z(n1329) );
  ANDN U2239 ( .A(n1258), .B(n983), .Z(n1395) );
  XNOR U2240 ( .A(n1335), .B(n1331), .Z(n1383) );
  XNOR U2241 ( .A(n1402), .B(n1403), .Z(n1335) );
  IV U2242 ( .A(n1334), .Z(n1403) );
  XNOR U2243 ( .A(n1346), .B(n1345), .Z(n1333) );
  XOR U2244 ( .A(n1409), .B(n1356), .Z(n1345) );
  XNOR U2245 ( .A(n1341), .B(n1343), .Z(n1356) );
  NANDN U2246 ( .B(n1001), .A(n1166), .Z(n1343) );
  XNOR U2247 ( .A(n1339), .B(n1410), .Z(n1341) );
  ANDN U2248 ( .A(n1042), .B(n1168), .Z(n1410) );
  XOR U2249 ( .A(n1411), .B(n1412), .Z(n1339) );
  AND U2250 ( .A(n1413), .B(n1414), .Z(n1412) );
  XOR U2251 ( .A(n1415), .B(n1411), .Z(n1414) );
  XNOR U2252 ( .A(n1355), .B(n1344), .Z(n1409) );
  XOR U2253 ( .A(n1419), .B(n1351), .Z(n1355) );
  XNOR U2254 ( .A(n1349), .B(n1420), .Z(n1351) );
  ANDN U2255 ( .A(n1149), .B(n1067), .Z(n1420) );
  XOR U2256 ( .A(n1421), .B(n1422), .Z(n1349) );
  AND U2257 ( .A(n1423), .B(n1424), .Z(n1422) );
  XNOR U2258 ( .A(n1425), .B(n1421), .Z(n1424) );
  AND U2259 ( .A(n1065), .B(n1095), .Z(n1353) );
  XNOR U2260 ( .A(n1364), .B(n1363), .Z(n1346) );
  XOR U2261 ( .A(n1429), .B(n1360), .Z(n1363) );
  XNOR U2262 ( .A(n1359), .B(n1430), .Z(n1360) );
  ANDN U2263 ( .A(n974), .B(n1300), .Z(n1430) );
  XOR U2264 ( .A(n1431), .B(n1432), .Z(n1359) );
  AND U2265 ( .A(n1433), .B(n1434), .Z(n1432) );
  XNOR U2266 ( .A(n1435), .B(n1431), .Z(n1434) );
  AND U2267 ( .A(n1298), .B(n933), .Z(n1361) );
  XNOR U2268 ( .A(n1370), .B(n1372), .Z(n1364) );
  NAND U2269 ( .A(n1439), .B(n877), .Z(n1372) );
  XNOR U2270 ( .A(n1368), .B(n1440), .Z(n1370) );
  ANDN U2271 ( .A(n908), .B(n1441), .Z(n1440) );
  NANDN U2272 ( .B(n1442), .A(n1443), .Z(n1368) );
  NAND U2273 ( .A(n1444), .B(n1445), .Z(n1443) );
  MUX U2274 ( .IN0(Y[17]), .IN1(n785), .SEL(n829), .F(n304) );
  XOR U2275 ( .A(n1450), .B(Y0[18]), .Z(n785) );
  XOR U2276 ( .A(n1451), .B(n1452), .Z(n1450) );
  AND U2277 ( .A(n841), .B(n1454), .Z(n1453) );
  XOR U2278 ( .A(n1448), .B(n1452), .Z(n1454) );
  XOR U2279 ( .A(n1447), .B(n1452), .Z(n1448) );
  XOR U2280 ( .A(n1382), .B(n1381), .Z(n1452) );
  XNOR U2281 ( .A(n1457), .B(n1406), .Z(n1400) );
  XNOR U2282 ( .A(n1394), .B(n1393), .Z(n1406) );
  XOR U2283 ( .A(n1458), .B(n1389), .Z(n1393) );
  XNOR U2284 ( .A(n1387), .B(n1459), .Z(n1389) );
  ANDN U2285 ( .A(n1386), .B(n939), .Z(n1459) );
  XOR U2286 ( .A(n1460), .B(n1461), .Z(n1387) );
  AND U2287 ( .A(n1462), .B(n1463), .Z(n1461) );
  XNOR U2288 ( .A(n1464), .B(n1460), .Z(n1463) );
  AND U2289 ( .A(n937), .B(n1323), .Z(n1391) );
  XNOR U2290 ( .A(n1397), .B(n1398), .Z(n1394) );
  NANDN U2291 ( .B(n1188), .A(n1021), .Z(n1398) );
  XNOR U2292 ( .A(n1396), .B(n1468), .Z(n1397) );
  ANDN U2293 ( .A(n1258), .B(n1023), .Z(n1468) );
  XOR U2294 ( .A(n1469), .B(n1470), .Z(n1396) );
  AND U2295 ( .A(n1471), .B(n1472), .Z(n1470) );
  XOR U2296 ( .A(n1473), .B(n1469), .Z(n1472) );
  XNOR U2297 ( .A(n1405), .B(n1399), .Z(n1457) );
  XOR U2298 ( .A(n1477), .B(n1407), .Z(n1405) );
  NAND U2299 ( .A(n1481), .B(n1482), .Z(n1408) );
  NANDN U2300 ( .B(n1483), .A(n876), .Z(n1482) );
  NANDN U2301 ( .B(n1484), .A(n1485), .Z(n1481) );
  XNOR U2302 ( .A(n1418), .B(n1417), .Z(n1401) );
  XOR U2303 ( .A(n1489), .B(n1428), .Z(n1417) );
  XNOR U2304 ( .A(n1413), .B(n1415), .Z(n1428) );
  NANDN U2305 ( .B(n1001), .A(n1230), .Z(n1415) );
  XNOR U2306 ( .A(n1411), .B(n1490), .Z(n1413) );
  ANDN U2307 ( .A(n1042), .B(n1232), .Z(n1490) );
  XOR U2308 ( .A(n1491), .B(n1492), .Z(n1411) );
  AND U2309 ( .A(n1493), .B(n1494), .Z(n1492) );
  XOR U2310 ( .A(n1495), .B(n1491), .Z(n1494) );
  XNOR U2311 ( .A(n1427), .B(n1416), .Z(n1489) );
  XOR U2312 ( .A(n1499), .B(n1423), .Z(n1427) );
  XNOR U2313 ( .A(n1421), .B(n1500), .Z(n1423) );
  ANDN U2314 ( .A(n1149), .B(n1109), .Z(n1500) );
  XOR U2315 ( .A(n1501), .B(n1502), .Z(n1421) );
  AND U2316 ( .A(n1503), .B(n1504), .Z(n1502) );
  XNOR U2317 ( .A(n1505), .B(n1501), .Z(n1504) );
  AND U2318 ( .A(n1107), .B(n1095), .Z(n1425) );
  XOR U2319 ( .A(n1438), .B(n1437), .Z(n1418) );
  XOR U2320 ( .A(n1509), .B(n1433), .Z(n1437) );
  XNOR U2321 ( .A(n1431), .B(n1510), .Z(n1433) );
  ANDN U2322 ( .A(n974), .B(n1367), .Z(n1510) );
  AND U2323 ( .A(n1365), .B(n933), .Z(n1435) );
  XOR U2324 ( .A(n1445), .B(n1444), .Z(n1438) );
  NAND U2325 ( .A(n1517), .B(n877), .Z(n1444) );
  XNOR U2326 ( .A(n1442), .B(n1518), .Z(n1445) );
  ANDN U2327 ( .A(n908), .B(n1519), .Z(n1518) );
  NANDN U2328 ( .B(n1520), .A(n1521), .Z(n1442) );
  NAND U2329 ( .A(n1522), .B(n1523), .Z(n1521) );
  IV U2330 ( .A(n1446), .Z(n1447) );
  MUX U2331 ( .IN0(Y[16]), .IN1(n782), .SEL(n829), .F(n303) );
  XOR U2332 ( .A(n1528), .B(Y0[17]), .Z(n782) );
  XOR U2333 ( .A(n1529), .B(n1530), .Z(n1528) );
  AND U2334 ( .A(n841), .B(n1532), .Z(n1531) );
  XOR U2335 ( .A(n1526), .B(n1530), .Z(n1532) );
  XOR U2336 ( .A(n1525), .B(n1530), .Z(n1526) );
  XOR U2337 ( .A(n1456), .B(n1455), .Z(n1530) );
  XNOR U2338 ( .A(n1535), .B(n1488), .Z(n1475) );
  XNOR U2339 ( .A(n1467), .B(n1466), .Z(n1488) );
  XOR U2340 ( .A(n1536), .B(n1462), .Z(n1466) );
  XNOR U2341 ( .A(n1460), .B(n1537), .Z(n1462) );
  ANDN U2342 ( .A(n1386), .B(n983), .Z(n1537) );
  XOR U2343 ( .A(n1538), .B(n1539), .Z(n1460) );
  AND U2344 ( .A(n1540), .B(n1541), .Z(n1539) );
  XNOR U2345 ( .A(n1542), .B(n1538), .Z(n1541) );
  AND U2346 ( .A(n981), .B(n1323), .Z(n1464) );
  XNOR U2347 ( .A(n1471), .B(n1473), .Z(n1467) );
  NANDN U2348 ( .B(n1188), .A(n1065), .Z(n1473) );
  XNOR U2349 ( .A(n1469), .B(n1546), .Z(n1471) );
  ANDN U2350 ( .A(n1258), .B(n1067), .Z(n1546) );
  XOR U2351 ( .A(n1547), .B(n1548), .Z(n1469) );
  AND U2352 ( .A(n1549), .B(n1550), .Z(n1548) );
  XOR U2353 ( .A(n1551), .B(n1547), .Z(n1550) );
  XOR U2354 ( .A(n1487), .B(n1474), .Z(n1535) );
  XNOR U2355 ( .A(n1555), .B(n1479), .Z(n1487) );
  XNOR U2356 ( .A(n1556), .B(n1485), .Z(n1479) );
  AND U2357 ( .A(n906), .B(n1557), .Z(n1485) );
  NAND U2358 ( .A(n1558), .B(n1484), .Z(n1556) );
  XOR U2359 ( .A(n1559), .B(n1560), .Z(n1484) );
  AND U2360 ( .A(n1561), .B(n1562), .Z(n1560) );
  XOR U2361 ( .A(n1563), .B(n1559), .Z(n1562) );
  NANDN U2362 ( .B(n909), .A(n1564), .Z(n1558) );
  XNOR U2363 ( .A(n1478), .B(n1486), .Z(n1555) );
  IV U2364 ( .A(n1480), .Z(n1478) );
  XNOR U2365 ( .A(n1498), .B(n1497), .Z(n1476) );
  XOR U2366 ( .A(n1570), .B(n1508), .Z(n1497) );
  XNOR U2367 ( .A(n1493), .B(n1495), .Z(n1508) );
  NANDN U2368 ( .B(n1001), .A(n1298), .Z(n1495) );
  XNOR U2369 ( .A(n1491), .B(n1571), .Z(n1493) );
  ANDN U2370 ( .A(n1042), .B(n1300), .Z(n1571) );
  XNOR U2371 ( .A(n1507), .B(n1496), .Z(n1570) );
  XOR U2372 ( .A(n1578), .B(n1503), .Z(n1507) );
  XNOR U2373 ( .A(n1501), .B(n1579), .Z(n1503) );
  ANDN U2374 ( .A(n1149), .B(n1168), .Z(n1579) );
  XOR U2375 ( .A(n1580), .B(n1581), .Z(n1501) );
  AND U2376 ( .A(n1582), .B(n1583), .Z(n1581) );
  XNOR U2377 ( .A(n1584), .B(n1580), .Z(n1583) );
  AND U2378 ( .A(n1166), .B(n1095), .Z(n1505) );
  XOR U2379 ( .A(n1516), .B(n1515), .Z(n1498) );
  XOR U2380 ( .A(n1588), .B(n1512), .Z(n1515) );
  XNOR U2381 ( .A(n1511), .B(n1589), .Z(n1512) );
  ANDN U2382 ( .A(n974), .B(n1441), .Z(n1589) );
  XOR U2383 ( .A(n1590), .B(n1591), .Z(n1511) );
  AND U2384 ( .A(n1592), .B(n1593), .Z(n1591) );
  XNOR U2385 ( .A(n1594), .B(n1590), .Z(n1593) );
  AND U2386 ( .A(n1439), .B(n933), .Z(n1513) );
  XOR U2387 ( .A(n1523), .B(n1522), .Z(n1516) );
  NAND U2388 ( .A(n1598), .B(n877), .Z(n1522) );
  XNOR U2389 ( .A(n1520), .B(n1599), .Z(n1523) );
  ANDN U2390 ( .A(n908), .B(n1600), .Z(n1599) );
  NAND U2391 ( .A(n1601), .B(n1602), .Z(n1520) );
  NAND U2392 ( .A(n1603), .B(n1604), .Z(n1601) );
  IV U2393 ( .A(n1524), .Z(n1525) );
  MUX U2394 ( .IN0(Y[15]), .IN1(n779), .SEL(n829), .F(n302) );
  XOR U2395 ( .A(n1609), .B(Y0[16]), .Z(n779) );
  XOR U2396 ( .A(n1610), .B(n1611), .Z(n1609) );
  AND U2397 ( .A(n841), .B(n1613), .Z(n1612) );
  XOR U2398 ( .A(n1607), .B(n1611), .Z(n1613) );
  XOR U2399 ( .A(n1606), .B(n1611), .Z(n1607) );
  XOR U2400 ( .A(n1534), .B(n1533), .Z(n1611) );
  XNOR U2401 ( .A(n1617), .B(n1567), .Z(n1553) );
  XNOR U2402 ( .A(n1545), .B(n1544), .Z(n1567) );
  XOR U2403 ( .A(n1618), .B(n1540), .Z(n1544) );
  XNOR U2404 ( .A(n1538), .B(n1619), .Z(n1540) );
  ANDN U2405 ( .A(n1386), .B(n1023), .Z(n1619) );
  XOR U2406 ( .A(n1620), .B(n1621), .Z(n1538) );
  AND U2407 ( .A(n1622), .B(n1623), .Z(n1621) );
  XNOR U2408 ( .A(n1624), .B(n1620), .Z(n1623) );
  AND U2409 ( .A(n1021), .B(n1323), .Z(n1542) );
  XNOR U2410 ( .A(n1549), .B(n1551), .Z(n1545) );
  NANDN U2411 ( .B(n1188), .A(n1107), .Z(n1551) );
  XNOR U2412 ( .A(n1547), .B(n1628), .Z(n1549) );
  ANDN U2413 ( .A(n1258), .B(n1109), .Z(n1628) );
  XNOR U2414 ( .A(n1566), .B(n1552), .Z(n1617) );
  XOR U2415 ( .A(n1635), .B(n1569), .Z(n1566) );
  XNOR U2416 ( .A(n1561), .B(n1563), .Z(n1569) );
  NAND U2417 ( .A(n937), .B(n1557), .Z(n1563) );
  XNOR U2418 ( .A(n1559), .B(n1636), .Z(n1561) );
  ANDN U2419 ( .A(n1564), .B(n939), .Z(n1636) );
  XOR U2420 ( .A(n1637), .B(n1638), .Z(n1559) );
  AND U2421 ( .A(n1639), .B(n1640), .Z(n1638) );
  XOR U2422 ( .A(n1641), .B(n1637), .Z(n1640) );
  XNOR U2423 ( .A(n1568), .B(n1565), .Z(n1635) );
  AND U2424 ( .A(n1646), .B(n1647), .Z(n1645) );
  NANDN U2425 ( .B(n1648), .A(n876), .Z(n1647) );
  NANDN U2426 ( .B(n1649), .A(n1650), .Z(n1646) );
  XNOR U2427 ( .A(n1577), .B(n1576), .Z(n1554) );
  XOR U2428 ( .A(n1654), .B(n1587), .Z(n1576) );
  XNOR U2429 ( .A(n1573), .B(n1574), .Z(n1587) );
  NANDN U2430 ( .B(n1001), .A(n1365), .Z(n1574) );
  XNOR U2431 ( .A(n1572), .B(n1655), .Z(n1573) );
  ANDN U2432 ( .A(n1042), .B(n1367), .Z(n1655) );
  XNOR U2433 ( .A(n1586), .B(n1575), .Z(n1654) );
  XOR U2434 ( .A(n1662), .B(n1582), .Z(n1586) );
  XNOR U2435 ( .A(n1580), .B(n1663), .Z(n1582) );
  ANDN U2436 ( .A(n1149), .B(n1232), .Z(n1663) );
  XOR U2437 ( .A(n1664), .B(n1665), .Z(n1580) );
  AND U2438 ( .A(n1666), .B(n1667), .Z(n1665) );
  XNOR U2439 ( .A(n1668), .B(n1664), .Z(n1667) );
  AND U2440 ( .A(n1230), .B(n1095), .Z(n1584) );
  XOR U2441 ( .A(n1597), .B(n1596), .Z(n1577) );
  XOR U2442 ( .A(n1672), .B(n1592), .Z(n1596) );
  XNOR U2443 ( .A(n1590), .B(n1673), .Z(n1592) );
  ANDN U2444 ( .A(n974), .B(n1519), .Z(n1673) );
  XOR U2445 ( .A(n1674), .B(n1675), .Z(n1590) );
  AND U2446 ( .A(n1676), .B(n1677), .Z(n1675) );
  XNOR U2447 ( .A(n1678), .B(n1674), .Z(n1677) );
  AND U2448 ( .A(n1517), .B(n933), .Z(n1594) );
  XOR U2449 ( .A(n1604), .B(n1603), .Z(n1597) );
  NAND U2450 ( .A(n1682), .B(n877), .Z(n1603) );
  XOR U2451 ( .A(n1602), .B(n1683), .Z(n1604) );
  ANDN U2452 ( .A(n908), .B(n1684), .Z(n1683) );
  ANDN U2453 ( .A(n1685), .B(n1686), .Z(n1602) );
  NAND U2454 ( .A(n1687), .B(n1688), .Z(n1685) );
  IV U2455 ( .A(n1605), .Z(n1606) );
  MUX U2456 ( .IN0(Y[14]), .IN1(n776), .SEL(n829), .F(n301) );
  XOR U2457 ( .A(n1693), .B(Y0[15]), .Z(n776) );
  XOR U2458 ( .A(n1694), .B(n1695), .Z(n1693) );
  AND U2459 ( .A(n841), .B(n1697), .Z(n1696) );
  XOR U2460 ( .A(n1691), .B(n1695), .Z(n1697) );
  XOR U2461 ( .A(n1690), .B(n1695), .Z(n1691) );
  XNOR U2462 ( .A(n1616), .B(n1615), .Z(n1695) );
  XOR U2463 ( .A(n1698), .B(n1699), .Z(n1615) );
  XOR U2464 ( .A(n1700), .B(n1701), .Z(n1699) );
  XOR U2465 ( .A(n1702), .B(n1700), .Z(n1701) );
  XNOR U2466 ( .A(n1708), .B(n1644), .Z(n1633) );
  XNOR U2467 ( .A(n1627), .B(n1626), .Z(n1644) );
  XOR U2468 ( .A(n1709), .B(n1622), .Z(n1626) );
  XNOR U2469 ( .A(n1620), .B(n1710), .Z(n1622) );
  ANDN U2470 ( .A(n1386), .B(n1067), .Z(n1710) );
  AND U2471 ( .A(n1065), .B(n1323), .Z(n1624) );
  XNOR U2472 ( .A(n1630), .B(n1631), .Z(n1627) );
  NANDN U2473 ( .B(n1188), .A(n1166), .Z(n1631) );
  XNOR U2474 ( .A(n1629), .B(n1717), .Z(n1630) );
  ANDN U2475 ( .A(n1258), .B(n1168), .Z(n1717) );
  XOR U2476 ( .A(n1718), .B(n1719), .Z(n1629) );
  AND U2477 ( .A(n1720), .B(n1721), .Z(n1719) );
  XOR U2478 ( .A(n1722), .B(n1718), .Z(n1721) );
  XNOR U2479 ( .A(n1643), .B(n1632), .Z(n1708) );
  XOR U2480 ( .A(n1726), .B(n1653), .Z(n1643) );
  XNOR U2481 ( .A(n1639), .B(n1641), .Z(n1653) );
  NAND U2482 ( .A(n981), .B(n1557), .Z(n1641) );
  XNOR U2483 ( .A(n1637), .B(n1727), .Z(n1639) );
  ANDN U2484 ( .A(n1564), .B(n983), .Z(n1727) );
  XOR U2485 ( .A(n1728), .B(n1729), .Z(n1637) );
  AND U2486 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U2487 ( .A(n1732), .B(n1728), .Z(n1731) );
  XNOR U2488 ( .A(n1652), .B(n1642), .Z(n1726) );
  XOR U2489 ( .A(n1740), .B(n1650), .Z(n1736) );
  AND U2490 ( .A(n906), .B(n1741), .Z(n1650) );
  NAND U2491 ( .A(n1742), .B(n1649), .Z(n1740) );
  XOR U2492 ( .A(n1743), .B(n1744), .Z(n1649) );
  AND U2493 ( .A(n1745), .B(n1746), .Z(n1744) );
  XNOR U2494 ( .A(n1747), .B(n1743), .Z(n1746) );
  NANDN U2495 ( .B(n909), .A(n1748), .Z(n1742) );
  XNOR U2496 ( .A(n1661), .B(n1660), .Z(n1634) );
  XOR U2497 ( .A(n1749), .B(n1671), .Z(n1660) );
  XNOR U2498 ( .A(n1657), .B(n1658), .Z(n1671) );
  NANDN U2499 ( .B(n1001), .A(n1439), .Z(n1658) );
  XNOR U2500 ( .A(n1656), .B(n1750), .Z(n1657) );
  ANDN U2501 ( .A(n1042), .B(n1441), .Z(n1750) );
  XNOR U2502 ( .A(n1670), .B(n1659), .Z(n1749) );
  XOR U2503 ( .A(n1757), .B(n1666), .Z(n1670) );
  XNOR U2504 ( .A(n1664), .B(n1758), .Z(n1666) );
  ANDN U2505 ( .A(n1149), .B(n1300), .Z(n1758) );
  AND U2506 ( .A(n1298), .B(n1095), .Z(n1668) );
  XOR U2507 ( .A(n1681), .B(n1680), .Z(n1661) );
  XOR U2508 ( .A(n1765), .B(n1676), .Z(n1680) );
  XNOR U2509 ( .A(n1674), .B(n1766), .Z(n1676) );
  ANDN U2510 ( .A(n974), .B(n1600), .Z(n1766) );
  AND U2511 ( .A(n1598), .B(n933), .Z(n1678) );
  XOR U2512 ( .A(n1688), .B(n1687), .Z(n1681) );
  NAND U2513 ( .A(n1773), .B(n877), .Z(n1687) );
  XNOR U2514 ( .A(n1686), .B(n1774), .Z(n1688) );
  ANDN U2515 ( .A(n908), .B(n1775), .Z(n1774) );
  NAND U2516 ( .A(n1776), .B(n1777), .Z(n1686) );
  NAND U2517 ( .A(n1778), .B(n1779), .Z(n1776) );
  IV U2518 ( .A(n1689), .Z(n1690) );
  MUX U2519 ( .IN0(Y[13]), .IN1(n773), .SEL(n829), .F(n300) );
  XOR U2520 ( .A(n1784), .B(Y0[14]), .Z(n773) );
  XOR U2521 ( .A(n1785), .B(n1786), .Z(n1784) );
  AND U2522 ( .A(n841), .B(n1788), .Z(n1787) );
  XOR U2523 ( .A(n1782), .B(n1786), .Z(n1788) );
  XOR U2524 ( .A(n1781), .B(n1786), .Z(n1782) );
  XOR U2525 ( .A(n1789), .B(n1703), .Z(n1706) );
  NAND U2526 ( .A(n1700), .B(n1793), .Z(n1704) );
  AND U2527 ( .A(n1794), .B(n1795), .Z(n1793) );
  NANDN U2528 ( .B(n1796), .A(n876), .Z(n1795) );
  NANDN U2529 ( .B(n1797), .A(n1798), .Z(n1794) );
  AND U2530 ( .A(n1799), .B(n1800), .Z(n1700) );
  NANDN U2531 ( .B(n1801), .A(n1802), .Z(n1800) );
  OR U2532 ( .A(n1803), .B(n1804), .Z(n1799) );
  XNOR U2533 ( .A(n1725), .B(n1724), .Z(n1707) );
  XOR U2534 ( .A(n1808), .B(n1735), .Z(n1724) );
  XNOR U2535 ( .A(n1716), .B(n1715), .Z(n1735) );
  XOR U2536 ( .A(n1809), .B(n1712), .Z(n1715) );
  XNOR U2537 ( .A(n1711), .B(n1810), .Z(n1712) );
  ANDN U2538 ( .A(n1386), .B(n1109), .Z(n1810) );
  XOR U2539 ( .A(n1811), .B(n1812), .Z(n1711) );
  AND U2540 ( .A(n1813), .B(n1814), .Z(n1812) );
  XNOR U2541 ( .A(n1815), .B(n1811), .Z(n1814) );
  AND U2542 ( .A(n1107), .B(n1323), .Z(n1713) );
  XNOR U2543 ( .A(n1720), .B(n1722), .Z(n1716) );
  NANDN U2544 ( .B(n1188), .A(n1230), .Z(n1722) );
  XNOR U2545 ( .A(n1718), .B(n1819), .Z(n1720) );
  ANDN U2546 ( .A(n1258), .B(n1232), .Z(n1819) );
  XNOR U2547 ( .A(n1734), .B(n1723), .Z(n1808) );
  XOR U2548 ( .A(n1826), .B(n1739), .Z(n1734) );
  XNOR U2549 ( .A(n1730), .B(n1732), .Z(n1739) );
  NAND U2550 ( .A(n1021), .B(n1557), .Z(n1732) );
  XNOR U2551 ( .A(n1728), .B(n1827), .Z(n1730) );
  ANDN U2552 ( .A(n1564), .B(n1023), .Z(n1827) );
  XOR U2553 ( .A(n1828), .B(n1829), .Z(n1728) );
  AND U2554 ( .A(n1830), .B(n1831), .Z(n1829) );
  XOR U2555 ( .A(n1832), .B(n1828), .Z(n1831) );
  XNOR U2556 ( .A(n1738), .B(n1733), .Z(n1826) );
  XOR U2557 ( .A(n1836), .B(n1745), .Z(n1738) );
  XNOR U2558 ( .A(n1743), .B(n1837), .Z(n1745) );
  ANDN U2559 ( .A(n1748), .B(n939), .Z(n1837) );
  XOR U2560 ( .A(n1838), .B(n1839), .Z(n1743) );
  AND U2561 ( .A(n1840), .B(n1841), .Z(n1839) );
  XNOR U2562 ( .A(n1842), .B(n1838), .Z(n1841) );
  AND U2563 ( .A(n937), .B(n1741), .Z(n1747) );
  XNOR U2564 ( .A(n1756), .B(n1755), .Z(n1725) );
  XOR U2565 ( .A(n1846), .B(n1764), .Z(n1755) );
  XNOR U2566 ( .A(n1752), .B(n1753), .Z(n1764) );
  NANDN U2567 ( .B(n1001), .A(n1517), .Z(n1753) );
  XNOR U2568 ( .A(n1751), .B(n1847), .Z(n1752) );
  ANDN U2569 ( .A(n1042), .B(n1519), .Z(n1847) );
  XNOR U2570 ( .A(n1763), .B(n1754), .Z(n1846) );
  XOR U2571 ( .A(n1854), .B(n1760), .Z(n1763) );
  XNOR U2572 ( .A(n1759), .B(n1855), .Z(n1760) );
  ANDN U2573 ( .A(n1149), .B(n1367), .Z(n1855) );
  AND U2574 ( .A(n1365), .B(n1095), .Z(n1761) );
  XOR U2575 ( .A(n1772), .B(n1771), .Z(n1756) );
  XOR U2576 ( .A(n1862), .B(n1768), .Z(n1771) );
  XNOR U2577 ( .A(n1767), .B(n1863), .Z(n1768) );
  ANDN U2578 ( .A(n974), .B(n1684), .Z(n1863) );
  AND U2579 ( .A(n1682), .B(n933), .Z(n1769) );
  XOR U2580 ( .A(n1779), .B(n1778), .Z(n1772) );
  NAND U2581 ( .A(n1870), .B(n877), .Z(n1778) );
  XOR U2582 ( .A(n1777), .B(n1871), .Z(n1779) );
  ANDN U2583 ( .A(n908), .B(n1872), .Z(n1871) );
  ANDN U2584 ( .A(n1873), .B(n1874), .Z(n1777) );
  NAND U2585 ( .A(n1875), .B(n1876), .Z(n1873) );
  IV U2586 ( .A(n1780), .Z(n1781) );
  MUX U2587 ( .IN0(Y[12]), .IN1(n770), .SEL(n829), .F(n299) );
  XOR U2588 ( .A(n1881), .B(Y0[13]), .Z(n770) );
  XNOR U2589 ( .A(n1882), .B(n1883), .Z(n1881) );
  AND U2590 ( .A(n841), .B(n1885), .Z(n1884) );
  XNOR U2591 ( .A(n1879), .B(n1883), .Z(n1885) );
  XNOR U2592 ( .A(n1878), .B(n1883), .Z(n1879) );
  XNOR U2593 ( .A(n1807), .B(n1806), .Z(n1883) );
  XOR U2594 ( .A(n1886), .B(n1791), .Z(n1806) );
  NANDN U2595 ( .B(n1887), .A(n1888), .Z(n1797) );
  XOR U2596 ( .A(n1891), .B(n1804), .Z(n1801) );
  NAND U2597 ( .A(n1892), .B(n906), .Z(n1804) );
  NAND U2598 ( .A(n1893), .B(n1803), .Z(n1891) );
  NANDN U2599 ( .B(n909), .A(n1897), .Z(n1893) );
  XNOR U2600 ( .A(n1790), .B(n1805), .Z(n1886) );
  IV U2601 ( .A(n1792), .Z(n1790) );
  XNOR U2602 ( .A(n1825), .B(n1824), .Z(n1807) );
  XOR U2603 ( .A(n1904), .B(n1835), .Z(n1824) );
  XNOR U2604 ( .A(n1818), .B(n1817), .Z(n1835) );
  XOR U2605 ( .A(n1905), .B(n1813), .Z(n1817) );
  XNOR U2606 ( .A(n1811), .B(n1906), .Z(n1813) );
  ANDN U2607 ( .A(n1386), .B(n1168), .Z(n1906) );
  XOR U2608 ( .A(n1907), .B(n1908), .Z(n1811) );
  AND U2609 ( .A(n1909), .B(n1910), .Z(n1908) );
  XNOR U2610 ( .A(n1911), .B(n1907), .Z(n1910) );
  AND U2611 ( .A(n1166), .B(n1323), .Z(n1815) );
  XNOR U2612 ( .A(n1821), .B(n1822), .Z(n1818) );
  NANDN U2613 ( .B(n1188), .A(n1298), .Z(n1822) );
  XNOR U2614 ( .A(n1820), .B(n1915), .Z(n1821) );
  ANDN U2615 ( .A(n1258), .B(n1300), .Z(n1915) );
  XNOR U2616 ( .A(n1834), .B(n1823), .Z(n1904) );
  XOR U2617 ( .A(n1922), .B(n1845), .Z(n1834) );
  XNOR U2618 ( .A(n1830), .B(n1832), .Z(n1845) );
  NAND U2619 ( .A(n1065), .B(n1557), .Z(n1832) );
  XNOR U2620 ( .A(n1828), .B(n1923), .Z(n1830) );
  ANDN U2621 ( .A(n1564), .B(n1067), .Z(n1923) );
  XOR U2622 ( .A(n1924), .B(n1925), .Z(n1828) );
  AND U2623 ( .A(n1926), .B(n1927), .Z(n1925) );
  XOR U2624 ( .A(n1928), .B(n1924), .Z(n1927) );
  XNOR U2625 ( .A(n1844), .B(n1833), .Z(n1922) );
  XOR U2626 ( .A(n1932), .B(n1840), .Z(n1844) );
  XNOR U2627 ( .A(n1838), .B(n1933), .Z(n1840) );
  ANDN U2628 ( .A(n1748), .B(n983), .Z(n1933) );
  XOR U2629 ( .A(n1934), .B(n1935), .Z(n1838) );
  AND U2630 ( .A(n1936), .B(n1937), .Z(n1935) );
  XNOR U2631 ( .A(n1938), .B(n1934), .Z(n1937) );
  AND U2632 ( .A(n981), .B(n1741), .Z(n1842) );
  XNOR U2633 ( .A(n1853), .B(n1852), .Z(n1825) );
  XOR U2634 ( .A(n1942), .B(n1861), .Z(n1852) );
  XNOR U2635 ( .A(n1849), .B(n1850), .Z(n1861) );
  NANDN U2636 ( .B(n1001), .A(n1598), .Z(n1850) );
  XNOR U2637 ( .A(n1848), .B(n1943), .Z(n1849) );
  ANDN U2638 ( .A(n1042), .B(n1600), .Z(n1943) );
  XNOR U2639 ( .A(n1860), .B(n1851), .Z(n1942) );
  XOR U2640 ( .A(n1950), .B(n1857), .Z(n1860) );
  XNOR U2641 ( .A(n1856), .B(n1951), .Z(n1857) );
  ANDN U2642 ( .A(n1149), .B(n1441), .Z(n1951) );
  AND U2643 ( .A(n1439), .B(n1095), .Z(n1858) );
  XOR U2644 ( .A(n1869), .B(n1868), .Z(n1853) );
  XOR U2645 ( .A(n1958), .B(n1865), .Z(n1868) );
  XNOR U2646 ( .A(n1864), .B(n1959), .Z(n1865) );
  ANDN U2647 ( .A(n974), .B(n1775), .Z(n1959) );
  AND U2648 ( .A(n1773), .B(n933), .Z(n1866) );
  XOR U2649 ( .A(n1876), .B(n1875), .Z(n1869) );
  NAND U2650 ( .A(n1966), .B(n877), .Z(n1875) );
  XNOR U2651 ( .A(n1874), .B(n1967), .Z(n1876) );
  ANDN U2652 ( .A(n908), .B(n1968), .Z(n1967) );
  NAND U2653 ( .A(n1969), .B(n1970), .Z(n1874) );
  NAND U2654 ( .A(n1971), .B(n1972), .Z(n1969) );
  IV U2655 ( .A(n1877), .Z(n1878) );
  MUX U2656 ( .IN0(Y[11]), .IN1(n767), .SEL(n829), .F(n298) );
  XOR U2657 ( .A(n1977), .B(Y0[12]), .Z(n767) );
  XOR U2658 ( .A(n1978), .B(n1979), .Z(n1977) );
  AND U2659 ( .A(n841), .B(n1981), .Z(n1980) );
  XOR U2660 ( .A(n1975), .B(n1979), .Z(n1981) );
  XOR U2661 ( .A(n1974), .B(n1979), .Z(n1975) );
  XNOR U2662 ( .A(n1982), .B(n1903), .Z(n1899) );
  XOR U2663 ( .A(n1888), .B(n1887), .Z(n1903) );
  NANDN U2664 ( .B(n1983), .A(n1984), .Z(n1887) );
  AND U2665 ( .A(n1986), .B(n1987), .Z(n1985) );
  NANDN U2666 ( .B(n1988), .A(n876), .Z(n1987) );
  NANDN U2667 ( .B(n1989), .A(n1990), .Z(n1986) );
  XNOR U2668 ( .A(n1895), .B(n1896), .Z(n1890) );
  NAND U2669 ( .A(n1892), .B(n937), .Z(n1896) );
  XNOR U2670 ( .A(n1894), .B(n1994), .Z(n1895) );
  ANDN U2671 ( .A(n1897), .B(n939), .Z(n1994) );
  XNOR U2672 ( .A(n1902), .B(n1898), .Z(n1982) );
  IV U2673 ( .A(n1901), .Z(n1902) );
  XNOR U2674 ( .A(n1921), .B(n1920), .Z(n1900) );
  XOR U2675 ( .A(n2004), .B(n1931), .Z(n1920) );
  XNOR U2676 ( .A(n1914), .B(n1913), .Z(n1931) );
  XOR U2677 ( .A(n2005), .B(n1909), .Z(n1913) );
  XNOR U2678 ( .A(n1907), .B(n2006), .Z(n1909) );
  ANDN U2679 ( .A(n1386), .B(n1232), .Z(n2006) );
  AND U2680 ( .A(n1230), .B(n1323), .Z(n1911) );
  XNOR U2681 ( .A(n1917), .B(n1918), .Z(n1914) );
  NANDN U2682 ( .B(n1188), .A(n1365), .Z(n1918) );
  XNOR U2683 ( .A(n1916), .B(n2013), .Z(n1917) );
  ANDN U2684 ( .A(n1258), .B(n1367), .Z(n2013) );
  XNOR U2685 ( .A(n1930), .B(n1919), .Z(n2004) );
  XOR U2686 ( .A(n2020), .B(n1941), .Z(n1930) );
  XNOR U2687 ( .A(n1926), .B(n1928), .Z(n1941) );
  NAND U2688 ( .A(n1107), .B(n1557), .Z(n1928) );
  XNOR U2689 ( .A(n1924), .B(n2021), .Z(n1926) );
  ANDN U2690 ( .A(n1564), .B(n1109), .Z(n2021) );
  XNOR U2691 ( .A(n1940), .B(n1929), .Z(n2020) );
  XOR U2692 ( .A(n2028), .B(n1936), .Z(n1940) );
  XNOR U2693 ( .A(n1934), .B(n2029), .Z(n1936) );
  ANDN U2694 ( .A(n1748), .B(n1023), .Z(n2029) );
  XOR U2695 ( .A(n2030), .B(n2031), .Z(n1934) );
  AND U2696 ( .A(n2032), .B(n2033), .Z(n2031) );
  XNOR U2697 ( .A(n2034), .B(n2030), .Z(n2033) );
  AND U2698 ( .A(n1021), .B(n1741), .Z(n1938) );
  XNOR U2699 ( .A(n1949), .B(n1948), .Z(n1921) );
  XOR U2700 ( .A(n2038), .B(n1957), .Z(n1948) );
  XNOR U2701 ( .A(n1945), .B(n1946), .Z(n1957) );
  NANDN U2702 ( .B(n1001), .A(n1682), .Z(n1946) );
  XNOR U2703 ( .A(n1944), .B(n2039), .Z(n1945) );
  ANDN U2704 ( .A(n1042), .B(n1684), .Z(n2039) );
  XNOR U2705 ( .A(n1956), .B(n1947), .Z(n2038) );
  XOR U2706 ( .A(n2046), .B(n1953), .Z(n1956) );
  XNOR U2707 ( .A(n1952), .B(n2047), .Z(n1953) );
  ANDN U2708 ( .A(n1149), .B(n1519), .Z(n2047) );
  AND U2709 ( .A(n1517), .B(n1095), .Z(n1954) );
  XOR U2710 ( .A(n1965), .B(n1964), .Z(n1949) );
  XOR U2711 ( .A(n2054), .B(n1961), .Z(n1964) );
  XNOR U2712 ( .A(n1960), .B(n2055), .Z(n1961) );
  ANDN U2713 ( .A(n974), .B(n1872), .Z(n2055) );
  AND U2714 ( .A(n1870), .B(n933), .Z(n1962) );
  XOR U2715 ( .A(n1972), .B(n1971), .Z(n1965) );
  NAND U2716 ( .A(n2062), .B(n877), .Z(n1971) );
  XOR U2717 ( .A(n1970), .B(n2063), .Z(n1972) );
  ANDN U2718 ( .A(n908), .B(n2064), .Z(n2063) );
  ANDN U2719 ( .A(n2065), .B(n2066), .Z(n1970) );
  NAND U2720 ( .A(n2067), .B(n2068), .Z(n2065) );
  IV U2721 ( .A(n1973), .Z(n1974) );
  MUX U2722 ( .IN0(Y[10]), .IN1(n764), .SEL(n829), .F(n297) );
  XOR U2723 ( .A(n2073), .B(Y0[11]), .Z(n764) );
  XNOR U2724 ( .A(n2074), .B(n2075), .Z(n2073) );
  AND U2725 ( .A(n841), .B(n2077), .Z(n2076) );
  XNOR U2726 ( .A(n2071), .B(n2075), .Z(n2077) );
  XNOR U2727 ( .A(n2070), .B(n2075), .Z(n2071) );
  XNOR U2728 ( .A(n2000), .B(n1999), .Z(n2075) );
  XOR U2729 ( .A(n2078), .B(n2003), .Z(n1999) );
  XOR U2730 ( .A(n1993), .B(n1992), .Z(n1983) );
  XOR U2731 ( .A(n2086), .B(n1990), .Z(n2082) );
  AND U2732 ( .A(n2087), .B(n906), .Z(n1990) );
  NAND U2733 ( .A(n2088), .B(n1989), .Z(n2086) );
  XOR U2734 ( .A(n2089), .B(n2090), .Z(n1989) );
  AND U2735 ( .A(n2091), .B(n2092), .Z(n2090) );
  XNOR U2736 ( .A(n2093), .B(n2089), .Z(n2092) );
  NANDN U2737 ( .B(n909), .A(n2094), .Z(n2088) );
  XNOR U2738 ( .A(n1996), .B(n1997), .Z(n1993) );
  NAND U2739 ( .A(n1892), .B(n981), .Z(n1997) );
  XNOR U2740 ( .A(n1995), .B(n2095), .Z(n1996) );
  ANDN U2741 ( .A(n1897), .B(n983), .Z(n2095) );
  XNOR U2742 ( .A(n2002), .B(n1998), .Z(n2078) );
  IV U2743 ( .A(n2001), .Z(n2002) );
  XNOR U2744 ( .A(n2019), .B(n2018), .Z(n2000) );
  XOR U2745 ( .A(n2105), .B(n2027), .Z(n2018) );
  XNOR U2746 ( .A(n2012), .B(n2011), .Z(n2027) );
  XOR U2747 ( .A(n2106), .B(n2008), .Z(n2011) );
  XNOR U2748 ( .A(n2007), .B(n2107), .Z(n2008) );
  ANDN U2749 ( .A(n1386), .B(n1300), .Z(n2107) );
  AND U2750 ( .A(n1298), .B(n1323), .Z(n2009) );
  XNOR U2751 ( .A(n2015), .B(n2016), .Z(n2012) );
  NANDN U2752 ( .B(n1188), .A(n1439), .Z(n2016) );
  XNOR U2753 ( .A(n2014), .B(n2114), .Z(n2015) );
  ANDN U2754 ( .A(n1258), .B(n1441), .Z(n2114) );
  XNOR U2755 ( .A(n2026), .B(n2017), .Z(n2105) );
  XOR U2756 ( .A(n2121), .B(n2037), .Z(n2026) );
  XNOR U2757 ( .A(n2023), .B(n2024), .Z(n2037) );
  NAND U2758 ( .A(n1166), .B(n1557), .Z(n2024) );
  XNOR U2759 ( .A(n2022), .B(n2122), .Z(n2023) );
  ANDN U2760 ( .A(n1564), .B(n1168), .Z(n2122) );
  XNOR U2761 ( .A(n2036), .B(n2025), .Z(n2121) );
  XOR U2762 ( .A(n2129), .B(n2032), .Z(n2036) );
  XNOR U2763 ( .A(n2030), .B(n2130), .Z(n2032) );
  ANDN U2764 ( .A(n1748), .B(n1067), .Z(n2130) );
  XOR U2765 ( .A(n2131), .B(n2132), .Z(n2030) );
  AND U2766 ( .A(n2133), .B(n2134), .Z(n2132) );
  XNOR U2767 ( .A(n2135), .B(n2131), .Z(n2134) );
  AND U2768 ( .A(n1065), .B(n1741), .Z(n2034) );
  XNOR U2769 ( .A(n2045), .B(n2044), .Z(n2019) );
  XOR U2770 ( .A(n2139), .B(n2053), .Z(n2044) );
  XNOR U2771 ( .A(n2041), .B(n2042), .Z(n2053) );
  NANDN U2772 ( .B(n1001), .A(n1773), .Z(n2042) );
  XNOR U2773 ( .A(n2040), .B(n2140), .Z(n2041) );
  ANDN U2774 ( .A(n1042), .B(n1775), .Z(n2140) );
  XNOR U2775 ( .A(n2052), .B(n2043), .Z(n2139) );
  XOR U2776 ( .A(n2147), .B(n2049), .Z(n2052) );
  XNOR U2777 ( .A(n2048), .B(n2148), .Z(n2049) );
  ANDN U2778 ( .A(n1149), .B(n1600), .Z(n2148) );
  AND U2779 ( .A(n1598), .B(n1095), .Z(n2050) );
  XOR U2780 ( .A(n2061), .B(n2060), .Z(n2045) );
  XOR U2781 ( .A(n2155), .B(n2057), .Z(n2060) );
  XNOR U2782 ( .A(n2056), .B(n2156), .Z(n2057) );
  ANDN U2783 ( .A(n974), .B(n1968), .Z(n2156) );
  AND U2784 ( .A(n1966), .B(n933), .Z(n2058) );
  XOR U2785 ( .A(n2068), .B(n2067), .Z(n2061) );
  NAND U2786 ( .A(n2163), .B(n877), .Z(n2067) );
  XNOR U2787 ( .A(n2066), .B(n2164), .Z(n2068) );
  ANDN U2788 ( .A(n908), .B(n2165), .Z(n2164) );
  NAND U2789 ( .A(n2166), .B(n2167), .Z(n2066) );
  NAND U2790 ( .A(n2168), .B(n2169), .Z(n2166) );
  IV U2791 ( .A(n2069), .Z(n2070) );
  MUX U2792 ( .IN0(Y[9]), .IN1(n761), .SEL(n829), .F(n296) );
  XOR U2793 ( .A(n2174), .B(Y0[10]), .Z(n761) );
  XOR U2794 ( .A(n2175), .B(n2176), .Z(n2174) );
  AND U2795 ( .A(n841), .B(n2178), .Z(n2177) );
  XOR U2796 ( .A(n2172), .B(n2176), .Z(n2178) );
  XOR U2797 ( .A(n2171), .B(n2176), .Z(n2172) );
  XNOR U2798 ( .A(n2179), .B(n2104), .Z(n2100) );
  XNOR U2799 ( .A(n2081), .B(n2080), .Z(n2104) );
  XOR U2800 ( .A(n2079), .B(n2180), .Z(n2080) );
  AND U2801 ( .A(n2181), .B(n2182), .Z(n2180) );
  NANDN U2802 ( .B(n2183), .A(n2184), .Z(n2182) );
  AND U2803 ( .A(n2185), .B(n2186), .Z(n2181) );
  NANDN U2804 ( .B(n2187), .A(n876), .Z(n2186) );
  OR U2805 ( .A(n2188), .B(n2189), .Z(n2185) );
  XNOR U2806 ( .A(n2085), .B(n2084), .Z(n2081) );
  XOR U2807 ( .A(n2193), .B(n2091), .Z(n2084) );
  XNOR U2808 ( .A(n2089), .B(n2194), .Z(n2091) );
  ANDN U2809 ( .A(n2094), .B(n939), .Z(n2194) );
  XOR U2810 ( .A(n2195), .B(n2196), .Z(n2089) );
  AND U2811 ( .A(n2197), .B(n2198), .Z(n2196) );
  XNOR U2812 ( .A(n2199), .B(n2195), .Z(n2198) );
  AND U2813 ( .A(n2087), .B(n937), .Z(n2093) );
  XNOR U2814 ( .A(n2097), .B(n2098), .Z(n2085) );
  NAND U2815 ( .A(n1892), .B(n1021), .Z(n2098) );
  XNOR U2816 ( .A(n2096), .B(n2203), .Z(n2097) );
  ANDN U2817 ( .A(n1897), .B(n1023), .Z(n2203) );
  XNOR U2818 ( .A(n2103), .B(n2099), .Z(n2179) );
  IV U2819 ( .A(n2102), .Z(n2103) );
  XNOR U2820 ( .A(n2120), .B(n2119), .Z(n2101) );
  XOR U2821 ( .A(n2213), .B(n2128), .Z(n2119) );
  XNOR U2822 ( .A(n2113), .B(n2112), .Z(n2128) );
  XOR U2823 ( .A(n2214), .B(n2109), .Z(n2112) );
  XNOR U2824 ( .A(n2108), .B(n2215), .Z(n2109) );
  ANDN U2825 ( .A(n1386), .B(n1367), .Z(n2215) );
  AND U2826 ( .A(n1365), .B(n1323), .Z(n2110) );
  XNOR U2827 ( .A(n2116), .B(n2117), .Z(n2113) );
  NANDN U2828 ( .B(n1188), .A(n1517), .Z(n2117) );
  XNOR U2829 ( .A(n2115), .B(n2222), .Z(n2116) );
  ANDN U2830 ( .A(n1258), .B(n1519), .Z(n2222) );
  XNOR U2831 ( .A(n2127), .B(n2118), .Z(n2213) );
  XOR U2832 ( .A(n2229), .B(n2138), .Z(n2127) );
  XNOR U2833 ( .A(n2124), .B(n2125), .Z(n2138) );
  NAND U2834 ( .A(n1230), .B(n1557), .Z(n2125) );
  XNOR U2835 ( .A(n2123), .B(n2230), .Z(n2124) );
  ANDN U2836 ( .A(n1564), .B(n1232), .Z(n2230) );
  XNOR U2837 ( .A(n2137), .B(n2126), .Z(n2229) );
  XOR U2838 ( .A(n2237), .B(n2133), .Z(n2137) );
  XNOR U2839 ( .A(n2131), .B(n2238), .Z(n2133) );
  ANDN U2840 ( .A(n1748), .B(n1109), .Z(n2238) );
  AND U2841 ( .A(n1107), .B(n1741), .Z(n2135) );
  XNOR U2842 ( .A(n2146), .B(n2145), .Z(n2120) );
  XOR U2843 ( .A(n2245), .B(n2154), .Z(n2145) );
  XNOR U2844 ( .A(n2142), .B(n2143), .Z(n2154) );
  NANDN U2845 ( .B(n1001), .A(n1870), .Z(n2143) );
  XNOR U2846 ( .A(n2141), .B(n2246), .Z(n2142) );
  ANDN U2847 ( .A(n1042), .B(n1872), .Z(n2246) );
  XNOR U2848 ( .A(n2153), .B(n2144), .Z(n2245) );
  XOR U2849 ( .A(n2253), .B(n2150), .Z(n2153) );
  XNOR U2850 ( .A(n2149), .B(n2254), .Z(n2150) );
  ANDN U2851 ( .A(n1149), .B(n1684), .Z(n2254) );
  AND U2852 ( .A(n1682), .B(n1095), .Z(n2151) );
  XOR U2853 ( .A(n2162), .B(n2161), .Z(n2146) );
  XOR U2854 ( .A(n2261), .B(n2158), .Z(n2161) );
  XNOR U2855 ( .A(n2157), .B(n2262), .Z(n2158) );
  ANDN U2856 ( .A(n974), .B(n2064), .Z(n2262) );
  AND U2857 ( .A(n2062), .B(n933), .Z(n2159) );
  XOR U2858 ( .A(n2169), .B(n2168), .Z(n2162) );
  NAND U2859 ( .A(n2269), .B(n877), .Z(n2168) );
  XOR U2860 ( .A(n2167), .B(n2270), .Z(n2169) );
  ANDN U2861 ( .A(n908), .B(n2271), .Z(n2270) );
  ANDN U2862 ( .A(n2272), .B(n2273), .Z(n2167) );
  NAND U2863 ( .A(n2274), .B(n2275), .Z(n2272) );
  IV U2864 ( .A(n2170), .Z(n2171) );
  MUX U2865 ( .IN0(Y[8]), .IN1(n758), .SEL(n829), .F(n295) );
  XOR U2866 ( .A(n2280), .B(Y0[9]), .Z(n758) );
  XOR U2867 ( .A(n2281), .B(n2282), .Z(n2280) );
  AND U2868 ( .A(n841), .B(n2284), .Z(n2283) );
  XOR U2869 ( .A(n2278), .B(n2282), .Z(n2284) );
  XOR U2870 ( .A(n2277), .B(n2282), .Z(n2278) );
  XNOR U2871 ( .A(n2285), .B(n2212), .Z(n2208) );
  XNOR U2872 ( .A(n2192), .B(n2191), .Z(n2212) );
  XOR U2873 ( .A(n2286), .B(n2188), .Z(n2191) );
  XNOR U2874 ( .A(n2287), .B(n2184), .Z(n2188) );
  AND U2875 ( .A(n2288), .B(n906), .Z(n2184) );
  NAND U2876 ( .A(n2289), .B(n2183), .Z(n2287) );
  NANDN U2877 ( .B(n909), .A(n2293), .Z(n2289) );
  XNOR U2878 ( .A(n2189), .B(n2190), .Z(n2286) );
  XNOR U2879 ( .A(n2297), .B(n2300), .Z(n2299) );
  XNOR U2880 ( .A(n2202), .B(n2201), .Z(n2192) );
  XOR U2881 ( .A(n2301), .B(n2197), .Z(n2201) );
  XNOR U2882 ( .A(n2195), .B(n2302), .Z(n2197) );
  ANDN U2883 ( .A(n2094), .B(n983), .Z(n2302) );
  XOR U2884 ( .A(n2303), .B(n2304), .Z(n2195) );
  AND U2885 ( .A(n2305), .B(n2306), .Z(n2304) );
  XNOR U2886 ( .A(n2307), .B(n2303), .Z(n2306) );
  AND U2887 ( .A(n2087), .B(n981), .Z(n2199) );
  XNOR U2888 ( .A(n2205), .B(n2206), .Z(n2202) );
  NAND U2889 ( .A(n1892), .B(n1065), .Z(n2206) );
  XNOR U2890 ( .A(n2204), .B(n2311), .Z(n2205) );
  ANDN U2891 ( .A(n1897), .B(n1067), .Z(n2311) );
  XNOR U2892 ( .A(n2211), .B(n2207), .Z(n2285) );
  IV U2893 ( .A(n2210), .Z(n2211) );
  XNOR U2894 ( .A(n2228), .B(n2227), .Z(n2209) );
  XOR U2895 ( .A(n2320), .B(n2236), .Z(n2227) );
  XNOR U2896 ( .A(n2221), .B(n2220), .Z(n2236) );
  XOR U2897 ( .A(n2321), .B(n2217), .Z(n2220) );
  XNOR U2898 ( .A(n2216), .B(n2322), .Z(n2217) );
  ANDN U2899 ( .A(n1386), .B(n1441), .Z(n2322) );
  AND U2900 ( .A(n1439), .B(n1323), .Z(n2218) );
  XNOR U2901 ( .A(n2224), .B(n2225), .Z(n2221) );
  NANDN U2902 ( .B(n1188), .A(n1598), .Z(n2225) );
  XNOR U2903 ( .A(n2223), .B(n2329), .Z(n2224) );
  ANDN U2904 ( .A(n1258), .B(n1600), .Z(n2329) );
  XNOR U2905 ( .A(n2235), .B(n2226), .Z(n2320) );
  XOR U2906 ( .A(n2336), .B(n2244), .Z(n2235) );
  XNOR U2907 ( .A(n2232), .B(n2233), .Z(n2244) );
  NAND U2908 ( .A(n1298), .B(n1557), .Z(n2233) );
  XNOR U2909 ( .A(n2231), .B(n2337), .Z(n2232) );
  ANDN U2910 ( .A(n1564), .B(n1300), .Z(n2337) );
  XNOR U2911 ( .A(n2243), .B(n2234), .Z(n2336) );
  XOR U2912 ( .A(n2344), .B(n2240), .Z(n2243) );
  XNOR U2913 ( .A(n2239), .B(n2345), .Z(n2240) );
  ANDN U2914 ( .A(n1748), .B(n1168), .Z(n2345) );
  AND U2915 ( .A(n1166), .B(n1741), .Z(n2241) );
  XNOR U2916 ( .A(n2252), .B(n2251), .Z(n2228) );
  XOR U2917 ( .A(n2352), .B(n2260), .Z(n2251) );
  XNOR U2918 ( .A(n2248), .B(n2249), .Z(n2260) );
  NANDN U2919 ( .B(n1001), .A(n1966), .Z(n2249) );
  XNOR U2920 ( .A(n2247), .B(n2353), .Z(n2248) );
  ANDN U2921 ( .A(n1042), .B(n1968), .Z(n2353) );
  XNOR U2922 ( .A(n2259), .B(n2250), .Z(n2352) );
  XOR U2923 ( .A(n2360), .B(n2256), .Z(n2259) );
  XNOR U2924 ( .A(n2255), .B(n2361), .Z(n2256) );
  ANDN U2925 ( .A(n1149), .B(n1775), .Z(n2361) );
  AND U2926 ( .A(n1773), .B(n1095), .Z(n2257) );
  XOR U2927 ( .A(n2268), .B(n2267), .Z(n2252) );
  XOR U2928 ( .A(n2368), .B(n2264), .Z(n2267) );
  XNOR U2929 ( .A(n2263), .B(n2369), .Z(n2264) );
  ANDN U2930 ( .A(n974), .B(n2165), .Z(n2369) );
  AND U2931 ( .A(n2163), .B(n933), .Z(n2265) );
  XOR U2932 ( .A(n2275), .B(n2274), .Z(n2268) );
  NAND U2933 ( .A(n2376), .B(n877), .Z(n2274) );
  XNOR U2934 ( .A(n2273), .B(n2377), .Z(n2275) );
  ANDN U2935 ( .A(n908), .B(n2378), .Z(n2377) );
  NAND U2936 ( .A(n2379), .B(n2380), .Z(n2273) );
  NAND U2937 ( .A(n2381), .B(n2382), .Z(n2379) );
  IV U2938 ( .A(n2276), .Z(n2277) );
  MUX U2939 ( .IN0(Y[7]), .IN1(n755), .SEL(n829), .F(n294) );
  XOR U2940 ( .A(n2387), .B(Y0[8]), .Z(n755) );
  XOR U2941 ( .A(n2388), .B(n2389), .Z(n2387) );
  AND U2942 ( .A(n841), .B(n2391), .Z(n2390) );
  XOR U2943 ( .A(n2385), .B(n2389), .Z(n2391) );
  XOR U2944 ( .A(n2384), .B(n2389), .Z(n2385) );
  XNOR U2945 ( .A(n2392), .B(n2319), .Z(n2316) );
  XNOR U2946 ( .A(n2296), .B(n2295), .Z(n2319) );
  XOR U2947 ( .A(n2393), .B(n2300), .Z(n2295) );
  XNOR U2948 ( .A(n2291), .B(n2292), .Z(n2300) );
  NAND U2949 ( .A(n2288), .B(n937), .Z(n2292) );
  XNOR U2950 ( .A(n2290), .B(n2394), .Z(n2291) );
  ANDN U2951 ( .A(n2293), .B(n939), .Z(n2394) );
  XNOR U2952 ( .A(n2298), .B(n2294), .Z(n2393) );
  XOR U2953 ( .A(n2297), .B(n2401), .Z(n2298) );
  AND U2954 ( .A(n2402), .B(n2403), .Z(n2401) );
  NANDN U2955 ( .B(n2404), .A(n876), .Z(n2403) );
  NANDN U2956 ( .B(n2405), .A(n2406), .Z(n2402) );
  XNOR U2957 ( .A(n2310), .B(n2309), .Z(n2296) );
  XOR U2958 ( .A(n2410), .B(n2305), .Z(n2309) );
  XNOR U2959 ( .A(n2303), .B(n2411), .Z(n2305) );
  ANDN U2960 ( .A(n2094), .B(n1023), .Z(n2411) );
  AND U2961 ( .A(n2087), .B(n1021), .Z(n2307) );
  XNOR U2962 ( .A(n2313), .B(n2314), .Z(n2310) );
  NAND U2963 ( .A(n1892), .B(n1107), .Z(n2314) );
  XNOR U2964 ( .A(n2312), .B(n2418), .Z(n2313) );
  ANDN U2965 ( .A(n1897), .B(n1109), .Z(n2418) );
  XNOR U2966 ( .A(n2335), .B(n2334), .Z(n2317) );
  XOR U2967 ( .A(n2428), .B(n2343), .Z(n2334) );
  XNOR U2968 ( .A(n2328), .B(n2327), .Z(n2343) );
  XOR U2969 ( .A(n2429), .B(n2324), .Z(n2327) );
  XNOR U2970 ( .A(n2323), .B(n2430), .Z(n2324) );
  ANDN U2971 ( .A(n1386), .B(n1519), .Z(n2430) );
  AND U2972 ( .A(n1517), .B(n1323), .Z(n2325) );
  XNOR U2973 ( .A(n2331), .B(n2332), .Z(n2328) );
  NANDN U2974 ( .B(n1188), .A(n1682), .Z(n2332) );
  XNOR U2975 ( .A(n2330), .B(n2437), .Z(n2331) );
  ANDN U2976 ( .A(n1258), .B(n1684), .Z(n2437) );
  XNOR U2977 ( .A(n2342), .B(n2333), .Z(n2428) );
  XOR U2978 ( .A(n2444), .B(n2351), .Z(n2342) );
  XNOR U2979 ( .A(n2339), .B(n2340), .Z(n2351) );
  NAND U2980 ( .A(n1365), .B(n1557), .Z(n2340) );
  XNOR U2981 ( .A(n2338), .B(n2445), .Z(n2339) );
  ANDN U2982 ( .A(n1564), .B(n1367), .Z(n2445) );
  XNOR U2983 ( .A(n2350), .B(n2341), .Z(n2444) );
  XOR U2984 ( .A(n2452), .B(n2347), .Z(n2350) );
  XNOR U2985 ( .A(n2346), .B(n2453), .Z(n2347) );
  ANDN U2986 ( .A(n1748), .B(n1232), .Z(n2453) );
  AND U2987 ( .A(n1230), .B(n1741), .Z(n2348) );
  XNOR U2988 ( .A(n2359), .B(n2358), .Z(n2335) );
  XOR U2989 ( .A(n2460), .B(n2367), .Z(n2358) );
  XNOR U2990 ( .A(n2355), .B(n2356), .Z(n2367) );
  NANDN U2991 ( .B(n1001), .A(n2062), .Z(n2356) );
  XNOR U2992 ( .A(n2354), .B(n2461), .Z(n2355) );
  ANDN U2993 ( .A(n1042), .B(n2064), .Z(n2461) );
  XNOR U2994 ( .A(n2366), .B(n2357), .Z(n2460) );
  XOR U2995 ( .A(n2468), .B(n2363), .Z(n2366) );
  XNOR U2996 ( .A(n2362), .B(n2469), .Z(n2363) );
  ANDN U2997 ( .A(n1149), .B(n1872), .Z(n2469) );
  AND U2998 ( .A(n1870), .B(n1095), .Z(n2364) );
  XOR U2999 ( .A(n2375), .B(n2374), .Z(n2359) );
  XOR U3000 ( .A(n2476), .B(n2371), .Z(n2374) );
  XNOR U3001 ( .A(n2370), .B(n2477), .Z(n2371) );
  ANDN U3002 ( .A(n974), .B(n2271), .Z(n2477) );
  AND U3003 ( .A(n2269), .B(n933), .Z(n2372) );
  XOR U3004 ( .A(n2382), .B(n2381), .Z(n2375) );
  NAND U3005 ( .A(n2484), .B(n877), .Z(n2381) );
  XOR U3006 ( .A(n2380), .B(n2485), .Z(n2382) );
  ANDN U3007 ( .A(n908), .B(n2486), .Z(n2485) );
  ANDN U3008 ( .A(n2487), .B(n2488), .Z(n2380) );
  NAND U3009 ( .A(n2489), .B(n2490), .Z(n2487) );
  IV U3010 ( .A(n2383), .Z(n2384) );
  MUX U3011 ( .IN0(Y[6]), .IN1(n752), .SEL(n829), .F(n293) );
  XOR U3012 ( .A(n2495), .B(Y0[7]), .Z(n752) );
  XOR U3013 ( .A(n2496), .B(n2497), .Z(n2495) );
  AND U3014 ( .A(n841), .B(n2499), .Z(n2498) );
  XOR U3015 ( .A(n2493), .B(n2497), .Z(n2499) );
  XOR U3016 ( .A(n2492), .B(n2497), .Z(n2493) );
  XNOR U3017 ( .A(n2500), .B(n2427), .Z(n2423) );
  XNOR U3018 ( .A(n2400), .B(n2399), .Z(n2427) );
  XOR U3019 ( .A(n2501), .B(n2409), .Z(n2399) );
  XNOR U3020 ( .A(n2396), .B(n2397), .Z(n2409) );
  NAND U3021 ( .A(n2288), .B(n981), .Z(n2397) );
  XNOR U3022 ( .A(n2395), .B(n2502), .Z(n2396) );
  ANDN U3023 ( .A(n2293), .B(n983), .Z(n2502) );
  XOR U3024 ( .A(n2503), .B(n2504), .Z(n2395) );
  AND U3025 ( .A(n2505), .B(n2506), .Z(n2504) );
  XOR U3026 ( .A(n2507), .B(n2503), .Z(n2506) );
  XNOR U3027 ( .A(n2408), .B(n2398), .Z(n2501) );
  XOR U3028 ( .A(n2515), .B(n2406), .Z(n2511) );
  AND U3029 ( .A(n2516), .B(n906), .Z(n2406) );
  NAND U3030 ( .A(n2517), .B(n2405), .Z(n2515) );
  XOR U3031 ( .A(n2518), .B(n2519), .Z(n2405) );
  AND U3032 ( .A(n2520), .B(n2521), .Z(n2519) );
  XNOR U3033 ( .A(n2522), .B(n2518), .Z(n2521) );
  NANDN U3034 ( .B(n909), .A(n2523), .Z(n2517) );
  XNOR U3035 ( .A(n2417), .B(n2416), .Z(n2400) );
  XOR U3036 ( .A(n2524), .B(n2413), .Z(n2416) );
  XNOR U3037 ( .A(n2412), .B(n2525), .Z(n2413) );
  ANDN U3038 ( .A(n2094), .B(n1067), .Z(n2525) );
  AND U3039 ( .A(n2087), .B(n1065), .Z(n2414) );
  XNOR U3040 ( .A(n2420), .B(n2421), .Z(n2417) );
  NAND U3041 ( .A(n1892), .B(n1166), .Z(n2421) );
  XNOR U3042 ( .A(n2419), .B(n2532), .Z(n2420) );
  ANDN U3043 ( .A(n1897), .B(n1168), .Z(n2532) );
  XNOR U3044 ( .A(n2426), .B(n2422), .Z(n2500) );
  XOR U3045 ( .A(n2543), .B(n2544), .Z(n2539) );
  NANDN U3046 ( .B(n2545), .A(n2546), .Z(n2543) );
  XNOR U3047 ( .A(n2443), .B(n2442), .Z(n2424) );
  XOR U3048 ( .A(n2547), .B(n2451), .Z(n2442) );
  XNOR U3049 ( .A(n2436), .B(n2435), .Z(n2451) );
  XOR U3050 ( .A(n2548), .B(n2432), .Z(n2435) );
  XNOR U3051 ( .A(n2431), .B(n2549), .Z(n2432) );
  ANDN U3052 ( .A(n1386), .B(n1600), .Z(n2549) );
  AND U3053 ( .A(n1598), .B(n1323), .Z(n2433) );
  XNOR U3054 ( .A(n2439), .B(n2440), .Z(n2436) );
  NANDN U3055 ( .B(n1188), .A(n1773), .Z(n2440) );
  XNOR U3056 ( .A(n2438), .B(n2556), .Z(n2439) );
  ANDN U3057 ( .A(n1258), .B(n1775), .Z(n2556) );
  XNOR U3058 ( .A(n2450), .B(n2441), .Z(n2547) );
  XOR U3059 ( .A(n2563), .B(n2459), .Z(n2450) );
  XNOR U3060 ( .A(n2447), .B(n2448), .Z(n2459) );
  NAND U3061 ( .A(n1439), .B(n1557), .Z(n2448) );
  XNOR U3062 ( .A(n2446), .B(n2564), .Z(n2447) );
  ANDN U3063 ( .A(n1564), .B(n1441), .Z(n2564) );
  XNOR U3064 ( .A(n2458), .B(n2449), .Z(n2563) );
  XOR U3065 ( .A(n2571), .B(n2455), .Z(n2458) );
  XNOR U3066 ( .A(n2454), .B(n2572), .Z(n2455) );
  ANDN U3067 ( .A(n1748), .B(n1300), .Z(n2572) );
  AND U3068 ( .A(n1298), .B(n1741), .Z(n2456) );
  XNOR U3069 ( .A(n2467), .B(n2466), .Z(n2443) );
  XOR U3070 ( .A(n2579), .B(n2475), .Z(n2466) );
  XNOR U3071 ( .A(n2463), .B(n2464), .Z(n2475) );
  NANDN U3072 ( .B(n1001), .A(n2163), .Z(n2464) );
  XNOR U3073 ( .A(n2462), .B(n2580), .Z(n2463) );
  ANDN U3074 ( .A(n1042), .B(n2165), .Z(n2580) );
  XNOR U3075 ( .A(n2474), .B(n2465), .Z(n2579) );
  XOR U3076 ( .A(n2587), .B(n2471), .Z(n2474) );
  XNOR U3077 ( .A(n2470), .B(n2588), .Z(n2471) );
  ANDN U3078 ( .A(n1149), .B(n1968), .Z(n2588) );
  AND U3079 ( .A(n1966), .B(n1095), .Z(n2472) );
  XOR U3080 ( .A(n2483), .B(n2482), .Z(n2467) );
  XOR U3081 ( .A(n2595), .B(n2479), .Z(n2482) );
  XNOR U3082 ( .A(n2478), .B(n2596), .Z(n2479) );
  ANDN U3083 ( .A(n974), .B(n2378), .Z(n2596) );
  AND U3084 ( .A(n2376), .B(n933), .Z(n2480) );
  XOR U3085 ( .A(n2490), .B(n2489), .Z(n2483) );
  NAND U3086 ( .A(n2603), .B(n877), .Z(n2489) );
  XNOR U3087 ( .A(n2488), .B(n2604), .Z(n2490) );
  ANDN U3088 ( .A(n908), .B(n2605), .Z(n2604) );
  NAND U3089 ( .A(n2606), .B(n2607), .Z(n2488) );
  NAND U3090 ( .A(n2608), .B(n2609), .Z(n2606) );
  IV U3091 ( .A(n2491), .Z(n2492) );
  MUX U3092 ( .IN0(Y[5]), .IN1(n749), .SEL(n829), .F(n292) );
  XOR U3093 ( .A(n2614), .B(Y0[6]), .Z(n749) );
  XOR U3094 ( .A(n2615), .B(n2616), .Z(n2614) );
  AND U3095 ( .A(n841), .B(n2618), .Z(n2617) );
  XOR U3096 ( .A(n2612), .B(n2616), .Z(n2618) );
  XOR U3097 ( .A(n2611), .B(n2616), .Z(n2612) );
  XNOR U3098 ( .A(n2619), .B(n2542), .Z(n2537) );
  XNOR U3099 ( .A(n2510), .B(n2509), .Z(n2542) );
  XOR U3100 ( .A(n2620), .B(n2514), .Z(n2509) );
  XNOR U3101 ( .A(n2505), .B(n2507), .Z(n2514) );
  NAND U3102 ( .A(n2288), .B(n1021), .Z(n2507) );
  XNOR U3103 ( .A(n2503), .B(n2621), .Z(n2505) );
  ANDN U3104 ( .A(n2293), .B(n1023), .Z(n2621) );
  XNOR U3105 ( .A(n2513), .B(n2508), .Z(n2620) );
  XOR U3106 ( .A(n2628), .B(n2520), .Z(n2513) );
  XNOR U3107 ( .A(n2518), .B(n2629), .Z(n2520) );
  ANDN U3108 ( .A(n2523), .B(n939), .Z(n2629) );
  XOR U3109 ( .A(n2630), .B(n2631), .Z(n2518) );
  AND U3110 ( .A(n2632), .B(n2633), .Z(n2631) );
  XNOR U3111 ( .A(n2634), .B(n2630), .Z(n2633) );
  AND U3112 ( .A(n2516), .B(n937), .Z(n2522) );
  XNOR U3113 ( .A(n2531), .B(n2530), .Z(n2510) );
  XOR U3114 ( .A(n2638), .B(n2527), .Z(n2530) );
  XNOR U3115 ( .A(n2526), .B(n2639), .Z(n2527) );
  ANDN U3116 ( .A(n2094), .B(n1109), .Z(n2639) );
  AND U3117 ( .A(n2087), .B(n1107), .Z(n2528) );
  XNOR U3118 ( .A(n2534), .B(n2535), .Z(n2531) );
  NAND U3119 ( .A(n1892), .B(n1230), .Z(n2535) );
  XNOR U3120 ( .A(n2533), .B(n2646), .Z(n2534) );
  ANDN U3121 ( .A(n1897), .B(n1232), .Z(n2646) );
  XNOR U3122 ( .A(n2541), .B(n2536), .Z(n2619) );
  XOR U3123 ( .A(n2540), .B(n2653), .Z(n2541) );
  AND U3124 ( .A(n2544), .B(n2654), .Z(n2653) );
  AND U3125 ( .A(n2655), .B(n2656), .Z(n2654) );
  NANDN U3126 ( .B(n2657), .A(n876), .Z(n2656) );
  NAND U3127 ( .A(n2658), .B(n2659), .Z(n2655) );
  ANDN U3128 ( .A(n2546), .B(n2545), .Z(n2544) );
  ANDN U3129 ( .A(n2660), .B(n2661), .Z(n2545) );
  OR U3130 ( .A(n2662), .B(n2663), .Z(n2546) );
  XNOR U3131 ( .A(n2562), .B(n2561), .Z(n2538) );
  XOR U3132 ( .A(n2667), .B(n2570), .Z(n2561) );
  XNOR U3133 ( .A(n2555), .B(n2554), .Z(n2570) );
  XOR U3134 ( .A(n2668), .B(n2551), .Z(n2554) );
  XNOR U3135 ( .A(n2550), .B(n2669), .Z(n2551) );
  ANDN U3136 ( .A(n1386), .B(n1684), .Z(n2669) );
  AND U3137 ( .A(n1682), .B(n1323), .Z(n2552) );
  XNOR U3138 ( .A(n2558), .B(n2559), .Z(n2555) );
  NANDN U3139 ( .B(n1188), .A(n1870), .Z(n2559) );
  XNOR U3140 ( .A(n2557), .B(n2676), .Z(n2558) );
  ANDN U3141 ( .A(n1258), .B(n1872), .Z(n2676) );
  XNOR U3142 ( .A(n2569), .B(n2560), .Z(n2667) );
  XOR U3143 ( .A(n2683), .B(n2578), .Z(n2569) );
  XNOR U3144 ( .A(n2566), .B(n2567), .Z(n2578) );
  NAND U3145 ( .A(n1517), .B(n1557), .Z(n2567) );
  XNOR U3146 ( .A(n2565), .B(n2684), .Z(n2566) );
  ANDN U3147 ( .A(n1564), .B(n1519), .Z(n2684) );
  XNOR U3148 ( .A(n2577), .B(n2568), .Z(n2683) );
  XOR U3149 ( .A(n2691), .B(n2574), .Z(n2577) );
  XNOR U3150 ( .A(n2573), .B(n2692), .Z(n2574) );
  ANDN U3151 ( .A(n1748), .B(n1367), .Z(n2692) );
  AND U3152 ( .A(n1365), .B(n1741), .Z(n2575) );
  XNOR U3153 ( .A(n2586), .B(n2585), .Z(n2562) );
  XOR U3154 ( .A(n2699), .B(n2594), .Z(n2585) );
  XNOR U3155 ( .A(n2582), .B(n2583), .Z(n2594) );
  NANDN U3156 ( .B(n1001), .A(n2269), .Z(n2583) );
  XNOR U3157 ( .A(n2581), .B(n2700), .Z(n2582) );
  ANDN U3158 ( .A(n1042), .B(n2271), .Z(n2700) );
  XNOR U3159 ( .A(n2593), .B(n2584), .Z(n2699) );
  XOR U3160 ( .A(n2707), .B(n2590), .Z(n2593) );
  XNOR U3161 ( .A(n2589), .B(n2708), .Z(n2590) );
  ANDN U3162 ( .A(n1149), .B(n2064), .Z(n2708) );
  AND U3163 ( .A(n2062), .B(n1095), .Z(n2591) );
  XOR U3164 ( .A(n2602), .B(n2601), .Z(n2586) );
  XOR U3165 ( .A(n2715), .B(n2598), .Z(n2601) );
  XNOR U3166 ( .A(n2597), .B(n2716), .Z(n2598) );
  ANDN U3167 ( .A(n974), .B(n2486), .Z(n2716) );
  AND U3168 ( .A(n2484), .B(n933), .Z(n2599) );
  XOR U3169 ( .A(n2609), .B(n2608), .Z(n2602) );
  NAND U3170 ( .A(n2723), .B(n877), .Z(n2608) );
  XOR U3171 ( .A(n2607), .B(n2724), .Z(n2609) );
  ANDN U3172 ( .A(n908), .B(n2725), .Z(n2724) );
  ANDN U3173 ( .A(n2726), .B(n2727), .Z(n2607) );
  NAND U3174 ( .A(n2728), .B(n2729), .Z(n2726) );
  IV U3175 ( .A(n2610), .Z(n2611) );
  MUX U3176 ( .IN0(Y[4]), .IN1(n746), .SEL(n829), .F(n291) );
  XOR U3177 ( .A(n2734), .B(Y0[5]), .Z(n746) );
  XOR U3178 ( .A(n2735), .B(n2736), .Z(n2734) );
  AND U3179 ( .A(n841), .B(n2738), .Z(n2737) );
  XOR U3180 ( .A(n2732), .B(n2736), .Z(n2738) );
  XOR U3181 ( .A(n2731), .B(n2736), .Z(n2732) );
  XNOR U3182 ( .A(n2739), .B(n2666), .Z(n2651) );
  XNOR U3183 ( .A(n2627), .B(n2626), .Z(n2666) );
  XOR U3184 ( .A(n2740), .B(n2637), .Z(n2626) );
  XNOR U3185 ( .A(n2623), .B(n2624), .Z(n2637) );
  NAND U3186 ( .A(n2288), .B(n1065), .Z(n2624) );
  XNOR U3187 ( .A(n2622), .B(n2741), .Z(n2623) );
  ANDN U3188 ( .A(n2293), .B(n1067), .Z(n2741) );
  XNOR U3189 ( .A(n2636), .B(n2625), .Z(n2740) );
  XOR U3190 ( .A(n2748), .B(n2632), .Z(n2636) );
  XNOR U3191 ( .A(n2630), .B(n2749), .Z(n2632) );
  ANDN U3192 ( .A(n2523), .B(n983), .Z(n2749) );
  XOR U3193 ( .A(n2750), .B(n2751), .Z(n2630) );
  AND U3194 ( .A(n2752), .B(n2753), .Z(n2751) );
  XNOR U3195 ( .A(n2754), .B(n2750), .Z(n2753) );
  AND U3196 ( .A(n2516), .B(n981), .Z(n2634) );
  XNOR U3197 ( .A(n2645), .B(n2644), .Z(n2627) );
  XOR U3198 ( .A(n2758), .B(n2641), .Z(n2644) );
  XNOR U3199 ( .A(n2640), .B(n2759), .Z(n2641) );
  ANDN U3200 ( .A(n2094), .B(n1168), .Z(n2759) );
  AND U3201 ( .A(n2087), .B(n1166), .Z(n2642) );
  XNOR U3202 ( .A(n2648), .B(n2649), .Z(n2645) );
  NAND U3203 ( .A(n1892), .B(n1298), .Z(n2649) );
  XNOR U3204 ( .A(n2647), .B(n2766), .Z(n2648) );
  ANDN U3205 ( .A(n1897), .B(n1300), .Z(n2766) );
  XOR U3206 ( .A(n2665), .B(n2650), .Z(n2739) );
  XOR U3207 ( .A(n2773), .B(n2658), .Z(n2665) );
  XOR U3208 ( .A(n2777), .B(n2663), .Z(n2661) );
  NAND U3209 ( .A(n2778), .B(n906), .Z(n2663) );
  NAND U3210 ( .A(n2779), .B(n2662), .Z(n2777) );
  NANDN U3211 ( .B(n909), .A(n2783), .Z(n2779) );
  ANDN U3212 ( .A(n2784), .B(n2785), .Z(n2659) );
  XNOR U3213 ( .A(n2682), .B(n2681), .Z(n2652) );
  XOR U3214 ( .A(n2789), .B(n2690), .Z(n2681) );
  XNOR U3215 ( .A(n2675), .B(n2674), .Z(n2690) );
  XOR U3216 ( .A(n2790), .B(n2671), .Z(n2674) );
  XNOR U3217 ( .A(n2670), .B(n2791), .Z(n2671) );
  ANDN U3218 ( .A(n1386), .B(n1775), .Z(n2791) );
  AND U3219 ( .A(n1773), .B(n1323), .Z(n2672) );
  XNOR U3220 ( .A(n2678), .B(n2679), .Z(n2675) );
  NANDN U3221 ( .B(n1188), .A(n1966), .Z(n2679) );
  XNOR U3222 ( .A(n2677), .B(n2798), .Z(n2678) );
  ANDN U3223 ( .A(n1258), .B(n1968), .Z(n2798) );
  XNOR U3224 ( .A(n2689), .B(n2680), .Z(n2789) );
  XOR U3225 ( .A(n2805), .B(n2698), .Z(n2689) );
  XNOR U3226 ( .A(n2686), .B(n2687), .Z(n2698) );
  NAND U3227 ( .A(n1598), .B(n1557), .Z(n2687) );
  XNOR U3228 ( .A(n2685), .B(n2806), .Z(n2686) );
  ANDN U3229 ( .A(n1564), .B(n1600), .Z(n2806) );
  XNOR U3230 ( .A(n2697), .B(n2688), .Z(n2805) );
  XOR U3231 ( .A(n2813), .B(n2694), .Z(n2697) );
  XNOR U3232 ( .A(n2693), .B(n2814), .Z(n2694) );
  ANDN U3233 ( .A(n1748), .B(n1441), .Z(n2814) );
  AND U3234 ( .A(n1439), .B(n1741), .Z(n2695) );
  XNOR U3235 ( .A(n2706), .B(n2705), .Z(n2682) );
  XOR U3236 ( .A(n2821), .B(n2714), .Z(n2705) );
  XNOR U3237 ( .A(n2702), .B(n2703), .Z(n2714) );
  NANDN U3238 ( .B(n1001), .A(n2376), .Z(n2703) );
  XNOR U3239 ( .A(n2701), .B(n2822), .Z(n2702) );
  ANDN U3240 ( .A(n1042), .B(n2378), .Z(n2822) );
  XNOR U3241 ( .A(n2713), .B(n2704), .Z(n2821) );
  XOR U3242 ( .A(n2829), .B(n2710), .Z(n2713) );
  XNOR U3243 ( .A(n2709), .B(n2830), .Z(n2710) );
  ANDN U3244 ( .A(n1149), .B(n2165), .Z(n2830) );
  AND U3245 ( .A(n2163), .B(n1095), .Z(n2711) );
  XOR U3246 ( .A(n2722), .B(n2721), .Z(n2706) );
  XOR U3247 ( .A(n2837), .B(n2718), .Z(n2721) );
  XNOR U3248 ( .A(n2717), .B(n2838), .Z(n2718) );
  ANDN U3249 ( .A(n974), .B(n2605), .Z(n2838) );
  AND U3250 ( .A(n2603), .B(n933), .Z(n2719) );
  XOR U3251 ( .A(n2729), .B(n2728), .Z(n2722) );
  NAND U3252 ( .A(n2845), .B(n877), .Z(n2728) );
  XNOR U3253 ( .A(n2727), .B(n2846), .Z(n2729) );
  ANDN U3254 ( .A(n908), .B(n2847), .Z(n2846) );
  NAND U3255 ( .A(n2848), .B(n2849), .Z(n2727) );
  NAND U3256 ( .A(n2850), .B(n2851), .Z(n2848) );
  IV U3257 ( .A(n2730), .Z(n2731) );
  MUX U3258 ( .IN0(Y[3]), .IN1(n743), .SEL(n829), .F(n290) );
  XNOR U3259 ( .A(n2855), .B(Y0[4]), .Z(n743) );
  XNOR U3260 ( .A(n2857), .B(n2858), .Z(n2855) );
  XOR U3261 ( .A(n2856), .B(n2859), .Z(n2857) );
  AND U3262 ( .A(n841), .B(n2860), .Z(n2859) );
  XNOR U3263 ( .A(n2853), .B(n2858), .Z(n2860) );
  XOR U3264 ( .A(n2858), .B(n2852), .Z(n2853) );
  NOR U3265 ( .A(n2861), .B(n2862), .Z(n2852) );
  XNOR U3266 ( .A(n2863), .B(n2788), .Z(n2771) );
  XNOR U3267 ( .A(n2747), .B(n2746), .Z(n2788) );
  XOR U3268 ( .A(n2864), .B(n2757), .Z(n2746) );
  XNOR U3269 ( .A(n2743), .B(n2744), .Z(n2757) );
  NAND U3270 ( .A(n2288), .B(n1107), .Z(n2744) );
  XNOR U3271 ( .A(n2742), .B(n2865), .Z(n2743) );
  ANDN U3272 ( .A(n2293), .B(n1109), .Z(n2865) );
  XNOR U3273 ( .A(n2756), .B(n2745), .Z(n2864) );
  XOR U3274 ( .A(n2872), .B(n2752), .Z(n2756) );
  XNOR U3275 ( .A(n2750), .B(n2873), .Z(n2752) );
  ANDN U3276 ( .A(n2523), .B(n1023), .Z(n2873) );
  AND U3277 ( .A(n2516), .B(n1021), .Z(n2754) );
  XNOR U3278 ( .A(n2765), .B(n2764), .Z(n2747) );
  XOR U3279 ( .A(n2880), .B(n2761), .Z(n2764) );
  XNOR U3280 ( .A(n2760), .B(n2881), .Z(n2761) );
  ANDN U3281 ( .A(n2094), .B(n1232), .Z(n2881) );
  AND U3282 ( .A(n2087), .B(n1230), .Z(n2762) );
  XNOR U3283 ( .A(n2768), .B(n2769), .Z(n2765) );
  NAND U3284 ( .A(n1892), .B(n1365), .Z(n2769) );
  XNOR U3285 ( .A(n2767), .B(n2888), .Z(n2768) );
  ANDN U3286 ( .A(n1897), .B(n1367), .Z(n2888) );
  XNOR U3287 ( .A(n2787), .B(n2770), .Z(n2863) );
  XOR U3288 ( .A(n2895), .B(n2785), .Z(n2787) );
  XOR U3289 ( .A(n2776), .B(n2775), .Z(n2785) );
  XNOR U3290 ( .A(n2774), .B(n2896), .Z(n2775) );
  AND U3291 ( .A(n2897), .B(n2898), .Z(n2896) );
  NANDN U3292 ( .B(n2899), .A(n876), .Z(n2898) );
  NANDN U3293 ( .B(n2900), .A(n2901), .Z(n2897) );
  XNOR U3294 ( .A(n2781), .B(n2782), .Z(n2776) );
  NAND U3295 ( .A(n2778), .B(n937), .Z(n2782) );
  XNOR U3296 ( .A(n2780), .B(n2905), .Z(n2781) );
  ANDN U3297 ( .A(n2783), .B(n939), .Z(n2905) );
  NOR U3298 ( .A(n2909), .B(n2910), .Z(n2784) );
  XNOR U3299 ( .A(n2804), .B(n2803), .Z(n2772) );
  XOR U3300 ( .A(n2914), .B(n2812), .Z(n2803) );
  XNOR U3301 ( .A(n2797), .B(n2796), .Z(n2812) );
  XOR U3302 ( .A(n2915), .B(n2793), .Z(n2796) );
  XNOR U3303 ( .A(n2792), .B(n2916), .Z(n2793) );
  ANDN U3304 ( .A(n1386), .B(n1872), .Z(n2916) );
  AND U3305 ( .A(n1870), .B(n1323), .Z(n2794) );
  XNOR U3306 ( .A(n2800), .B(n2801), .Z(n2797) );
  NANDN U3307 ( .B(n1188), .A(n2062), .Z(n2801) );
  XNOR U3308 ( .A(n2799), .B(n2923), .Z(n2800) );
  ANDN U3309 ( .A(n1258), .B(n2064), .Z(n2923) );
  XNOR U3310 ( .A(n2811), .B(n2802), .Z(n2914) );
  XOR U3311 ( .A(n2930), .B(n2820), .Z(n2811) );
  XNOR U3312 ( .A(n2808), .B(n2809), .Z(n2820) );
  NAND U3313 ( .A(n1682), .B(n1557), .Z(n2809) );
  XNOR U3314 ( .A(n2807), .B(n2931), .Z(n2808) );
  ANDN U3315 ( .A(n1564), .B(n1684), .Z(n2931) );
  XNOR U3316 ( .A(n2819), .B(n2810), .Z(n2930) );
  XOR U3317 ( .A(n2938), .B(n2816), .Z(n2819) );
  XNOR U3318 ( .A(n2815), .B(n2939), .Z(n2816) );
  ANDN U3319 ( .A(n1748), .B(n1519), .Z(n2939) );
  AND U3320 ( .A(n1517), .B(n1741), .Z(n2817) );
  XNOR U3321 ( .A(n2828), .B(n2827), .Z(n2804) );
  XOR U3322 ( .A(n2946), .B(n2836), .Z(n2827) );
  XNOR U3323 ( .A(n2824), .B(n2825), .Z(n2836) );
  NANDN U3324 ( .B(n1001), .A(n2484), .Z(n2825) );
  XNOR U3325 ( .A(n2823), .B(n2947), .Z(n2824) );
  ANDN U3326 ( .A(n1042), .B(n2486), .Z(n2947) );
  XNOR U3327 ( .A(n2835), .B(n2826), .Z(n2946) );
  XOR U3328 ( .A(n2954), .B(n2832), .Z(n2835) );
  XNOR U3329 ( .A(n2831), .B(n2955), .Z(n2832) );
  ANDN U3330 ( .A(n1149), .B(n2271), .Z(n2955) );
  AND U3331 ( .A(n2269), .B(n1095), .Z(n2833) );
  XOR U3332 ( .A(n2844), .B(n2843), .Z(n2828) );
  XOR U3333 ( .A(n2962), .B(n2840), .Z(n2843) );
  XNOR U3334 ( .A(n2839), .B(n2963), .Z(n2840) );
  ANDN U3335 ( .A(n974), .B(n2725), .Z(n2963) );
  AND U3336 ( .A(n2723), .B(n933), .Z(n2841) );
  XOR U3337 ( .A(n2851), .B(n2850), .Z(n2844) );
  NAND U3338 ( .A(n2970), .B(n877), .Z(n2850) );
  XOR U3339 ( .A(n2849), .B(n2971), .Z(n2851) );
  ANDN U3340 ( .A(n908), .B(n2972), .Z(n2971) );
  ANDN U3341 ( .A(n2973), .B(n2974), .Z(n2849) );
  NAND U3342 ( .A(n2975), .B(n2976), .Z(n2973) );
  IV U3343 ( .A(n2854), .Z(n2856) );
  MUX U3344 ( .IN0(Y[2]), .IN1(n740), .SEL(n829), .F(n289) );
  IV U3345 ( .A(n2980), .Z(n829) );
  XNOR U3346 ( .A(n2978), .B(Y0[3]), .Z(n740) );
  XNOR U3347 ( .A(n2981), .B(n2982), .Z(n2978) );
  XOR U3348 ( .A(n2979), .B(n2983), .Z(n2981) );
  AND U3349 ( .A(n841), .B(n2984), .Z(n2983) );
  XNOR U3350 ( .A(n2862), .B(n2982), .Z(n2984) );
  NANDN U3351 ( .B(n2985), .A(n2986), .Z(n2861) );
  XNOR U3352 ( .A(n2987), .B(n2913), .Z(n2893) );
  XNOR U3353 ( .A(n2871), .B(n2870), .Z(n2913) );
  XOR U3354 ( .A(n2988), .B(n2879), .Z(n2870) );
  XNOR U3355 ( .A(n2867), .B(n2868), .Z(n2879) );
  NAND U3356 ( .A(n2288), .B(n1166), .Z(n2868) );
  XNOR U3357 ( .A(n2866), .B(n2989), .Z(n2867) );
  ANDN U3358 ( .A(n2293), .B(n1168), .Z(n2989) );
  XNOR U3359 ( .A(n2878), .B(n2869), .Z(n2988) );
  XOR U3360 ( .A(n2996), .B(n2875), .Z(n2878) );
  XNOR U3361 ( .A(n2874), .B(n2997), .Z(n2875) );
  ANDN U3362 ( .A(n2523), .B(n1067), .Z(n2997) );
  AND U3363 ( .A(n2516), .B(n1065), .Z(n2876) );
  XNOR U3364 ( .A(n2887), .B(n2886), .Z(n2871) );
  XOR U3365 ( .A(n3004), .B(n2883), .Z(n2886) );
  XNOR U3366 ( .A(n2882), .B(n3005), .Z(n2883) );
  ANDN U3367 ( .A(n2094), .B(n1300), .Z(n3005) );
  AND U3368 ( .A(n2087), .B(n1298), .Z(n2884) );
  XNOR U3369 ( .A(n2890), .B(n2891), .Z(n2887) );
  NAND U3370 ( .A(n1892), .B(n1439), .Z(n2891) );
  XNOR U3371 ( .A(n2889), .B(n3012), .Z(n2890) );
  ANDN U3372 ( .A(n1897), .B(n1441), .Z(n3012) );
  XNOR U3373 ( .A(n2912), .B(n2892), .Z(n2987) );
  XOR U3374 ( .A(n3019), .B(n2910), .Z(n2912) );
  XOR U3375 ( .A(n2904), .B(n2903), .Z(n2910) );
  XOR U3376 ( .A(n3024), .B(n2901), .Z(n3020) );
  AND U3377 ( .A(n3025), .B(n906), .Z(n2901) );
  NAND U3378 ( .A(n3026), .B(n2900), .Z(n3024) );
  XOR U3379 ( .A(n3027), .B(n3028), .Z(n2900) );
  AND U3380 ( .A(n3029), .B(n3030), .Z(n3028) );
  XNOR U3381 ( .A(n3031), .B(n3027), .Z(n3030) );
  NANDN U3382 ( .B(n909), .A(n3032), .Z(n3026) );
  XNOR U3383 ( .A(n2907), .B(n2908), .Z(n2904) );
  NAND U3384 ( .A(n2778), .B(n981), .Z(n2908) );
  XNOR U3385 ( .A(n2906), .B(n3033), .Z(n2907) );
  ANDN U3386 ( .A(n2783), .B(n983), .Z(n3033) );
  XOR U3387 ( .A(n3034), .B(n3035), .Z(n2906) );
  AND U3388 ( .A(n3036), .B(n3037), .Z(n3035) );
  XOR U3389 ( .A(n3038), .B(n3034), .Z(n3037) );
  XNOR U3390 ( .A(n2909), .B(n2911), .Z(n3019) );
  XNOR U3391 ( .A(n3042), .B(n3045), .Z(n3044) );
  XNOR U3392 ( .A(n2929), .B(n2928), .Z(n2894) );
  XOR U3393 ( .A(n3046), .B(n2937), .Z(n2928) );
  XNOR U3394 ( .A(n2922), .B(n2921), .Z(n2937) );
  XOR U3395 ( .A(n3047), .B(n2918), .Z(n2921) );
  XNOR U3396 ( .A(n2917), .B(n3048), .Z(n2918) );
  ANDN U3397 ( .A(n1386), .B(n1968), .Z(n3048) );
  AND U3398 ( .A(n1966), .B(n1323), .Z(n2919) );
  XNOR U3399 ( .A(n2925), .B(n2926), .Z(n2922) );
  NANDN U3400 ( .B(n1188), .A(n2163), .Z(n2926) );
  XNOR U3401 ( .A(n2924), .B(n3055), .Z(n2925) );
  ANDN U3402 ( .A(n1258), .B(n2165), .Z(n3055) );
  XNOR U3403 ( .A(n2936), .B(n2927), .Z(n3046) );
  XOR U3404 ( .A(n3062), .B(n2945), .Z(n2936) );
  XNOR U3405 ( .A(n2933), .B(n2934), .Z(n2945) );
  NAND U3406 ( .A(n1773), .B(n1557), .Z(n2934) );
  XNOR U3407 ( .A(n2932), .B(n3063), .Z(n2933) );
  ANDN U3408 ( .A(n1564), .B(n1775), .Z(n3063) );
  XNOR U3409 ( .A(n2944), .B(n2935), .Z(n3062) );
  XOR U3410 ( .A(n3070), .B(n2941), .Z(n2944) );
  XNOR U3411 ( .A(n2940), .B(n3071), .Z(n2941) );
  ANDN U3412 ( .A(n1748), .B(n1600), .Z(n3071) );
  AND U3413 ( .A(n1598), .B(n1741), .Z(n2942) );
  XNOR U3414 ( .A(n2953), .B(n2952), .Z(n2929) );
  XOR U3415 ( .A(n3078), .B(n2961), .Z(n2952) );
  XNOR U3416 ( .A(n2949), .B(n2950), .Z(n2961) );
  NANDN U3417 ( .B(n1001), .A(n2603), .Z(n2950) );
  XNOR U3418 ( .A(n2948), .B(n3079), .Z(n2949) );
  ANDN U3419 ( .A(n1042), .B(n2605), .Z(n3079) );
  XNOR U3420 ( .A(n2960), .B(n2951), .Z(n3078) );
  XOR U3421 ( .A(n3086), .B(n2957), .Z(n2960) );
  XNOR U3422 ( .A(n2956), .B(n3087), .Z(n2957) );
  ANDN U3423 ( .A(n1149), .B(n2378), .Z(n3087) );
  AND U3424 ( .A(n2376), .B(n1095), .Z(n2958) );
  XOR U3425 ( .A(n2969), .B(n2968), .Z(n2953) );
  XOR U3426 ( .A(n3094), .B(n2965), .Z(n2968) );
  XNOR U3427 ( .A(n2964), .B(n3095), .Z(n2965) );
  ANDN U3428 ( .A(n974), .B(n2847), .Z(n3095) );
  AND U3429 ( .A(n2845), .B(n933), .Z(n2966) );
  XOR U3430 ( .A(n2976), .B(n2975), .Z(n2969) );
  NAND U3431 ( .A(n3102), .B(n877), .Z(n2975) );
  XNOR U3432 ( .A(n2974), .B(n3103), .Z(n2976) );
  ANDN U3433 ( .A(n908), .B(n3104), .Z(n3103) );
  NAND U3434 ( .A(n3105), .B(n3106), .Z(n2974) );
  NAND U3435 ( .A(n3107), .B(n3108), .Z(n3105) );
  IV U3436 ( .A(n2977), .Z(n2979) );
  MUX U3437 ( .IN0(n737), .IN1(Y[1]), .SEL(n2980), .F(n288) );
  XNOR U3438 ( .A(n3110), .B(Y0[2]), .Z(n737) );
  XNOR U3439 ( .A(n3111), .B(n3112), .Z(n3110) );
  XNOR U3440 ( .A(n3109), .B(n3113), .Z(n3111) );
  AND U3441 ( .A(n841), .B(n3114), .Z(n3113) );
  XNOR U3442 ( .A(n2985), .B(n3112), .Z(n3114) );
  XOR U3443 ( .A(n3112), .B(n2986), .Z(n2985) );
  ANDN U3444 ( .A(n3115), .B(n3116), .Z(n2986) );
  XNOR U3445 ( .A(n3117), .B(n3041), .Z(n3017) );
  XNOR U3446 ( .A(n2995), .B(n2994), .Z(n3041) );
  XOR U3447 ( .A(n3118), .B(n3003), .Z(n2994) );
  XNOR U3448 ( .A(n2991), .B(n2992), .Z(n3003) );
  NAND U3449 ( .A(n2288), .B(n1230), .Z(n2992) );
  XNOR U3450 ( .A(n2990), .B(n3119), .Z(n2991) );
  ANDN U3451 ( .A(n2293), .B(n1232), .Z(n3119) );
  XNOR U3452 ( .A(n3002), .B(n2993), .Z(n3118) );
  XOR U3453 ( .A(n3126), .B(n2999), .Z(n3002) );
  XNOR U3454 ( .A(n2998), .B(n3127), .Z(n2999) );
  ANDN U3455 ( .A(n2523), .B(n1109), .Z(n3127) );
  AND U3456 ( .A(n2516), .B(n1107), .Z(n3000) );
  XNOR U3457 ( .A(n3011), .B(n3010), .Z(n2995) );
  XOR U3458 ( .A(n3134), .B(n3007), .Z(n3010) );
  XNOR U3459 ( .A(n3006), .B(n3135), .Z(n3007) );
  ANDN U3460 ( .A(n2094), .B(n1367), .Z(n3135) );
  AND U3461 ( .A(n2087), .B(n1365), .Z(n3008) );
  XNOR U3462 ( .A(n3014), .B(n3015), .Z(n3011) );
  NAND U3463 ( .A(n1892), .B(n1517), .Z(n3015) );
  XNOR U3464 ( .A(n3013), .B(n3142), .Z(n3014) );
  ANDN U3465 ( .A(n1897), .B(n1519), .Z(n3142) );
  XOR U3466 ( .A(n3040), .B(n3016), .Z(n3117) );
  XNOR U3467 ( .A(n3149), .B(n3045), .Z(n3040) );
  XNOR U3468 ( .A(n3023), .B(n3022), .Z(n3045) );
  XOR U3469 ( .A(n3150), .B(n3029), .Z(n3022) );
  XNOR U3470 ( .A(n3027), .B(n3151), .Z(n3029) );
  ANDN U3471 ( .A(n3032), .B(n939), .Z(n3151) );
  AND U3472 ( .A(n3025), .B(n937), .Z(n3031) );
  XNOR U3473 ( .A(n3036), .B(n3038), .Z(n3023) );
  NAND U3474 ( .A(n2778), .B(n1021), .Z(n3038) );
  XNOR U3475 ( .A(n3034), .B(n3158), .Z(n3036) );
  ANDN U3476 ( .A(n2783), .B(n1023), .Z(n3158) );
  XNOR U3477 ( .A(n3043), .B(n3039), .Z(n3149) );
  XOR U3478 ( .A(n3042), .B(n3165), .Z(n3043) );
  AND U3479 ( .A(n3166), .B(n3167), .Z(n3165) );
  NANDN U3480 ( .B(n3168), .A(n3169), .Z(n3167) );
  AND U3481 ( .A(n3170), .B(n3171), .Z(n3166) );
  NANDN U3482 ( .B(n3172), .A(n876), .Z(n3171) );
  OR U3483 ( .A(n3173), .B(n3174), .Z(n3170) );
  XNOR U3484 ( .A(n3061), .B(n3060), .Z(n3018) );
  XOR U3485 ( .A(n3178), .B(n3069), .Z(n3060) );
  XNOR U3486 ( .A(n3054), .B(n3053), .Z(n3069) );
  XOR U3487 ( .A(n3179), .B(n3050), .Z(n3053) );
  XNOR U3488 ( .A(n3049), .B(n3180), .Z(n3050) );
  ANDN U3489 ( .A(n1386), .B(n2064), .Z(n3180) );
  AND U3490 ( .A(n2062), .B(n1323), .Z(n3051) );
  XNOR U3491 ( .A(n3057), .B(n3058), .Z(n3054) );
  NANDN U3492 ( .B(n1188), .A(n2269), .Z(n3058) );
  XNOR U3493 ( .A(n3056), .B(n3187), .Z(n3057) );
  ANDN U3494 ( .A(n1258), .B(n2271), .Z(n3187) );
  XNOR U3495 ( .A(n3068), .B(n3059), .Z(n3178) );
  XOR U3496 ( .A(n3194), .B(n3077), .Z(n3068) );
  XNOR U3497 ( .A(n3065), .B(n3066), .Z(n3077) );
  NAND U3498 ( .A(n1870), .B(n1557), .Z(n3066) );
  XNOR U3499 ( .A(n3064), .B(n3195), .Z(n3065) );
  ANDN U3500 ( .A(n1564), .B(n1872), .Z(n3195) );
  XNOR U3501 ( .A(n3076), .B(n3067), .Z(n3194) );
  XOR U3502 ( .A(n3202), .B(n3073), .Z(n3076) );
  XNOR U3503 ( .A(n3072), .B(n3203), .Z(n3073) );
  ANDN U3504 ( .A(n1748), .B(n1684), .Z(n3203) );
  AND U3505 ( .A(n1682), .B(n1741), .Z(n3074) );
  XNOR U3506 ( .A(n3085), .B(n3084), .Z(n3061) );
  XOR U3507 ( .A(n3210), .B(n3093), .Z(n3084) );
  XNOR U3508 ( .A(n3081), .B(n3082), .Z(n3093) );
  NANDN U3509 ( .B(n1001), .A(n2723), .Z(n3082) );
  XNOR U3510 ( .A(n3080), .B(n3211), .Z(n3081) );
  ANDN U3511 ( .A(n1042), .B(n2725), .Z(n3211) );
  XNOR U3512 ( .A(n3092), .B(n3083), .Z(n3210) );
  XOR U3513 ( .A(n3218), .B(n3089), .Z(n3092) );
  XNOR U3514 ( .A(n3088), .B(n3219), .Z(n3089) );
  ANDN U3515 ( .A(n1149), .B(n2486), .Z(n3219) );
  AND U3516 ( .A(n2484), .B(n1095), .Z(n3090) );
  XOR U3517 ( .A(n3101), .B(n3100), .Z(n3085) );
  XOR U3518 ( .A(n3226), .B(n3097), .Z(n3100) );
  XNOR U3519 ( .A(n3096), .B(n3227), .Z(n3097) );
  ANDN U3520 ( .A(n974), .B(n2972), .Z(n3227) );
  AND U3521 ( .A(n2970), .B(n933), .Z(n3098) );
  XOR U3522 ( .A(n3108), .B(n3107), .Z(n3101) );
  NAND U3523 ( .A(n3234), .B(n877), .Z(n3107) );
  XOR U3524 ( .A(n3106), .B(n3235), .Z(n3108) );
  ANDN U3525 ( .A(n908), .B(n3236), .Z(n3235) );
  ANDN U3526 ( .A(n3237), .B(n3238), .Z(n3106) );
  NAND U3527 ( .A(n3239), .B(n3240), .Z(n3237) );
  MUX U3528 ( .IN0(n733), .IN1(Y[0]), .SEL(n2980), .F(n287) );
  NANDN U3529 ( .B(rst), .A(n828), .Z(n2980) );
  AND U3530 ( .A(n3243), .B(n3244), .Z(n828) );
  ANDN U3531 ( .A(n3245), .B(n[2]), .Z(n3244) );
  NOR U3532 ( .A(n[5]), .B(n[6]), .Z(n3245) );
  AND U3533 ( .A(n729), .B(n3246), .Z(n3243) );
  NOR U3534 ( .A(n[0]), .B(n[1]), .Z(n3246) );
  NOR U3535 ( .A(n[4]), .B(n[3]), .Z(n729) );
  XOR U3536 ( .A(n3242), .B(Y0[1]), .Z(n733) );
  XOR U3537 ( .A(n3247), .B(n3248), .Z(n3242) );
  XOR U3538 ( .A(n3249), .B(n3241), .Z(n3247) );
  NAND U3539 ( .A(n3250), .B(n841), .Z(n3249) );
  XOR U3540 ( .A(A[31]), .B(X[31]), .Z(n841) );
  XOR U3541 ( .A(n3115), .B(n3248), .Z(n3250) );
  XOR U3542 ( .A(n3116), .B(n3248), .Z(n3115) );
  XNOR U3543 ( .A(n3251), .B(n3164), .Z(n3147) );
  XNOR U3544 ( .A(n3125), .B(n3124), .Z(n3164) );
  XOR U3545 ( .A(n3252), .B(n3133), .Z(n3124) );
  XNOR U3546 ( .A(n3121), .B(n3122), .Z(n3133) );
  NAND U3547 ( .A(n2288), .B(n1298), .Z(n3122) );
  XNOR U3548 ( .A(n3120), .B(n3253), .Z(n3121) );
  ANDN U3549 ( .A(n2293), .B(n1300), .Z(n3253) );
  XNOR U3550 ( .A(n3132), .B(n3123), .Z(n3252) );
  XOR U3551 ( .A(n3260), .B(n3129), .Z(n3132) );
  XNOR U3552 ( .A(n3128), .B(n3261), .Z(n3129) );
  ANDN U3553 ( .A(n2523), .B(n1168), .Z(n3261) );
  AND U3554 ( .A(n2516), .B(n1166), .Z(n3130) );
  XNOR U3555 ( .A(n3141), .B(n3140), .Z(n3125) );
  XOR U3556 ( .A(n3268), .B(n3137), .Z(n3140) );
  XNOR U3557 ( .A(n3136), .B(n3269), .Z(n3137) );
  ANDN U3558 ( .A(n2094), .B(n1441), .Z(n3269) );
  AND U3559 ( .A(n2087), .B(n1439), .Z(n3138) );
  XNOR U3560 ( .A(n3144), .B(n3145), .Z(n3141) );
  NAND U3561 ( .A(n1892), .B(n1598), .Z(n3145) );
  XNOR U3562 ( .A(n3143), .B(n3276), .Z(n3144) );
  ANDN U3563 ( .A(n1897), .B(n1600), .Z(n3276) );
  XOR U3564 ( .A(n3163), .B(n3146), .Z(n3251) );
  XNOR U3565 ( .A(n3283), .B(n3177), .Z(n3163) );
  XNOR U3566 ( .A(n3157), .B(n3156), .Z(n3177) );
  XOR U3567 ( .A(n3284), .B(n3153), .Z(n3156) );
  XNOR U3568 ( .A(n3152), .B(n3285), .Z(n3153) );
  ANDN U3569 ( .A(n3032), .B(n983), .Z(n3285) );
  AND U3570 ( .A(n3025), .B(n981), .Z(n3154) );
  XNOR U3571 ( .A(n3160), .B(n3161), .Z(n3157) );
  NAND U3572 ( .A(n2778), .B(n1065), .Z(n3161) );
  XNOR U3573 ( .A(n3159), .B(n3292), .Z(n3160) );
  ANDN U3574 ( .A(n2783), .B(n1067), .Z(n3292) );
  XOR U3575 ( .A(n3176), .B(n3162), .Z(n3283) );
  XNOR U3576 ( .A(n3299), .B(n3173), .Z(n3176) );
  XNOR U3577 ( .A(n3300), .B(n3169), .Z(n3173) );
  AND U3578 ( .A(n3301), .B(n906), .Z(n3169) );
  NAND U3579 ( .A(n3302), .B(n3168), .Z(n3300) );
  NANDN U3580 ( .B(n909), .A(n3306), .Z(n3302) );
  XNOR U3581 ( .A(n3174), .B(n3175), .Z(n3299) );
  XNOR U3582 ( .A(n3310), .B(n3313), .Z(n3312) );
  XNOR U3583 ( .A(n3193), .B(n3192), .Z(n3148) );
  XOR U3584 ( .A(n3314), .B(n3201), .Z(n3192) );
  XNOR U3585 ( .A(n3186), .B(n3185), .Z(n3201) );
  XOR U3586 ( .A(n3315), .B(n3182), .Z(n3185) );
  XNOR U3587 ( .A(n3181), .B(n3316), .Z(n3182) );
  ANDN U3588 ( .A(n1386), .B(n2165), .Z(n3316) );
  AND U3589 ( .A(n2163), .B(n1323), .Z(n3183) );
  XNOR U3590 ( .A(n3189), .B(n3190), .Z(n3186) );
  NANDN U3591 ( .B(n1188), .A(n2376), .Z(n3190) );
  XNOR U3592 ( .A(n3188), .B(n3323), .Z(n3189) );
  ANDN U3593 ( .A(n1258), .B(n2378), .Z(n3323) );
  XNOR U3594 ( .A(n3200), .B(n3191), .Z(n3314) );
  XOR U3595 ( .A(n3330), .B(n3209), .Z(n3200) );
  XNOR U3596 ( .A(n3197), .B(n3198), .Z(n3209) );
  NAND U3597 ( .A(n1966), .B(n1557), .Z(n3198) );
  XNOR U3598 ( .A(n3196), .B(n3331), .Z(n3197) );
  ANDN U3599 ( .A(n1564), .B(n1968), .Z(n3331) );
  XNOR U3600 ( .A(n3208), .B(n3199), .Z(n3330) );
  XOR U3601 ( .A(n3338), .B(n3205), .Z(n3208) );
  XNOR U3602 ( .A(n3204), .B(n3339), .Z(n3205) );
  ANDN U3603 ( .A(n1748), .B(n1775), .Z(n3339) );
  AND U3604 ( .A(n1773), .B(n1741), .Z(n3206) );
  XNOR U3605 ( .A(n3217), .B(n3216), .Z(n3193) );
  XOR U3606 ( .A(n3346), .B(n3225), .Z(n3216) );
  XNOR U3607 ( .A(n3213), .B(n3214), .Z(n3225) );
  NANDN U3608 ( .B(n1001), .A(n2845), .Z(n3214) );
  XNOR U3609 ( .A(n3212), .B(n3347), .Z(n3213) );
  ANDN U3610 ( .A(n1042), .B(n2847), .Z(n3347) );
  XNOR U3611 ( .A(n3224), .B(n3215), .Z(n3346) );
  XOR U3612 ( .A(n3354), .B(n3221), .Z(n3224) );
  XNOR U3613 ( .A(n3220), .B(n3355), .Z(n3221) );
  ANDN U3614 ( .A(n1149), .B(n2605), .Z(n3355) );
  AND U3615 ( .A(n2603), .B(n1095), .Z(n3222) );
  XOR U3616 ( .A(n3233), .B(n3232), .Z(n3217) );
  XOR U3617 ( .A(n3362), .B(n3229), .Z(n3232) );
  XNOR U3618 ( .A(n3228), .B(n3363), .Z(n3229) );
  ANDN U3619 ( .A(n974), .B(n3104), .Z(n3363) );
  AND U3620 ( .A(n3102), .B(n933), .Z(n3230) );
  XOR U3621 ( .A(n3240), .B(n3239), .Z(n3233) );
  NAND U3622 ( .A(n3370), .B(n877), .Z(n3239) );
  XNOR U3623 ( .A(n3238), .B(n3371), .Z(n3240) );
  ANDN U3624 ( .A(n908), .B(n3372), .Z(n3371) );
  NAND U3625 ( .A(n3373), .B(n3374), .Z(n3238) );
  NAND U3626 ( .A(n3375), .B(n3376), .Z(n3373) );
  XNOR U3627 ( .A(n3377), .B(n3298), .Z(n3281) );
  XNOR U3628 ( .A(n3259), .B(n3258), .Z(n3298) );
  XOR U3629 ( .A(n3378), .B(n3267), .Z(n3258) );
  XNOR U3630 ( .A(n3255), .B(n3256), .Z(n3267) );
  NAND U3631 ( .A(n2288), .B(n1365), .Z(n3256) );
  XNOR U3632 ( .A(n3254), .B(n3379), .Z(n3255) );
  ANDN U3633 ( .A(n2293), .B(n1367), .Z(n3379) );
  XOR U3634 ( .A(n3380), .B(n3381), .Z(n3254) );
  AND U3635 ( .A(n3382), .B(n3383), .Z(n3381) );
  XOR U3636 ( .A(n3384), .B(n3380), .Z(n3383) );
  XNOR U3637 ( .A(n3266), .B(n3257), .Z(n3378) );
  XOR U3638 ( .A(n3388), .B(n3263), .Z(n3266) );
  XNOR U3639 ( .A(n3262), .B(n3389), .Z(n3263) );
  ANDN U3640 ( .A(n2523), .B(n1232), .Z(n3389) );
  XOR U3641 ( .A(n3390), .B(n3391), .Z(n3262) );
  AND U3642 ( .A(n3392), .B(n3393), .Z(n3391) );
  XNOR U3643 ( .A(n3394), .B(n3390), .Z(n3393) );
  AND U3644 ( .A(n2516), .B(n1230), .Z(n3264) );
  XNOR U3645 ( .A(n3275), .B(n3274), .Z(n3259) );
  XOR U3646 ( .A(n3398), .B(n3271), .Z(n3274) );
  XNOR U3647 ( .A(n3270), .B(n3399), .Z(n3271) );
  ANDN U3648 ( .A(n2094), .B(n1519), .Z(n3399) );
  AND U3649 ( .A(n2087), .B(n1517), .Z(n3272) );
  XNOR U3650 ( .A(n3278), .B(n3279), .Z(n3275) );
  NAND U3651 ( .A(n1892), .B(n1682), .Z(n3279) );
  XNOR U3652 ( .A(n3277), .B(n3406), .Z(n3278) );
  ANDN U3653 ( .A(n1897), .B(n1684), .Z(n3406) );
  XNOR U3654 ( .A(n3297), .B(n3280), .Z(n3377) );
  XNOR U3655 ( .A(n3410), .B(n3411), .Z(n3280) );
  XNOR U3656 ( .A(n3412), .B(n3309), .Z(n3297) );
  XNOR U3657 ( .A(n3291), .B(n3290), .Z(n3309) );
  XOR U3658 ( .A(n3413), .B(n3287), .Z(n3290) );
  XNOR U3659 ( .A(n3286), .B(n3414), .Z(n3287) );
  ANDN U3660 ( .A(n3032), .B(n1023), .Z(n3414) );
  XOR U3661 ( .A(n3415), .B(n3416), .Z(n3286) );
  AND U3662 ( .A(n3417), .B(n3418), .Z(n3416) );
  XNOR U3663 ( .A(n3419), .B(n3415), .Z(n3418) );
  AND U3664 ( .A(n3025), .B(n1021), .Z(n3288) );
  XNOR U3665 ( .A(n3294), .B(n3295), .Z(n3291) );
  NAND U3666 ( .A(n2778), .B(n1107), .Z(n3295) );
  XNOR U3667 ( .A(n3293), .B(n3423), .Z(n3294) );
  ANDN U3668 ( .A(n2783), .B(n1109), .Z(n3423) );
  XOR U3669 ( .A(n3424), .B(n3425), .Z(n3293) );
  AND U3670 ( .A(n3426), .B(n3427), .Z(n3425) );
  XOR U3671 ( .A(n3428), .B(n3424), .Z(n3427) );
  XNOR U3672 ( .A(n3308), .B(n3296), .Z(n3412) );
  XOR U3673 ( .A(n3429), .B(n3430), .Z(n3296) );
  AND U3674 ( .A(n3431), .B(n3432), .Z(n3430) );
  XOR U3675 ( .A(n3433), .B(n3434), .Z(n3432) );
  XNOR U3676 ( .A(n3435), .B(n3429), .Z(n3433) );
  XNOR U3677 ( .A(n3386), .B(n3436), .Z(n3431) );
  XNOR U3678 ( .A(n3429), .B(n3387), .Z(n3436) );
  XNOR U3679 ( .A(n3405), .B(n3404), .Z(n3387) );
  XOR U3680 ( .A(n3437), .B(n3401), .Z(n3404) );
  XNOR U3681 ( .A(n3400), .B(n3438), .Z(n3401) );
  ANDN U3682 ( .A(n2094), .B(n1600), .Z(n3438) );
  AND U3683 ( .A(n2087), .B(n1598), .Z(n3402) );
  XNOR U3684 ( .A(n3408), .B(n3409), .Z(n3405) );
  NAND U3685 ( .A(n1773), .B(n1892), .Z(n3409) );
  XNOR U3686 ( .A(n3407), .B(n3445), .Z(n3408) );
  ANDN U3687 ( .A(n1897), .B(n1775), .Z(n3445) );
  XOR U3688 ( .A(n3449), .B(n3397), .Z(n3386) );
  XNOR U3689 ( .A(n3382), .B(n3384), .Z(n3397) );
  NAND U3690 ( .A(n2288), .B(n1439), .Z(n3384) );
  XNOR U3691 ( .A(n3380), .B(n3450), .Z(n3382) );
  ANDN U3692 ( .A(n2293), .B(n1441), .Z(n3450) );
  XNOR U3693 ( .A(n3396), .B(n3385), .Z(n3449) );
  XOR U3694 ( .A(n3457), .B(n3392), .Z(n3396) );
  XNOR U3695 ( .A(n3390), .B(n3458), .Z(n3392) );
  ANDN U3696 ( .A(n2523), .B(n1300), .Z(n3458) );
  XOR U3697 ( .A(n3459), .B(n3460), .Z(n3390) );
  AND U3698 ( .A(n3461), .B(n3462), .Z(n3460) );
  XNOR U3699 ( .A(n3463), .B(n3459), .Z(n3462) );
  AND U3700 ( .A(n2516), .B(n1298), .Z(n3394) );
  XOR U3701 ( .A(n3467), .B(n3468), .Z(n3429) );
  AND U3702 ( .A(n3469), .B(n3470), .Z(n3468) );
  XOR U3703 ( .A(n3471), .B(n3472), .Z(n3470) );
  XOR U3704 ( .A(n3467), .B(n3473), .Z(n3472) );
  XNOR U3705 ( .A(n3455), .B(n3474), .Z(n3469) );
  XNOR U3706 ( .A(n3467), .B(n3456), .Z(n3474) );
  XNOR U3707 ( .A(n3444), .B(n3443), .Z(n3456) );
  XOR U3708 ( .A(n3475), .B(n3440), .Z(n3443) );
  XNOR U3709 ( .A(n3439), .B(n3476), .Z(n3440) );
  ANDN U3710 ( .A(n2094), .B(n1684), .Z(n3476) );
  XOR U3711 ( .A(n3477), .B(n3478), .Z(n3439) );
  AND U3712 ( .A(n3479), .B(n3480), .Z(n3478) );
  XNOR U3713 ( .A(n3481), .B(n3477), .Z(n3480) );
  AND U3714 ( .A(n2087), .B(n1682), .Z(n3441) );
  XNOR U3715 ( .A(n3447), .B(n3448), .Z(n3444) );
  NAND U3716 ( .A(n1870), .B(n1892), .Z(n3448) );
  XNOR U3717 ( .A(n3446), .B(n3485), .Z(n3447) );
  ANDN U3718 ( .A(n1897), .B(n1872), .Z(n3485) );
  XOR U3719 ( .A(n3486), .B(n3487), .Z(n3446) );
  AND U3720 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR U3721 ( .A(n3490), .B(n3486), .Z(n3489) );
  XOR U3722 ( .A(n3491), .B(n3466), .Z(n3455) );
  XNOR U3723 ( .A(n3452), .B(n3453), .Z(n3466) );
  NAND U3724 ( .A(n2288), .B(n1517), .Z(n3453) );
  XNOR U3725 ( .A(n3451), .B(n3492), .Z(n3452) );
  ANDN U3726 ( .A(n2293), .B(n1519), .Z(n3492) );
  XOR U3727 ( .A(n3493), .B(n3494), .Z(n3451) );
  AND U3728 ( .A(n3495), .B(n3496), .Z(n3494) );
  XOR U3729 ( .A(n3497), .B(n3493), .Z(n3496) );
  XNOR U3730 ( .A(n3465), .B(n3454), .Z(n3491) );
  XOR U3731 ( .A(n3501), .B(n3461), .Z(n3465) );
  XNOR U3732 ( .A(n3459), .B(n3502), .Z(n3461) );
  ANDN U3733 ( .A(n2523), .B(n1367), .Z(n3502) );
  XOR U3734 ( .A(n3503), .B(n3504), .Z(n3459) );
  AND U3735 ( .A(n3505), .B(n3506), .Z(n3504) );
  XNOR U3736 ( .A(n3507), .B(n3503), .Z(n3506) );
  XOR U3737 ( .A(n3508), .B(n3463), .Z(n3501) );
  AND U3738 ( .A(n2516), .B(n1365), .Z(n3463) );
  IV U3739 ( .A(n3464), .Z(n3508) );
  XOR U3740 ( .A(n3512), .B(n3513), .Z(n3467) );
  AND U3741 ( .A(n3514), .B(n3515), .Z(n3513) );
  XOR U3742 ( .A(n3516), .B(n3517), .Z(n3515) );
  XOR U3743 ( .A(n3512), .B(n3518), .Z(n3517) );
  XNOR U3744 ( .A(n3499), .B(n3519), .Z(n3514) );
  XNOR U3745 ( .A(n3512), .B(n3500), .Z(n3519) );
  XNOR U3746 ( .A(n3484), .B(n3483), .Z(n3500) );
  XOR U3747 ( .A(n3520), .B(n3479), .Z(n3483) );
  XNOR U3748 ( .A(n3477), .B(n3521), .Z(n3479) );
  ANDN U3749 ( .A(n2094), .B(n1775), .Z(n3521) );
  XOR U3750 ( .A(n3522), .B(n3523), .Z(n3477) );
  AND U3751 ( .A(n3524), .B(n3525), .Z(n3523) );
  XNOR U3752 ( .A(n3526), .B(n3522), .Z(n3525) );
  AND U3753 ( .A(n1773), .B(n2087), .Z(n3481) );
  XNOR U3754 ( .A(n3488), .B(n3490), .Z(n3484) );
  NAND U3755 ( .A(n1966), .B(n1892), .Z(n3490) );
  XNOR U3756 ( .A(n3486), .B(n3530), .Z(n3488) );
  ANDN U3757 ( .A(n1897), .B(n1968), .Z(n3530) );
  XOR U3758 ( .A(n3534), .B(n3511), .Z(n3499) );
  XNOR U3759 ( .A(n3495), .B(n3497), .Z(n3511) );
  NAND U3760 ( .A(n2288), .B(n1598), .Z(n3497) );
  XNOR U3761 ( .A(n3493), .B(n3535), .Z(n3495) );
  ANDN U3762 ( .A(n2293), .B(n1600), .Z(n3535) );
  XOR U3763 ( .A(n3536), .B(n3537), .Z(n3493) );
  AND U3764 ( .A(n3538), .B(n3539), .Z(n3537) );
  XOR U3765 ( .A(n3540), .B(n3536), .Z(n3539) );
  XNOR U3766 ( .A(n3510), .B(n3498), .Z(n3534) );
  XOR U3767 ( .A(n3544), .B(n3505), .Z(n3510) );
  XNOR U3768 ( .A(n3503), .B(n3545), .Z(n3505) );
  ANDN U3769 ( .A(n2523), .B(n1441), .Z(n3545) );
  XOR U3770 ( .A(n3546), .B(n3547), .Z(n3503) );
  AND U3771 ( .A(n3548), .B(n3549), .Z(n3547) );
  XNOR U3772 ( .A(n3550), .B(n3546), .Z(n3549) );
  AND U3773 ( .A(n2516), .B(n1439), .Z(n3507) );
  XOR U3774 ( .A(n3554), .B(n3555), .Z(n3512) );
  AND U3775 ( .A(n3556), .B(n3557), .Z(n3555) );
  XOR U3776 ( .A(n3558), .B(n3559), .Z(n3557) );
  XOR U3777 ( .A(n3554), .B(n3560), .Z(n3559) );
  XNOR U3778 ( .A(n3542), .B(n3561), .Z(n3556) );
  XNOR U3779 ( .A(n3554), .B(n3543), .Z(n3561) );
  XNOR U3780 ( .A(n3529), .B(n3528), .Z(n3543) );
  XOR U3781 ( .A(n3562), .B(n3524), .Z(n3528) );
  XNOR U3782 ( .A(n3522), .B(n3563), .Z(n3524) );
  ANDN U3783 ( .A(n2094), .B(n1872), .Z(n3563) );
  XOR U3784 ( .A(n3564), .B(n3565), .Z(n3522) );
  AND U3785 ( .A(n3566), .B(n3567), .Z(n3565) );
  XNOR U3786 ( .A(n3568), .B(n3564), .Z(n3567) );
  AND U3787 ( .A(n1870), .B(n2087), .Z(n3526) );
  XNOR U3788 ( .A(n3532), .B(n3533), .Z(n3529) );
  NAND U3789 ( .A(n2062), .B(n1892), .Z(n3533) );
  XNOR U3790 ( .A(n3531), .B(n3572), .Z(n3532) );
  ANDN U3791 ( .A(n1897), .B(n2064), .Z(n3572) );
  XOR U3792 ( .A(n3573), .B(n3574), .Z(n3531) );
  AND U3793 ( .A(n3575), .B(n3576), .Z(n3574) );
  XOR U3794 ( .A(n3577), .B(n3573), .Z(n3576) );
  XOR U3795 ( .A(n3578), .B(n3553), .Z(n3542) );
  XNOR U3796 ( .A(n3538), .B(n3540), .Z(n3553) );
  NAND U3797 ( .A(n2288), .B(n1682), .Z(n3540) );
  XNOR U3798 ( .A(n3536), .B(n3579), .Z(n3538) );
  ANDN U3799 ( .A(n2293), .B(n1684), .Z(n3579) );
  XNOR U3800 ( .A(n3552), .B(n3541), .Z(n3578) );
  XOR U3801 ( .A(n3586), .B(n3548), .Z(n3552) );
  XNOR U3802 ( .A(n3546), .B(n3587), .Z(n3548) );
  ANDN U3803 ( .A(n2523), .B(n1519), .Z(n3587) );
  XOR U3804 ( .A(n3588), .B(n3589), .Z(n3546) );
  AND U3805 ( .A(n3590), .B(n3591), .Z(n3589) );
  XNOR U3806 ( .A(n3592), .B(n3588), .Z(n3591) );
  XOR U3807 ( .A(n3593), .B(n3550), .Z(n3586) );
  AND U3808 ( .A(n2516), .B(n1517), .Z(n3550) );
  IV U3809 ( .A(n3551), .Z(n3593) );
  XOR U3810 ( .A(n3597), .B(n3598), .Z(n3554) );
  AND U3811 ( .A(n3599), .B(n3600), .Z(n3598) );
  XOR U3812 ( .A(n3601), .B(n3602), .Z(n3600) );
  XOR U3813 ( .A(n3597), .B(n3603), .Z(n3602) );
  XNOR U3814 ( .A(n3584), .B(n3604), .Z(n3599) );
  XNOR U3815 ( .A(n3597), .B(n3585), .Z(n3604) );
  XNOR U3816 ( .A(n3571), .B(n3570), .Z(n3585) );
  XOR U3817 ( .A(n3605), .B(n3566), .Z(n3570) );
  XNOR U3818 ( .A(n3564), .B(n3606), .Z(n3566) );
  ANDN U3819 ( .A(n2094), .B(n1968), .Z(n3606) );
  XOR U3820 ( .A(n3607), .B(n3608), .Z(n3564) );
  AND U3821 ( .A(n3609), .B(n3610), .Z(n3608) );
  XNOR U3822 ( .A(n3611), .B(n3607), .Z(n3610) );
  AND U3823 ( .A(n1966), .B(n2087), .Z(n3568) );
  XNOR U3824 ( .A(n3575), .B(n3577), .Z(n3571) );
  NAND U3825 ( .A(n2163), .B(n1892), .Z(n3577) );
  XNOR U3826 ( .A(n3573), .B(n3615), .Z(n3575) );
  ANDN U3827 ( .A(n1897), .B(n2165), .Z(n3615) );
  XOR U3828 ( .A(n3619), .B(n3596), .Z(n3584) );
  XNOR U3829 ( .A(n3581), .B(n3582), .Z(n3596) );
  NAND U3830 ( .A(n1773), .B(n2288), .Z(n3582) );
  XNOR U3831 ( .A(n3580), .B(n3620), .Z(n3581) );
  ANDN U3832 ( .A(n2293), .B(n1775), .Z(n3620) );
  XOR U3833 ( .A(n3621), .B(n3622), .Z(n3580) );
  AND U3834 ( .A(n3623), .B(n3624), .Z(n3622) );
  XOR U3835 ( .A(n3625), .B(n3621), .Z(n3624) );
  XNOR U3836 ( .A(n3595), .B(n3583), .Z(n3619) );
  XOR U3837 ( .A(n3629), .B(n3590), .Z(n3595) );
  XNOR U3838 ( .A(n3588), .B(n3630), .Z(n3590) );
  ANDN U3839 ( .A(n2523), .B(n1600), .Z(n3630) );
  XOR U3840 ( .A(n3631), .B(n3632), .Z(n3588) );
  AND U3841 ( .A(n3633), .B(n3634), .Z(n3632) );
  XNOR U3842 ( .A(n3635), .B(n3631), .Z(n3634) );
  AND U3843 ( .A(n2516), .B(n1598), .Z(n3592) );
  XOR U3844 ( .A(n3639), .B(n3640), .Z(n3597) );
  AND U3845 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U3846 ( .A(n3643), .B(n3644), .Z(n3642) );
  XOR U3847 ( .A(n3639), .B(n3645), .Z(n3644) );
  XNOR U3848 ( .A(n3627), .B(n3646), .Z(n3641) );
  XNOR U3849 ( .A(n3639), .B(n3628), .Z(n3646) );
  XNOR U3850 ( .A(n3614), .B(n3613), .Z(n3628) );
  XOR U3851 ( .A(n3647), .B(n3609), .Z(n3613) );
  XNOR U3852 ( .A(n3607), .B(n3648), .Z(n3609) );
  ANDN U3853 ( .A(n2094), .B(n2064), .Z(n3648) );
  XOR U3854 ( .A(n3649), .B(n3650), .Z(n3607) );
  AND U3855 ( .A(n3651), .B(n3652), .Z(n3650) );
  XNOR U3856 ( .A(n3653), .B(n3649), .Z(n3652) );
  XOR U3857 ( .A(n3654), .B(n3611), .Z(n3647) );
  AND U3858 ( .A(n2062), .B(n2087), .Z(n3611) );
  IV U3859 ( .A(n3612), .Z(n3654) );
  XNOR U3860 ( .A(n3617), .B(n3618), .Z(n3614) );
  NAND U3861 ( .A(n2269), .B(n1892), .Z(n3618) );
  XNOR U3862 ( .A(n3616), .B(n3658), .Z(n3617) );
  ANDN U3863 ( .A(n1897), .B(n2271), .Z(n3658) );
  XOR U3864 ( .A(n3659), .B(n3660), .Z(n3616) );
  AND U3865 ( .A(n3661), .B(n3662), .Z(n3660) );
  XOR U3866 ( .A(n3663), .B(n3659), .Z(n3662) );
  XOR U3867 ( .A(n3664), .B(n3638), .Z(n3627) );
  XNOR U3868 ( .A(n3623), .B(n3625), .Z(n3638) );
  NAND U3869 ( .A(n1870), .B(n2288), .Z(n3625) );
  XNOR U3870 ( .A(n3621), .B(n3665), .Z(n3623) );
  ANDN U3871 ( .A(n2293), .B(n1872), .Z(n3665) );
  XOR U3872 ( .A(n3666), .B(n3667), .Z(n3621) );
  AND U3873 ( .A(n3668), .B(n3669), .Z(n3667) );
  XOR U3874 ( .A(n3670), .B(n3666), .Z(n3669) );
  XNOR U3875 ( .A(n3637), .B(n3626), .Z(n3664) );
  XOR U3876 ( .A(n3674), .B(n3633), .Z(n3637) );
  XNOR U3877 ( .A(n3631), .B(n3675), .Z(n3633) );
  ANDN U3878 ( .A(n2523), .B(n1684), .Z(n3675) );
  XOR U3879 ( .A(n3676), .B(n3677), .Z(n3631) );
  AND U3880 ( .A(n3678), .B(n3679), .Z(n3677) );
  XNOR U3881 ( .A(n3680), .B(n3676), .Z(n3679) );
  XOR U3882 ( .A(n3681), .B(n3635), .Z(n3674) );
  AND U3883 ( .A(n2516), .B(n1682), .Z(n3635) );
  IV U3884 ( .A(n3636), .Z(n3681) );
  XOR U3885 ( .A(n3685), .B(n3686), .Z(n3639) );
  AND U3886 ( .A(n3687), .B(n3688), .Z(n3686) );
  XOR U3887 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR U3888 ( .A(n3685), .B(n3691), .Z(n3690) );
  XNOR U3889 ( .A(n3672), .B(n3692), .Z(n3687) );
  XNOR U3890 ( .A(n3685), .B(n3673), .Z(n3692) );
  XNOR U3891 ( .A(n3657), .B(n3656), .Z(n3673) );
  XOR U3892 ( .A(n3693), .B(n3651), .Z(n3656) );
  XNOR U3893 ( .A(n3649), .B(n3694), .Z(n3651) );
  ANDN U3894 ( .A(n2094), .B(n2165), .Z(n3694) );
  XOR U3895 ( .A(n3695), .B(n3696), .Z(n3649) );
  AND U3896 ( .A(n3697), .B(n3698), .Z(n3696) );
  XNOR U3897 ( .A(n3699), .B(n3695), .Z(n3698) );
  XOR U3898 ( .A(n3700), .B(n3653), .Z(n3693) );
  AND U3899 ( .A(n2163), .B(n2087), .Z(n3653) );
  IV U3900 ( .A(n3655), .Z(n3700) );
  XNOR U3901 ( .A(n3661), .B(n3663), .Z(n3657) );
  NAND U3902 ( .A(n2376), .B(n1892), .Z(n3663) );
  XNOR U3903 ( .A(n3659), .B(n3704), .Z(n3661) );
  ANDN U3904 ( .A(n1897), .B(n2378), .Z(n3704) );
  XOR U3905 ( .A(n3705), .B(n3706), .Z(n3659) );
  AND U3906 ( .A(n3707), .B(n3708), .Z(n3706) );
  XOR U3907 ( .A(n3709), .B(n3705), .Z(n3708) );
  XOR U3908 ( .A(n3710), .B(n3684), .Z(n3672) );
  XNOR U3909 ( .A(n3668), .B(n3670), .Z(n3684) );
  NAND U3910 ( .A(n1966), .B(n2288), .Z(n3670) );
  XNOR U3911 ( .A(n3666), .B(n3711), .Z(n3668) );
  ANDN U3912 ( .A(n2293), .B(n1968), .Z(n3711) );
  XNOR U3913 ( .A(n3683), .B(n3671), .Z(n3710) );
  XOR U3914 ( .A(n3718), .B(n3678), .Z(n3683) );
  XNOR U3915 ( .A(n3676), .B(n3719), .Z(n3678) );
  ANDN U3916 ( .A(n2523), .B(n1775), .Z(n3719) );
  XOR U3917 ( .A(n3720), .B(n3721), .Z(n3676) );
  AND U3918 ( .A(n3722), .B(n3723), .Z(n3721) );
  XNOR U3919 ( .A(n3724), .B(n3720), .Z(n3723) );
  XOR U3920 ( .A(n3725), .B(n3680), .Z(n3718) );
  AND U3921 ( .A(n1773), .B(n2516), .Z(n3680) );
  IV U3922 ( .A(n3682), .Z(n3725) );
  XOR U3923 ( .A(n3729), .B(n3730), .Z(n3685) );
  AND U3924 ( .A(n3731), .B(n3732), .Z(n3730) );
  XOR U3925 ( .A(n3733), .B(n3734), .Z(n3732) );
  XOR U3926 ( .A(n3729), .B(n3735), .Z(n3734) );
  XNOR U3927 ( .A(n3716), .B(n3736), .Z(n3731) );
  XNOR U3928 ( .A(n3729), .B(n3717), .Z(n3736) );
  XNOR U3929 ( .A(n3703), .B(n3702), .Z(n3717) );
  XOR U3930 ( .A(n3737), .B(n3697), .Z(n3702) );
  XNOR U3931 ( .A(n3695), .B(n3738), .Z(n3697) );
  ANDN U3932 ( .A(n2094), .B(n2271), .Z(n3738) );
  XOR U3933 ( .A(n3739), .B(n3740), .Z(n3695) );
  AND U3934 ( .A(n3741), .B(n3742), .Z(n3740) );
  XNOR U3935 ( .A(n3743), .B(n3739), .Z(n3742) );
  XOR U3936 ( .A(n3744), .B(n3699), .Z(n3737) );
  AND U3937 ( .A(n2269), .B(n2087), .Z(n3699) );
  IV U3938 ( .A(n3701), .Z(n3744) );
  XNOR U3939 ( .A(n3707), .B(n3709), .Z(n3703) );
  NAND U3940 ( .A(n2484), .B(n1892), .Z(n3709) );
  XNOR U3941 ( .A(n3705), .B(n3748), .Z(n3707) );
  ANDN U3942 ( .A(n1897), .B(n2486), .Z(n3748) );
  XOR U3943 ( .A(n3749), .B(n3750), .Z(n3705) );
  AND U3944 ( .A(n3751), .B(n3752), .Z(n3750) );
  XOR U3945 ( .A(n3753), .B(n3749), .Z(n3752) );
  XOR U3946 ( .A(n3754), .B(n3728), .Z(n3716) );
  XNOR U3947 ( .A(n3713), .B(n3714), .Z(n3728) );
  NAND U3948 ( .A(n2062), .B(n2288), .Z(n3714) );
  XNOR U3949 ( .A(n3712), .B(n3755), .Z(n3713) );
  ANDN U3950 ( .A(n2293), .B(n2064), .Z(n3755) );
  XOR U3951 ( .A(n3756), .B(n3757), .Z(n3712) );
  AND U3952 ( .A(n3758), .B(n3759), .Z(n3757) );
  XOR U3953 ( .A(n3760), .B(n3756), .Z(n3759) );
  XNOR U3954 ( .A(n3727), .B(n3715), .Z(n3754) );
  XOR U3955 ( .A(n3764), .B(n3722), .Z(n3727) );
  XNOR U3956 ( .A(n3720), .B(n3765), .Z(n3722) );
  ANDN U3957 ( .A(n2523), .B(n1872), .Z(n3765) );
  XOR U3958 ( .A(n3766), .B(n3767), .Z(n3720) );
  AND U3959 ( .A(n3768), .B(n3769), .Z(n3767) );
  XNOR U3960 ( .A(n3770), .B(n3766), .Z(n3769) );
  XOR U3961 ( .A(n3771), .B(n3724), .Z(n3764) );
  AND U3962 ( .A(n1870), .B(n2516), .Z(n3724) );
  IV U3963 ( .A(n3726), .Z(n3771) );
  XOR U3964 ( .A(n3775), .B(n3776), .Z(n3729) );
  AND U3965 ( .A(n3777), .B(n3778), .Z(n3776) );
  XOR U3966 ( .A(n3779), .B(n3780), .Z(n3778) );
  XOR U3967 ( .A(n3775), .B(n3781), .Z(n3780) );
  XNOR U3968 ( .A(n3762), .B(n3782), .Z(n3777) );
  XNOR U3969 ( .A(n3775), .B(n3763), .Z(n3782) );
  XNOR U3970 ( .A(n3747), .B(n3746), .Z(n3763) );
  XOR U3971 ( .A(n3783), .B(n3741), .Z(n3746) );
  XNOR U3972 ( .A(n3739), .B(n3784), .Z(n3741) );
  ANDN U3973 ( .A(n2094), .B(n2378), .Z(n3784) );
  XOR U3974 ( .A(n3785), .B(n3786), .Z(n3739) );
  AND U3975 ( .A(n3787), .B(n3788), .Z(n3786) );
  XNOR U3976 ( .A(n3789), .B(n3785), .Z(n3788) );
  XOR U3977 ( .A(n3790), .B(n3743), .Z(n3783) );
  AND U3978 ( .A(n2376), .B(n2087), .Z(n3743) );
  IV U3979 ( .A(n3745), .Z(n3790) );
  XNOR U3980 ( .A(n3751), .B(n3753), .Z(n3747) );
  NAND U3981 ( .A(n2603), .B(n1892), .Z(n3753) );
  XNOR U3982 ( .A(n3749), .B(n3794), .Z(n3751) );
  ANDN U3983 ( .A(n1897), .B(n2605), .Z(n3794) );
  XOR U3984 ( .A(n3795), .B(n3796), .Z(n3749) );
  AND U3985 ( .A(n3797), .B(n3798), .Z(n3796) );
  XOR U3986 ( .A(n3799), .B(n3795), .Z(n3798) );
  XOR U3987 ( .A(n3800), .B(n3774), .Z(n3762) );
  XNOR U3988 ( .A(n3758), .B(n3760), .Z(n3774) );
  NAND U3989 ( .A(n2163), .B(n2288), .Z(n3760) );
  XNOR U3990 ( .A(n3756), .B(n3801), .Z(n3758) );
  ANDN U3991 ( .A(n2293), .B(n2165), .Z(n3801) );
  XOR U3992 ( .A(n3802), .B(n3803), .Z(n3756) );
  AND U3993 ( .A(n3804), .B(n3805), .Z(n3803) );
  XOR U3994 ( .A(n3806), .B(n3802), .Z(n3805) );
  XNOR U3995 ( .A(n3773), .B(n3761), .Z(n3800) );
  XOR U3996 ( .A(n3810), .B(n3768), .Z(n3773) );
  XNOR U3997 ( .A(n3766), .B(n3811), .Z(n3768) );
  ANDN U3998 ( .A(n2523), .B(n1968), .Z(n3811) );
  XOR U3999 ( .A(n3812), .B(n3813), .Z(n3766) );
  AND U4000 ( .A(n3814), .B(n3815), .Z(n3813) );
  XNOR U4001 ( .A(n3816), .B(n3812), .Z(n3815) );
  XOR U4002 ( .A(n3817), .B(n3770), .Z(n3810) );
  AND U4003 ( .A(n1966), .B(n2516), .Z(n3770) );
  IV U4004 ( .A(n3772), .Z(n3817) );
  XOR U4005 ( .A(n3821), .B(n3822), .Z(n3775) );
  AND U4006 ( .A(n3823), .B(n3824), .Z(n3822) );
  XOR U4007 ( .A(n3825), .B(n3826), .Z(n3824) );
  XOR U4008 ( .A(n3821), .B(n3827), .Z(n3826) );
  XNOR U4009 ( .A(n3808), .B(n3828), .Z(n3823) );
  XNOR U4010 ( .A(n3821), .B(n3809), .Z(n3828) );
  XNOR U4011 ( .A(n3793), .B(n3792), .Z(n3809) );
  XOR U4012 ( .A(n3829), .B(n3787), .Z(n3792) );
  XNOR U4013 ( .A(n3785), .B(n3830), .Z(n3787) );
  ANDN U4014 ( .A(n2094), .B(n2486), .Z(n3830) );
  XOR U4015 ( .A(n3831), .B(n3832), .Z(n3785) );
  AND U4016 ( .A(n3833), .B(n3834), .Z(n3832) );
  XNOR U4017 ( .A(n3835), .B(n3831), .Z(n3834) );
  XOR U4018 ( .A(n3836), .B(n3789), .Z(n3829) );
  AND U4019 ( .A(n2484), .B(n2087), .Z(n3789) );
  IV U4020 ( .A(n3791), .Z(n3836) );
  XNOR U4021 ( .A(n3797), .B(n3799), .Z(n3793) );
  NAND U4022 ( .A(n2723), .B(n1892), .Z(n3799) );
  XNOR U4023 ( .A(n3795), .B(n3840), .Z(n3797) );
  ANDN U4024 ( .A(n1897), .B(n2725), .Z(n3840) );
  XOR U4025 ( .A(n3841), .B(n3842), .Z(n3795) );
  AND U4026 ( .A(n3843), .B(n3844), .Z(n3842) );
  XOR U4027 ( .A(n3845), .B(n3841), .Z(n3844) );
  XOR U4028 ( .A(n3846), .B(n3820), .Z(n3808) );
  XNOR U4029 ( .A(n3804), .B(n3806), .Z(n3820) );
  NAND U4030 ( .A(n2269), .B(n2288), .Z(n3806) );
  XNOR U4031 ( .A(n3802), .B(n3847), .Z(n3804) );
  ANDN U4032 ( .A(n2293), .B(n2271), .Z(n3847) );
  XOR U4033 ( .A(n3848), .B(n3849), .Z(n3802) );
  AND U4034 ( .A(n3850), .B(n3851), .Z(n3849) );
  XOR U4035 ( .A(n3852), .B(n3848), .Z(n3851) );
  XNOR U4036 ( .A(n3819), .B(n3807), .Z(n3846) );
  XOR U4037 ( .A(n3856), .B(n3814), .Z(n3819) );
  XNOR U4038 ( .A(n3812), .B(n3857), .Z(n3814) );
  ANDN U4039 ( .A(n2523), .B(n2064), .Z(n3857) );
  XOR U4040 ( .A(n3858), .B(n3859), .Z(n3812) );
  AND U4041 ( .A(n3860), .B(n3861), .Z(n3859) );
  XNOR U4042 ( .A(n3862), .B(n3858), .Z(n3861) );
  XOR U4043 ( .A(n3863), .B(n3816), .Z(n3856) );
  AND U4044 ( .A(n2062), .B(n2516), .Z(n3816) );
  IV U4045 ( .A(n3818), .Z(n3863) );
  XOR U4046 ( .A(n3867), .B(n3868), .Z(n3821) );
  AND U4047 ( .A(n3869), .B(n3870), .Z(n3868) );
  XOR U4048 ( .A(n3871), .B(n3872), .Z(n3870) );
  XOR U4049 ( .A(n3867), .B(n3873), .Z(n3872) );
  XNOR U4050 ( .A(n3854), .B(n3874), .Z(n3869) );
  XNOR U4051 ( .A(n3867), .B(n3855), .Z(n3874) );
  XNOR U4052 ( .A(n3839), .B(n3838), .Z(n3855) );
  XOR U4053 ( .A(n3875), .B(n3833), .Z(n3838) );
  XNOR U4054 ( .A(n3831), .B(n3876), .Z(n3833) );
  ANDN U4055 ( .A(n2094), .B(n2605), .Z(n3876) );
  XOR U4056 ( .A(n3877), .B(n3878), .Z(n3831) );
  AND U4057 ( .A(n3879), .B(n3880), .Z(n3878) );
  XNOR U4058 ( .A(n3881), .B(n3877), .Z(n3880) );
  XOR U4059 ( .A(n3882), .B(n3835), .Z(n3875) );
  AND U4060 ( .A(n2603), .B(n2087), .Z(n3835) );
  IV U4061 ( .A(n3837), .Z(n3882) );
  XNOR U4062 ( .A(n3843), .B(n3845), .Z(n3839) );
  NAND U4063 ( .A(n2845), .B(n1892), .Z(n3845) );
  XNOR U4064 ( .A(n3841), .B(n3886), .Z(n3843) );
  ANDN U4065 ( .A(n1897), .B(n2847), .Z(n3886) );
  XOR U4066 ( .A(n3890), .B(n3866), .Z(n3854) );
  XNOR U4067 ( .A(n3850), .B(n3852), .Z(n3866) );
  NAND U4068 ( .A(n2376), .B(n2288), .Z(n3852) );
  XNOR U4069 ( .A(n3848), .B(n3891), .Z(n3850) );
  ANDN U4070 ( .A(n2293), .B(n2378), .Z(n3891) );
  XOR U4071 ( .A(n3892), .B(n3893), .Z(n3848) );
  AND U4072 ( .A(n3894), .B(n3895), .Z(n3893) );
  XOR U4073 ( .A(n3896), .B(n3892), .Z(n3895) );
  XNOR U4074 ( .A(n3865), .B(n3853), .Z(n3890) );
  XOR U4075 ( .A(n3900), .B(n3860), .Z(n3865) );
  XNOR U4076 ( .A(n3858), .B(n3901), .Z(n3860) );
  ANDN U4077 ( .A(n2523), .B(n2165), .Z(n3901) );
  XOR U4078 ( .A(n3902), .B(n3903), .Z(n3858) );
  AND U4079 ( .A(n3904), .B(n3905), .Z(n3903) );
  XNOR U4080 ( .A(n3906), .B(n3902), .Z(n3905) );
  XOR U4081 ( .A(n3907), .B(n3862), .Z(n3900) );
  AND U4082 ( .A(n2163), .B(n2516), .Z(n3862) );
  IV U4083 ( .A(n3864), .Z(n3907) );
  XOR U4084 ( .A(n3911), .B(n3912), .Z(n3867) );
  AND U4085 ( .A(n3913), .B(n3914), .Z(n3912) );
  XOR U4086 ( .A(n3915), .B(n3916), .Z(n3914) );
  XOR U4087 ( .A(n3911), .B(n3917), .Z(n3916) );
  XNOR U4088 ( .A(n3898), .B(n3918), .Z(n3913) );
  XNOR U4089 ( .A(n3911), .B(n3899), .Z(n3918) );
  XNOR U4090 ( .A(n3885), .B(n3884), .Z(n3899) );
  XOR U4091 ( .A(n3919), .B(n3879), .Z(n3884) );
  XNOR U4092 ( .A(n3877), .B(n3920), .Z(n3879) );
  ANDN U4093 ( .A(n2094), .B(n2725), .Z(n3920) );
  XOR U4094 ( .A(n3921), .B(n3922), .Z(n3877) );
  AND U4095 ( .A(n3923), .B(n3924), .Z(n3922) );
  XNOR U4096 ( .A(n3925), .B(n3921), .Z(n3924) );
  XOR U4097 ( .A(n3926), .B(n3881), .Z(n3919) );
  AND U4098 ( .A(n2723), .B(n2087), .Z(n3881) );
  IV U4099 ( .A(n3883), .Z(n3926) );
  XNOR U4100 ( .A(n3888), .B(n3889), .Z(n3885) );
  NAND U4101 ( .A(n2970), .B(n1892), .Z(n3889) );
  XNOR U4102 ( .A(n3887), .B(n3930), .Z(n3888) );
  ANDN U4103 ( .A(n1897), .B(n2972), .Z(n3930) );
  XOR U4104 ( .A(n3931), .B(n3932), .Z(n3887) );
  AND U4105 ( .A(n3933), .B(n3934), .Z(n3932) );
  XOR U4106 ( .A(n3935), .B(n3931), .Z(n3934) );
  XOR U4107 ( .A(n3936), .B(n3910), .Z(n3898) );
  XNOR U4108 ( .A(n3894), .B(n3896), .Z(n3910) );
  NAND U4109 ( .A(n2484), .B(n2288), .Z(n3896) );
  XNOR U4110 ( .A(n3892), .B(n3937), .Z(n3894) );
  ANDN U4111 ( .A(n2293), .B(n2486), .Z(n3937) );
  XOR U4112 ( .A(n3938), .B(n3939), .Z(n3892) );
  AND U4113 ( .A(n3940), .B(n3941), .Z(n3939) );
  XOR U4114 ( .A(n3942), .B(n3938), .Z(n3941) );
  XNOR U4115 ( .A(n3909), .B(n3897), .Z(n3936) );
  XOR U4116 ( .A(n3946), .B(n3904), .Z(n3909) );
  XNOR U4117 ( .A(n3902), .B(n3947), .Z(n3904) );
  ANDN U4118 ( .A(n2523), .B(n2271), .Z(n3947) );
  XOR U4119 ( .A(n3948), .B(n3949), .Z(n3902) );
  AND U4120 ( .A(n3950), .B(n3951), .Z(n3949) );
  XNOR U4121 ( .A(n3952), .B(n3948), .Z(n3951) );
  XOR U4122 ( .A(n3953), .B(n3906), .Z(n3946) );
  AND U4123 ( .A(n2269), .B(n2516), .Z(n3906) );
  IV U4124 ( .A(n3908), .Z(n3953) );
  XOR U4125 ( .A(n3957), .B(n3958), .Z(n3911) );
  AND U4126 ( .A(n3959), .B(n3960), .Z(n3958) );
  XOR U4127 ( .A(n3961), .B(n3962), .Z(n3960) );
  XOR U4128 ( .A(n3957), .B(n3963), .Z(n3962) );
  XNOR U4129 ( .A(n3944), .B(n3964), .Z(n3959) );
  XNOR U4130 ( .A(n3957), .B(n3945), .Z(n3964) );
  XNOR U4131 ( .A(n3929), .B(n3928), .Z(n3945) );
  XOR U4132 ( .A(n3965), .B(n3923), .Z(n3928) );
  XNOR U4133 ( .A(n3921), .B(n3966), .Z(n3923) );
  ANDN U4134 ( .A(n2094), .B(n2847), .Z(n3966) );
  XOR U4135 ( .A(n3967), .B(n3968), .Z(n3921) );
  AND U4136 ( .A(n3969), .B(n3970), .Z(n3968) );
  XNOR U4137 ( .A(n3971), .B(n3967), .Z(n3970) );
  XOR U4138 ( .A(n3972), .B(n3925), .Z(n3965) );
  AND U4139 ( .A(n2845), .B(n2087), .Z(n3925) );
  IV U4140 ( .A(n3927), .Z(n3972) );
  XNOR U4141 ( .A(n3933), .B(n3935), .Z(n3929) );
  NAND U4142 ( .A(n3102), .B(n1892), .Z(n3935) );
  XNOR U4143 ( .A(n3931), .B(n3976), .Z(n3933) );
  ANDN U4144 ( .A(n1897), .B(n3104), .Z(n3976) );
  XOR U4145 ( .A(n3977), .B(n3978), .Z(n3931) );
  AND U4146 ( .A(n3979), .B(n3980), .Z(n3978) );
  XOR U4147 ( .A(n3981), .B(n3977), .Z(n3980) );
  XOR U4148 ( .A(n3982), .B(n3956), .Z(n3944) );
  XNOR U4149 ( .A(n3940), .B(n3942), .Z(n3956) );
  NAND U4150 ( .A(n2603), .B(n2288), .Z(n3942) );
  XNOR U4151 ( .A(n3938), .B(n3983), .Z(n3940) );
  ANDN U4152 ( .A(n2293), .B(n2605), .Z(n3983) );
  XOR U4153 ( .A(n3984), .B(n3985), .Z(n3938) );
  AND U4154 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U4155 ( .A(n3988), .B(n3984), .Z(n3987) );
  XNOR U4156 ( .A(n3955), .B(n3943), .Z(n3982) );
  XOR U4157 ( .A(n3992), .B(n3950), .Z(n3955) );
  XNOR U4158 ( .A(n3948), .B(n3993), .Z(n3950) );
  ANDN U4159 ( .A(n2523), .B(n2378), .Z(n3993) );
  XOR U4160 ( .A(n3994), .B(n3995), .Z(n3948) );
  AND U4161 ( .A(n3996), .B(n3997), .Z(n3995) );
  XNOR U4162 ( .A(n3998), .B(n3994), .Z(n3997) );
  XOR U4163 ( .A(n3999), .B(n3952), .Z(n3992) );
  AND U4164 ( .A(n2376), .B(n2516), .Z(n3952) );
  IV U4165 ( .A(n3954), .Z(n3999) );
  XOR U4166 ( .A(n4003), .B(n4004), .Z(n3957) );
  AND U4167 ( .A(n4005), .B(n4006), .Z(n4004) );
  XOR U4168 ( .A(n4007), .B(n4008), .Z(n4006) );
  XOR U4169 ( .A(n4003), .B(n4009), .Z(n4008) );
  XNOR U4170 ( .A(n3990), .B(n4010), .Z(n4005) );
  XNOR U4171 ( .A(n4003), .B(n3991), .Z(n4010) );
  XNOR U4172 ( .A(n3975), .B(n3974), .Z(n3991) );
  XOR U4173 ( .A(n4011), .B(n3969), .Z(n3974) );
  XNOR U4174 ( .A(n3967), .B(n4012), .Z(n3969) );
  ANDN U4175 ( .A(n2094), .B(n2972), .Z(n4012) );
  XOR U4176 ( .A(n4013), .B(n4014), .Z(n3967) );
  AND U4177 ( .A(n4015), .B(n4016), .Z(n4014) );
  XNOR U4178 ( .A(n4017), .B(n4013), .Z(n4016) );
  XOR U4179 ( .A(n4018), .B(n3971), .Z(n4011) );
  AND U4180 ( .A(n2970), .B(n2087), .Z(n3971) );
  IV U4181 ( .A(n3973), .Z(n4018) );
  XNOR U4182 ( .A(n3979), .B(n3981), .Z(n3975) );
  NAND U4183 ( .A(n3234), .B(n1892), .Z(n3981) );
  XNOR U4184 ( .A(n3977), .B(n4022), .Z(n3979) );
  ANDN U4185 ( .A(n1897), .B(n3236), .Z(n4022) );
  XOR U4186 ( .A(n4023), .B(n4024), .Z(n3977) );
  AND U4187 ( .A(n4025), .B(n4026), .Z(n4024) );
  XOR U4188 ( .A(n4027), .B(n4023), .Z(n4026) );
  XOR U4189 ( .A(n4028), .B(n4002), .Z(n3990) );
  XNOR U4190 ( .A(n3986), .B(n3988), .Z(n4002) );
  NAND U4191 ( .A(n2723), .B(n2288), .Z(n3988) );
  XNOR U4192 ( .A(n3984), .B(n4029), .Z(n3986) );
  ANDN U4193 ( .A(n2293), .B(n2725), .Z(n4029) );
  XOR U4194 ( .A(n4030), .B(n4031), .Z(n3984) );
  AND U4195 ( .A(n4032), .B(n4033), .Z(n4031) );
  XOR U4196 ( .A(n4034), .B(n4030), .Z(n4033) );
  XNOR U4197 ( .A(n4001), .B(n3989), .Z(n4028) );
  XOR U4198 ( .A(n4038), .B(n3996), .Z(n4001) );
  XNOR U4199 ( .A(n3994), .B(n4039), .Z(n3996) );
  ANDN U4200 ( .A(n2523), .B(n2486), .Z(n4039) );
  XOR U4201 ( .A(n4040), .B(n4041), .Z(n3994) );
  AND U4202 ( .A(n4042), .B(n4043), .Z(n4041) );
  XNOR U4203 ( .A(n4044), .B(n4040), .Z(n4043) );
  XOR U4204 ( .A(n4045), .B(n3998), .Z(n4038) );
  AND U4205 ( .A(n2484), .B(n2516), .Z(n3998) );
  IV U4206 ( .A(n4000), .Z(n4045) );
  XOR U4207 ( .A(n4049), .B(n4050), .Z(n4003) );
  AND U4208 ( .A(n4051), .B(n4052), .Z(n4050) );
  XOR U4209 ( .A(n4053), .B(n4054), .Z(n4052) );
  XOR U4210 ( .A(n4049), .B(n4055), .Z(n4054) );
  XNOR U4211 ( .A(n4036), .B(n4056), .Z(n4051) );
  XNOR U4212 ( .A(n4049), .B(n4037), .Z(n4056) );
  XNOR U4213 ( .A(n4021), .B(n4020), .Z(n4037) );
  XOR U4214 ( .A(n4057), .B(n4015), .Z(n4020) );
  XNOR U4215 ( .A(n4013), .B(n4058), .Z(n4015) );
  ANDN U4216 ( .A(n2094), .B(n3104), .Z(n4058) );
  XOR U4217 ( .A(n4062), .B(n4017), .Z(n4057) );
  AND U4218 ( .A(n3102), .B(n2087), .Z(n4017) );
  IV U4219 ( .A(n4019), .Z(n4062) );
  XNOR U4220 ( .A(n4025), .B(n4027), .Z(n4021) );
  NAND U4221 ( .A(n3370), .B(n1892), .Z(n4027) );
  XNOR U4222 ( .A(n4023), .B(n4066), .Z(n4025) );
  ANDN U4223 ( .A(n1897), .B(n3372), .Z(n4066) );
  XOR U4224 ( .A(n4070), .B(n4048), .Z(n4036) );
  XNOR U4225 ( .A(n4032), .B(n4034), .Z(n4048) );
  NAND U4226 ( .A(n2845), .B(n2288), .Z(n4034) );
  XNOR U4227 ( .A(n4030), .B(n4071), .Z(n4032) );
  ANDN U4228 ( .A(n2293), .B(n2847), .Z(n4071) );
  XOR U4229 ( .A(n4072), .B(n4073), .Z(n4030) );
  AND U4230 ( .A(n4074), .B(n4075), .Z(n4073) );
  XOR U4231 ( .A(n4076), .B(n4072), .Z(n4075) );
  XNOR U4232 ( .A(n4047), .B(n4035), .Z(n4070) );
  XOR U4233 ( .A(n4080), .B(n4042), .Z(n4047) );
  XNOR U4234 ( .A(n4040), .B(n4081), .Z(n4042) );
  ANDN U4235 ( .A(n2523), .B(n2605), .Z(n4081) );
  XOR U4236 ( .A(n4082), .B(n4083), .Z(n4040) );
  AND U4237 ( .A(n4084), .B(n4085), .Z(n4083) );
  XNOR U4238 ( .A(n4086), .B(n4082), .Z(n4085) );
  XOR U4239 ( .A(n4087), .B(n4044), .Z(n4080) );
  AND U4240 ( .A(n2603), .B(n2516), .Z(n4044) );
  IV U4241 ( .A(n4046), .Z(n4087) );
  XOR U4242 ( .A(n4092), .B(n4093), .Z(n3411) );
  XOR U4243 ( .A(n4094), .B(n4091), .Z(n4092) );
  XNOR U4244 ( .A(n4079), .B(n4078), .Z(n3410) );
  XOR U4245 ( .A(n4095), .B(n4090), .Z(n4078) );
  XNOR U4246 ( .A(n4074), .B(n4076), .Z(n4090) );
  NAND U4247 ( .A(n2970), .B(n2288), .Z(n4076) );
  XNOR U4248 ( .A(n4072), .B(n4096), .Z(n4074) );
  ANDN U4249 ( .A(n2293), .B(n2972), .Z(n4096) );
  XOR U4250 ( .A(n4089), .B(n4077), .Z(n4095) );
  XOR U4251 ( .A(n4100), .B(n4101), .Z(n4077) );
  XOR U4252 ( .A(n4102), .B(n4084), .Z(n4089) );
  XNOR U4253 ( .A(n4082), .B(n4103), .Z(n4084) );
  ANDN U4254 ( .A(n2523), .B(n2725), .Z(n4103) );
  AND U4255 ( .A(n2723), .B(n2516), .Z(n4086) );
  XNOR U4256 ( .A(n4107), .B(n4108), .Z(n4088) );
  AND U4257 ( .A(n4109), .B(n4110), .Z(n4108) );
  XNOR U4258 ( .A(n4105), .B(n4111), .Z(n4110) );
  XNOR U4259 ( .A(n4106), .B(n4107), .Z(n4111) );
  AND U4260 ( .A(n2845), .B(n2516), .Z(n4106) );
  XOR U4261 ( .A(n4104), .B(n4112), .Z(n4105) );
  ANDN U4262 ( .A(n2523), .B(n2847), .Z(n4112) );
  XNOR U4263 ( .A(n4098), .B(n4116), .Z(n4109) );
  XNOR U4264 ( .A(n4099), .B(n4107), .Z(n4116) );
  AND U4265 ( .A(n3102), .B(n2288), .Z(n4099) );
  XOR U4266 ( .A(n4097), .B(n4117), .Z(n4098) );
  ANDN U4267 ( .A(n2293), .B(n3104), .Z(n4117) );
  XOR U4268 ( .A(n4121), .B(n4122), .Z(n4107) );
  AND U4269 ( .A(n4123), .B(n4124), .Z(n4122) );
  XNOR U4270 ( .A(n4114), .B(n4125), .Z(n4124) );
  XNOR U4271 ( .A(n4115), .B(n4121), .Z(n4125) );
  AND U4272 ( .A(n2970), .B(n2516), .Z(n4115) );
  XOR U4273 ( .A(n4113), .B(n4126), .Z(n4114) );
  ANDN U4274 ( .A(n2523), .B(n2972), .Z(n4126) );
  XNOR U4275 ( .A(n4119), .B(n4130), .Z(n4123) );
  XNOR U4276 ( .A(n4120), .B(n4121), .Z(n4130) );
  AND U4277 ( .A(n3234), .B(n2288), .Z(n4120) );
  XOR U4278 ( .A(n4118), .B(n4131), .Z(n4119) );
  ANDN U4279 ( .A(n2293), .B(n3236), .Z(n4131) );
  XOR U4280 ( .A(n4135), .B(n4136), .Z(n4121) );
  AND U4281 ( .A(n4137), .B(n4138), .Z(n4136) );
  XNOR U4282 ( .A(n4128), .B(n4139), .Z(n4138) );
  XNOR U4283 ( .A(n4129), .B(n4135), .Z(n4139) );
  AND U4284 ( .A(n3102), .B(n2516), .Z(n4129) );
  XOR U4285 ( .A(n4127), .B(n4140), .Z(n4128) );
  ANDN U4286 ( .A(n2523), .B(n3104), .Z(n4140) );
  XNOR U4287 ( .A(n4133), .B(n4144), .Z(n4137) );
  XNOR U4288 ( .A(n4134), .B(n4135), .Z(n4144) );
  AND U4289 ( .A(n3370), .B(n2288), .Z(n4134) );
  XOR U4290 ( .A(n4132), .B(n4145), .Z(n4133) );
  ANDN U4291 ( .A(n2293), .B(n3372), .Z(n4145) );
  XNOR U4292 ( .A(n4150), .B(n4142), .Z(n4101) );
  XNOR U4293 ( .A(n4141), .B(n4151), .Z(n4142) );
  ANDN U4294 ( .A(n2523), .B(n3236), .Z(n4151) );
  XNOR U4295 ( .A(n4154), .B(n4152), .Z(n4153) );
  ANDN U4296 ( .A(n2523), .B(n3372), .Z(n4154) );
  XNOR U4297 ( .A(n4149), .B(n4143), .Z(n4150) );
  AND U4298 ( .A(n3234), .B(n2516), .Z(n4143) );
  XNOR U4299 ( .A(n4147), .B(n4148), .Z(n4100) );
  NAND U4300 ( .A(n4158), .B(n2288), .Z(n4148) );
  XNOR U4301 ( .A(n4146), .B(n4159), .Z(n4147) );
  ANDN U4302 ( .A(n2293), .B(n4160), .Z(n4159) );
  NAND U4303 ( .A(A[0]), .B(n4161), .Z(n4146) );
  NANDN U4304 ( .B(n2288), .A(n4162), .Z(n4161) );
  NANDN U4305 ( .B(n4163), .A(n2293), .Z(n4162) );
  IV U4306 ( .A(n2187), .Z(n2288) );
  XNOR U4307 ( .A(n4156), .B(n4157), .Z(n4149) );
  NAND U4308 ( .A(n4158), .B(n2516), .Z(n4157) );
  XNOR U4309 ( .A(n4155), .B(n4166), .Z(n4156) );
  ANDN U4310 ( .A(n2523), .B(n4160), .Z(n4166) );
  NAND U4311 ( .A(A[0]), .B(n4167), .Z(n4155) );
  NANDN U4312 ( .B(n2516), .A(n4168), .Z(n4167) );
  NANDN U4313 ( .B(n4163), .A(n2523), .Z(n4168) );
  IV U4314 ( .A(n2404), .Z(n2516) );
  XNOR U4315 ( .A(n4065), .B(n4064), .Z(n4079) );
  XOR U4316 ( .A(n4171), .B(n4060), .Z(n4064) );
  XNOR U4317 ( .A(n4059), .B(n4172), .Z(n4060) );
  ANDN U4318 ( .A(n2094), .B(n3236), .Z(n4172) );
  XNOR U4319 ( .A(n4175), .B(n4173), .Z(n4174) );
  ANDN U4320 ( .A(n2094), .B(n3372), .Z(n4175) );
  XNOR U4321 ( .A(n4063), .B(n4061), .Z(n4171) );
  AND U4322 ( .A(n3234), .B(n2087), .Z(n4061) );
  XNOR U4323 ( .A(n4177), .B(n4178), .Z(n4063) );
  NAND U4324 ( .A(n4158), .B(n2087), .Z(n4178) );
  XNOR U4325 ( .A(n4176), .B(n4179), .Z(n4177) );
  ANDN U4326 ( .A(n2094), .B(n4160), .Z(n4179) );
  NAND U4327 ( .A(A[0]), .B(n4180), .Z(n4176) );
  NANDN U4328 ( .B(n2087), .A(n4181), .Z(n4180) );
  NANDN U4329 ( .B(n4163), .A(n2094), .Z(n4181) );
  IV U4330 ( .A(n1988), .Z(n2087) );
  XNOR U4331 ( .A(n4068), .B(n4069), .Z(n4065) );
  NAND U4332 ( .A(n4158), .B(n1892), .Z(n4069) );
  XNOR U4333 ( .A(n4067), .B(n4184), .Z(n4068) );
  ANDN U4334 ( .A(n1897), .B(n4160), .Z(n4184) );
  NAND U4335 ( .A(A[0]), .B(n4185), .Z(n4067) );
  NANDN U4336 ( .B(n1892), .A(n4186), .Z(n4185) );
  NANDN U4337 ( .B(n4163), .A(n1897), .Z(n4186) );
  IV U4338 ( .A(n1796), .Z(n1892) );
  XNOR U4339 ( .A(n4189), .B(n4190), .Z(n4091) );
  XOR U4340 ( .A(n4191), .B(n3313), .Z(n3308) );
  XNOR U4341 ( .A(n3304), .B(n3305), .Z(n3313) );
  NAND U4342 ( .A(n3301), .B(n937), .Z(n3305) );
  XNOR U4343 ( .A(n3303), .B(n4192), .Z(n3304) );
  ANDN U4344 ( .A(n3306), .B(n939), .Z(n4192) );
  XOR U4345 ( .A(n4193), .B(n4194), .Z(n3303) );
  AND U4346 ( .A(n4195), .B(n4196), .Z(n4194) );
  XOR U4347 ( .A(n4197), .B(n4193), .Z(n4196) );
  XNOR U4348 ( .A(n3311), .B(n3307), .Z(n4191) );
  XNOR U4349 ( .A(n3422), .B(n3421), .Z(n3434) );
  XOR U4350 ( .A(n4199), .B(n3417), .Z(n3421) );
  XNOR U4351 ( .A(n3415), .B(n4200), .Z(n3417) );
  ANDN U4352 ( .A(n3032), .B(n1067), .Z(n4200) );
  XOR U4353 ( .A(n4201), .B(n4202), .Z(n3415) );
  AND U4354 ( .A(n4203), .B(n4204), .Z(n4202) );
  XNOR U4355 ( .A(n4205), .B(n4201), .Z(n4204) );
  AND U4356 ( .A(n3025), .B(n1065), .Z(n3419) );
  XNOR U4357 ( .A(n3426), .B(n3428), .Z(n3422) );
  NAND U4358 ( .A(n2778), .B(n1166), .Z(n3428) );
  XNOR U4359 ( .A(n3424), .B(n4209), .Z(n3426) );
  ANDN U4360 ( .A(n2783), .B(n1168), .Z(n4209) );
  XOR U4361 ( .A(n4210), .B(n4211), .Z(n3424) );
  AND U4362 ( .A(n4212), .B(n4213), .Z(n4211) );
  XOR U4363 ( .A(n4214), .B(n4210), .Z(n4213) );
  XOR U4364 ( .A(n4215), .B(n4216), .Z(n3435) );
  XNOR U4365 ( .A(n4217), .B(n4198), .Z(n4215) );
  XOR U4366 ( .A(n4219), .B(n4220), .Z(n3473) );
  XOR U4367 ( .A(n4221), .B(n4218), .Z(n4219) );
  XNOR U4368 ( .A(n4208), .B(n4207), .Z(n3471) );
  XOR U4369 ( .A(n4222), .B(n4203), .Z(n4207) );
  XNOR U4370 ( .A(n4201), .B(n4223), .Z(n4203) );
  ANDN U4371 ( .A(n3032), .B(n1109), .Z(n4223) );
  XOR U4372 ( .A(n4224), .B(n4225), .Z(n4201) );
  AND U4373 ( .A(n4226), .B(n4227), .Z(n4225) );
  XNOR U4374 ( .A(n4228), .B(n4224), .Z(n4227) );
  XOR U4375 ( .A(n4229), .B(n4205), .Z(n4222) );
  AND U4376 ( .A(n3025), .B(n1107), .Z(n4205) );
  IV U4377 ( .A(n4206), .Z(n4229) );
  XNOR U4378 ( .A(n4212), .B(n4214), .Z(n4208) );
  NAND U4379 ( .A(n2778), .B(n1230), .Z(n4214) );
  XNOR U4380 ( .A(n4210), .B(n4233), .Z(n4212) );
  ANDN U4381 ( .A(n2783), .B(n1232), .Z(n4233) );
  XOR U4382 ( .A(n4234), .B(n4235), .Z(n4210) );
  AND U4383 ( .A(n4236), .B(n4237), .Z(n4235) );
  XOR U4384 ( .A(n4238), .B(n4234), .Z(n4237) );
  XOR U4385 ( .A(n4240), .B(n4241), .Z(n3518) );
  XOR U4386 ( .A(n4242), .B(n4239), .Z(n4240) );
  XNOR U4387 ( .A(n4232), .B(n4231), .Z(n3516) );
  XOR U4388 ( .A(n4243), .B(n4226), .Z(n4231) );
  XNOR U4389 ( .A(n4224), .B(n4244), .Z(n4226) );
  ANDN U4390 ( .A(n3032), .B(n1168), .Z(n4244) );
  XOR U4391 ( .A(n4245), .B(n4246), .Z(n4224) );
  AND U4392 ( .A(n4247), .B(n4248), .Z(n4246) );
  XNOR U4393 ( .A(n4249), .B(n4245), .Z(n4248) );
  XOR U4394 ( .A(n4250), .B(n4228), .Z(n4243) );
  AND U4395 ( .A(n3025), .B(n1166), .Z(n4228) );
  IV U4396 ( .A(n4230), .Z(n4250) );
  XNOR U4397 ( .A(n4236), .B(n4238), .Z(n4232) );
  NAND U4398 ( .A(n2778), .B(n1298), .Z(n4238) );
  XNOR U4399 ( .A(n4234), .B(n4254), .Z(n4236) );
  ANDN U4400 ( .A(n2783), .B(n1300), .Z(n4254) );
  XOR U4401 ( .A(n4255), .B(n4256), .Z(n4234) );
  AND U4402 ( .A(n4257), .B(n4258), .Z(n4256) );
  XOR U4403 ( .A(n4259), .B(n4255), .Z(n4258) );
  XOR U4404 ( .A(n4261), .B(n4262), .Z(n3560) );
  XOR U4405 ( .A(n4263), .B(n4260), .Z(n4261) );
  XNOR U4406 ( .A(n4253), .B(n4252), .Z(n3558) );
  XOR U4407 ( .A(n4264), .B(n4247), .Z(n4252) );
  XNOR U4408 ( .A(n4245), .B(n4265), .Z(n4247) );
  ANDN U4409 ( .A(n3032), .B(n1232), .Z(n4265) );
  XOR U4410 ( .A(n4266), .B(n4267), .Z(n4245) );
  AND U4411 ( .A(n4268), .B(n4269), .Z(n4267) );
  XNOR U4412 ( .A(n4270), .B(n4266), .Z(n4269) );
  AND U4413 ( .A(n3025), .B(n1230), .Z(n4249) );
  XNOR U4414 ( .A(n4257), .B(n4259), .Z(n4253) );
  NAND U4415 ( .A(n2778), .B(n1365), .Z(n4259) );
  XNOR U4416 ( .A(n4255), .B(n4274), .Z(n4257) );
  ANDN U4417 ( .A(n2783), .B(n1367), .Z(n4274) );
  XOR U4418 ( .A(n4275), .B(n4276), .Z(n4255) );
  AND U4419 ( .A(n4277), .B(n4278), .Z(n4276) );
  XOR U4420 ( .A(n4279), .B(n4275), .Z(n4278) );
  XOR U4421 ( .A(n4281), .B(n4282), .Z(n3603) );
  XOR U4422 ( .A(n4283), .B(n4280), .Z(n4281) );
  XNOR U4423 ( .A(n4273), .B(n4272), .Z(n3601) );
  XOR U4424 ( .A(n4284), .B(n4268), .Z(n4272) );
  XNOR U4425 ( .A(n4266), .B(n4285), .Z(n4268) );
  ANDN U4426 ( .A(n3032), .B(n1300), .Z(n4285) );
  XOR U4427 ( .A(n4286), .B(n4287), .Z(n4266) );
  AND U4428 ( .A(n4288), .B(n4289), .Z(n4287) );
  XNOR U4429 ( .A(n4290), .B(n4286), .Z(n4289) );
  XOR U4430 ( .A(n4291), .B(n4270), .Z(n4284) );
  AND U4431 ( .A(n3025), .B(n1298), .Z(n4270) );
  IV U4432 ( .A(n4271), .Z(n4291) );
  XNOR U4433 ( .A(n4277), .B(n4279), .Z(n4273) );
  NAND U4434 ( .A(n2778), .B(n1439), .Z(n4279) );
  XNOR U4435 ( .A(n4275), .B(n4295), .Z(n4277) );
  ANDN U4436 ( .A(n2783), .B(n1441), .Z(n4295) );
  XOR U4437 ( .A(n4296), .B(n4297), .Z(n4275) );
  AND U4438 ( .A(n4298), .B(n4299), .Z(n4297) );
  XOR U4439 ( .A(n4300), .B(n4296), .Z(n4299) );
  XOR U4440 ( .A(n4302), .B(n4303), .Z(n3645) );
  XOR U4441 ( .A(n4304), .B(n4301), .Z(n4302) );
  XNOR U4442 ( .A(n4294), .B(n4293), .Z(n3643) );
  XOR U4443 ( .A(n4305), .B(n4288), .Z(n4293) );
  XNOR U4444 ( .A(n4286), .B(n4306), .Z(n4288) );
  ANDN U4445 ( .A(n3032), .B(n1367), .Z(n4306) );
  XOR U4446 ( .A(n4307), .B(n4308), .Z(n4286) );
  AND U4447 ( .A(n4309), .B(n4310), .Z(n4308) );
  XNOR U4448 ( .A(n4311), .B(n4307), .Z(n4310) );
  XOR U4449 ( .A(n4312), .B(n4290), .Z(n4305) );
  AND U4450 ( .A(n3025), .B(n1365), .Z(n4290) );
  IV U4451 ( .A(n4292), .Z(n4312) );
  XNOR U4452 ( .A(n4298), .B(n4300), .Z(n4294) );
  NAND U4453 ( .A(n2778), .B(n1517), .Z(n4300) );
  XNOR U4454 ( .A(n4296), .B(n4316), .Z(n4298) );
  ANDN U4455 ( .A(n2783), .B(n1519), .Z(n4316) );
  XOR U4456 ( .A(n4317), .B(n4318), .Z(n4296) );
  AND U4457 ( .A(n4319), .B(n4320), .Z(n4318) );
  XOR U4458 ( .A(n4321), .B(n4317), .Z(n4320) );
  XOR U4459 ( .A(n4323), .B(n4324), .Z(n3691) );
  XOR U4460 ( .A(n4325), .B(n4322), .Z(n4323) );
  XNOR U4461 ( .A(n4315), .B(n4314), .Z(n3689) );
  XOR U4462 ( .A(n4326), .B(n4309), .Z(n4314) );
  XNOR U4463 ( .A(n4307), .B(n4327), .Z(n4309) );
  ANDN U4464 ( .A(n3032), .B(n1441), .Z(n4327) );
  XOR U4465 ( .A(n4328), .B(n4329), .Z(n4307) );
  AND U4466 ( .A(n4330), .B(n4331), .Z(n4329) );
  XNOR U4467 ( .A(n4332), .B(n4328), .Z(n4331) );
  XOR U4468 ( .A(n4333), .B(n4311), .Z(n4326) );
  AND U4469 ( .A(n3025), .B(n1439), .Z(n4311) );
  IV U4470 ( .A(n4313), .Z(n4333) );
  XNOR U4471 ( .A(n4319), .B(n4321), .Z(n4315) );
  NAND U4472 ( .A(n2778), .B(n1598), .Z(n4321) );
  XNOR U4473 ( .A(n4317), .B(n4337), .Z(n4319) );
  ANDN U4474 ( .A(n2783), .B(n1600), .Z(n4337) );
  XOR U4475 ( .A(n4338), .B(n4339), .Z(n4317) );
  AND U4476 ( .A(n4340), .B(n4341), .Z(n4339) );
  XOR U4477 ( .A(n4342), .B(n4338), .Z(n4341) );
  XOR U4478 ( .A(n4344), .B(n4345), .Z(n3735) );
  XOR U4479 ( .A(n4346), .B(n4343), .Z(n4344) );
  XNOR U4480 ( .A(n4336), .B(n4335), .Z(n3733) );
  XOR U4481 ( .A(n4347), .B(n4330), .Z(n4335) );
  XNOR U4482 ( .A(n4328), .B(n4348), .Z(n4330) );
  ANDN U4483 ( .A(n3032), .B(n1519), .Z(n4348) );
  XOR U4484 ( .A(n4349), .B(n4350), .Z(n4328) );
  AND U4485 ( .A(n4351), .B(n4352), .Z(n4350) );
  XNOR U4486 ( .A(n4353), .B(n4349), .Z(n4352) );
  XOR U4487 ( .A(n4354), .B(n4332), .Z(n4347) );
  AND U4488 ( .A(n3025), .B(n1517), .Z(n4332) );
  IV U4489 ( .A(n4334), .Z(n4354) );
  XNOR U4490 ( .A(n4340), .B(n4342), .Z(n4336) );
  NAND U4491 ( .A(n2778), .B(n1682), .Z(n4342) );
  XNOR U4492 ( .A(n4338), .B(n4358), .Z(n4340) );
  ANDN U4493 ( .A(n2783), .B(n1684), .Z(n4358) );
  XOR U4494 ( .A(n4359), .B(n4360), .Z(n4338) );
  AND U4495 ( .A(n4361), .B(n4362), .Z(n4360) );
  XOR U4496 ( .A(n4363), .B(n4359), .Z(n4362) );
  XOR U4497 ( .A(n4365), .B(n4366), .Z(n3781) );
  XOR U4498 ( .A(n4367), .B(n4364), .Z(n4365) );
  XNOR U4499 ( .A(n4357), .B(n4356), .Z(n3779) );
  XOR U4500 ( .A(n4368), .B(n4351), .Z(n4356) );
  XNOR U4501 ( .A(n4349), .B(n4369), .Z(n4351) );
  ANDN U4502 ( .A(n3032), .B(n1600), .Z(n4369) );
  XOR U4503 ( .A(n4370), .B(n4371), .Z(n4349) );
  AND U4504 ( .A(n4372), .B(n4373), .Z(n4371) );
  XNOR U4505 ( .A(n4374), .B(n4370), .Z(n4373) );
  XOR U4506 ( .A(n4375), .B(n4353), .Z(n4368) );
  AND U4507 ( .A(n3025), .B(n1598), .Z(n4353) );
  IV U4508 ( .A(n4355), .Z(n4375) );
  XNOR U4509 ( .A(n4361), .B(n4363), .Z(n4357) );
  NAND U4510 ( .A(n2778), .B(n1773), .Z(n4363) );
  XNOR U4511 ( .A(n4359), .B(n4379), .Z(n4361) );
  ANDN U4512 ( .A(n2783), .B(n1775), .Z(n4379) );
  XOR U4513 ( .A(n4380), .B(n4381), .Z(n4359) );
  AND U4514 ( .A(n4382), .B(n4383), .Z(n4381) );
  XOR U4515 ( .A(n4384), .B(n4380), .Z(n4383) );
  XOR U4516 ( .A(n4386), .B(n4387), .Z(n3827) );
  XOR U4517 ( .A(n4388), .B(n4385), .Z(n4386) );
  XNOR U4518 ( .A(n4378), .B(n4377), .Z(n3825) );
  XOR U4519 ( .A(n4389), .B(n4372), .Z(n4377) );
  XNOR U4520 ( .A(n4370), .B(n4390), .Z(n4372) );
  ANDN U4521 ( .A(n3032), .B(n1684), .Z(n4390) );
  XOR U4522 ( .A(n4391), .B(n4392), .Z(n4370) );
  AND U4523 ( .A(n4393), .B(n4394), .Z(n4392) );
  XNOR U4524 ( .A(n4395), .B(n4391), .Z(n4394) );
  XOR U4525 ( .A(n4396), .B(n4374), .Z(n4389) );
  AND U4526 ( .A(n3025), .B(n1682), .Z(n4374) );
  IV U4527 ( .A(n4376), .Z(n4396) );
  XNOR U4528 ( .A(n4382), .B(n4384), .Z(n4378) );
  NAND U4529 ( .A(n2778), .B(n1870), .Z(n4384) );
  XNOR U4530 ( .A(n4380), .B(n4400), .Z(n4382) );
  ANDN U4531 ( .A(n2783), .B(n1872), .Z(n4400) );
  XOR U4532 ( .A(n4401), .B(n4402), .Z(n4380) );
  AND U4533 ( .A(n4403), .B(n4404), .Z(n4402) );
  XOR U4534 ( .A(n4405), .B(n4401), .Z(n4404) );
  XOR U4535 ( .A(n4407), .B(n4408), .Z(n3873) );
  XOR U4536 ( .A(n4409), .B(n4406), .Z(n4407) );
  XNOR U4537 ( .A(n4399), .B(n4398), .Z(n3871) );
  XOR U4538 ( .A(n4410), .B(n4393), .Z(n4398) );
  XNOR U4539 ( .A(n4391), .B(n4411), .Z(n4393) );
  ANDN U4540 ( .A(n3032), .B(n1775), .Z(n4411) );
  XOR U4541 ( .A(n4412), .B(n4413), .Z(n4391) );
  AND U4542 ( .A(n4414), .B(n4415), .Z(n4413) );
  XNOR U4543 ( .A(n4416), .B(n4412), .Z(n4415) );
  XOR U4544 ( .A(n4417), .B(n4395), .Z(n4410) );
  AND U4545 ( .A(n3025), .B(n1773), .Z(n4395) );
  IV U4546 ( .A(n4397), .Z(n4417) );
  XNOR U4547 ( .A(n4403), .B(n4405), .Z(n4399) );
  NAND U4548 ( .A(n2778), .B(n1966), .Z(n4405) );
  XNOR U4549 ( .A(n4401), .B(n4421), .Z(n4403) );
  ANDN U4550 ( .A(n2783), .B(n1968), .Z(n4421) );
  XOR U4551 ( .A(n4422), .B(n4423), .Z(n4401) );
  AND U4552 ( .A(n4424), .B(n4425), .Z(n4423) );
  XOR U4553 ( .A(n4426), .B(n4422), .Z(n4425) );
  XOR U4554 ( .A(n4428), .B(n4429), .Z(n3917) );
  XOR U4555 ( .A(n4430), .B(n4427), .Z(n4428) );
  XNOR U4556 ( .A(n4420), .B(n4419), .Z(n3915) );
  XOR U4557 ( .A(n4431), .B(n4414), .Z(n4419) );
  XNOR U4558 ( .A(n4412), .B(n4432), .Z(n4414) );
  ANDN U4559 ( .A(n3032), .B(n1872), .Z(n4432) );
  XOR U4560 ( .A(n4433), .B(n4434), .Z(n4412) );
  AND U4561 ( .A(n4435), .B(n4436), .Z(n4434) );
  XNOR U4562 ( .A(n4437), .B(n4433), .Z(n4436) );
  XOR U4563 ( .A(n4438), .B(n4416), .Z(n4431) );
  AND U4564 ( .A(n3025), .B(n1870), .Z(n4416) );
  IV U4565 ( .A(n4418), .Z(n4438) );
  XNOR U4566 ( .A(n4424), .B(n4426), .Z(n4420) );
  NAND U4567 ( .A(n2778), .B(n2062), .Z(n4426) );
  XNOR U4568 ( .A(n4422), .B(n4442), .Z(n4424) );
  ANDN U4569 ( .A(n2783), .B(n2064), .Z(n4442) );
  XOR U4570 ( .A(n4443), .B(n4444), .Z(n4422) );
  AND U4571 ( .A(n4445), .B(n4446), .Z(n4444) );
  XOR U4572 ( .A(n4447), .B(n4443), .Z(n4446) );
  XOR U4573 ( .A(n4449), .B(n4450), .Z(n3963) );
  XOR U4574 ( .A(n4451), .B(n4448), .Z(n4449) );
  XNOR U4575 ( .A(n4441), .B(n4440), .Z(n3961) );
  XOR U4576 ( .A(n4452), .B(n4435), .Z(n4440) );
  XNOR U4577 ( .A(n4433), .B(n4453), .Z(n4435) );
  ANDN U4578 ( .A(n3032), .B(n1968), .Z(n4453) );
  XOR U4579 ( .A(n4454), .B(n4455), .Z(n4433) );
  AND U4580 ( .A(n4456), .B(n4457), .Z(n4455) );
  XNOR U4581 ( .A(n4458), .B(n4454), .Z(n4457) );
  XOR U4582 ( .A(n4459), .B(n4437), .Z(n4452) );
  AND U4583 ( .A(n3025), .B(n1966), .Z(n4437) );
  IV U4584 ( .A(n4439), .Z(n4459) );
  XNOR U4585 ( .A(n4445), .B(n4447), .Z(n4441) );
  NAND U4586 ( .A(n2778), .B(n2163), .Z(n4447) );
  XNOR U4587 ( .A(n4443), .B(n4463), .Z(n4445) );
  ANDN U4588 ( .A(n2783), .B(n2165), .Z(n4463) );
  XOR U4589 ( .A(n4464), .B(n4465), .Z(n4443) );
  AND U4590 ( .A(n4466), .B(n4467), .Z(n4465) );
  XOR U4591 ( .A(n4468), .B(n4464), .Z(n4467) );
  XOR U4592 ( .A(n4470), .B(n4471), .Z(n4009) );
  XOR U4593 ( .A(n4472), .B(n4469), .Z(n4470) );
  XNOR U4594 ( .A(n4462), .B(n4461), .Z(n4007) );
  XOR U4595 ( .A(n4473), .B(n4456), .Z(n4461) );
  XNOR U4596 ( .A(n4454), .B(n4474), .Z(n4456) );
  ANDN U4597 ( .A(n3032), .B(n2064), .Z(n4474) );
  XOR U4598 ( .A(n4475), .B(n4476), .Z(n4454) );
  AND U4599 ( .A(n4477), .B(n4478), .Z(n4476) );
  XNOR U4600 ( .A(n4479), .B(n4475), .Z(n4478) );
  XOR U4601 ( .A(n4480), .B(n4458), .Z(n4473) );
  AND U4602 ( .A(n3025), .B(n2062), .Z(n4458) );
  IV U4603 ( .A(n4460), .Z(n4480) );
  XNOR U4604 ( .A(n4466), .B(n4468), .Z(n4462) );
  NAND U4605 ( .A(n2778), .B(n2269), .Z(n4468) );
  XNOR U4606 ( .A(n4464), .B(n4484), .Z(n4466) );
  ANDN U4607 ( .A(n2783), .B(n2271), .Z(n4484) );
  XOR U4608 ( .A(n4485), .B(n4486), .Z(n4464) );
  AND U4609 ( .A(n4487), .B(n4488), .Z(n4486) );
  XOR U4610 ( .A(n4489), .B(n4485), .Z(n4488) );
  XOR U4611 ( .A(n4491), .B(n4492), .Z(n4055) );
  XOR U4612 ( .A(n4493), .B(n4490), .Z(n4491) );
  XNOR U4613 ( .A(n4483), .B(n4482), .Z(n4053) );
  XOR U4614 ( .A(n4494), .B(n4477), .Z(n4482) );
  XNOR U4615 ( .A(n4475), .B(n4495), .Z(n4477) );
  ANDN U4616 ( .A(n3032), .B(n2165), .Z(n4495) );
  XOR U4617 ( .A(n4496), .B(n4497), .Z(n4475) );
  AND U4618 ( .A(n4498), .B(n4499), .Z(n4497) );
  XNOR U4619 ( .A(n4500), .B(n4496), .Z(n4499) );
  XOR U4620 ( .A(n4501), .B(n4479), .Z(n4494) );
  AND U4621 ( .A(n3025), .B(n2163), .Z(n4479) );
  IV U4622 ( .A(n4481), .Z(n4501) );
  XNOR U4623 ( .A(n4487), .B(n4489), .Z(n4483) );
  NAND U4624 ( .A(n2778), .B(n2376), .Z(n4489) );
  XNOR U4625 ( .A(n4485), .B(n4505), .Z(n4487) );
  ANDN U4626 ( .A(n2783), .B(n2378), .Z(n4505) );
  XOR U4627 ( .A(n4506), .B(n4507), .Z(n4485) );
  AND U4628 ( .A(n4508), .B(n4509), .Z(n4507) );
  XOR U4629 ( .A(n4510), .B(n4506), .Z(n4509) );
  XOR U4630 ( .A(n4512), .B(n4513), .Z(n4094) );
  XOR U4631 ( .A(n4514), .B(n4511), .Z(n4512) );
  XNOR U4632 ( .A(n4504), .B(n4503), .Z(n4093) );
  XOR U4633 ( .A(n4515), .B(n4498), .Z(n4503) );
  XNOR U4634 ( .A(n4496), .B(n4516), .Z(n4498) );
  ANDN U4635 ( .A(n3032), .B(n2271), .Z(n4516) );
  AND U4636 ( .A(n3025), .B(n2269), .Z(n4500) );
  XNOR U4637 ( .A(n4508), .B(n4510), .Z(n4504) );
  NAND U4638 ( .A(n2778), .B(n2484), .Z(n4510) );
  XNOR U4639 ( .A(n4506), .B(n4523), .Z(n4508) );
  ANDN U4640 ( .A(n2783), .B(n2486), .Z(n4523) );
  XOR U4641 ( .A(n4527), .B(n4528), .Z(n4511) );
  AND U4642 ( .A(n4529), .B(n4530), .Z(n4528) );
  XOR U4643 ( .A(n4531), .B(n4532), .Z(n4530) );
  XNOR U4644 ( .A(n4527), .B(n4533), .Z(n4532) );
  XNOR U4645 ( .A(n4521), .B(n4534), .Z(n4529) );
  XNOR U4646 ( .A(n4527), .B(n4522), .Z(n4534) );
  XNOR U4647 ( .A(n4525), .B(n4526), .Z(n4522) );
  NAND U4648 ( .A(n2603), .B(n2778), .Z(n4526) );
  XNOR U4649 ( .A(n4524), .B(n4535), .Z(n4525) );
  ANDN U4650 ( .A(n2783), .B(n2605), .Z(n4535) );
  XOR U4651 ( .A(n4539), .B(n4518), .Z(n4521) );
  XNOR U4652 ( .A(n4517), .B(n4540), .Z(n4518) );
  ANDN U4653 ( .A(n3032), .B(n2378), .Z(n4540) );
  AND U4654 ( .A(n3025), .B(n2376), .Z(n4519) );
  XOR U4655 ( .A(n4547), .B(n4548), .Z(n4527) );
  AND U4656 ( .A(n4549), .B(n4550), .Z(n4548) );
  XOR U4657 ( .A(n4551), .B(n4552), .Z(n4550) );
  XNOR U4658 ( .A(n4547), .B(n4553), .Z(n4552) );
  XNOR U4659 ( .A(n4545), .B(n4554), .Z(n4549) );
  XNOR U4660 ( .A(n4547), .B(n4546), .Z(n4554) );
  XNOR U4661 ( .A(n4537), .B(n4538), .Z(n4546) );
  NAND U4662 ( .A(n2723), .B(n2778), .Z(n4538) );
  XNOR U4663 ( .A(n4536), .B(n4555), .Z(n4537) );
  ANDN U4664 ( .A(n2783), .B(n2725), .Z(n4555) );
  XOR U4665 ( .A(n4559), .B(n4542), .Z(n4545) );
  XNOR U4666 ( .A(n4541), .B(n4560), .Z(n4542) );
  ANDN U4667 ( .A(n3032), .B(n2486), .Z(n4560) );
  AND U4668 ( .A(n3025), .B(n2484), .Z(n4543) );
  XOR U4669 ( .A(n4567), .B(n4568), .Z(n4547) );
  AND U4670 ( .A(n4569), .B(n4570), .Z(n4568) );
  XOR U4671 ( .A(n4571), .B(n4572), .Z(n4570) );
  XNOR U4672 ( .A(n4567), .B(n4573), .Z(n4572) );
  XNOR U4673 ( .A(n4565), .B(n4574), .Z(n4569) );
  XNOR U4674 ( .A(n4567), .B(n4566), .Z(n4574) );
  XNOR U4675 ( .A(n4557), .B(n4558), .Z(n4566) );
  NAND U4676 ( .A(n2845), .B(n2778), .Z(n4558) );
  XNOR U4677 ( .A(n4556), .B(n4575), .Z(n4557) );
  ANDN U4678 ( .A(n2783), .B(n2847), .Z(n4575) );
  XOR U4679 ( .A(n4579), .B(n4562), .Z(n4565) );
  XNOR U4680 ( .A(n4561), .B(n4580), .Z(n4562) );
  ANDN U4681 ( .A(n3032), .B(n2605), .Z(n4580) );
  AND U4682 ( .A(n2603), .B(n3025), .Z(n4563) );
  XOR U4683 ( .A(n4587), .B(n4588), .Z(n4567) );
  AND U4684 ( .A(n4589), .B(n4590), .Z(n4588) );
  XOR U4685 ( .A(n4591), .B(n4592), .Z(n4590) );
  XNOR U4686 ( .A(n4587), .B(n4593), .Z(n4592) );
  XNOR U4687 ( .A(n4585), .B(n4594), .Z(n4589) );
  XNOR U4688 ( .A(n4587), .B(n4586), .Z(n4594) );
  XNOR U4689 ( .A(n4577), .B(n4578), .Z(n4586) );
  NAND U4690 ( .A(n2970), .B(n2778), .Z(n4578) );
  XNOR U4691 ( .A(n4576), .B(n4595), .Z(n4577) );
  ANDN U4692 ( .A(n2783), .B(n2972), .Z(n4595) );
  XOR U4693 ( .A(n4599), .B(n4582), .Z(n4585) );
  XNOR U4694 ( .A(n4581), .B(n4600), .Z(n4582) );
  ANDN U4695 ( .A(n3032), .B(n2725), .Z(n4600) );
  AND U4696 ( .A(n2723), .B(n3025), .Z(n4583) );
  XOR U4697 ( .A(n4607), .B(n4608), .Z(n4587) );
  AND U4698 ( .A(n4609), .B(n4610), .Z(n4608) );
  XOR U4699 ( .A(n4611), .B(n4612), .Z(n4610) );
  XNOR U4700 ( .A(n4607), .B(n4613), .Z(n4612) );
  XNOR U4701 ( .A(n4605), .B(n4614), .Z(n4609) );
  XNOR U4702 ( .A(n4607), .B(n4606), .Z(n4614) );
  XNOR U4703 ( .A(n4597), .B(n4598), .Z(n4606) );
  NAND U4704 ( .A(n3102), .B(n2778), .Z(n4598) );
  XNOR U4705 ( .A(n4596), .B(n4615), .Z(n4597) );
  ANDN U4706 ( .A(n2783), .B(n3104), .Z(n4615) );
  XOR U4707 ( .A(n4619), .B(n4602), .Z(n4605) );
  XNOR U4708 ( .A(n4601), .B(n4620), .Z(n4602) );
  ANDN U4709 ( .A(n3032), .B(n2847), .Z(n4620) );
  AND U4710 ( .A(n2845), .B(n3025), .Z(n4603) );
  XOR U4711 ( .A(n4627), .B(n4628), .Z(n4607) );
  AND U4712 ( .A(n4629), .B(n4630), .Z(n4628) );
  XOR U4713 ( .A(n4631), .B(n4632), .Z(n4630) );
  XNOR U4714 ( .A(n4627), .B(n4633), .Z(n4632) );
  XNOR U4715 ( .A(n4625), .B(n4634), .Z(n4629) );
  XNOR U4716 ( .A(n4627), .B(n4626), .Z(n4634) );
  XNOR U4717 ( .A(n4617), .B(n4618), .Z(n4626) );
  NAND U4718 ( .A(n3234), .B(n2778), .Z(n4618) );
  XNOR U4719 ( .A(n4616), .B(n4635), .Z(n4617) );
  ANDN U4720 ( .A(n2783), .B(n3236), .Z(n4635) );
  XOR U4721 ( .A(n4636), .B(n4637), .Z(n4616) );
  AND U4722 ( .A(n4638), .B(n4639), .Z(n4637) );
  XOR U4723 ( .A(n4640), .B(n4636), .Z(n4639) );
  XOR U4724 ( .A(n4641), .B(n4622), .Z(n4625) );
  XNOR U4725 ( .A(n4621), .B(n4642), .Z(n4622) );
  ANDN U4726 ( .A(n3032), .B(n2972), .Z(n4642) );
  XOR U4727 ( .A(n4643), .B(n4644), .Z(n4621) );
  AND U4728 ( .A(n4645), .B(n4646), .Z(n4644) );
  XNOR U4729 ( .A(n4647), .B(n4643), .Z(n4646) );
  AND U4730 ( .A(n2970), .B(n3025), .Z(n4623) );
  XOR U4731 ( .A(n4651), .B(n4652), .Z(n4627) );
  AND U4732 ( .A(n4653), .B(n4654), .Z(n4652) );
  XOR U4733 ( .A(n4655), .B(n4656), .Z(n4654) );
  XNOR U4734 ( .A(n4651), .B(n4657), .Z(n4656) );
  XNOR U4735 ( .A(n4649), .B(n4658), .Z(n4653) );
  XNOR U4736 ( .A(n4651), .B(n4650), .Z(n4658) );
  XNOR U4737 ( .A(n4638), .B(n4640), .Z(n4650) );
  NAND U4738 ( .A(n3370), .B(n2778), .Z(n4640) );
  XNOR U4739 ( .A(n4636), .B(n4659), .Z(n4638) );
  ANDN U4740 ( .A(n2783), .B(n3372), .Z(n4659) );
  XOR U4741 ( .A(n4663), .B(n4645), .Z(n4649) );
  XNOR U4742 ( .A(n4643), .B(n4664), .Z(n4645) );
  ANDN U4743 ( .A(n3032), .B(n3104), .Z(n4664) );
  XOR U4744 ( .A(n4665), .B(n4666), .Z(n4643) );
  AND U4745 ( .A(n4667), .B(n4668), .Z(n4666) );
  XNOR U4746 ( .A(n4669), .B(n4665), .Z(n4668) );
  AND U4747 ( .A(n3102), .B(n3025), .Z(n4647) );
  XOR U4748 ( .A(n4674), .B(n4675), .Z(n4190) );
  XNOR U4749 ( .A(n4672), .B(n4671), .Z(n4189) );
  XOR U4750 ( .A(n4677), .B(n4667), .Z(n4671) );
  XNOR U4751 ( .A(n4665), .B(n4678), .Z(n4667) );
  ANDN U4752 ( .A(n3032), .B(n3236), .Z(n4678) );
  XNOR U4753 ( .A(n4681), .B(n4679), .Z(n4680) );
  ANDN U4754 ( .A(n3032), .B(n3372), .Z(n4681) );
  XNOR U4755 ( .A(n4670), .B(n4669), .Z(n4677) );
  AND U4756 ( .A(n3234), .B(n3025), .Z(n4669) );
  XNOR U4757 ( .A(n4683), .B(n4684), .Z(n4670) );
  NAND U4758 ( .A(n4158), .B(n3025), .Z(n4684) );
  XNOR U4759 ( .A(n4682), .B(n4685), .Z(n4683) );
  ANDN U4760 ( .A(n3032), .B(n4160), .Z(n4685) );
  NAND U4761 ( .A(A[0]), .B(n4686), .Z(n4682) );
  NANDN U4762 ( .B(n3025), .A(n4687), .Z(n4686) );
  NANDN U4763 ( .B(n4163), .A(n3032), .Z(n4687) );
  IV U4764 ( .A(n2899), .Z(n3025) );
  XNOR U4765 ( .A(n4661), .B(n4662), .Z(n4672) );
  NAND U4766 ( .A(n4158), .B(n2778), .Z(n4662) );
  XNOR U4767 ( .A(n4660), .B(n4690), .Z(n4661) );
  ANDN U4768 ( .A(n2783), .B(n4160), .Z(n4690) );
  NAND U4769 ( .A(A[0]), .B(n4691), .Z(n4660) );
  NANDN U4770 ( .B(n2778), .A(n4692), .Z(n4691) );
  NANDN U4771 ( .B(n4163), .A(n2783), .Z(n4692) );
  IV U4772 ( .A(n2657), .Z(n2778) );
  XOR U4773 ( .A(n4695), .B(n4696), .Z(n4673) );
  XOR U4774 ( .A(n3310), .B(n4697), .Z(n3311) );
  AND U4775 ( .A(n4698), .B(n4699), .Z(n4697) );
  NANDN U4776 ( .B(n4700), .A(n876), .Z(n4699) );
  NANDN U4777 ( .B(n4701), .A(n4702), .Z(n4698) );
  XNOR U4778 ( .A(n4195), .B(n4197), .Z(n4216) );
  NAND U4779 ( .A(n3301), .B(n981), .Z(n4197) );
  XNOR U4780 ( .A(n4193), .B(n4704), .Z(n4195) );
  ANDN U4781 ( .A(n3306), .B(n983), .Z(n4704) );
  XOR U4782 ( .A(n4705), .B(n4706), .Z(n4193) );
  AND U4783 ( .A(n4707), .B(n4708), .Z(n4706) );
  XOR U4784 ( .A(n4709), .B(n4705), .Z(n4708) );
  XNOR U4785 ( .A(n4710), .B(n4711), .Z(n4217) );
  IV U4786 ( .A(n4703), .Z(n4711) );
  XOR U4787 ( .A(n4712), .B(n4702), .Z(n4710) );
  AND U4788 ( .A(n4713), .B(n906), .Z(n4702) );
  IV U4789 ( .A(n939), .Z(n906) );
  NAND U4790 ( .A(n4714), .B(n4701), .Z(n4712) );
  XOR U4791 ( .A(n4715), .B(n4716), .Z(n4701) );
  AND U4792 ( .A(n4717), .B(n4718), .Z(n4716) );
  XNOR U4793 ( .A(n4719), .B(n4715), .Z(n4718) );
  NANDN U4794 ( .B(n909), .A(X[0]), .Z(n4714) );
  IV U4795 ( .A(n876), .Z(n909) );
  AND U4796 ( .A(n4720), .B(n4721), .Z(n876) );
  AND U4797 ( .A(A[31]), .B(n4722), .Z(n4720) );
  XNOR U4798 ( .A(n4707), .B(n4709), .Z(n4220) );
  NAND U4799 ( .A(n3301), .B(n1021), .Z(n4709) );
  XNOR U4800 ( .A(n4705), .B(n4724), .Z(n4707) );
  ANDN U4801 ( .A(n3306), .B(n1023), .Z(n4724) );
  XOR U4802 ( .A(n4725), .B(n4726), .Z(n4705) );
  AND U4803 ( .A(n4727), .B(n4728), .Z(n4726) );
  XOR U4804 ( .A(n4729), .B(n4725), .Z(n4728) );
  XNOR U4805 ( .A(n4730), .B(n4717), .Z(n4221) );
  XNOR U4806 ( .A(n4715), .B(n4731), .Z(n4717) );
  ANDN U4807 ( .A(X[0]), .B(n939), .Z(n4731) );
  XOR U4808 ( .A(n4722), .B(A[30]), .Z(n4721) );
  ANDN U4809 ( .A(n4732), .B(n4733), .Z(n4722) );
  XOR U4810 ( .A(n4734), .B(n4735), .Z(n4715) );
  AND U4811 ( .A(n4736), .B(n4737), .Z(n4735) );
  XNOR U4812 ( .A(n4738), .B(n4734), .Z(n4737) );
  XOR U4813 ( .A(n4739), .B(n4719), .Z(n4730) );
  AND U4814 ( .A(n4713), .B(n937), .Z(n4719) );
  IV U4815 ( .A(n983), .Z(n937) );
  IV U4816 ( .A(n4723), .Z(n4739) );
  XNOR U4817 ( .A(n4727), .B(n4729), .Z(n4241) );
  NAND U4818 ( .A(n3301), .B(n1065), .Z(n4729) );
  XNOR U4819 ( .A(n4725), .B(n4741), .Z(n4727) );
  ANDN U4820 ( .A(n3306), .B(n1067), .Z(n4741) );
  XOR U4821 ( .A(n4742), .B(n4743), .Z(n4725) );
  AND U4822 ( .A(n4744), .B(n4745), .Z(n4743) );
  XOR U4823 ( .A(n4746), .B(n4742), .Z(n4745) );
  XNOR U4824 ( .A(n4747), .B(n4736), .Z(n4242) );
  XNOR U4825 ( .A(n4734), .B(n4748), .Z(n4736) );
  ANDN U4826 ( .A(X[0]), .B(n983), .Z(n4748) );
  ANDN U4827 ( .A(n4749), .B(n4750), .Z(n4732) );
  XOR U4828 ( .A(n4751), .B(n4752), .Z(n4734) );
  AND U4829 ( .A(n4753), .B(n4754), .Z(n4752) );
  XNOR U4830 ( .A(n4755), .B(n4751), .Z(n4754) );
  XOR U4831 ( .A(n4756), .B(n4738), .Z(n4747) );
  AND U4832 ( .A(n4713), .B(n981), .Z(n4738) );
  IV U4833 ( .A(n1023), .Z(n981) );
  IV U4834 ( .A(n4740), .Z(n4756) );
  XNOR U4835 ( .A(n4744), .B(n4746), .Z(n4262) );
  NAND U4836 ( .A(n3301), .B(n1107), .Z(n4746) );
  XNOR U4837 ( .A(n4742), .B(n4758), .Z(n4744) );
  ANDN U4838 ( .A(n3306), .B(n1109), .Z(n4758) );
  XOR U4839 ( .A(n4759), .B(n4760), .Z(n4742) );
  AND U4840 ( .A(n4761), .B(n4762), .Z(n4760) );
  XOR U4841 ( .A(n4763), .B(n4759), .Z(n4762) );
  XNOR U4842 ( .A(n4764), .B(n4753), .Z(n4263) );
  XNOR U4843 ( .A(n4751), .B(n4765), .Z(n4753) );
  ANDN U4844 ( .A(X[0]), .B(n1023), .Z(n4765) );
  XNOR U4845 ( .A(n4749), .B(A[28]), .Z(n4750) );
  ANDN U4846 ( .A(n4766), .B(n4767), .Z(n4749) );
  XOR U4847 ( .A(n4768), .B(n4769), .Z(n4751) );
  AND U4848 ( .A(n4770), .B(n4771), .Z(n4769) );
  XNOR U4849 ( .A(n4772), .B(n4768), .Z(n4771) );
  AND U4850 ( .A(n4713), .B(n1021), .Z(n4755) );
  IV U4851 ( .A(n1067), .Z(n1021) );
  XNOR U4852 ( .A(n4761), .B(n4763), .Z(n4282) );
  NAND U4853 ( .A(n3301), .B(n1166), .Z(n4763) );
  XNOR U4854 ( .A(n4759), .B(n4774), .Z(n4761) );
  ANDN U4855 ( .A(n3306), .B(n1168), .Z(n4774) );
  XOR U4856 ( .A(n4775), .B(n4776), .Z(n4759) );
  AND U4857 ( .A(n4777), .B(n4778), .Z(n4776) );
  XOR U4858 ( .A(n4779), .B(n4775), .Z(n4778) );
  XNOR U4859 ( .A(n4780), .B(n4770), .Z(n4283) );
  XNOR U4860 ( .A(n4768), .B(n4781), .Z(n4770) );
  ANDN U4861 ( .A(X[0]), .B(n1067), .Z(n4781) );
  ANDN U4862 ( .A(n4782), .B(n4783), .Z(n4766) );
  XOR U4863 ( .A(n4784), .B(n4785), .Z(n4768) );
  AND U4864 ( .A(n4786), .B(n4787), .Z(n4785) );
  XNOR U4865 ( .A(n4788), .B(n4784), .Z(n4787) );
  AND U4866 ( .A(n4713), .B(n1065), .Z(n4772) );
  IV U4867 ( .A(n1109), .Z(n1065) );
  XNOR U4868 ( .A(n4777), .B(n4779), .Z(n4303) );
  NAND U4869 ( .A(n3301), .B(n1230), .Z(n4779) );
  XNOR U4870 ( .A(n4775), .B(n4790), .Z(n4777) );
  ANDN U4871 ( .A(n3306), .B(n1232), .Z(n4790) );
  XOR U4872 ( .A(n4791), .B(n4792), .Z(n4775) );
  AND U4873 ( .A(n4793), .B(n4794), .Z(n4792) );
  XOR U4874 ( .A(n4795), .B(n4791), .Z(n4794) );
  XNOR U4875 ( .A(n4796), .B(n4786), .Z(n4304) );
  XNOR U4876 ( .A(n4784), .B(n4797), .Z(n4786) );
  ANDN U4877 ( .A(X[0]), .B(n1109), .Z(n4797) );
  XNOR U4878 ( .A(n4782), .B(A[26]), .Z(n4783) );
  ANDN U4879 ( .A(n4798), .B(n4799), .Z(n4782) );
  XOR U4880 ( .A(n4800), .B(n4801), .Z(n4784) );
  AND U4881 ( .A(n4802), .B(n4803), .Z(n4801) );
  XNOR U4882 ( .A(n4804), .B(n4800), .Z(n4803) );
  XOR U4883 ( .A(n4805), .B(n4788), .Z(n4796) );
  AND U4884 ( .A(n4713), .B(n1107), .Z(n4788) );
  IV U4885 ( .A(n1168), .Z(n1107) );
  IV U4886 ( .A(n4789), .Z(n4805) );
  XNOR U4887 ( .A(n4793), .B(n4795), .Z(n4324) );
  NAND U4888 ( .A(n3301), .B(n1298), .Z(n4795) );
  XNOR U4889 ( .A(n4791), .B(n4807), .Z(n4793) );
  ANDN U4890 ( .A(n3306), .B(n1300), .Z(n4807) );
  XOR U4891 ( .A(n4808), .B(n4809), .Z(n4791) );
  AND U4892 ( .A(n4810), .B(n4811), .Z(n4809) );
  XOR U4893 ( .A(n4812), .B(n4808), .Z(n4811) );
  XNOR U4894 ( .A(n4813), .B(n4802), .Z(n4325) );
  XNOR U4895 ( .A(n4800), .B(n4814), .Z(n4802) );
  ANDN U4896 ( .A(X[0]), .B(n1168), .Z(n4814) );
  ANDN U4897 ( .A(n4815), .B(n4816), .Z(n4798) );
  XOR U4898 ( .A(n4817), .B(n4818), .Z(n4800) );
  AND U4899 ( .A(n4819), .B(n4820), .Z(n4818) );
  XNOR U4900 ( .A(n4821), .B(n4817), .Z(n4820) );
  XOR U4901 ( .A(n4822), .B(n4804), .Z(n4813) );
  AND U4902 ( .A(n4713), .B(n1166), .Z(n4804) );
  IV U4903 ( .A(n1232), .Z(n1166) );
  IV U4904 ( .A(n4806), .Z(n4822) );
  XNOR U4905 ( .A(n4810), .B(n4812), .Z(n4345) );
  NAND U4906 ( .A(n3301), .B(n1365), .Z(n4812) );
  XNOR U4907 ( .A(n4808), .B(n4824), .Z(n4810) );
  ANDN U4908 ( .A(n3306), .B(n1367), .Z(n4824) );
  XOR U4909 ( .A(n4825), .B(n4826), .Z(n4808) );
  AND U4910 ( .A(n4827), .B(n4828), .Z(n4826) );
  XOR U4911 ( .A(n4829), .B(n4825), .Z(n4828) );
  XNOR U4912 ( .A(n4830), .B(n4819), .Z(n4346) );
  XNOR U4913 ( .A(n4817), .B(n4831), .Z(n4819) );
  ANDN U4914 ( .A(X[0]), .B(n1232), .Z(n4831) );
  XNOR U4915 ( .A(n4815), .B(A[24]), .Z(n4816) );
  ANDN U4916 ( .A(n4832), .B(n4833), .Z(n4815) );
  XOR U4917 ( .A(n4834), .B(n4835), .Z(n4817) );
  AND U4918 ( .A(n4836), .B(n4837), .Z(n4835) );
  XNOR U4919 ( .A(n4838), .B(n4834), .Z(n4837) );
  XOR U4920 ( .A(n4839), .B(n4821), .Z(n4830) );
  AND U4921 ( .A(n4713), .B(n1230), .Z(n4821) );
  IV U4922 ( .A(n1300), .Z(n1230) );
  IV U4923 ( .A(n4823), .Z(n4839) );
  XNOR U4924 ( .A(n4827), .B(n4829), .Z(n4366) );
  NAND U4925 ( .A(n3301), .B(n1439), .Z(n4829) );
  XNOR U4926 ( .A(n4825), .B(n4841), .Z(n4827) );
  ANDN U4927 ( .A(n3306), .B(n1441), .Z(n4841) );
  XOR U4928 ( .A(n4842), .B(n4843), .Z(n4825) );
  AND U4929 ( .A(n4844), .B(n4845), .Z(n4843) );
  XOR U4930 ( .A(n4846), .B(n4842), .Z(n4845) );
  XNOR U4931 ( .A(n4847), .B(n4836), .Z(n4367) );
  XNOR U4932 ( .A(n4834), .B(n4848), .Z(n4836) );
  ANDN U4933 ( .A(X[0]), .B(n1300), .Z(n4848) );
  ANDN U4934 ( .A(n4849), .B(n4850), .Z(n4832) );
  XOR U4935 ( .A(n4851), .B(n4852), .Z(n4834) );
  AND U4936 ( .A(n4853), .B(n4854), .Z(n4852) );
  XNOR U4937 ( .A(n4855), .B(n4851), .Z(n4854) );
  XOR U4938 ( .A(n4856), .B(n4838), .Z(n4847) );
  AND U4939 ( .A(n4713), .B(n1298), .Z(n4838) );
  IV U4940 ( .A(n1367), .Z(n1298) );
  IV U4941 ( .A(n4840), .Z(n4856) );
  XNOR U4942 ( .A(n4844), .B(n4846), .Z(n4387) );
  NAND U4943 ( .A(n3301), .B(n1517), .Z(n4846) );
  XNOR U4944 ( .A(n4842), .B(n4858), .Z(n4844) );
  ANDN U4945 ( .A(n3306), .B(n1519), .Z(n4858) );
  XOR U4946 ( .A(n4859), .B(n4860), .Z(n4842) );
  AND U4947 ( .A(n4861), .B(n4862), .Z(n4860) );
  XOR U4948 ( .A(n4863), .B(n4859), .Z(n4862) );
  XNOR U4949 ( .A(n4864), .B(n4853), .Z(n4388) );
  XNOR U4950 ( .A(n4851), .B(n4865), .Z(n4853) );
  ANDN U4951 ( .A(X[0]), .B(n1367), .Z(n4865) );
  XNOR U4952 ( .A(n4849), .B(A[22]), .Z(n4850) );
  ANDN U4953 ( .A(n4866), .B(n4867), .Z(n4849) );
  XOR U4954 ( .A(n4868), .B(n4869), .Z(n4851) );
  AND U4955 ( .A(n4870), .B(n4871), .Z(n4869) );
  XNOR U4956 ( .A(n4872), .B(n4868), .Z(n4871) );
  XOR U4957 ( .A(n4873), .B(n4855), .Z(n4864) );
  AND U4958 ( .A(n4713), .B(n1365), .Z(n4855) );
  IV U4959 ( .A(n1441), .Z(n1365) );
  IV U4960 ( .A(n4857), .Z(n4873) );
  XNOR U4961 ( .A(n4861), .B(n4863), .Z(n4408) );
  NAND U4962 ( .A(n3301), .B(n1598), .Z(n4863) );
  XNOR U4963 ( .A(n4859), .B(n4875), .Z(n4861) );
  ANDN U4964 ( .A(n3306), .B(n1600), .Z(n4875) );
  XOR U4965 ( .A(n4876), .B(n4877), .Z(n4859) );
  AND U4966 ( .A(n4878), .B(n4879), .Z(n4877) );
  XOR U4967 ( .A(n4880), .B(n4876), .Z(n4879) );
  XNOR U4968 ( .A(n4881), .B(n4870), .Z(n4409) );
  XNOR U4969 ( .A(n4868), .B(n4882), .Z(n4870) );
  ANDN U4970 ( .A(X[0]), .B(n1441), .Z(n4882) );
  ANDN U4971 ( .A(n4883), .B(n4884), .Z(n4866) );
  XOR U4972 ( .A(n4885), .B(n4886), .Z(n4868) );
  AND U4973 ( .A(n4887), .B(n4888), .Z(n4886) );
  XNOR U4974 ( .A(n4889), .B(n4885), .Z(n4888) );
  XOR U4975 ( .A(n4890), .B(n4872), .Z(n4881) );
  AND U4976 ( .A(n4713), .B(n1439), .Z(n4872) );
  IV U4977 ( .A(n1519), .Z(n1439) );
  IV U4978 ( .A(n4874), .Z(n4890) );
  XNOR U4979 ( .A(n4878), .B(n4880), .Z(n4429) );
  NAND U4980 ( .A(n3301), .B(n1682), .Z(n4880) );
  XNOR U4981 ( .A(n4876), .B(n4892), .Z(n4878) );
  ANDN U4982 ( .A(n3306), .B(n1684), .Z(n4892) );
  XOR U4983 ( .A(n4893), .B(n4894), .Z(n4876) );
  AND U4984 ( .A(n4895), .B(n4896), .Z(n4894) );
  XOR U4985 ( .A(n4897), .B(n4893), .Z(n4896) );
  XNOR U4986 ( .A(n4898), .B(n4887), .Z(n4430) );
  XNOR U4987 ( .A(n4885), .B(n4899), .Z(n4887) );
  ANDN U4988 ( .A(X[0]), .B(n1519), .Z(n4899) );
  XNOR U4989 ( .A(n4883), .B(A[20]), .Z(n4884) );
  ANDN U4990 ( .A(n4900), .B(n4901), .Z(n4883) );
  XOR U4991 ( .A(n4902), .B(n4903), .Z(n4885) );
  AND U4992 ( .A(n4904), .B(n4905), .Z(n4903) );
  XNOR U4993 ( .A(n4906), .B(n4902), .Z(n4905) );
  XOR U4994 ( .A(n4907), .B(n4889), .Z(n4898) );
  AND U4995 ( .A(n4713), .B(n1517), .Z(n4889) );
  IV U4996 ( .A(n1600), .Z(n1517) );
  IV U4997 ( .A(n4891), .Z(n4907) );
  XNOR U4998 ( .A(n4895), .B(n4897), .Z(n4450) );
  NAND U4999 ( .A(n3301), .B(n1773), .Z(n4897) );
  XNOR U5000 ( .A(n4893), .B(n4909), .Z(n4895) );
  ANDN U5001 ( .A(n3306), .B(n1775), .Z(n4909) );
  XOR U5002 ( .A(n4910), .B(n4911), .Z(n4893) );
  AND U5003 ( .A(n4912), .B(n4913), .Z(n4911) );
  XOR U5004 ( .A(n4914), .B(n4910), .Z(n4913) );
  XNOR U5005 ( .A(n4915), .B(n4904), .Z(n4451) );
  XNOR U5006 ( .A(n4902), .B(n4916), .Z(n4904) );
  ANDN U5007 ( .A(X[0]), .B(n1600), .Z(n4916) );
  ANDN U5008 ( .A(n4917), .B(n4918), .Z(n4900) );
  XOR U5009 ( .A(n4919), .B(n4920), .Z(n4902) );
  AND U5010 ( .A(n4921), .B(n4922), .Z(n4920) );
  XNOR U5011 ( .A(n4923), .B(n4919), .Z(n4922) );
  XOR U5012 ( .A(n4924), .B(n4906), .Z(n4915) );
  AND U5013 ( .A(n4713), .B(n1598), .Z(n4906) );
  IV U5014 ( .A(n1684), .Z(n1598) );
  IV U5015 ( .A(n4908), .Z(n4924) );
  XNOR U5016 ( .A(n4912), .B(n4914), .Z(n4471) );
  NAND U5017 ( .A(n3301), .B(n1870), .Z(n4914) );
  XNOR U5018 ( .A(n4910), .B(n4926), .Z(n4912) );
  ANDN U5019 ( .A(n3306), .B(n1872), .Z(n4926) );
  XOR U5020 ( .A(n4927), .B(n4928), .Z(n4910) );
  AND U5021 ( .A(n4929), .B(n4930), .Z(n4928) );
  XOR U5022 ( .A(n4931), .B(n4927), .Z(n4930) );
  XNOR U5023 ( .A(n4932), .B(n4921), .Z(n4472) );
  XNOR U5024 ( .A(n4919), .B(n4933), .Z(n4921) );
  ANDN U5025 ( .A(X[0]), .B(n1684), .Z(n4933) );
  XNOR U5026 ( .A(n4917), .B(A[18]), .Z(n4918) );
  ANDN U5027 ( .A(n4934), .B(n4935), .Z(n4917) );
  XOR U5028 ( .A(n4936), .B(n4937), .Z(n4919) );
  AND U5029 ( .A(n4938), .B(n4939), .Z(n4937) );
  XNOR U5030 ( .A(n4940), .B(n4936), .Z(n4939) );
  XOR U5031 ( .A(n4941), .B(n4923), .Z(n4932) );
  AND U5032 ( .A(n4713), .B(n1682), .Z(n4923) );
  IV U5033 ( .A(n1775), .Z(n1682) );
  IV U5034 ( .A(n4925), .Z(n4941) );
  XNOR U5035 ( .A(n4929), .B(n4931), .Z(n4492) );
  NAND U5036 ( .A(n3301), .B(n1966), .Z(n4931) );
  XNOR U5037 ( .A(n4927), .B(n4943), .Z(n4929) );
  ANDN U5038 ( .A(n3306), .B(n1968), .Z(n4943) );
  XOR U5039 ( .A(n4944), .B(n4945), .Z(n4927) );
  AND U5040 ( .A(n4946), .B(n4947), .Z(n4945) );
  XOR U5041 ( .A(n4948), .B(n4944), .Z(n4947) );
  XNOR U5042 ( .A(n4949), .B(n4938), .Z(n4493) );
  XNOR U5043 ( .A(n4936), .B(n4950), .Z(n4938) );
  ANDN U5044 ( .A(X[0]), .B(n1775), .Z(n4950) );
  ANDN U5045 ( .A(n4951), .B(n4952), .Z(n4934) );
  XOR U5046 ( .A(n4953), .B(n4954), .Z(n4936) );
  AND U5047 ( .A(n4955), .B(n4956), .Z(n4954) );
  XNOR U5048 ( .A(n4957), .B(n4953), .Z(n4956) );
  XOR U5049 ( .A(n4958), .B(n4940), .Z(n4949) );
  AND U5050 ( .A(n4713), .B(n1773), .Z(n4940) );
  IV U5051 ( .A(n1872), .Z(n1773) );
  IV U5052 ( .A(n4942), .Z(n4958) );
  XNOR U5053 ( .A(n4946), .B(n4948), .Z(n4513) );
  NAND U5054 ( .A(n3301), .B(n2062), .Z(n4948) );
  XNOR U5055 ( .A(n4944), .B(n4960), .Z(n4946) );
  ANDN U5056 ( .A(n3306), .B(n2064), .Z(n4960) );
  XNOR U5057 ( .A(n4964), .B(n4955), .Z(n4514) );
  XNOR U5058 ( .A(n4953), .B(n4965), .Z(n4955) );
  ANDN U5059 ( .A(X[0]), .B(n1872), .Z(n4965) );
  AND U5060 ( .A(n4713), .B(n1870), .Z(n4957) );
  XNOR U5061 ( .A(n4962), .B(n4963), .Z(n4531) );
  NAND U5062 ( .A(n3301), .B(n2163), .Z(n4963) );
  XNOR U5063 ( .A(n4961), .B(n4970), .Z(n4962) );
  ANDN U5064 ( .A(n3306), .B(n2165), .Z(n4970) );
  XNOR U5065 ( .A(n4974), .B(n4967), .Z(n4533) );
  XNOR U5066 ( .A(n4966), .B(n4975), .Z(n4967) );
  ANDN U5067 ( .A(X[0]), .B(n1968), .Z(n4975) );
  AND U5068 ( .A(n4713), .B(n1966), .Z(n4968) );
  XNOR U5069 ( .A(n4972), .B(n4973), .Z(n4551) );
  NAND U5070 ( .A(n3301), .B(n2269), .Z(n4973) );
  XNOR U5071 ( .A(n4971), .B(n4980), .Z(n4972) );
  ANDN U5072 ( .A(n3306), .B(n2271), .Z(n4980) );
  XNOR U5073 ( .A(n4984), .B(n4977), .Z(n4553) );
  XNOR U5074 ( .A(n4976), .B(n4985), .Z(n4977) );
  ANDN U5075 ( .A(X[0]), .B(n2064), .Z(n4985) );
  AND U5076 ( .A(n4713), .B(n2062), .Z(n4978) );
  XNOR U5077 ( .A(n4982), .B(n4983), .Z(n4571) );
  NAND U5078 ( .A(n3301), .B(n2376), .Z(n4983) );
  XNOR U5079 ( .A(n4981), .B(n4990), .Z(n4982) );
  ANDN U5080 ( .A(n3306), .B(n2378), .Z(n4990) );
  XNOR U5081 ( .A(n4994), .B(n4987), .Z(n4573) );
  XNOR U5082 ( .A(n4986), .B(n4995), .Z(n4987) );
  ANDN U5083 ( .A(X[0]), .B(n2165), .Z(n4995) );
  XOR U5084 ( .A(n4996), .B(n4997), .Z(n4986) );
  AND U5085 ( .A(n4998), .B(n4999), .Z(n4997) );
  XNOR U5086 ( .A(n5000), .B(n4996), .Z(n4999) );
  AND U5087 ( .A(n4713), .B(n2163), .Z(n4988) );
  XNOR U5088 ( .A(n4992), .B(n4993), .Z(n4591) );
  NAND U5089 ( .A(n3301), .B(n2484), .Z(n4993) );
  XNOR U5090 ( .A(n4991), .B(n5002), .Z(n4992) );
  ANDN U5091 ( .A(n3306), .B(n2486), .Z(n5002) );
  XOR U5092 ( .A(n5003), .B(n5004), .Z(n4991) );
  AND U5093 ( .A(n5005), .B(n5006), .Z(n5004) );
  XOR U5094 ( .A(n5007), .B(n5003), .Z(n5006) );
  XNOR U5095 ( .A(n5008), .B(n4998), .Z(n4593) );
  XNOR U5096 ( .A(n4996), .B(n5009), .Z(n4998) );
  ANDN U5097 ( .A(X[0]), .B(n2271), .Z(n5009) );
  XOR U5098 ( .A(n5010), .B(n5011), .Z(n4996) );
  AND U5099 ( .A(n5012), .B(n5013), .Z(n5011) );
  XNOR U5100 ( .A(n5014), .B(n5010), .Z(n5013) );
  XOR U5101 ( .A(n5015), .B(n5000), .Z(n5008) );
  AND U5102 ( .A(n4713), .B(n2269), .Z(n5000) );
  IV U5103 ( .A(n5001), .Z(n5015) );
  XNOR U5104 ( .A(n5005), .B(n5007), .Z(n4611) );
  NAND U5105 ( .A(n3301), .B(n2603), .Z(n5007) );
  XNOR U5106 ( .A(n5003), .B(n5017), .Z(n5005) );
  ANDN U5107 ( .A(n3306), .B(n2605), .Z(n5017) );
  XOR U5108 ( .A(n5018), .B(n5019), .Z(n5003) );
  AND U5109 ( .A(n5020), .B(n5021), .Z(n5019) );
  XOR U5110 ( .A(n5022), .B(n5018), .Z(n5021) );
  XNOR U5111 ( .A(n5023), .B(n5012), .Z(n4613) );
  XNOR U5112 ( .A(n5010), .B(n5024), .Z(n5012) );
  ANDN U5113 ( .A(X[0]), .B(n2378), .Z(n5024) );
  XOR U5114 ( .A(n5025), .B(n5026), .Z(n5010) );
  AND U5115 ( .A(n5027), .B(n5028), .Z(n5026) );
  XNOR U5116 ( .A(n5029), .B(n5025), .Z(n5028) );
  XOR U5117 ( .A(n5030), .B(n5014), .Z(n5023) );
  AND U5118 ( .A(n4713), .B(n2376), .Z(n5014) );
  IV U5119 ( .A(n5016), .Z(n5030) );
  XNOR U5120 ( .A(n5020), .B(n5022), .Z(n4631) );
  NAND U5121 ( .A(n3301), .B(n2723), .Z(n5022) );
  XNOR U5122 ( .A(n5018), .B(n5032), .Z(n5020) );
  ANDN U5123 ( .A(n3306), .B(n2725), .Z(n5032) );
  XNOR U5124 ( .A(n5036), .B(n5027), .Z(n4633) );
  XNOR U5125 ( .A(n5025), .B(n5037), .Z(n5027) );
  ANDN U5126 ( .A(X[0]), .B(n2486), .Z(n5037) );
  XOR U5127 ( .A(n5038), .B(n5039), .Z(n5025) );
  AND U5128 ( .A(n5040), .B(n5041), .Z(n5039) );
  XNOR U5129 ( .A(n5042), .B(n5038), .Z(n5041) );
  AND U5130 ( .A(n4713), .B(n2484), .Z(n5029) );
  XNOR U5131 ( .A(n5034), .B(n5035), .Z(n4655) );
  NAND U5132 ( .A(n3301), .B(n2845), .Z(n5035) );
  XNOR U5133 ( .A(n5033), .B(n5044), .Z(n5034) );
  ANDN U5134 ( .A(n3306), .B(n2847), .Z(n5044) );
  XNOR U5135 ( .A(n5048), .B(n5040), .Z(n4657) );
  XNOR U5136 ( .A(n5038), .B(n5049), .Z(n5040) );
  ANDN U5137 ( .A(X[0]), .B(n2605), .Z(n5049) );
  XOR U5138 ( .A(n5050), .B(n5051), .Z(n5038) );
  AND U5139 ( .A(n5052), .B(n5053), .Z(n5051) );
  XNOR U5140 ( .A(n5054), .B(n5050), .Z(n5053) );
  AND U5141 ( .A(n4713), .B(n2603), .Z(n5042) );
  XNOR U5142 ( .A(n5046), .B(n5047), .Z(n4675) );
  NAND U5143 ( .A(n3301), .B(n2970), .Z(n5047) );
  XNOR U5144 ( .A(n5045), .B(n5056), .Z(n5046) );
  ANDN U5145 ( .A(n3306), .B(n2972), .Z(n5056) );
  XNOR U5146 ( .A(n5060), .B(n5052), .Z(n4676) );
  XNOR U5147 ( .A(n5050), .B(n5061), .Z(n5052) );
  ANDN U5148 ( .A(X[0]), .B(n2725), .Z(n5061) );
  AND U5149 ( .A(n4713), .B(n2723), .Z(n5054) );
  XNOR U5150 ( .A(n5065), .B(n5066), .Z(n5055) );
  AND U5151 ( .A(n5067), .B(n5068), .Z(n5066) );
  XNOR U5152 ( .A(n5063), .B(n5069), .Z(n5068) );
  XNOR U5153 ( .A(n5064), .B(n5065), .Z(n5069) );
  AND U5154 ( .A(n4713), .B(n2845), .Z(n5064) );
  XOR U5155 ( .A(n5062), .B(n5070), .Z(n5063) );
  ANDN U5156 ( .A(X[0]), .B(n2847), .Z(n5070) );
  XNOR U5157 ( .A(n5058), .B(n5074), .Z(n5067) );
  XNOR U5158 ( .A(n5059), .B(n5065), .Z(n5074) );
  AND U5159 ( .A(n3102), .B(n3301), .Z(n5059) );
  XOR U5160 ( .A(n5057), .B(n5075), .Z(n5058) );
  ANDN U5161 ( .A(n3306), .B(n3104), .Z(n5075) );
  XOR U5162 ( .A(n5079), .B(n5080), .Z(n5065) );
  AND U5163 ( .A(n5081), .B(n5082), .Z(n5080) );
  XNOR U5164 ( .A(n5072), .B(n5083), .Z(n5082) );
  XNOR U5165 ( .A(n5073), .B(n5079), .Z(n5083) );
  AND U5166 ( .A(n4713), .B(n2970), .Z(n5073) );
  XOR U5167 ( .A(n5071), .B(n5084), .Z(n5072) );
  ANDN U5168 ( .A(X[0]), .B(n2972), .Z(n5084) );
  XNOR U5169 ( .A(n5077), .B(n5088), .Z(n5081) );
  XNOR U5170 ( .A(n5078), .B(n5079), .Z(n5088) );
  AND U5171 ( .A(n3234), .B(n3301), .Z(n5078) );
  XOR U5172 ( .A(n5076), .B(n5089), .Z(n5077) );
  ANDN U5173 ( .A(n3306), .B(n3236), .Z(n5089) );
  XOR U5174 ( .A(n5090), .B(n5091), .Z(n5076) );
  ANDN U5175 ( .A(n5092), .B(n5093), .Z(n5091) );
  XNOR U5176 ( .A(n5094), .B(n5090), .Z(n5092) );
  XOR U5177 ( .A(n5095), .B(n5096), .Z(n5079) );
  AND U5178 ( .A(n5097), .B(n5098), .Z(n5096) );
  XNOR U5179 ( .A(n5086), .B(n5099), .Z(n5098) );
  XNOR U5180 ( .A(n5087), .B(n5095), .Z(n5099) );
  AND U5181 ( .A(n4713), .B(n3102), .Z(n5087) );
  XOR U5182 ( .A(n5085), .B(n5100), .Z(n5086) );
  ANDN U5183 ( .A(X[0]), .B(n3104), .Z(n5100) );
  XNOR U5184 ( .A(n5093), .B(n5104), .Z(n5097) );
  XNOR U5185 ( .A(n5094), .B(n5095), .Z(n5104) );
  AND U5186 ( .A(n3370), .B(n3301), .Z(n5094) );
  XOR U5187 ( .A(n5090), .B(n5105), .Z(n5093) );
  ANDN U5188 ( .A(n3306), .B(n3372), .Z(n5105) );
  XNOR U5189 ( .A(n5110), .B(n5102), .Z(n4696) );
  XNOR U5190 ( .A(n5101), .B(n5111), .Z(n5102) );
  ANDN U5191 ( .A(X[0]), .B(n3236), .Z(n5111) );
  XNOR U5192 ( .A(n5114), .B(n5112), .Z(n5113) );
  ANDN U5193 ( .A(X[0]), .B(n3372), .Z(n5114) );
  ANDN U5194 ( .A(n4713), .B(n4160), .Z(n5115) );
  XNOR U5195 ( .A(n5109), .B(n5103), .Z(n5110) );
  AND U5196 ( .A(n4713), .B(n3234), .Z(n5103) );
  XNOR U5197 ( .A(n5107), .B(n5108), .Z(n4695) );
  NAND U5198 ( .A(n4158), .B(n3301), .Z(n5108) );
  XNOR U5199 ( .A(n5106), .B(n5119), .Z(n5107) );
  ANDN U5200 ( .A(n3306), .B(n4160), .Z(n5119) );
  NAND U5201 ( .A(A[0]), .B(n5120), .Z(n5106) );
  NANDN U5202 ( .B(n3301), .A(n5121), .Z(n5120) );
  NANDN U5203 ( .B(n4163), .A(n3306), .Z(n5121) );
  IV U5204 ( .A(n3172), .Z(n3301) );
  XNOR U5205 ( .A(n5117), .B(n5118), .Z(n5109) );
  NAND U5206 ( .A(n4158), .B(n4713), .Z(n5118) );
  XNOR U5207 ( .A(n5116), .B(n5124), .Z(n5117) );
  ANDN U5208 ( .A(X[0]), .B(n4160), .Z(n5124) );
  NAND U5209 ( .A(A[0]), .B(n5125), .Z(n5116) );
  NANDN U5210 ( .B(n4713), .A(n5126), .Z(n5125) );
  NANDN U5211 ( .B(n4163), .A(X[0]), .Z(n5126) );
  IV U5212 ( .A(n4700), .Z(n4713) );
  XNOR U5213 ( .A(n3329), .B(n3328), .Z(n3282) );
  XOR U5214 ( .A(n5128), .B(n3337), .Z(n3328) );
  XNOR U5215 ( .A(n3322), .B(n3321), .Z(n3337) );
  XOR U5216 ( .A(n5129), .B(n3318), .Z(n3321) );
  XNOR U5217 ( .A(n3317), .B(n5130), .Z(n3318) );
  ANDN U5218 ( .A(n1386), .B(n2271), .Z(n5130) );
  AND U5219 ( .A(n2269), .B(n1323), .Z(n3319) );
  XNOR U5220 ( .A(n3325), .B(n3326), .Z(n3322) );
  NANDN U5221 ( .B(n1188), .A(n2484), .Z(n3326) );
  XNOR U5222 ( .A(n3324), .B(n5137), .Z(n3325) );
  ANDN U5223 ( .A(n1258), .B(n2486), .Z(n5137) );
  XOR U5224 ( .A(n3336), .B(n3327), .Z(n5128) );
  XNOR U5225 ( .A(n5141), .B(n5142), .Z(n3327) );
  XOR U5226 ( .A(n5143), .B(n3345), .Z(n3336) );
  XNOR U5227 ( .A(n3333), .B(n3334), .Z(n3345) );
  NAND U5228 ( .A(n2062), .B(n1557), .Z(n3334) );
  XNOR U5229 ( .A(n3332), .B(n5144), .Z(n3333) );
  ANDN U5230 ( .A(n1564), .B(n2064), .Z(n5144) );
  XNOR U5231 ( .A(n3344), .B(n3335), .Z(n5143) );
  XOR U5232 ( .A(n5148), .B(n5149), .Z(n3335) );
  AND U5233 ( .A(n5150), .B(n5151), .Z(n5149) );
  XOR U5234 ( .A(n5152), .B(n5153), .Z(n5151) );
  XNOR U5235 ( .A(n5148), .B(n5154), .Z(n5153) );
  XNOR U5236 ( .A(n5135), .B(n5155), .Z(n5150) );
  XNOR U5237 ( .A(n5148), .B(n5136), .Z(n5155) );
  XNOR U5238 ( .A(n5139), .B(n5140), .Z(n5136) );
  NANDN U5239 ( .B(n1188), .A(n2603), .Z(n5140) );
  XNOR U5240 ( .A(n5138), .B(n5156), .Z(n5139) );
  ANDN U5241 ( .A(n1258), .B(n2605), .Z(n5156) );
  XOR U5242 ( .A(n5160), .B(n5132), .Z(n5135) );
  XNOR U5243 ( .A(n5131), .B(n5161), .Z(n5132) );
  ANDN U5244 ( .A(n1386), .B(n2378), .Z(n5161) );
  AND U5245 ( .A(n2376), .B(n1323), .Z(n5133) );
  XOR U5246 ( .A(n5168), .B(n5169), .Z(n5148) );
  AND U5247 ( .A(n5170), .B(n5171), .Z(n5169) );
  XOR U5248 ( .A(n5172), .B(n5173), .Z(n5171) );
  XNOR U5249 ( .A(n5168), .B(n5174), .Z(n5173) );
  XNOR U5250 ( .A(n5166), .B(n5175), .Z(n5170) );
  XNOR U5251 ( .A(n5168), .B(n5167), .Z(n5175) );
  XNOR U5252 ( .A(n5158), .B(n5159), .Z(n5167) );
  NANDN U5253 ( .B(n1188), .A(n2723), .Z(n5159) );
  XNOR U5254 ( .A(n5157), .B(n5176), .Z(n5158) );
  ANDN U5255 ( .A(n1258), .B(n2725), .Z(n5176) );
  XOR U5256 ( .A(n5180), .B(n5163), .Z(n5166) );
  XNOR U5257 ( .A(n5162), .B(n5181), .Z(n5163) );
  ANDN U5258 ( .A(n1386), .B(n2486), .Z(n5181) );
  AND U5259 ( .A(n2484), .B(n1323), .Z(n5164) );
  XOR U5260 ( .A(n5188), .B(n5189), .Z(n5168) );
  AND U5261 ( .A(n5190), .B(n5191), .Z(n5189) );
  XOR U5262 ( .A(n5192), .B(n5193), .Z(n5191) );
  XNOR U5263 ( .A(n5188), .B(n5194), .Z(n5193) );
  XNOR U5264 ( .A(n5186), .B(n5195), .Z(n5190) );
  XNOR U5265 ( .A(n5188), .B(n5187), .Z(n5195) );
  XNOR U5266 ( .A(n5178), .B(n5179), .Z(n5187) );
  NANDN U5267 ( .B(n1188), .A(n2845), .Z(n5179) );
  XNOR U5268 ( .A(n5177), .B(n5196), .Z(n5178) );
  ANDN U5269 ( .A(n1258), .B(n2847), .Z(n5196) );
  XOR U5270 ( .A(n5200), .B(n5183), .Z(n5186) );
  XNOR U5271 ( .A(n5182), .B(n5201), .Z(n5183) );
  ANDN U5272 ( .A(n1386), .B(n2605), .Z(n5201) );
  AND U5273 ( .A(n2603), .B(n1323), .Z(n5184) );
  XOR U5274 ( .A(n5208), .B(n5209), .Z(n5188) );
  AND U5275 ( .A(n5210), .B(n5211), .Z(n5209) );
  XOR U5276 ( .A(n5212), .B(n5213), .Z(n5211) );
  XNOR U5277 ( .A(n5208), .B(n5214), .Z(n5213) );
  XNOR U5278 ( .A(n5206), .B(n5215), .Z(n5210) );
  XNOR U5279 ( .A(n5208), .B(n5207), .Z(n5215) );
  XNOR U5280 ( .A(n5198), .B(n5199), .Z(n5207) );
  NANDN U5281 ( .B(n1188), .A(n2970), .Z(n5199) );
  XNOR U5282 ( .A(n5197), .B(n5216), .Z(n5198) );
  ANDN U5283 ( .A(n1258), .B(n2972), .Z(n5216) );
  XOR U5284 ( .A(n5220), .B(n5203), .Z(n5206) );
  XNOR U5285 ( .A(n5202), .B(n5221), .Z(n5203) );
  ANDN U5286 ( .A(n1386), .B(n2725), .Z(n5221) );
  AND U5287 ( .A(n2723), .B(n1323), .Z(n5204) );
  XOR U5288 ( .A(n5228), .B(n5229), .Z(n5208) );
  AND U5289 ( .A(n5230), .B(n5231), .Z(n5229) );
  XOR U5290 ( .A(n5232), .B(n5233), .Z(n5231) );
  XNOR U5291 ( .A(n5228), .B(n5234), .Z(n5233) );
  XNOR U5292 ( .A(n5226), .B(n5235), .Z(n5230) );
  XNOR U5293 ( .A(n5228), .B(n5227), .Z(n5235) );
  XNOR U5294 ( .A(n5218), .B(n5219), .Z(n5227) );
  NANDN U5295 ( .B(n1188), .A(n3102), .Z(n5219) );
  XNOR U5296 ( .A(n5217), .B(n5236), .Z(n5218) );
  ANDN U5297 ( .A(n1258), .B(n3104), .Z(n5236) );
  XOR U5298 ( .A(n5240), .B(n5223), .Z(n5226) );
  XNOR U5299 ( .A(n5222), .B(n5241), .Z(n5223) );
  ANDN U5300 ( .A(n1386), .B(n2847), .Z(n5241) );
  XOR U5301 ( .A(n5242), .B(n5243), .Z(n5222) );
  AND U5302 ( .A(n5244), .B(n5245), .Z(n5243) );
  XNOR U5303 ( .A(n5246), .B(n5242), .Z(n5245) );
  AND U5304 ( .A(n2845), .B(n1323), .Z(n5224) );
  XOR U5305 ( .A(n5250), .B(n5251), .Z(n5228) );
  AND U5306 ( .A(n5252), .B(n5253), .Z(n5251) );
  XOR U5307 ( .A(n5254), .B(n5255), .Z(n5253) );
  XNOR U5308 ( .A(n5250), .B(n5256), .Z(n5255) );
  XNOR U5309 ( .A(n5248), .B(n5257), .Z(n5252) );
  XNOR U5310 ( .A(n5250), .B(n5249), .Z(n5257) );
  XNOR U5311 ( .A(n5238), .B(n5239), .Z(n5249) );
  NANDN U5312 ( .B(n1188), .A(n3234), .Z(n5239) );
  XNOR U5313 ( .A(n5237), .B(n5258), .Z(n5238) );
  ANDN U5314 ( .A(n1258), .B(n3236), .Z(n5258) );
  XOR U5315 ( .A(n5259), .B(n5260), .Z(n5237) );
  AND U5316 ( .A(n5261), .B(n5262), .Z(n5260) );
  XOR U5317 ( .A(n5263), .B(n5259), .Z(n5262) );
  XOR U5318 ( .A(n5264), .B(n5244), .Z(n5248) );
  XNOR U5319 ( .A(n5242), .B(n5265), .Z(n5244) );
  ANDN U5320 ( .A(n1386), .B(n2972), .Z(n5265) );
  XOR U5321 ( .A(n5266), .B(n5267), .Z(n5242) );
  AND U5322 ( .A(n5268), .B(n5269), .Z(n5267) );
  XNOR U5323 ( .A(n5270), .B(n5266), .Z(n5269) );
  AND U5324 ( .A(n2970), .B(n1323), .Z(n5246) );
  XOR U5325 ( .A(n5274), .B(n5275), .Z(n5250) );
  AND U5326 ( .A(n5276), .B(n5277), .Z(n5275) );
  XOR U5327 ( .A(n5278), .B(n5279), .Z(n5277) );
  XNOR U5328 ( .A(n5274), .B(n5280), .Z(n5279) );
  XNOR U5329 ( .A(n5272), .B(n5281), .Z(n5276) );
  XNOR U5330 ( .A(n5274), .B(n5273), .Z(n5281) );
  XNOR U5331 ( .A(n5261), .B(n5263), .Z(n5273) );
  NANDN U5332 ( .B(n1188), .A(n3370), .Z(n5263) );
  XNOR U5333 ( .A(n5259), .B(n5282), .Z(n5261) );
  ANDN U5334 ( .A(n1258), .B(n3372), .Z(n5282) );
  XOR U5335 ( .A(n5286), .B(n5268), .Z(n5272) );
  XNOR U5336 ( .A(n5266), .B(n5287), .Z(n5268) );
  ANDN U5337 ( .A(n1386), .B(n3104), .Z(n5287) );
  AND U5338 ( .A(n3102), .B(n1323), .Z(n5270) );
  XOR U5339 ( .A(n5295), .B(n5296), .Z(n5142) );
  XNOR U5340 ( .A(n5293), .B(n5292), .Z(n5141) );
  XOR U5341 ( .A(n5298), .B(n5289), .Z(n5292) );
  XNOR U5342 ( .A(n5288), .B(n5299), .Z(n5289) );
  ANDN U5343 ( .A(n1386), .B(n3236), .Z(n5299) );
  XNOR U5344 ( .A(n5302), .B(n5300), .Z(n5301) );
  ANDN U5345 ( .A(n1386), .B(n3372), .Z(n5302) );
  XNOR U5346 ( .A(n5291), .B(n5290), .Z(n5298) );
  AND U5347 ( .A(n3234), .B(n1323), .Z(n5290) );
  XNOR U5348 ( .A(n5305), .B(n5306), .Z(n5291) );
  NAND U5349 ( .A(n4158), .B(n1323), .Z(n5306) );
  XNOR U5350 ( .A(n5304), .B(n5307), .Z(n5305) );
  ANDN U5351 ( .A(n1386), .B(n4160), .Z(n5307) );
  NAND U5352 ( .A(A[0]), .B(n5308), .Z(n5304) );
  NANDN U5353 ( .B(n1323), .A(n5309), .Z(n5308) );
  NANDN U5354 ( .B(n4163), .A(n1386), .Z(n5309) );
  IV U5355 ( .A(n5303), .Z(n1323) );
  XNOR U5356 ( .A(n5284), .B(n5285), .Z(n5293) );
  NANDN U5357 ( .B(n1188), .A(n4158), .Z(n5285) );
  XNOR U5358 ( .A(n5283), .B(n5312), .Z(n5284) );
  ANDN U5359 ( .A(n1258), .B(n4160), .Z(n5312) );
  NAND U5360 ( .A(A[0]), .B(n5313), .Z(n5283) );
  NAND U5361 ( .A(n5314), .B(n1188), .Z(n5313) );
  NANDN U5362 ( .B(n4163), .A(n1258), .Z(n5314) );
  XOR U5363 ( .A(n5317), .B(n5318), .Z(n5294) );
  XOR U5364 ( .A(n5319), .B(n3341), .Z(n3344) );
  XNOR U5365 ( .A(n3340), .B(n5320), .Z(n3341) );
  ANDN U5366 ( .A(n1748), .B(n1872), .Z(n5320) );
  XNOR U5367 ( .A(n4951), .B(A[16]), .Z(n4952) );
  ANDN U5368 ( .A(n5321), .B(n5322), .Z(n4951) );
  AND U5369 ( .A(n1870), .B(n1741), .Z(n3342) );
  IV U5370 ( .A(n1968), .Z(n1870) );
  XNOR U5371 ( .A(n5146), .B(n5147), .Z(n5152) );
  NAND U5372 ( .A(n2163), .B(n1557), .Z(n5147) );
  XNOR U5373 ( .A(n5145), .B(n5327), .Z(n5146) );
  ANDN U5374 ( .A(n1564), .B(n2165), .Z(n5327) );
  XNOR U5375 ( .A(n5331), .B(n5324), .Z(n5154) );
  XNOR U5376 ( .A(n5323), .B(n5332), .Z(n5324) );
  ANDN U5377 ( .A(n1748), .B(n1968), .Z(n5332) );
  ANDN U5378 ( .A(n5333), .B(n5334), .Z(n5321) );
  AND U5379 ( .A(n1966), .B(n1741), .Z(n5325) );
  IV U5380 ( .A(n2064), .Z(n1966) );
  XNOR U5381 ( .A(n5329), .B(n5330), .Z(n5172) );
  NAND U5382 ( .A(n2269), .B(n1557), .Z(n5330) );
  XNOR U5383 ( .A(n5328), .B(n5339), .Z(n5329) );
  ANDN U5384 ( .A(n1564), .B(n2271), .Z(n5339) );
  XNOR U5385 ( .A(n5343), .B(n5336), .Z(n5174) );
  XNOR U5386 ( .A(n5335), .B(n5344), .Z(n5336) );
  ANDN U5387 ( .A(n1748), .B(n2064), .Z(n5344) );
  XNOR U5388 ( .A(n5333), .B(A[14]), .Z(n5334) );
  ANDN U5389 ( .A(n5345), .B(n5346), .Z(n5333) );
  AND U5390 ( .A(n2062), .B(n1741), .Z(n5337) );
  IV U5391 ( .A(n2165), .Z(n2062) );
  XNOR U5392 ( .A(n5341), .B(n5342), .Z(n5192) );
  NAND U5393 ( .A(n2376), .B(n1557), .Z(n5342) );
  XNOR U5394 ( .A(n5340), .B(n5351), .Z(n5341) );
  ANDN U5395 ( .A(n1564), .B(n2378), .Z(n5351) );
  XNOR U5396 ( .A(n5355), .B(n5348), .Z(n5194) );
  XNOR U5397 ( .A(n5347), .B(n5356), .Z(n5348) );
  ANDN U5398 ( .A(n1748), .B(n2165), .Z(n5356) );
  ANDN U5399 ( .A(n5357), .B(n5358), .Z(n5345) );
  AND U5400 ( .A(n2163), .B(n1741), .Z(n5349) );
  IV U5401 ( .A(n2271), .Z(n2163) );
  XNOR U5402 ( .A(n5353), .B(n5354), .Z(n5212) );
  NAND U5403 ( .A(n2484), .B(n1557), .Z(n5354) );
  XNOR U5404 ( .A(n5352), .B(n5363), .Z(n5353) );
  ANDN U5405 ( .A(n1564), .B(n2486), .Z(n5363) );
  XNOR U5406 ( .A(n5367), .B(n5360), .Z(n5214) );
  XNOR U5407 ( .A(n5359), .B(n5368), .Z(n5360) );
  ANDN U5408 ( .A(n1748), .B(n2271), .Z(n5368) );
  XNOR U5409 ( .A(n5357), .B(A[12]), .Z(n5358) );
  ANDN U5410 ( .A(n5369), .B(n5370), .Z(n5357) );
  AND U5411 ( .A(n2269), .B(n1741), .Z(n5361) );
  IV U5412 ( .A(n2378), .Z(n2269) );
  XNOR U5413 ( .A(n5365), .B(n5366), .Z(n5232) );
  NAND U5414 ( .A(n2603), .B(n1557), .Z(n5366) );
  XNOR U5415 ( .A(n5364), .B(n5375), .Z(n5365) );
  ANDN U5416 ( .A(n1564), .B(n2605), .Z(n5375) );
  XOR U5417 ( .A(n5376), .B(n5377), .Z(n5364) );
  AND U5418 ( .A(n5378), .B(n5379), .Z(n5377) );
  XOR U5419 ( .A(n5380), .B(n5376), .Z(n5379) );
  XNOR U5420 ( .A(n5381), .B(n5372), .Z(n5234) );
  XNOR U5421 ( .A(n5371), .B(n5382), .Z(n5372) );
  ANDN U5422 ( .A(n1748), .B(n2378), .Z(n5382) );
  ANDN U5423 ( .A(n5383), .B(n5384), .Z(n5369) );
  AND U5424 ( .A(n2376), .B(n1741), .Z(n5373) );
  IV U5425 ( .A(n2486), .Z(n2376) );
  XNOR U5426 ( .A(n5378), .B(n5380), .Z(n5254) );
  NAND U5427 ( .A(n2723), .B(n1557), .Z(n5380) );
  XNOR U5428 ( .A(n5376), .B(n5389), .Z(n5378) );
  ANDN U5429 ( .A(n1564), .B(n2725), .Z(n5389) );
  XOR U5430 ( .A(n5390), .B(n5391), .Z(n5376) );
  AND U5431 ( .A(n5392), .B(n5393), .Z(n5391) );
  XOR U5432 ( .A(n5394), .B(n5390), .Z(n5393) );
  XNOR U5433 ( .A(n5395), .B(n5386), .Z(n5256) );
  XNOR U5434 ( .A(n5385), .B(n5396), .Z(n5386) );
  ANDN U5435 ( .A(n1748), .B(n2486), .Z(n5396) );
  XNOR U5436 ( .A(n5383), .B(A[10]), .Z(n5384) );
  ANDN U5437 ( .A(n5397), .B(n5398), .Z(n5383) );
  XOR U5438 ( .A(n5399), .B(n5400), .Z(n5385) );
  AND U5439 ( .A(n5401), .B(n5402), .Z(n5400) );
  XNOR U5440 ( .A(n5403), .B(n5399), .Z(n5402) );
  XOR U5441 ( .A(n5404), .B(n5387), .Z(n5395) );
  AND U5442 ( .A(n2484), .B(n1741), .Z(n5387) );
  IV U5443 ( .A(n2605), .Z(n2484) );
  IV U5444 ( .A(n5388), .Z(n5404) );
  XNOR U5445 ( .A(n5392), .B(n5394), .Z(n5278) );
  NAND U5446 ( .A(n2845), .B(n1557), .Z(n5394) );
  XNOR U5447 ( .A(n5390), .B(n5406), .Z(n5392) );
  ANDN U5448 ( .A(n1564), .B(n2847), .Z(n5406) );
  XNOR U5449 ( .A(n5410), .B(n5401), .Z(n5280) );
  XNOR U5450 ( .A(n5399), .B(n5411), .Z(n5401) );
  ANDN U5451 ( .A(n1748), .B(n2605), .Z(n5411) );
  ANDN U5452 ( .A(n5412), .B(n5413), .Z(n5397) );
  XOR U5453 ( .A(n5414), .B(n5415), .Z(n5399) );
  AND U5454 ( .A(n5416), .B(n5417), .Z(n5415) );
  XNOR U5455 ( .A(n5418), .B(n5414), .Z(n5417) );
  AND U5456 ( .A(n2603), .B(n1741), .Z(n5403) );
  IV U5457 ( .A(n2725), .Z(n2603) );
  XNOR U5458 ( .A(n5408), .B(n5409), .Z(n5296) );
  NAND U5459 ( .A(n2970), .B(n1557), .Z(n5409) );
  XNOR U5460 ( .A(n5407), .B(n5420), .Z(n5408) );
  ANDN U5461 ( .A(n1564), .B(n2972), .Z(n5420) );
  XNOR U5462 ( .A(n5424), .B(n5416), .Z(n5297) );
  XNOR U5463 ( .A(n5414), .B(n5425), .Z(n5416) );
  ANDN U5464 ( .A(n1748), .B(n2725), .Z(n5425) );
  AND U5465 ( .A(n2723), .B(n1741), .Z(n5418) );
  XNOR U5466 ( .A(n5429), .B(n5430), .Z(n5419) );
  AND U5467 ( .A(n5431), .B(n5432), .Z(n5430) );
  XNOR U5468 ( .A(n5427), .B(n5433), .Z(n5432) );
  XNOR U5469 ( .A(n5428), .B(n5429), .Z(n5433) );
  AND U5470 ( .A(n2845), .B(n1741), .Z(n5428) );
  XOR U5471 ( .A(n5426), .B(n5434), .Z(n5427) );
  ANDN U5472 ( .A(n1748), .B(n2847), .Z(n5434) );
  XNOR U5473 ( .A(n5422), .B(n5438), .Z(n5431) );
  XNOR U5474 ( .A(n5423), .B(n5429), .Z(n5438) );
  AND U5475 ( .A(n3102), .B(n1557), .Z(n5423) );
  XOR U5476 ( .A(n5421), .B(n5439), .Z(n5422) );
  ANDN U5477 ( .A(n1564), .B(n3104), .Z(n5439) );
  XOR U5478 ( .A(n5443), .B(n5444), .Z(n5429) );
  AND U5479 ( .A(n5445), .B(n5446), .Z(n5444) );
  XNOR U5480 ( .A(n5436), .B(n5447), .Z(n5446) );
  XNOR U5481 ( .A(n5437), .B(n5443), .Z(n5447) );
  AND U5482 ( .A(n2970), .B(n1741), .Z(n5437) );
  XOR U5483 ( .A(n5435), .B(n5448), .Z(n5436) );
  ANDN U5484 ( .A(n1748), .B(n2972), .Z(n5448) );
  XNOR U5485 ( .A(n5441), .B(n5452), .Z(n5445) );
  XNOR U5486 ( .A(n5442), .B(n5443), .Z(n5452) );
  AND U5487 ( .A(n3234), .B(n1557), .Z(n5442) );
  XOR U5488 ( .A(n5440), .B(n5453), .Z(n5441) );
  ANDN U5489 ( .A(n1564), .B(n3236), .Z(n5453) );
  XOR U5490 ( .A(n5454), .B(n5455), .Z(n5440) );
  ANDN U5491 ( .A(n5456), .B(n5457), .Z(n5455) );
  XNOR U5492 ( .A(n5458), .B(n5454), .Z(n5456) );
  XOR U5493 ( .A(n5459), .B(n5460), .Z(n5443) );
  AND U5494 ( .A(n5461), .B(n5462), .Z(n5460) );
  XNOR U5495 ( .A(n5450), .B(n5463), .Z(n5462) );
  XNOR U5496 ( .A(n5451), .B(n5459), .Z(n5463) );
  AND U5497 ( .A(n3102), .B(n1741), .Z(n5451) );
  XOR U5498 ( .A(n5449), .B(n5464), .Z(n5450) );
  ANDN U5499 ( .A(n1748), .B(n3104), .Z(n5464) );
  XNOR U5500 ( .A(n5457), .B(n5468), .Z(n5461) );
  XNOR U5501 ( .A(n5458), .B(n5459), .Z(n5468) );
  AND U5502 ( .A(n3370), .B(n1557), .Z(n5458) );
  XOR U5503 ( .A(n5454), .B(n5469), .Z(n5457) );
  ANDN U5504 ( .A(n1564), .B(n3372), .Z(n5469) );
  XNOR U5505 ( .A(n5474), .B(n5466), .Z(n5318) );
  XNOR U5506 ( .A(n5465), .B(n5475), .Z(n5466) );
  ANDN U5507 ( .A(n1748), .B(n3236), .Z(n5475) );
  XNOR U5508 ( .A(n5478), .B(n5476), .Z(n5477) );
  ANDN U5509 ( .A(n1748), .B(n3372), .Z(n5478) );
  XNOR U5510 ( .A(n5473), .B(n5467), .Z(n5474) );
  AND U5511 ( .A(n3234), .B(n1741), .Z(n5467) );
  XNOR U5512 ( .A(n5471), .B(n5472), .Z(n5317) );
  NAND U5513 ( .A(n4158), .B(n1557), .Z(n5472) );
  XNOR U5514 ( .A(n5470), .B(n5482), .Z(n5471) );
  ANDN U5515 ( .A(n1564), .B(n4160), .Z(n5482) );
  NAND U5516 ( .A(A[0]), .B(n5483), .Z(n5470) );
  NANDN U5517 ( .B(n1557), .A(n5484), .Z(n5483) );
  NANDN U5518 ( .B(n4163), .A(n1564), .Z(n5484) );
  IV U5519 ( .A(n1483), .Z(n1557) );
  XNOR U5520 ( .A(n5480), .B(n5481), .Z(n5473) );
  NAND U5521 ( .A(n4158), .B(n1741), .Z(n5481) );
  XNOR U5522 ( .A(n5479), .B(n5487), .Z(n5480) );
  ANDN U5523 ( .A(n1748), .B(n4160), .Z(n5487) );
  NAND U5524 ( .A(A[0]), .B(n5488), .Z(n5479) );
  NANDN U5525 ( .B(n1741), .A(n5489), .Z(n5488) );
  NANDN U5526 ( .B(n4163), .A(n1748), .Z(n5489) );
  IV U5527 ( .A(n1648), .Z(n1741) );
  XNOR U5528 ( .A(n3353), .B(n3352), .Z(n3329) );
  XOR U5529 ( .A(n5492), .B(n3361), .Z(n3352) );
  XNOR U5530 ( .A(n3349), .B(n3350), .Z(n3361) );
  NANDN U5531 ( .B(n1001), .A(n2970), .Z(n3350) );
  XNOR U5532 ( .A(n3348), .B(n5493), .Z(n3349) );
  ANDN U5533 ( .A(n1042), .B(n2972), .Z(n5493) );
  XOR U5534 ( .A(n3360), .B(n3351), .Z(n5492) );
  XOR U5535 ( .A(n5497), .B(n5498), .Z(n3351) );
  XOR U5536 ( .A(n5499), .B(n3357), .Z(n3360) );
  XNOR U5537 ( .A(n3356), .B(n5500), .Z(n3357) );
  ANDN U5538 ( .A(n1149), .B(n2725), .Z(n5500) );
  XNOR U5539 ( .A(n5412), .B(A[8]), .Z(n5413) );
  ANDN U5540 ( .A(n5501), .B(n5502), .Z(n5412) );
  AND U5541 ( .A(n2723), .B(n1095), .Z(n3358) );
  IV U5542 ( .A(n2847), .Z(n2723) );
  XNOR U5543 ( .A(n5506), .B(n5507), .Z(n3359) );
  AND U5544 ( .A(n5508), .B(n5509), .Z(n5507) );
  XNOR U5545 ( .A(n5504), .B(n5510), .Z(n5509) );
  XNOR U5546 ( .A(n5505), .B(n5506), .Z(n5510) );
  AND U5547 ( .A(n2845), .B(n1095), .Z(n5505) );
  IV U5548 ( .A(n2972), .Z(n2845) );
  XOR U5549 ( .A(n5503), .B(n5511), .Z(n5504) );
  ANDN U5550 ( .A(n1149), .B(n2847), .Z(n5511) );
  ANDN U5551 ( .A(n5512), .B(n5513), .Z(n5501) );
  XNOR U5552 ( .A(n5495), .B(n5517), .Z(n5508) );
  XNOR U5553 ( .A(n5496), .B(n5506), .Z(n5517) );
  ANDN U5554 ( .A(n3102), .B(n1001), .Z(n5496) );
  XOR U5555 ( .A(n5494), .B(n5518), .Z(n5495) );
  ANDN U5556 ( .A(n1042), .B(n3104), .Z(n5518) );
  XOR U5557 ( .A(n5522), .B(n5523), .Z(n5506) );
  AND U5558 ( .A(n5524), .B(n5525), .Z(n5523) );
  XNOR U5559 ( .A(n5515), .B(n5526), .Z(n5525) );
  XNOR U5560 ( .A(n5516), .B(n5522), .Z(n5526) );
  AND U5561 ( .A(n2970), .B(n1095), .Z(n5516) );
  IV U5562 ( .A(n3104), .Z(n2970) );
  XOR U5563 ( .A(n5514), .B(n5527), .Z(n5515) );
  ANDN U5564 ( .A(n1149), .B(n2972), .Z(n5527) );
  XNOR U5565 ( .A(n5512), .B(A[6]), .Z(n5513) );
  ANDN U5566 ( .A(n5528), .B(n5529), .Z(n5512) );
  XNOR U5567 ( .A(n5520), .B(n5533), .Z(n5524) );
  XNOR U5568 ( .A(n5521), .B(n5522), .Z(n5533) );
  ANDN U5569 ( .A(n3234), .B(n1001), .Z(n5521) );
  XOR U5570 ( .A(n5519), .B(n5534), .Z(n5520) );
  ANDN U5571 ( .A(n1042), .B(n3236), .Z(n5534) );
  XOR U5572 ( .A(n5535), .B(n5536), .Z(n5519) );
  ANDN U5573 ( .A(n5537), .B(n5538), .Z(n5536) );
  XNOR U5574 ( .A(n5539), .B(n5535), .Z(n5537) );
  XOR U5575 ( .A(n5540), .B(n5541), .Z(n5522) );
  AND U5576 ( .A(n5542), .B(n5543), .Z(n5541) );
  XNOR U5577 ( .A(n5531), .B(n5544), .Z(n5543) );
  XNOR U5578 ( .A(n5532), .B(n5540), .Z(n5544) );
  AND U5579 ( .A(n3102), .B(n1095), .Z(n5532) );
  XOR U5580 ( .A(n5530), .B(n5545), .Z(n5531) );
  ANDN U5581 ( .A(n1149), .B(n3104), .Z(n5545) );
  ANDN U5582 ( .A(n5546), .B(n5547), .Z(n5528) );
  XNOR U5583 ( .A(n5538), .B(n5551), .Z(n5542) );
  XNOR U5584 ( .A(n5539), .B(n5540), .Z(n5551) );
  ANDN U5585 ( .A(n3370), .B(n1001), .Z(n5539) );
  XOR U5586 ( .A(n5535), .B(n5552), .Z(n5538) );
  ANDN U5587 ( .A(n1042), .B(n3372), .Z(n5552) );
  XNOR U5588 ( .A(n5557), .B(n5549), .Z(n5498) );
  XNOR U5589 ( .A(n5548), .B(n5558), .Z(n5549) );
  ANDN U5590 ( .A(n1149), .B(n3236), .Z(n5558) );
  XNOR U5591 ( .A(n5561), .B(n5559), .Z(n5560) );
  ANDN U5592 ( .A(n1149), .B(n3372), .Z(n5561) );
  XNOR U5593 ( .A(n5556), .B(n5550), .Z(n5557) );
  AND U5594 ( .A(n3234), .B(n1095), .Z(n5550) );
  XNOR U5595 ( .A(n5554), .B(n5555), .Z(n5497) );
  NANDN U5596 ( .B(n1001), .A(n4158), .Z(n5555) );
  XNOR U5597 ( .A(n5553), .B(n5566), .Z(n5554) );
  ANDN U5598 ( .A(n1042), .B(n4160), .Z(n5566) );
  NAND U5599 ( .A(A[0]), .B(n5567), .Z(n5553) );
  NAND U5600 ( .A(n5568), .B(n1001), .Z(n5567) );
  NANDN U5601 ( .B(n4163), .A(n1042), .Z(n5568) );
  XNOR U5602 ( .A(n5564), .B(n5565), .Z(n5556) );
  NAND U5603 ( .A(n4158), .B(n1095), .Z(n5565) );
  XNOR U5604 ( .A(n5563), .B(n5571), .Z(n5564) );
  ANDN U5605 ( .A(n1149), .B(n4160), .Z(n5571) );
  NAND U5606 ( .A(A[0]), .B(n5572), .Z(n5563) );
  NANDN U5607 ( .B(n1095), .A(n5573), .Z(n5572) );
  NANDN U5608 ( .B(n4163), .A(n1149), .Z(n5573) );
  IV U5609 ( .A(n5562), .Z(n1095) );
  XOR U5610 ( .A(n3369), .B(n3368), .Z(n3353) );
  XOR U5611 ( .A(n5576), .B(n3365), .Z(n3368) );
  XNOR U5612 ( .A(n3364), .B(n5577), .Z(n3365) );
  ANDN U5613 ( .A(n974), .B(n3236), .Z(n5577) );
  IV U5614 ( .A(n3102), .Z(n3236) );
  XNOR U5615 ( .A(n5546), .B(A[4]), .Z(n5547) );
  ANDN U5616 ( .A(n5578), .B(n5579), .Z(n5546) );
  XNOR U5617 ( .A(n5582), .B(n5580), .Z(n5581) );
  ANDN U5618 ( .A(n974), .B(n3372), .Z(n5582) );
  IV U5619 ( .A(n3234), .Z(n3372) );
  IV U5620 ( .A(n4160), .Z(n3370) );
  XNOR U5621 ( .A(n3367), .B(n3366), .Z(n5576) );
  AND U5622 ( .A(n3234), .B(n933), .Z(n3366) );
  ANDN U5623 ( .A(n5587), .B(n5588), .Z(n5578) );
  XNOR U5624 ( .A(n5585), .B(n5586), .Z(n3367) );
  NAND U5625 ( .A(n4158), .B(n933), .Z(n5586) );
  XNOR U5626 ( .A(n5584), .B(n5589), .Z(n5585) );
  ANDN U5627 ( .A(n974), .B(n4160), .Z(n5589) );
  NAND U5628 ( .A(A[0]), .B(n5590), .Z(n5584) );
  NANDN U5629 ( .B(n933), .A(n5591), .Z(n5590) );
  NANDN U5630 ( .B(n4163), .A(n974), .Z(n5591) );
  IV U5631 ( .A(n5583), .Z(n933) );
  XOR U5632 ( .A(n3376), .B(n3375), .Z(n3369) );
  NAND U5633 ( .A(n4158), .B(n877), .Z(n3375) );
  IV U5634 ( .A(n4163), .Z(n4158) );
  XOR U5635 ( .A(n3374), .B(n5594), .Z(n3376) );
  ANDN U5636 ( .A(n908), .B(n4160), .Z(n5594) );
  XNOR U5637 ( .A(n5587), .B(A[2]), .Z(n5588) );
  NOR U5638 ( .A(A[0]), .B(n5595), .Z(n5587) );
  NANDN U5639 ( .B(n877), .A(n5597), .Z(n5596) );
  NANDN U5640 ( .B(n4163), .A(n908), .Z(n5597) );
  XOR U5641 ( .A(A[0]), .B(A[1]), .Z(n5595) );
  AND U5642 ( .A(n5599), .B(n5598), .Z(n877) );
  ANDN U5643 ( .A(X[31]), .B(n5600), .Z(n5599) );
  NANDN U5644 ( .B(n5601), .A(n5593), .Z(n5600) );
  XNOR U5645 ( .A(n5601), .B(X[29]), .Z(n5593) );
  NAND U5646 ( .A(n5592), .B(n5602), .Z(n5601) );
  XOR U5647 ( .A(n5602), .B(X[28]), .Z(n5592) );
  ANDN U5648 ( .A(n5569), .B(n5603), .Z(n5602) );
  XNOR U5649 ( .A(n5603), .B(X[27]), .Z(n5569) );
  NAND U5650 ( .A(n5570), .B(n5604), .Z(n5603) );
  XOR U5651 ( .A(n5604), .B(X[26]), .Z(n5570) );
  ANDN U5652 ( .A(n5575), .B(n5605), .Z(n5604) );
  XNOR U5653 ( .A(n5605), .B(X[25]), .Z(n5575) );
  NAND U5654 ( .A(n5574), .B(n5606), .Z(n5605) );
  XOR U5655 ( .A(n5606), .B(X[24]), .Z(n5574) );
  ANDN U5656 ( .A(n5315), .B(n5607), .Z(n5606) );
  XNOR U5657 ( .A(n5607), .B(X[23]), .Z(n5315) );
  NAND U5658 ( .A(n5316), .B(n5608), .Z(n5607) );
  XOR U5659 ( .A(n5608), .B(X[22]), .Z(n5316) );
  ANDN U5660 ( .A(n5311), .B(n5609), .Z(n5608) );
  XNOR U5661 ( .A(n5609), .B(X[21]), .Z(n5311) );
  NAND U5662 ( .A(n5310), .B(n5610), .Z(n5609) );
  XOR U5663 ( .A(n5610), .B(X[20]), .Z(n5310) );
  ANDN U5664 ( .A(n5486), .B(n5611), .Z(n5610) );
  XNOR U5665 ( .A(n5611), .B(X[19]), .Z(n5486) );
  NAND U5666 ( .A(n5485), .B(n5612), .Z(n5611) );
  XOR U5667 ( .A(n5612), .B(X[18]), .Z(n5485) );
  ANDN U5668 ( .A(n5491), .B(n5613), .Z(n5612) );
  XNOR U5669 ( .A(n5613), .B(X[17]), .Z(n5491) );
  NAND U5670 ( .A(n5490), .B(n5614), .Z(n5613) );
  XOR U5671 ( .A(n5614), .B(X[16]), .Z(n5490) );
  ANDN U5672 ( .A(n4188), .B(n5615), .Z(n5614) );
  XNOR U5673 ( .A(n5615), .B(X[15]), .Z(n4188) );
  NAND U5674 ( .A(n4187), .B(n5616), .Z(n5615) );
  XOR U5675 ( .A(n5616), .B(X[14]), .Z(n4187) );
  ANDN U5676 ( .A(n4183), .B(n5617), .Z(n5616) );
  XNOR U5677 ( .A(n5617), .B(X[13]), .Z(n4183) );
  NAND U5678 ( .A(n4182), .B(n5618), .Z(n5617) );
  XOR U5679 ( .A(n5618), .B(X[12]), .Z(n4182) );
  ANDN U5680 ( .A(n4165), .B(n5619), .Z(n5618) );
  XNOR U5681 ( .A(n5619), .B(X[11]), .Z(n4165) );
  NAND U5682 ( .A(n4164), .B(n5620), .Z(n5619) );
  XOR U5683 ( .A(n5620), .B(X[10]), .Z(n4164) );
  ANDN U5684 ( .A(n4170), .B(n5621), .Z(n5620) );
  XNOR U5685 ( .A(n5621), .B(X[9]), .Z(n4170) );
  NAND U5686 ( .A(n4169), .B(n5622), .Z(n5621) );
  XOR U5687 ( .A(n5622), .B(X[8]), .Z(n4169) );
  ANDN U5688 ( .A(n4694), .B(n5623), .Z(n5622) );
  XNOR U5689 ( .A(n5623), .B(X[7]), .Z(n4694) );
  NAND U5690 ( .A(n4693), .B(n5624), .Z(n5623) );
  XOR U5691 ( .A(n5624), .B(X[6]), .Z(n4693) );
  ANDN U5692 ( .A(n4689), .B(n5625), .Z(n5624) );
  XNOR U5693 ( .A(n5625), .B(X[5]), .Z(n4689) );
  NAND U5694 ( .A(n4688), .B(n5626), .Z(n5625) );
  XOR U5695 ( .A(n5626), .B(X[4]), .Z(n4688) );
  ANDN U5696 ( .A(n5123), .B(n5627), .Z(n5626) );
  XNOR U5697 ( .A(n5627), .B(X[3]), .Z(n5123) );
  NAND U5698 ( .A(n5122), .B(n5628), .Z(n5627) );
  XOR U5699 ( .A(n5628), .B(X[2]), .Z(n5122) );
  NOR U5700 ( .A(n5127), .B(X[0]), .Z(n5628) );
  XOR U5701 ( .A(X[0]), .B(X[1]), .Z(n5127) );
endmodule

