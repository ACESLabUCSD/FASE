
module MxM_TG_W16_N100 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MxM/n229 , \_MxM/n228 , \_MxM/n227 , \_MxM/n226 , \_MxM/n225 ,
         \_MxM/n224 , \_MxM/n223 , \_MxM/n222 , \_MxM/n221 , \_MxM/n220 ,
         \_MxM/n219 , \_MxM/n218 , \_MxM/n217 , \_MxM/n216 , \_MxM/n215 ,
         \_MxM/n214 , \_MxM/n213 , \_MxM/n212 , \_MxM/n211 , \_MxM/n210 ,
         \_MxM/n209 , \_MxM/n208 , \_MxM/n207 , \_MxM/n206 , \_MxM/n205 ,
         \_MxM/n204 , \_MxM/n203 , \_MxM/n202 , \_MxM/n201 , \_MxM/n200 ,
         \_MxM/n199 , \_MxM/n198 , \_MxM/n197 , \_MxM/n196 , \_MxM/n195 ,
         \_MxM/n194 , \_MxM/n193 , \_MxM/n192 , \_MxM/n191 , \_MxM/N12 ,
         \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/n[0] ,
         \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] ,
         \_MxM/n[6] , \_MxM/Y0[0] , \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] ,
         \_MxM/Y0[4] , \_MxM/Y0[5] , \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/Y0[8] ,
         \_MxM/Y0[9] , \_MxM/Y0[10] , \_MxM/Y0[11] , \_MxM/Y0[12] ,
         \_MxM/Y0[13] , \_MxM/Y0[14] , \_MxM/Y0[15] , \_MxM/add_39/carry[6] ,
         \_MxM/add_39/carry[5] , \_MxM/add_39/carry[4] ,
         \_MxM/add_39/carry[3] , \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n191 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n192 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n193 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n194 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n195 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n196 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n197 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n198 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n199 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n200 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n201 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n202 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n203 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n204 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n205 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n206 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/n207 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/n208 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/n209 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/n210 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/n211 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/n212 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/n213 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/n214 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n215 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n216 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n217 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n218 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n219 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n220 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n221 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n222 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n223 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n224 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n225 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n226 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n227 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n228 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n229 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  MUX U1 ( .IN0(n1), .IN1(n1314), .SEL(n1315), .F(n1298) );
  IV U2 ( .A(n1316), .Z(n1) );
  MUX U3 ( .IN0(n2), .IN1(n981), .SEL(n982), .F(n958) );
  IV U4 ( .A(n983), .Z(n2) );
  MUX U5 ( .IN0(n1389), .IN1(n1407), .SEL(n1391), .F(n1370) );
  XOR U6 ( .A(n1172), .B(n1162), .Z(n978) );
  XOR U7 ( .A(n984), .B(n966), .Z(n970) );
  MUX U8 ( .IN0(n3), .IN1(n731), .SEL(n732), .F(n661) );
  IV U9 ( .A(n733), .Z(n3) );
  MUX U10 ( .IN0(n4), .IN1(n892), .SEL(n893), .F(n817) );
  IV U11 ( .A(n894), .Z(n4) );
  MUX U12 ( .IN0(n5), .IN1(n958), .SEL(n959), .F(n935) );
  IV U13 ( .A(n960), .Z(n5) );
  MUX U14 ( .IN0(n6), .IN1(n1154), .SEL(n1155), .F(n1144) );
  IV U15 ( .A(n1156), .Z(n6) );
  XOR U16 ( .A(n1157), .B(n1149), .Z(n955) );
  MUX U17 ( .IN0(n1109), .IN1(n1112), .SEL(n1110), .F(n1094) );
  MUX U18 ( .IN0(n7), .IN1(n456), .SEL(n457), .F(n405) );
  IV U19 ( .A(n458), .Z(n7) );
  MUX U20 ( .IN0(n8), .IN1(n808), .SEL(n809), .F(n731) );
  IV U21 ( .A(n810), .Z(n8) );
  XNOR U22 ( .A(n1452), .B(n1453), .Z(n896) );
  XOR U23 ( .A(n959), .B(n960), .Z(n971) );
  MUX U24 ( .IN0(n9), .IN1(n908), .SEL(n909), .F(n846) );
  IV U25 ( .A(n910), .Z(n9) );
  XOR U26 ( .A(n1145), .B(n1146), .Z(n953) );
  MUX U27 ( .IN0(n10), .IN1(n585), .SEL(n586), .F(n520) );
  IV U28 ( .A(n587), .Z(n10) );
  MUX U29 ( .IN0(e_input[8]), .IN1(n1437), .SEL(e_input[15]), .F(n468) );
  MUX U30 ( .IN0(n1150), .IN1(n11), .SEL(n1149), .F(n1141) );
  IV U31 ( .A(n1148), .Z(n11) );
  MUX U32 ( .IN0(e_input[13]), .IN1(n1463), .SEL(e_input[15]), .F(n250) );
  MUX U33 ( .IN0(n1325), .IN1(n1328), .SEL(n1326), .F(n1309) );
  MUX U34 ( .IN0(n12), .IN1(n935), .SEL(n936), .F(n916) );
  IV U35 ( .A(n937), .Z(n12) );
  MUX U36 ( .IN0(n13), .IN1(n1144), .SEL(n1145), .F(n923) );
  IV U37 ( .A(n1146), .Z(n13) );
  XOR U38 ( .A(n961), .B(n943), .Z(n947) );
  MUX U39 ( .IN0(e_input[9]), .IN1(n1438), .SEL(e_input[15]), .F(n414) );
  MUX U40 ( .IN0(n291), .IN1(n14), .SEL(n290), .F(n252) );
  IV U41 ( .A(n289), .Z(n14) );
  MUX U42 ( .IN0(e_input[11]), .IN1(n1418), .SEL(e_input[15]), .F(n320) );
  MUX U43 ( .IN0(n381), .IN1(n379), .SEL(n380), .F(n334) );
  MUX U44 ( .IN0(n15), .IN1(n174), .SEL(n173), .F(n182) );
  IV U45 ( .A(n185), .Z(n15) );
  MUX U46 ( .IN0(n16), .IN1(n1329), .SEL(n1330), .F(n1325) );
  IV U47 ( .A(n1331), .Z(n16) );
  XOR U48 ( .A(n1155), .B(n1156), .Z(n976) );
  MUX U49 ( .IN0(n17), .IN1(n712), .SEL(n713), .F(n643) );
  IV U50 ( .A(n714), .Z(n17) );
  MUX U51 ( .IN0(n18), .IN1(n771), .SEL(n772), .F(n708) );
  IV U52 ( .A(n773), .Z(n18) );
  MUX U53 ( .IN0(e_input[10]), .IN1(n1417), .SEL(e_input[15]), .F(n361) );
  MUX U54 ( .IN0(n471), .IN1(n19), .SEL(n470), .F(n416) );
  IV U55 ( .A(n469), .Z(n19) );
  MUX U56 ( .IN0(n547), .IN1(n545), .SEL(n546), .F(n480) );
  XNOR U57 ( .A(n1439), .B(n893), .Z(n897) );
  XOR U58 ( .A(n183), .B(n204), .Z(n202) );
  MUX U59 ( .IN0(n1370), .IN1(n1388), .SEL(n1372), .F(n1339) );
  MUX U60 ( .IN0(n1258), .IN1(n1280), .SEL(n1260), .F(n1240) );
  MUX U61 ( .IN0(n20), .IN1(n916), .SEL(n917), .F(n854) );
  IV U62 ( .A(n918), .Z(n20) );
  MUX U63 ( .IN0(n21), .IN1(n1161), .SEL(n1162), .F(n1148) );
  IV U64 ( .A(n1163), .Z(n21) );
  MUX U65 ( .IN0(n22), .IN1(n883), .SEL(n884), .F(n808) );
  IV U66 ( .A(n885), .Z(n22) );
  MUX U67 ( .IN0(g_input[11]), .IN1(n1192), .SEL(g_input[15]), .F(n337) );
  MUX U68 ( .IN0(n419), .IN1(n27), .SEL(n418), .F(n368) );
  MUX U69 ( .IN0(n680), .IN1(n678), .SEL(n679), .F(n610) );
  MUX U70 ( .IN0(n710), .IN1(n23), .SEL(n709), .F(n638) );
  IV U71 ( .A(n708), .Z(n23) );
  NAND U72 ( .A(n252), .B(n287), .Z(n286) );
  XOR U73 ( .A(n230), .B(n238), .Z(n236) );
  MUX U74 ( .IN0(n24), .IN1(n1176), .SEL(n1177), .F(n1161) );
  IV U75 ( .A(n1178), .Z(n24) );
  MUX U76 ( .IN0(n25), .IN1(n723), .SEL(n724), .F(n653) );
  IV U77 ( .A(n725), .Z(n25) );
  MUX U78 ( .IN0(n26), .IN1(n779), .SEL(n780), .F(n712) );
  IV U79 ( .A(n781), .Z(n26) );
  MUX U80 ( .IN0(e_input[4]), .IN1(n1123), .SEL(e_input[15]), .F(n707) );
  XOR U81 ( .A(n1419), .B(n1404), .Z(n1344) );
  MUX U82 ( .IN0(n463), .IN1(n465), .SEL(n464), .F(n27) );
  IV U83 ( .A(n27), .Z(n417) );
  MUX U84 ( .IN0(n641), .IN1(n28), .SEL(n640), .F(n568) );
  IV U85 ( .A(n639), .Z(n28) );
  MUX U86 ( .IN0(n748), .IN1(n746), .SEL(n747), .F(n678) );
  MUX U87 ( .IN0(n866), .IN1(n29), .SEL(n865), .F(n789) );
  IV U88 ( .A(n864), .Z(n29) );
  XNOR U89 ( .A(n371), .B(n331), .Z(n335) );
  XOR U90 ( .A(n261), .B(n269), .Z(n267) );
  XOR U91 ( .A(n936), .B(n937), .Z(n948) );
  MUX U92 ( .IN0(n1264), .IN1(n1274), .SEL(n1266), .F(n1250) );
  MUX U93 ( .IN0(n1339), .IN1(n1369), .SEL(n1341), .F(n875) );
  XNOR U94 ( .A(n1116), .B(n1117), .Z(n1100) );
  MUX U95 ( .IN0(g_input[9]), .IN1(n1230), .SEL(g_input[15]), .F(n431) );
  MUX U96 ( .IN0(g_input[12]), .IN1(n1174), .SEL(g_input[15]), .F(n292) );
  XOR U97 ( .A(n340), .B(n383), .Z(n341) );
  MUX U98 ( .IN0(n735), .IN1(n737), .SEL(n736), .F(n667) );
  MUX U99 ( .IN0(n777), .IN1(n775), .SEL(n776), .F(n702) );
  XOR U100 ( .A(n865), .B(n866), .Z(n872) );
  XNOR U101 ( .A(n368), .B(n411), .Z(n369) );
  XNOR U102 ( .A(n472), .B(n425), .Z(n429) );
  MUX U103 ( .IN0(n30), .IN1(n656), .SEL(n657), .F(n588) );
  IV U104 ( .A(n658), .Z(n30) );
  MUX U105 ( .IN0(n515), .IN1(n517), .SEL(n516), .F(n31) );
  IV U106 ( .A(n31), .Z(n451) );
  XOR U107 ( .A(n298), .B(n306), .Z(n304) );
  MUX U108 ( .IN0(n1256), .IN1(n32), .SEL(n1106), .F(n1237) );
  IV U109 ( .A(n1105), .Z(n32) );
  MUX U110 ( .IN0(n1102), .IN1(n1100), .SEL(n1101), .F(n1073) );
  XOR U111 ( .A(n1147), .B(n1141), .Z(n932) );
  MUX U112 ( .IN0(n33), .IN1(n875), .SEL(n876), .F(n800) );
  IV U113 ( .A(n877), .Z(n33) );
  MUX U114 ( .IN0(n34), .IN1(n923), .SEL(n924), .F(n864) );
  IV U115 ( .A(n925), .Z(n34) );
  XOR U116 ( .A(n938), .B(n909), .Z(n913) );
  MUX U117 ( .IN0(n599), .IN1(n601), .SEL(n600), .F(n534) );
  MUX U118 ( .IN0(n825), .IN1(n823), .SEL(n824), .F(n746) );
  XOR U119 ( .A(n1345), .B(n884), .Z(n888) );
  XNOR U120 ( .A(n420), .B(n376), .Z(n380) );
  MUX U121 ( .IN0(n35), .IN1(n459), .SEL(n460), .F(n408) );
  IV U122 ( .A(n461), .Z(n35) );
  MUX U123 ( .IN0(n36), .IN1(n574), .SEL(n575), .F(n514) );
  IV U124 ( .A(n576), .Z(n36) );
  NAND U125 ( .A(n638), .B(n706), .Z(n705) );
  MUX U126 ( .IN0(n580), .IN1(n582), .SEL(n581), .F(n515) );
  MUX U127 ( .IN0(n37), .IN1(n554), .SEL(n555), .F(n489) );
  IV U128 ( .A(\_MxM/Y0[5] ), .Z(n37) );
  XOR U129 ( .A(n343), .B(n351), .Z(n349) );
  MUX U130 ( .IN0(n38), .IN1(n1309), .SEL(n1310), .F(n1292) );
  IV U131 ( .A(n1311), .Z(n38) );
  MUX U132 ( .IN0(g_input[1]), .IN1(n1465), .SEL(g_input[15]), .F(n1119) );
  MUX U133 ( .IN0(n39), .IN1(n520), .SEL(n521), .F(n456) );
  IV U134 ( .A(n522), .Z(n39) );
  MUX U135 ( .IN0(g_input[6]), .IN1(n1361), .SEL(g_input[15]), .F(n613) );
  MUX U136 ( .IN0(g_input[7]), .IN1(n1348), .SEL(g_input[15]), .F(n548) );
  MUX U137 ( .IN0(g_input[5]), .IN1(n1381), .SEL(g_input[15]), .F(n681) );
  MUX U138 ( .IN0(n40), .IN1(n854), .SEL(n855), .F(n779) );
  IV U139 ( .A(n856), .Z(n40) );
  XOR U140 ( .A(n924), .B(n925), .Z(n930) );
  MUX U141 ( .IN0(n667), .IN1(n669), .SEL(n668), .F(n599) );
  XNOR U142 ( .A(n906), .B(n847), .Z(n851) );
  XOR U143 ( .A(n258), .B(n293), .Z(n259) );
  MUX U144 ( .IN0(n41), .IN1(n323), .SEL(n324), .F(n276) );
  IV U145 ( .A(n325), .Z(n41) );
  NAND U146 ( .A(n416), .B(n467), .Z(n466) );
  MUX U147 ( .IN0(n570), .IN1(n568), .SEL(n569), .F(n512) );
  XNOR U148 ( .A(n602), .B(n542), .Z(n546) );
  MUX U149 ( .IN0(n42), .IN1(n803), .SEL(n804), .F(n726) );
  IV U150 ( .A(n805), .Z(n42) );
  MUX U151 ( .IN0(n43), .IN1(n650), .SEL(n649), .F(n580) );
  IV U152 ( .A(n648), .Z(n43) );
  MUX U153 ( .IN0(n44), .IN1(n619), .SEL(n620), .F(n554) );
  IV U154 ( .A(\_MxM/Y0[4] ), .Z(n44) );
  XOR U155 ( .A(n388), .B(n396), .Z(n394) );
  MUX U156 ( .IN0(n1073), .IN1(n45), .SEL(n1074), .F(n1046) );
  IV U157 ( .A(n1075), .Z(n45) );
  MUX U158 ( .IN0(n1165), .IN1(n46), .SEL(n978), .F(n1152) );
  IV U159 ( .A(n976), .Z(n46) );
  XNOR U160 ( .A(n1330), .B(n1331), .Z(n1317) );
  MUX U161 ( .IN0(n47), .IN1(n653), .SEL(n654), .F(n585) );
  IV U162 ( .A(n655), .Z(n47) );
  MUX U163 ( .IN0(g_input[3]), .IN1(n1442), .SEL(g_input[15]), .F(n48) );
  IV U164 ( .A(n48), .Z(n826) );
  MUX U165 ( .IN0(g_input[4]), .IN1(n1399), .SEL(g_input[15]), .F(n49) );
  IV U166 ( .A(n49), .Z(n749) );
  MUX U167 ( .IN0(n912), .IN1(n50), .SEL(n913), .F(n850) );
  IV U168 ( .A(n914), .Z(n50) );
  XOR U169 ( .A(n1243), .B(n1244), .Z(n1105) );
  MUX U170 ( .IN0(n336), .IN1(n334), .SEL(n335), .F(n281) );
  MUX U171 ( .IN0(n51), .IN1(n643), .SEL(n644), .F(n574) );
  IV U172 ( .A(n645), .Z(n51) );
  XOR U173 ( .A(n551), .B(n614), .Z(n552) );
  MUX U174 ( .IN0(n812), .IN1(n814), .SEL(n813), .F(n735) );
  MUX U175 ( .IN0(n898), .IN1(n896), .SEL(n897), .F(n823) );
  MUX U176 ( .IN0(n52), .IN1(n365), .SEL(n366), .F(n323) );
  IV U177 ( .A(n367), .Z(n52) );
  XOR U178 ( .A(n526), .B(n470), .Z(n464) );
  XNOR U179 ( .A(n537), .B(n477), .Z(n481) );
  MUX U180 ( .IN0(n53), .IN1(n588), .SEL(n589), .F(n523) );
  IV U181 ( .A(n590), .Z(n53) );
  XOR U182 ( .A(n701), .B(n639), .Z(n640) );
  MUX U183 ( .IN0(n797), .IN1(n54), .SEL(n796), .F(n718) );
  IV U184 ( .A(n795), .Z(n54) );
  MUX U185 ( .IN0(n715), .IN1(n55), .SEL(n716), .F(n648) );
  IV U186 ( .A(n717), .Z(n55) );
  MUX U187 ( .IN0(n56), .IN1(n687), .SEL(n688), .F(n619) );
  IV U188 ( .A(\_MxM/Y0[3] ), .Z(n56) );
  XOR U189 ( .A(n443), .B(n449), .Z(n438) );
  MUX U190 ( .IN0(n57), .IN1(n1103), .SEL(n920), .F(n1076) );
  IV U191 ( .A(n919), .Z(n57) );
  MUX U192 ( .IN0(n1019), .IN1(n58), .SEL(n1020), .F(n992) );
  IV U193 ( .A(n1021), .Z(n58) );
  MUX U194 ( .IN0(e_input[1]), .IN1(n59), .SEL(e_input[15]), .F(n1136) );
  IV U195 ( .A(n1336), .Z(n59) );
  MUX U196 ( .IN0(e_input[6]), .IN1(n1128), .SEL(e_input[15]), .F(n573) );
  MUX U197 ( .IN0(e_input[3]), .IN1(n1322), .SEL(e_input[15]), .F(n792) );
  MUX U198 ( .IN0(n887), .IN1(n889), .SEL(n888), .F(n812) );
  MUX U199 ( .IN0(e_input[14]), .IN1(n1468), .SEL(e_input[15]), .F(n219) );
  NAND U200 ( .A(n317), .B(n360), .Z(n359) );
  XOR U201 ( .A(n591), .B(n531), .Z(n535) );
  XNOR U202 ( .A(n670), .B(n607), .Z(n611) );
  MUX U203 ( .IN0(n60), .IN1(n726), .SEL(n727), .F(n656) );
  IV U204 ( .A(n728), .Z(n60) );
  XNOR U205 ( .A(n769), .B(n709), .Z(n703) );
  MUX U206 ( .IN0(n782), .IN1(n61), .SEL(n783), .F(n715) );
  IV U207 ( .A(n784), .Z(n61) );
  MUX U208 ( .IN0(n62), .IN1(n261), .SEL(n262), .F(n230) );
  IV U209 ( .A(\_MxM/Y0[11] ), .Z(n62) );
  XOR U210 ( .A(n489), .B(n497), .Z(n495) );
  MUX U211 ( .IN0(n1237), .IN1(n63), .SEL(n1082), .F(n1218) );
  IV U212 ( .A(n1080), .Z(n63) );
  MUX U213 ( .IN0(n1292), .IN1(n1308), .SEL(n1294), .F(n1275) );
  MUX U214 ( .IN0(n969), .IN1(n64), .SEL(n970), .F(n946) );
  IV U215 ( .A(n971), .Z(n64) );
  XOR U216 ( .A(n917), .B(n918), .Z(n914) );
  XOR U217 ( .A(n1315), .B(n1316), .Z(n1130) );
  MUX U218 ( .IN0(n65), .IN1(n800), .SEL(n801), .F(n723) );
  IV U219 ( .A(n802), .Z(n65) );
  MUX U220 ( .IN0(g_input[10]), .IN1(n1210), .SEL(g_input[15]), .F(n382) );
  XNOR U221 ( .A(n1107), .B(n1097), .Z(n1101) );
  XOR U222 ( .A(n434), .B(n484), .Z(n435) );
  MUX U223 ( .IN0(n482), .IN1(n480), .SEL(n481), .F(n428) );
  MUX U224 ( .IN0(n704), .IN1(n702), .SEL(n703), .F(n639) );
  MUX U225 ( .IN0(g_input[13]), .IN1(n1160), .SEL(g_input[15]), .F(n255) );
  MUX U226 ( .IN0(n66), .IN1(n523), .SEL(n524), .F(n459) );
  IV U227 ( .A(n525), .Z(n66) );
  XOR U228 ( .A(n659), .B(n596), .Z(n600) );
  XNOR U229 ( .A(n815), .B(n743), .Z(n747) );
  MUX U230 ( .IN0(n67), .IN1(n878), .SEL(n879), .F(n803) );
  IV U231 ( .A(n880), .Z(n67) );
  MUX U232 ( .IN0(n68), .IN1(n867), .SEL(n868), .F(n795) );
  IV U233 ( .A(n869), .Z(n68) );
  MUX U234 ( .IN0(g_input[14]), .IN1(n1137), .SEL(g_input[15]), .F(n220) );
  MUX U235 ( .IN0(n278), .IN1(n69), .SEL(n277), .F(n246) );
  IV U236 ( .A(n276), .Z(n69) );
  XNOR U237 ( .A(n580), .B(n579), .Z(n632) );
  MUX U238 ( .IN0(\_MxM/Y0[13] ), .IN1(n70), .SEL(n184), .F(n176) );
  IV U239 ( .A(n183), .Z(n70) );
  MUX U240 ( .IN0(n71), .IN1(n343), .SEL(n344), .F(n298) );
  IV U241 ( .A(\_MxM/Y0[9] ), .Z(n71) );
  MUX U242 ( .IN0(n72), .IN1(n832), .SEL(n833), .F(n755) );
  IV U243 ( .A(\_MxM/Y0[1] ), .Z(n72) );
  XOR U244 ( .A(n554), .B(n562), .Z(n560) );
  MUX U245 ( .IN0(n1218), .IN1(n73), .SEL(n1055), .F(n1199) );
  IV U246 ( .A(n1053), .Z(n73) );
  MUX U247 ( .IN0(n992), .IN1(n74), .SEL(n993), .F(n969) );
  IV U248 ( .A(n994), .Z(n74) );
  MUX U249 ( .IN0(n1275), .IN1(n1291), .SEL(n1277), .F(n1264) );
  MUX U250 ( .IN0(n1152), .IN1(n75), .SEL(n955), .F(n1142) );
  IV U251 ( .A(n953), .Z(n75) );
  MUX U252 ( .IN0(g_input[8]), .IN1(n1248), .SEL(g_input[15]), .F(n483) );
  MUX U253 ( .IN0(g_input[2]), .IN1(n1455), .SEL(g_input[15]), .F(n899) );
  MUX U254 ( .IN0(n76), .IN1(n846), .SEL(n847), .F(n771) );
  IV U255 ( .A(n848), .Z(n76) );
  MUX U256 ( .IN0(n77), .IN1(n405), .SEL(n406), .F(n362) );
  IV U257 ( .A(n407), .Z(n77) );
  MUX U258 ( .IN0(n534), .IN1(n536), .SEL(n535), .F(n463) );
  MUX U259 ( .IN0(n612), .IN1(n610), .SEL(n611), .F(n545) );
  XOR U260 ( .A(n829), .B(n900), .Z(n830) );
  MUX U261 ( .IN0(n852), .IN1(n850), .SEL(n851), .F(n775) );
  XNOR U262 ( .A(n281), .B(n282), .Z(n280) );
  MUX U263 ( .IN0(n78), .IN1(n408), .SEL(n409), .F(n365) );
  IV U264 ( .A(n410), .Z(n78) );
  XOR U265 ( .A(n575), .B(n576), .Z(n570) );
  XOR U266 ( .A(n806), .B(n732), .Z(n736) );
  XNOR U267 ( .A(n890), .B(n820), .Z(n824) );
  NAND U268 ( .A(n789), .B(n862), .Z(n861) );
  XNOR U269 ( .A(n285), .B(n284), .Z(n278) );
  XNOR U270 ( .A(n680), .B(n679), .Z(n658) );
  MUX U271 ( .IN0(n720), .IN1(n718), .SEL(n719), .F(n79) );
  IV U272 ( .A(n79), .Z(n647) );
  MUX U273 ( .IN0(n857), .IN1(n80), .SEL(n858), .F(n782) );
  IV U274 ( .A(n859), .Z(n80) );
  MUX U275 ( .IN0(n451), .IN1(n81), .SEL(n452), .F(n402) );
  IV U276 ( .A(n453), .Z(n81) );
  MUX U277 ( .IN0(n82), .IN1(n230), .SEL(n231), .F(n183) );
  IV U278 ( .A(\_MxM/Y0[12] ), .Z(n82) );
  MUX U279 ( .IN0(n83), .IN1(n388), .SEL(n389), .F(n343) );
  IV U280 ( .A(\_MxM/Y0[8] ), .Z(n83) );
  XOR U281 ( .A(n619), .B(n627), .Z(n625) );
  MUX U282 ( .IN0(n1199), .IN1(n84), .SEL(n1028), .F(n1180) );
  IV U283 ( .A(n1026), .Z(n84) );
  MUX U284 ( .IN0(n85), .IN1(n1343), .SEL(n1344), .F(n1393) );
  IV U285 ( .A(n1413), .Z(n85) );
  NOR U286 ( .A(g_input[0]), .B(n1465), .Z(n1456) );
  XOR U287 ( .A(n1323), .B(n1310), .Z(n1131) );
  MUX U288 ( .IN0(n1142), .IN1(n86), .SEL(n932), .F(n870) );
  IV U289 ( .A(n930), .Z(n86) );
  MUX U290 ( .IN0(n430), .IN1(n428), .SEL(n429), .F(n379) );
  XOR U291 ( .A(n684), .B(n750), .Z(n685) );
  MUX U292 ( .IN0(n364), .IN1(n87), .SEL(n363), .F(n317) );
  IV U293 ( .A(n362), .Z(n87) );
  MUX U294 ( .IN0(e_input[7]), .IN1(n1129), .SEL(e_input[15]), .F(n506) );
  XNOR U295 ( .A(n738), .B(n675), .Z(n679) );
  XOR U296 ( .A(n729), .B(n664), .Z(n668) );
  XNOR U297 ( .A(n844), .B(n772), .Z(n776) );
  XNOR U298 ( .A(n898), .B(n897), .Z(n880) );
  MUX U299 ( .IN0(n254), .IN1(n280), .SEL(n253), .F(n225) );
  XNOR U300 ( .A(n336), .B(n335), .Z(n325) );
  XNOR U301 ( .A(n547), .B(n546), .Z(n525) );
  XNOR U302 ( .A(n612), .B(n611), .Z(n590) );
  XNOR U303 ( .A(n718), .B(n785), .Z(n719) );
  XNOR U304 ( .A(n461), .B(n460), .Z(n453) );
  XOR U305 ( .A(n567), .B(n508), .Z(n516) );
  XNOR U306 ( .A(n728), .B(n727), .Z(n717) );
  XNOR U307 ( .A(n805), .B(n804), .Z(n784) );
  XNOR U308 ( .A(n244), .B(n243), .Z(n268) );
  MUX U309 ( .IN0(n88), .IN1(n437), .SEL(n438), .F(n388) );
  IV U310 ( .A(\_MxM/Y0[7] ), .Z(n88) );
  MUX U311 ( .IN0(\_MxM/Y0[14] ), .IN1(n176), .SEL(n177), .F(n166) );
  XOR U312 ( .A(n687), .B(n695), .Z(n693) );
  MUX U313 ( .IN0(n1046), .IN1(n89), .SEL(n1047), .F(n1019) );
  IV U314 ( .A(n1048), .Z(n89) );
  MUX U315 ( .IN0(n90), .IN1(n1130), .SEL(n1131), .F(n1303) );
  IV U316 ( .A(n1317), .Z(n90) );
  MUX U317 ( .IN0(n1180), .IN1(n91), .SEL(n1001), .F(n1165) );
  IV U318 ( .A(n999), .Z(n91) );
  XOR U319 ( .A(n1441), .B(g_input[3]), .Z(n1442) );
  MUX U320 ( .IN0(n946), .IN1(n92), .SEL(n947), .F(n912) );
  IV U321 ( .A(n948), .Z(n92) );
  XOR U322 ( .A(n1411), .B(n1412), .Z(n1343) );
  XOR U323 ( .A(n1262), .B(n1253), .Z(n1106) );
  MUX U324 ( .IN0(e_input[5]), .IN1(n1124), .SEL(e_input[15]), .F(n636) );
  MUX U325 ( .IN0(e_input[2]), .IN1(n1321), .SEL(e_input[15]), .F(n863) );
  XNOR U326 ( .A(n1102), .B(n1101), .Z(n919) );
  XNOR U327 ( .A(n326), .B(n290), .Z(n284) );
  MUX U328 ( .IN0(n370), .IN1(n368), .SEL(n369), .F(n93) );
  IV U329 ( .A(n93), .Z(n322) );
  XOR U330 ( .A(n644), .B(n645), .Z(n641) );
  XOR U331 ( .A(n881), .B(n809), .Z(n813) );
  MUX U332 ( .IN0(n872), .IN1(n1132), .SEL(n871), .F(n794) );
  XNOR U333 ( .A(n852), .B(n851), .Z(n869) );
  AND U334 ( .A(n214), .B(n191), .Z(n213) );
  XNOR U335 ( .A(n381), .B(n380), .Z(n367) );
  XNOR U336 ( .A(n430), .B(n429), .Z(n410) );
  XNOR U337 ( .A(n482), .B(n481), .Z(n461) );
  XNOR U338 ( .A(n704), .B(n703), .Z(n720) );
  XNOR U339 ( .A(n748), .B(n747), .Z(n728) );
  XNOR U340 ( .A(n825), .B(n824), .Z(n805) );
  XNOR U341 ( .A(n777), .B(n776), .Z(n797) );
  XNOR U342 ( .A(n880), .B(n879), .Z(n859) );
  XNOR U343 ( .A(n245), .B(n246), .Z(n244) );
  XNOR U344 ( .A(n525), .B(n524), .Z(n517) );
  XNOR U345 ( .A(n590), .B(n589), .Z(n582) );
  XNOR U346 ( .A(n658), .B(n657), .Z(n650) );
  MUX U347 ( .IN0(n94), .IN1(n298), .SEL(n299), .F(n261) );
  IV U348 ( .A(\_MxM/Y0[10] ), .Z(n94) );
  MUX U349 ( .IN0(n95), .IN1(n489), .SEL(n490), .F(n437) );
  IV U350 ( .A(\_MxM/Y0[6] ), .Z(n95) );
  MUX U351 ( .IN0(n96), .IN1(n755), .SEL(n756), .F(n687) );
  IV U352 ( .A(\_MxM/Y0[2] ), .Z(n96) );
  MUX U353 ( .IN0(\_MxM/Y0[15] ), .IN1(n166), .SEL(n167), .F(n97) );
  IV U354 ( .A(n97), .Z(n163) );
  XOR U355 ( .A(n833), .B(\_MxM/Y0[1] ), .Z(n108) );
  ANDN U356 ( .A(n98), .B(\_MxM/n[0] ), .Z(\_MxM/n229 ) );
  AND U357 ( .A(\_MxM/N8 ), .B(n98), .Z(\_MxM/n228 ) );
  AND U358 ( .A(\_MxM/N9 ), .B(n98), .Z(\_MxM/n227 ) );
  AND U359 ( .A(\_MxM/N10 ), .B(n98), .Z(\_MxM/n226 ) );
  AND U360 ( .A(\_MxM/N11 ), .B(n98), .Z(\_MxM/n225 ) );
  AND U361 ( .A(\_MxM/N12 ), .B(n98), .Z(\_MxM/n224 ) );
  AND U362 ( .A(n98), .B(n99), .Z(\_MxM/n223 ) );
  XOR U363 ( .A(\_MxM/n[6] ), .B(\_MxM/add_39/carry[6] ), .Z(n99) );
  ANDN U364 ( .A(n100), .B(rst), .Z(n98) );
  NAND U365 ( .A(n101), .B(n102), .Z(n100) );
  AND U366 ( .A(\_MxM/n[0] ), .B(n103), .Z(n102) );
  NOR U367 ( .A(n104), .B(\_MxM/n[2] ), .Z(n103) );
  AND U368 ( .A(n105), .B(\_MxM/n[6] ), .Z(n101) );
  AND U369 ( .A(\_MxM/n[5] ), .B(\_MxM/n[1] ), .Z(n105) );
  NAND U370 ( .A(n106), .B(n107), .Z(\_MxM/n222 ) );
  OR U371 ( .A(n108), .B(n109), .Z(n107) );
  NANDN U372 ( .B(n110), .A(\_MxM/Y0[0] ), .Z(n106) );
  NAND U373 ( .A(n111), .B(n112), .Z(\_MxM/n221 ) );
  NANDN U374 ( .B(n109), .A(n113), .Z(n112) );
  NANDN U375 ( .B(n114), .A(rst), .Z(n111) );
  NAND U376 ( .A(n115), .B(n116), .Z(\_MxM/n220 ) );
  NANDN U377 ( .B(n109), .A(n117), .Z(n116) );
  NANDN U378 ( .B(n110), .A(\_MxM/Y0[2] ), .Z(n115) );
  NAND U379 ( .A(n118), .B(n119), .Z(\_MxM/n219 ) );
  NANDN U380 ( .B(n109), .A(n120), .Z(n119) );
  NANDN U381 ( .B(n110), .A(\_MxM/Y0[3] ), .Z(n118) );
  NAND U382 ( .A(n121), .B(n122), .Z(\_MxM/n218 ) );
  NANDN U383 ( .B(n109), .A(n123), .Z(n122) );
  NANDN U384 ( .B(n110), .A(\_MxM/Y0[4] ), .Z(n121) );
  NAND U385 ( .A(n124), .B(n125), .Z(\_MxM/n217 ) );
  NANDN U386 ( .B(n109), .A(n126), .Z(n125) );
  NANDN U387 ( .B(n110), .A(\_MxM/Y0[5] ), .Z(n124) );
  NAND U388 ( .A(n127), .B(n128), .Z(\_MxM/n216 ) );
  NANDN U389 ( .B(n109), .A(n129), .Z(n128) );
  NANDN U390 ( .B(n110), .A(\_MxM/Y0[6] ), .Z(n127) );
  NAND U391 ( .A(n130), .B(n131), .Z(\_MxM/n215 ) );
  NANDN U392 ( .B(n109), .A(n132), .Z(n131) );
  NANDN U393 ( .B(n110), .A(\_MxM/Y0[7] ), .Z(n130) );
  NAND U394 ( .A(n133), .B(n134), .Z(\_MxM/n214 ) );
  NANDN U395 ( .B(n109), .A(n135), .Z(n134) );
  NANDN U396 ( .B(n110), .A(\_MxM/Y0[8] ), .Z(n133) );
  NAND U397 ( .A(n136), .B(n137), .Z(\_MxM/n213 ) );
  NANDN U398 ( .B(n109), .A(n138), .Z(n137) );
  NANDN U399 ( .B(n110), .A(\_MxM/Y0[9] ), .Z(n136) );
  NAND U400 ( .A(n139), .B(n140), .Z(\_MxM/n212 ) );
  NANDN U401 ( .B(n109), .A(n141), .Z(n140) );
  NANDN U402 ( .B(n110), .A(\_MxM/Y0[10] ), .Z(n139) );
  NAND U403 ( .A(n142), .B(n143), .Z(\_MxM/n211 ) );
  NANDN U404 ( .B(n109), .A(n144), .Z(n143) );
  NANDN U405 ( .B(n110), .A(\_MxM/Y0[11] ), .Z(n142) );
  NAND U406 ( .A(n145), .B(n146), .Z(\_MxM/n210 ) );
  NANDN U407 ( .B(n109), .A(n147), .Z(n146) );
  NANDN U408 ( .B(n110), .A(\_MxM/Y0[12] ), .Z(n145) );
  NAND U409 ( .A(n148), .B(n149), .Z(\_MxM/n209 ) );
  NANDN U410 ( .B(n109), .A(n150), .Z(n149) );
  NANDN U411 ( .B(n110), .A(\_MxM/Y0[13] ), .Z(n148) );
  NAND U412 ( .A(n151), .B(n152), .Z(\_MxM/n208 ) );
  OR U413 ( .A(n153), .B(n109), .Z(n152) );
  NANDN U414 ( .B(n110), .A(\_MxM/Y0[14] ), .Z(n151) );
  NAND U415 ( .A(n154), .B(n155), .Z(\_MxM/n207 ) );
  OR U416 ( .A(n109), .B(n156), .Z(n155) );
  NANDN U417 ( .B(n157), .A(n110), .Z(n109) );
  NANDN U418 ( .B(n110), .A(\_MxM/Y0[15] ), .Z(n154) );
  NAND U419 ( .A(n158), .B(n159), .Z(\_MxM/n206 ) );
  NANDN U420 ( .B(n110), .A(o[15]), .Z(n159) );
  AND U421 ( .A(n160), .B(n161), .Z(n158) );
  NANDN U422 ( .B(n157), .A(o[15]), .Z(n161) );
  OR U423 ( .A(n156), .B(n162), .Z(n160) );
  XOR U424 ( .A(n163), .B(n164), .Z(n156) );
  XNOR U425 ( .A(\_MxM/Y0[15] ), .B(n165), .Z(n164) );
  NAND U426 ( .A(n168), .B(n169), .Z(\_MxM/n205 ) );
  NANDN U427 ( .B(n110), .A(o[14]), .Z(n169) );
  AND U428 ( .A(n170), .B(n171), .Z(n168) );
  NANDN U429 ( .B(n157), .A(o[14]), .Z(n171) );
  OR U430 ( .A(n153), .B(n162), .Z(n170) );
  XOR U431 ( .A(n167), .B(\_MxM/Y0[15] ), .Z(n153) );
  XOR U432 ( .A(n166), .B(n165), .Z(n167) );
  NAND U433 ( .A(n172), .B(n173), .Z(n165) );
  OR U434 ( .A(n174), .B(n175), .Z(n172) );
  NAND U435 ( .A(n178), .B(n179), .Z(\_MxM/n204 ) );
  NANDN U436 ( .B(n110), .A(o[13]), .Z(n179) );
  AND U437 ( .A(n180), .B(n181), .Z(n178) );
  NANDN U438 ( .B(n157), .A(o[13]), .Z(n181) );
  NANDN U439 ( .B(n162), .A(n150), .Z(n180) );
  XNOR U440 ( .A(n177), .B(\_MxM/Y0[14] ), .Z(n150) );
  XNOR U441 ( .A(n182), .B(n176), .Z(n177) );
  XNOR U442 ( .A(n175), .B(n185), .Z(n174) );
  OR U443 ( .A(n186), .B(n187), .Z(n175) );
  AND U444 ( .A(n188), .B(n189), .Z(n185) );
  OR U445 ( .A(n190), .B(n191), .Z(n189) );
  AND U446 ( .A(n192), .B(n193), .Z(n188) );
  OR U447 ( .A(n194), .B(n195), .Z(n193) );
  OR U448 ( .A(n196), .B(n197), .Z(n192) );
  NAND U449 ( .A(n198), .B(n199), .Z(\_MxM/n203 ) );
  NANDN U450 ( .B(n110), .A(o[12]), .Z(n199) );
  AND U451 ( .A(n200), .B(n201), .Z(n198) );
  NANDN U452 ( .B(n157), .A(o[12]), .Z(n201) );
  NANDN U453 ( .B(n162), .A(n147), .Z(n200) );
  XNOR U454 ( .A(n184), .B(\_MxM/Y0[13] ), .Z(n147) );
  XNOR U455 ( .A(n202), .B(n203), .Z(n184) );
  AND U456 ( .A(n173), .B(n205), .Z(n204) );
  XOR U457 ( .A(n186), .B(n206), .Z(n205) );
  XOR U458 ( .A(n206), .B(n187), .Z(n186) );
  OR U459 ( .A(n207), .B(n208), .Z(n187) );
  IV U460 ( .A(n203), .Z(n206) );
  XNOR U461 ( .A(n197), .B(n196), .Z(n203) );
  OR U462 ( .A(n209), .B(n210), .Z(n196) );
  AND U463 ( .A(n211), .B(n212), .Z(n197) );
  XNOR U464 ( .A(n190), .B(n213), .Z(n212) );
  NAND U465 ( .A(n215), .B(n216), .Z(n191) );
  NANDN U466 ( .B(n217), .A(n218), .Z(n215) );
  NANDN U467 ( .B(n194), .A(n219), .Z(n214) );
  NANDN U468 ( .B(n195), .A(n220), .Z(n190) );
  AND U469 ( .A(n221), .B(n222), .Z(n211) );
  OR U470 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U471 ( .A(n225), .B(n226), .Z(n221) );
  ANDN U472 ( .A(n227), .B(n228), .Z(n226) );
  XOR U473 ( .A(n225), .B(n229), .Z(n227) );
  NAND U474 ( .A(n232), .B(n233), .Z(\_MxM/n202 ) );
  NANDN U475 ( .B(n110), .A(o[11]), .Z(n233) );
  AND U476 ( .A(n234), .B(n235), .Z(n232) );
  NANDN U477 ( .B(n157), .A(o[11]), .Z(n235) );
  NANDN U478 ( .B(n162), .A(n144), .Z(n234) );
  XNOR U479 ( .A(n231), .B(\_MxM/Y0[12] ), .Z(n144) );
  XNOR U480 ( .A(n236), .B(n237), .Z(n231) );
  AND U481 ( .A(n173), .B(n239), .Z(n238) );
  XOR U482 ( .A(n207), .B(n240), .Z(n239) );
  XOR U483 ( .A(n240), .B(n208), .Z(n207) );
  OR U484 ( .A(n241), .B(n242), .Z(n208) );
  IV U485 ( .A(n237), .Z(n240) );
  XNOR U486 ( .A(n210), .B(n209), .Z(n237) );
  OR U487 ( .A(n243), .B(n244), .Z(n209) );
  XNOR U488 ( .A(n224), .B(n223), .Z(n210) );
  OR U489 ( .A(n245), .B(n246), .Z(n223) );
  XOR U490 ( .A(n229), .B(n228), .Z(n224) );
  XOR U491 ( .A(n225), .B(n247), .Z(n228) );
  AND U492 ( .A(n248), .B(n249), .Z(n247) );
  NANDN U493 ( .B(n194), .A(n250), .Z(n249) );
  OR U494 ( .A(n251), .B(n252), .Z(n248) );
  XOR U495 ( .A(n217), .B(n218), .Z(n229) );
  NANDN U496 ( .B(n195), .A(n255), .Z(n218) );
  XNOR U497 ( .A(n216), .B(n256), .Z(n217) );
  AND U498 ( .A(n220), .B(n219), .Z(n256) );
  ANDN U499 ( .A(n257), .B(n258), .Z(n216) );
  NANDN U500 ( .B(n259), .A(n260), .Z(n257) );
  NAND U501 ( .A(n263), .B(n264), .Z(\_MxM/n201 ) );
  NANDN U502 ( .B(n110), .A(o[10]), .Z(n264) );
  AND U503 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U504 ( .B(n157), .A(o[10]), .Z(n266) );
  NANDN U505 ( .B(n162), .A(n141), .Z(n265) );
  XNOR U506 ( .A(n262), .B(\_MxM/Y0[11] ), .Z(n141) );
  XNOR U507 ( .A(n267), .B(n268), .Z(n262) );
  AND U508 ( .A(n173), .B(n270), .Z(n269) );
  XOR U509 ( .A(n241), .B(n271), .Z(n270) );
  XOR U510 ( .A(n271), .B(n242), .Z(n241) );
  OR U511 ( .A(n272), .B(n273), .Z(n242) );
  IV U512 ( .A(n268), .Z(n271) );
  OR U513 ( .A(n274), .B(n275), .Z(n243) );
  XOR U514 ( .A(n254), .B(n253), .Z(n245) );
  XNOR U515 ( .A(n279), .B(n280), .Z(n253) );
  ANDN U516 ( .A(n283), .B(n284), .Z(n282) );
  XOR U517 ( .A(n281), .B(n285), .Z(n283) );
  XNOR U518 ( .A(n286), .B(n251), .Z(n279) );
  NAND U519 ( .A(n250), .B(n220), .Z(n251) );
  NANDN U520 ( .B(n194), .A(n288), .Z(n287) );
  XOR U521 ( .A(n259), .B(n260), .Z(n254) );
  NANDN U522 ( .B(n195), .A(n292), .Z(n260) );
  AND U523 ( .A(n255), .B(n219), .Z(n293) );
  NAND U524 ( .A(n294), .B(n295), .Z(n258) );
  NANDN U525 ( .B(n296), .A(n297), .Z(n294) );
  NAND U526 ( .A(n300), .B(n301), .Z(\_MxM/n200 ) );
  NANDN U527 ( .B(n110), .A(o[9]), .Z(n301) );
  AND U528 ( .A(n302), .B(n303), .Z(n300) );
  NANDN U529 ( .B(n157), .A(o[9]), .Z(n303) );
  NANDN U530 ( .B(n162), .A(n138), .Z(n302) );
  XNOR U531 ( .A(n299), .B(\_MxM/Y0[10] ), .Z(n138) );
  XNOR U532 ( .A(n304), .B(n305), .Z(n299) );
  AND U533 ( .A(n173), .B(n307), .Z(n306) );
  XOR U534 ( .A(n272), .B(n308), .Z(n307) );
  XOR U535 ( .A(n308), .B(n273), .Z(n272) );
  OR U536 ( .A(n309), .B(n310), .Z(n273) );
  IV U537 ( .A(n305), .Z(n308) );
  XNOR U538 ( .A(n275), .B(n274), .Z(n305) );
  OR U539 ( .A(n311), .B(n312), .Z(n274) );
  XNOR U540 ( .A(n278), .B(n277), .Z(n275) );
  XOR U541 ( .A(n276), .B(n313), .Z(n277) );
  AND U542 ( .A(n314), .B(n315), .Z(n313) );
  OR U543 ( .A(n316), .B(n317), .Z(n315) );
  AND U544 ( .A(n318), .B(n319), .Z(n314) );
  NANDN U545 ( .B(n194), .A(n320), .Z(n319) );
  NAND U546 ( .A(n321), .B(n322), .Z(n318) );
  XNOR U547 ( .A(n289), .B(n327), .Z(n290) );
  AND U548 ( .A(n220), .B(n288), .Z(n327) );
  XOR U549 ( .A(n328), .B(n329), .Z(n289) );
  ANDN U550 ( .A(n330), .B(n331), .Z(n329) );
  XNOR U551 ( .A(n332), .B(n328), .Z(n330) );
  XOR U552 ( .A(n333), .B(n291), .Z(n326) );
  NAND U553 ( .A(n250), .B(n255), .Z(n291) );
  IV U554 ( .A(n281), .Z(n333) );
  XNOR U555 ( .A(n296), .B(n297), .Z(n285) );
  NANDN U556 ( .B(n195), .A(n337), .Z(n297) );
  XNOR U557 ( .A(n295), .B(n338), .Z(n296) );
  AND U558 ( .A(n292), .B(n219), .Z(n338) );
  ANDN U559 ( .A(n339), .B(n340), .Z(n295) );
  NANDN U560 ( .B(n341), .A(n342), .Z(n339) );
  NAND U561 ( .A(n345), .B(n346), .Z(\_MxM/n199 ) );
  NANDN U562 ( .B(n110), .A(o[8]), .Z(n346) );
  AND U563 ( .A(n347), .B(n348), .Z(n345) );
  NANDN U564 ( .B(n157), .A(o[8]), .Z(n348) );
  NANDN U565 ( .B(n162), .A(n135), .Z(n347) );
  XNOR U566 ( .A(n344), .B(\_MxM/Y0[9] ), .Z(n135) );
  XNOR U567 ( .A(n349), .B(n350), .Z(n344) );
  AND U568 ( .A(n173), .B(n352), .Z(n351) );
  XOR U569 ( .A(n309), .B(n353), .Z(n352) );
  XOR U570 ( .A(n353), .B(n310), .Z(n309) );
  OR U571 ( .A(n354), .B(n355), .Z(n310) );
  IV U572 ( .A(n350), .Z(n353) );
  XNOR U573 ( .A(n312), .B(n311), .Z(n350) );
  OR U574 ( .A(n356), .B(n357), .Z(n311) );
  XNOR U575 ( .A(n325), .B(n324), .Z(n312) );
  XOR U576 ( .A(n358), .B(n321), .Z(n324) );
  XNOR U577 ( .A(n359), .B(n316), .Z(n321) );
  NAND U578 ( .A(n320), .B(n220), .Z(n316) );
  NANDN U579 ( .B(n194), .A(n361), .Z(n360) );
  XNOR U580 ( .A(n322), .B(n323), .Z(n358) );
  XNOR U581 ( .A(n328), .B(n372), .Z(n331) );
  AND U582 ( .A(n255), .B(n288), .Z(n372) );
  XOR U583 ( .A(n373), .B(n374), .Z(n328) );
  ANDN U584 ( .A(n375), .B(n376), .Z(n374) );
  XNOR U585 ( .A(n377), .B(n373), .Z(n375) );
  XOR U586 ( .A(n378), .B(n332), .Z(n371) );
  NAND U587 ( .A(n250), .B(n292), .Z(n332) );
  IV U588 ( .A(n334), .Z(n378) );
  XNOR U589 ( .A(n341), .B(n342), .Z(n336) );
  NANDN U590 ( .B(n195), .A(n382), .Z(n342) );
  AND U591 ( .A(n337), .B(n219), .Z(n383) );
  NAND U592 ( .A(n384), .B(n385), .Z(n340) );
  NANDN U593 ( .B(n386), .A(n387), .Z(n384) );
  NAND U594 ( .A(n390), .B(n391), .Z(\_MxM/n198 ) );
  NANDN U595 ( .B(n110), .A(o[7]), .Z(n391) );
  AND U596 ( .A(n392), .B(n393), .Z(n390) );
  NANDN U597 ( .B(n157), .A(o[7]), .Z(n393) );
  NANDN U598 ( .B(n162), .A(n132), .Z(n392) );
  XNOR U599 ( .A(n389), .B(\_MxM/Y0[8] ), .Z(n132) );
  XNOR U600 ( .A(n394), .B(n395), .Z(n389) );
  AND U601 ( .A(n173), .B(n397), .Z(n396) );
  XOR U602 ( .A(n354), .B(n398), .Z(n397) );
  XOR U603 ( .A(n398), .B(n355), .Z(n354) );
  OR U604 ( .A(n399), .B(n400), .Z(n355) );
  IV U605 ( .A(n395), .Z(n398) );
  XNOR U606 ( .A(n357), .B(n356), .Z(n395) );
  NANDN U607 ( .B(n401), .A(n402), .Z(n356) );
  XNOR U608 ( .A(n367), .B(n366), .Z(n357) );
  XOR U609 ( .A(n403), .B(n370), .Z(n366) );
  XNOR U610 ( .A(n363), .B(n364), .Z(n370) );
  NAND U611 ( .A(n320), .B(n255), .Z(n364) );
  XNOR U612 ( .A(n362), .B(n404), .Z(n363) );
  AND U613 ( .A(n220), .B(n361), .Z(n404) );
  XNOR U614 ( .A(n369), .B(n365), .Z(n403) );
  AND U615 ( .A(n412), .B(n413), .Z(n411) );
  NANDN U616 ( .B(n194), .A(n414), .Z(n413) );
  OR U617 ( .A(n415), .B(n416), .Z(n412) );
  XNOR U618 ( .A(n373), .B(n421), .Z(n376) );
  AND U619 ( .A(n292), .B(n288), .Z(n421) );
  XOR U620 ( .A(n422), .B(n423), .Z(n373) );
  ANDN U621 ( .A(n424), .B(n425), .Z(n423) );
  XNOR U622 ( .A(n426), .B(n422), .Z(n424) );
  XOR U623 ( .A(n427), .B(n377), .Z(n420) );
  NAND U624 ( .A(n250), .B(n337), .Z(n377) );
  IV U625 ( .A(n379), .Z(n427) );
  XNOR U626 ( .A(n386), .B(n387), .Z(n381) );
  NANDN U627 ( .B(n195), .A(n431), .Z(n387) );
  XNOR U628 ( .A(n385), .B(n432), .Z(n386) );
  AND U629 ( .A(n382), .B(n219), .Z(n432) );
  ANDN U630 ( .A(n433), .B(n434), .Z(n385) );
  NANDN U631 ( .B(n435), .A(n436), .Z(n433) );
  NAND U632 ( .A(n439), .B(n440), .Z(\_MxM/n197 ) );
  NANDN U633 ( .B(n110), .A(o[6]), .Z(n440) );
  AND U634 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U635 ( .B(n157), .A(o[6]), .Z(n442) );
  NANDN U636 ( .B(n162), .A(n129), .Z(n441) );
  XNOR U637 ( .A(n438), .B(\_MxM/Y0[7] ), .Z(n129) );
  XNOR U638 ( .A(n444), .B(n445), .Z(n443) );
  AND U639 ( .A(n173), .B(n446), .Z(n445) );
  XOR U640 ( .A(n399), .B(n449), .Z(n446) );
  XOR U641 ( .A(n449), .B(n400), .Z(n399) );
  OR U642 ( .A(n447), .B(n448), .Z(n400) );
  XNOR U643 ( .A(n401), .B(n402), .Z(n449) );
  XNOR U644 ( .A(n410), .B(n409), .Z(n401) );
  XOR U645 ( .A(n454), .B(n419), .Z(n409) );
  XNOR U646 ( .A(n406), .B(n407), .Z(n419) );
  NAND U647 ( .A(n320), .B(n292), .Z(n407) );
  XNOR U648 ( .A(n405), .B(n455), .Z(n406) );
  AND U649 ( .A(n255), .B(n361), .Z(n455) );
  XNOR U650 ( .A(n418), .B(n408), .Z(n454) );
  XNOR U651 ( .A(n462), .B(n417), .Z(n418) );
  XNOR U652 ( .A(n466), .B(n415), .Z(n462) );
  NAND U653 ( .A(n414), .B(n220), .Z(n415) );
  NANDN U654 ( .B(n194), .A(n468), .Z(n467) );
  XNOR U655 ( .A(n422), .B(n473), .Z(n425) );
  AND U656 ( .A(n337), .B(n288), .Z(n473) );
  XOR U657 ( .A(n474), .B(n475), .Z(n422) );
  ANDN U658 ( .A(n476), .B(n477), .Z(n475) );
  XNOR U659 ( .A(n478), .B(n474), .Z(n476) );
  XOR U660 ( .A(n479), .B(n426), .Z(n472) );
  NAND U661 ( .A(n250), .B(n382), .Z(n426) );
  IV U662 ( .A(n428), .Z(n479) );
  XNOR U663 ( .A(n435), .B(n436), .Z(n430) );
  NANDN U664 ( .B(n195), .A(n483), .Z(n436) );
  AND U665 ( .A(n431), .B(n219), .Z(n484) );
  NAND U666 ( .A(n485), .B(n486), .Z(n434) );
  NANDN U667 ( .B(n487), .A(n488), .Z(n485) );
  IV U668 ( .A(n437), .Z(n444) );
  NAND U669 ( .A(n491), .B(n492), .Z(\_MxM/n196 ) );
  NANDN U670 ( .B(n110), .A(o[5]), .Z(n492) );
  AND U671 ( .A(n493), .B(n494), .Z(n491) );
  NANDN U672 ( .B(n157), .A(o[5]), .Z(n494) );
  NANDN U673 ( .B(n162), .A(n126), .Z(n493) );
  XNOR U674 ( .A(n490), .B(\_MxM/Y0[6] ), .Z(n126) );
  XNOR U675 ( .A(n495), .B(n496), .Z(n490) );
  AND U676 ( .A(n173), .B(n498), .Z(n497) );
  XOR U677 ( .A(n447), .B(n499), .Z(n498) );
  XOR U678 ( .A(n499), .B(n448), .Z(n447) );
  OR U679 ( .A(n500), .B(n501), .Z(n448) );
  IV U680 ( .A(n496), .Z(n499) );
  XOR U681 ( .A(n453), .B(n452), .Z(n496) );
  XNOR U682 ( .A(n451), .B(n502), .Z(n452) );
  AND U683 ( .A(n450), .B(n503), .Z(n502) );
  AND U684 ( .A(n504), .B(n505), .Z(n503) );
  NANDN U685 ( .B(n194), .A(n506), .Z(n505) );
  OR U686 ( .A(n507), .B(n508), .Z(n504) );
  AND U687 ( .A(n509), .B(n510), .Z(n450) );
  NANDN U688 ( .B(n511), .A(n512), .Z(n510) );
  NANDN U689 ( .B(n513), .A(n514), .Z(n509) );
  XNOR U690 ( .A(n518), .B(n465), .Z(n460) );
  XNOR U691 ( .A(n457), .B(n458), .Z(n465) );
  NAND U692 ( .A(n320), .B(n337), .Z(n458) );
  XNOR U693 ( .A(n456), .B(n519), .Z(n457) );
  AND U694 ( .A(n292), .B(n361), .Z(n519) );
  XNOR U695 ( .A(n464), .B(n459), .Z(n518) );
  XNOR U696 ( .A(n469), .B(n527), .Z(n470) );
  AND U697 ( .A(n220), .B(n468), .Z(n527) );
  XOR U698 ( .A(n528), .B(n529), .Z(n469) );
  ANDN U699 ( .A(n530), .B(n531), .Z(n529) );
  XNOR U700 ( .A(n532), .B(n528), .Z(n530) );
  XOR U701 ( .A(n533), .B(n471), .Z(n526) );
  NAND U702 ( .A(n414), .B(n255), .Z(n471) );
  IV U703 ( .A(n463), .Z(n533) );
  XNOR U704 ( .A(n474), .B(n538), .Z(n477) );
  AND U705 ( .A(n382), .B(n288), .Z(n538) );
  XOR U706 ( .A(n539), .B(n540), .Z(n474) );
  ANDN U707 ( .A(n541), .B(n542), .Z(n540) );
  XNOR U708 ( .A(n543), .B(n539), .Z(n541) );
  XOR U709 ( .A(n544), .B(n478), .Z(n537) );
  NAND U710 ( .A(n250), .B(n431), .Z(n478) );
  IV U711 ( .A(n480), .Z(n544) );
  XNOR U712 ( .A(n487), .B(n488), .Z(n482) );
  NANDN U713 ( .B(n195), .A(n548), .Z(n488) );
  XNOR U714 ( .A(n486), .B(n549), .Z(n487) );
  AND U715 ( .A(n483), .B(n219), .Z(n549) );
  ANDN U716 ( .A(n550), .B(n551), .Z(n486) );
  NANDN U717 ( .B(n552), .A(n553), .Z(n550) );
  NAND U718 ( .A(n556), .B(n557), .Z(\_MxM/n195 ) );
  NANDN U719 ( .B(n110), .A(o[4]), .Z(n557) );
  AND U720 ( .A(n558), .B(n559), .Z(n556) );
  NANDN U721 ( .B(n157), .A(o[4]), .Z(n559) );
  NANDN U722 ( .B(n162), .A(n123), .Z(n558) );
  XNOR U723 ( .A(n555), .B(\_MxM/Y0[5] ), .Z(n123) );
  XNOR U724 ( .A(n560), .B(n561), .Z(n555) );
  AND U725 ( .A(n173), .B(n563), .Z(n562) );
  XOR U726 ( .A(n500), .B(n564), .Z(n563) );
  XOR U727 ( .A(n564), .B(n501), .Z(n500) );
  OR U728 ( .A(n565), .B(n566), .Z(n501) );
  IV U729 ( .A(n561), .Z(n564) );
  XOR U730 ( .A(n517), .B(n516), .Z(n561) );
  XOR U731 ( .A(n511), .B(n512), .Z(n508) );
  XOR U732 ( .A(n571), .B(n513), .Z(n511) );
  NAND U733 ( .A(n220), .B(n506), .Z(n513) );
  NANDN U734 ( .B(n514), .A(n572), .Z(n571) );
  NANDN U735 ( .B(n194), .A(n573), .Z(n572) );
  XOR U736 ( .A(n577), .B(n507), .Z(n567) );
  OR U737 ( .A(n578), .B(n579), .Z(n507) );
  IV U738 ( .A(n515), .Z(n577) );
  XNOR U739 ( .A(n583), .B(n536), .Z(n524) );
  XNOR U740 ( .A(n521), .B(n522), .Z(n536) );
  NAND U741 ( .A(n320), .B(n382), .Z(n522) );
  XNOR U742 ( .A(n520), .B(n584), .Z(n521) );
  AND U743 ( .A(n337), .B(n361), .Z(n584) );
  XNOR U744 ( .A(n535), .B(n523), .Z(n583) );
  XNOR U745 ( .A(n528), .B(n592), .Z(n531) );
  AND U746 ( .A(n255), .B(n468), .Z(n592) );
  XOR U747 ( .A(n593), .B(n594), .Z(n528) );
  ANDN U748 ( .A(n595), .B(n596), .Z(n594) );
  XNOR U749 ( .A(n597), .B(n593), .Z(n595) );
  XOR U750 ( .A(n598), .B(n532), .Z(n591) );
  NAND U751 ( .A(n414), .B(n292), .Z(n532) );
  IV U752 ( .A(n534), .Z(n598) );
  XNOR U753 ( .A(n539), .B(n603), .Z(n542) );
  AND U754 ( .A(n431), .B(n288), .Z(n603) );
  XOR U755 ( .A(n604), .B(n605), .Z(n539) );
  ANDN U756 ( .A(n606), .B(n607), .Z(n605) );
  XNOR U757 ( .A(n608), .B(n604), .Z(n606) );
  XOR U758 ( .A(n609), .B(n543), .Z(n602) );
  NAND U759 ( .A(n250), .B(n483), .Z(n543) );
  IV U760 ( .A(n545), .Z(n609) );
  XNOR U761 ( .A(n552), .B(n553), .Z(n547) );
  NANDN U762 ( .B(n195), .A(n613), .Z(n553) );
  AND U763 ( .A(n548), .B(n219), .Z(n614) );
  NAND U764 ( .A(n615), .B(n616), .Z(n551) );
  NANDN U765 ( .B(n617), .A(n618), .Z(n615) );
  NAND U766 ( .A(n621), .B(n622), .Z(\_MxM/n194 ) );
  NANDN U767 ( .B(n110), .A(o[3]), .Z(n622) );
  AND U768 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U769 ( .B(n157), .A(o[3]), .Z(n624) );
  NANDN U770 ( .B(n162), .A(n120), .Z(n623) );
  XNOR U771 ( .A(n620), .B(\_MxM/Y0[4] ), .Z(n120) );
  XNOR U772 ( .A(n625), .B(n626), .Z(n620) );
  AND U773 ( .A(n173), .B(n628), .Z(n627) );
  XOR U774 ( .A(n565), .B(n629), .Z(n628) );
  XOR U775 ( .A(n629), .B(n566), .Z(n565) );
  OR U776 ( .A(n630), .B(n631), .Z(n566) );
  IV U777 ( .A(n626), .Z(n629) );
  XOR U778 ( .A(n582), .B(n581), .Z(n626) );
  XOR U779 ( .A(n632), .B(n578), .Z(n581) );
  XOR U780 ( .A(n570), .B(n569), .Z(n578) );
  XOR U781 ( .A(n568), .B(n633), .Z(n569) );
  AND U782 ( .A(n634), .B(n635), .Z(n633) );
  NANDN U783 ( .B(n194), .A(n636), .Z(n635) );
  OR U784 ( .A(n637), .B(n638), .Z(n634) );
  NAND U785 ( .A(n255), .B(n506), .Z(n576) );
  XNOR U786 ( .A(n574), .B(n642), .Z(n575) );
  AND U787 ( .A(n573), .B(n220), .Z(n642) );
  NANDN U788 ( .B(n646), .A(n647), .Z(n579) );
  XNOR U789 ( .A(n651), .B(n601), .Z(n589) );
  XNOR U790 ( .A(n586), .B(n587), .Z(n601) );
  NAND U791 ( .A(n320), .B(n431), .Z(n587) );
  XNOR U792 ( .A(n585), .B(n652), .Z(n586) );
  AND U793 ( .A(n382), .B(n361), .Z(n652) );
  XNOR U794 ( .A(n600), .B(n588), .Z(n651) );
  XNOR U795 ( .A(n593), .B(n660), .Z(n596) );
  AND U796 ( .A(n292), .B(n468), .Z(n660) );
  XOR U797 ( .A(n661), .B(n662), .Z(n593) );
  ANDN U798 ( .A(n663), .B(n664), .Z(n662) );
  XNOR U799 ( .A(n665), .B(n661), .Z(n663) );
  XOR U800 ( .A(n666), .B(n597), .Z(n659) );
  NAND U801 ( .A(n414), .B(n337), .Z(n597) );
  IV U802 ( .A(n599), .Z(n666) );
  XNOR U803 ( .A(n604), .B(n671), .Z(n607) );
  AND U804 ( .A(n483), .B(n288), .Z(n671) );
  XOR U805 ( .A(n672), .B(n673), .Z(n604) );
  ANDN U806 ( .A(n674), .B(n675), .Z(n673) );
  XNOR U807 ( .A(n676), .B(n672), .Z(n674) );
  XOR U808 ( .A(n677), .B(n608), .Z(n670) );
  NAND U809 ( .A(n250), .B(n548), .Z(n608) );
  IV U810 ( .A(n610), .Z(n677) );
  XNOR U811 ( .A(n617), .B(n618), .Z(n612) );
  NANDN U812 ( .B(n195), .A(n681), .Z(n618) );
  XNOR U813 ( .A(n616), .B(n682), .Z(n617) );
  AND U814 ( .A(n613), .B(n219), .Z(n682) );
  ANDN U815 ( .A(n683), .B(n684), .Z(n616) );
  NANDN U816 ( .B(n685), .A(n686), .Z(n683) );
  NAND U817 ( .A(n689), .B(n690), .Z(\_MxM/n193 ) );
  NANDN U818 ( .B(n110), .A(o[2]), .Z(n690) );
  AND U819 ( .A(n691), .B(n692), .Z(n689) );
  NANDN U820 ( .B(n157), .A(o[2]), .Z(n692) );
  NANDN U821 ( .B(n162), .A(n117), .Z(n691) );
  XNOR U822 ( .A(n688), .B(\_MxM/Y0[3] ), .Z(n117) );
  XNOR U823 ( .A(n693), .B(n694), .Z(n688) );
  AND U824 ( .A(n173), .B(n696), .Z(n695) );
  XOR U825 ( .A(n630), .B(n697), .Z(n696) );
  XOR U826 ( .A(n697), .B(n631), .Z(n630) );
  OR U827 ( .A(n698), .B(n699), .Z(n631) );
  IV U828 ( .A(n694), .Z(n697) );
  XOR U829 ( .A(n650), .B(n649), .Z(n694) );
  XOR U830 ( .A(n700), .B(n646), .Z(n649) );
  XOR U831 ( .A(n641), .B(n640), .Z(n646) );
  XNOR U832 ( .A(n705), .B(n637), .Z(n701) );
  NAND U833 ( .A(n220), .B(n636), .Z(n637) );
  NANDN U834 ( .B(n194), .A(n707), .Z(n706) );
  NAND U835 ( .A(n292), .B(n506), .Z(n645) );
  XNOR U836 ( .A(n643), .B(n711), .Z(n644) );
  AND U837 ( .A(n573), .B(n255), .Z(n711) );
  XNOR U838 ( .A(n647), .B(n648), .Z(n700) );
  XNOR U839 ( .A(n721), .B(n669), .Z(n657) );
  XNOR U840 ( .A(n654), .B(n655), .Z(n669) );
  NAND U841 ( .A(n320), .B(n483), .Z(n655) );
  XNOR U842 ( .A(n653), .B(n722), .Z(n654) );
  AND U843 ( .A(n431), .B(n361), .Z(n722) );
  XNOR U844 ( .A(n668), .B(n656), .Z(n721) );
  XNOR U845 ( .A(n661), .B(n730), .Z(n664) );
  AND U846 ( .A(n337), .B(n468), .Z(n730) );
  XOR U847 ( .A(n734), .B(n665), .Z(n729) );
  NAND U848 ( .A(n414), .B(n382), .Z(n665) );
  IV U849 ( .A(n667), .Z(n734) );
  XNOR U850 ( .A(n672), .B(n739), .Z(n675) );
  AND U851 ( .A(n548), .B(n288), .Z(n739) );
  XOR U852 ( .A(n740), .B(n741), .Z(n672) );
  ANDN U853 ( .A(n742), .B(n743), .Z(n741) );
  XNOR U854 ( .A(n744), .B(n740), .Z(n742) );
  XOR U855 ( .A(n745), .B(n676), .Z(n738) );
  NAND U856 ( .A(n250), .B(n613), .Z(n676) );
  IV U857 ( .A(n678), .Z(n745) );
  XNOR U858 ( .A(n685), .B(n686), .Z(n680) );
  OR U859 ( .A(n749), .B(n195), .Z(n686) );
  AND U860 ( .A(n681), .B(n219), .Z(n750) );
  NAND U861 ( .A(n751), .B(n752), .Z(n684) );
  NANDN U862 ( .B(n753), .A(n754), .Z(n751) );
  NAND U863 ( .A(n757), .B(n758), .Z(\_MxM/n192 ) );
  NANDN U864 ( .B(n110), .A(o[1]), .Z(n758) );
  AND U865 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U866 ( .B(n157), .A(o[1]), .Z(n760) );
  NANDN U867 ( .B(n162), .A(n113), .Z(n759) );
  XNOR U868 ( .A(n756), .B(\_MxM/Y0[2] ), .Z(n113) );
  XNOR U869 ( .A(n761), .B(n762), .Z(n756) );
  XOR U870 ( .A(n755), .B(n763), .Z(n761) );
  AND U871 ( .A(n173), .B(n764), .Z(n763) );
  XOR U872 ( .A(n698), .B(n765), .Z(n764) );
  XOR U873 ( .A(n765), .B(n699), .Z(n698) );
  NANDN U874 ( .B(n766), .A(n767), .Z(n699) );
  IV U875 ( .A(n762), .Z(n765) );
  XOR U876 ( .A(n717), .B(n716), .Z(n762) );
  XNOR U877 ( .A(n768), .B(n720), .Z(n716) );
  XNOR U878 ( .A(n708), .B(n770), .Z(n709) );
  AND U879 ( .A(n707), .B(n220), .Z(n770) );
  XOR U880 ( .A(n774), .B(n710), .Z(n769) );
  NAND U881 ( .A(n255), .B(n636), .Z(n710) );
  IV U882 ( .A(n702), .Z(n774) );
  XNOR U883 ( .A(n713), .B(n714), .Z(n704) );
  NAND U884 ( .A(n337), .B(n506), .Z(n714) );
  XNOR U885 ( .A(n712), .B(n778), .Z(n713) );
  AND U886 ( .A(n573), .B(n292), .Z(n778) );
  XNOR U887 ( .A(n719), .B(n715), .Z(n768) );
  AND U888 ( .A(n786), .B(n787), .Z(n785) );
  OR U889 ( .A(n788), .B(n789), .Z(n787) );
  AND U890 ( .A(n790), .B(n791), .Z(n786) );
  NANDN U891 ( .B(n194), .A(n792), .Z(n791) );
  NANDN U892 ( .B(n793), .A(n794), .Z(n790) );
  XNOR U893 ( .A(n798), .B(n737), .Z(n727) );
  XNOR U894 ( .A(n724), .B(n725), .Z(n737) );
  NAND U895 ( .A(n320), .B(n548), .Z(n725) );
  XNOR U896 ( .A(n723), .B(n799), .Z(n724) );
  AND U897 ( .A(n483), .B(n361), .Z(n799) );
  XNOR U898 ( .A(n736), .B(n726), .Z(n798) );
  XNOR U899 ( .A(n731), .B(n807), .Z(n732) );
  AND U900 ( .A(n382), .B(n468), .Z(n807) );
  XOR U901 ( .A(n811), .B(n733), .Z(n806) );
  NAND U902 ( .A(n414), .B(n431), .Z(n733) );
  IV U903 ( .A(n735), .Z(n811) );
  XNOR U904 ( .A(n740), .B(n816), .Z(n743) );
  AND U905 ( .A(n613), .B(n288), .Z(n816) );
  XOR U906 ( .A(n817), .B(n818), .Z(n740) );
  ANDN U907 ( .A(n819), .B(n820), .Z(n818) );
  XNOR U908 ( .A(n821), .B(n817), .Z(n819) );
  XOR U909 ( .A(n822), .B(n744), .Z(n815) );
  NAND U910 ( .A(n250), .B(n681), .Z(n744) );
  IV U911 ( .A(n746), .Z(n822) );
  XNOR U912 ( .A(n753), .B(n754), .Z(n748) );
  OR U913 ( .A(n826), .B(n195), .Z(n754) );
  XNOR U914 ( .A(n752), .B(n827), .Z(n753) );
  ANDN U915 ( .A(n219), .B(n749), .Z(n827) );
  ANDN U916 ( .A(n828), .B(n829), .Z(n752) );
  NANDN U917 ( .B(n830), .A(n831), .Z(n828) );
  NAND U918 ( .A(n834), .B(n835), .Z(\_MxM/n191 ) );
  NANDN U919 ( .B(n110), .A(o[0]), .Z(n835) );
  AND U920 ( .A(n836), .B(n837), .Z(n834) );
  NANDN U921 ( .B(n157), .A(o[0]), .Z(n837) );
  IV U922 ( .A(n838), .Z(n157) );
  OR U923 ( .A(n162), .B(n108), .Z(n836) );
  IV U924 ( .A(\_MxM/Y0[1] ), .Z(n114) );
  XOR U925 ( .A(n839), .B(n840), .Z(n833) );
  XNOR U926 ( .A(n841), .B(n832), .Z(n839) );
  NAND U927 ( .A(\_MxM/Y0[0] ), .B(n766), .Z(n832) );
  NAND U928 ( .A(n842), .B(n173), .Z(n841) );
  XOR U929 ( .A(e_input[15]), .B(g_input[15]), .Z(n173) );
  XNOR U930 ( .A(n767), .B(n840), .Z(n842) );
  XNOR U931 ( .A(n766), .B(n840), .Z(n767) );
  XNOR U932 ( .A(n784), .B(n783), .Z(n840) );
  XNOR U933 ( .A(n843), .B(n797), .Z(n783) );
  XNOR U934 ( .A(n771), .B(n845), .Z(n772) );
  AND U935 ( .A(n707), .B(n255), .Z(n845) );
  XOR U936 ( .A(n849), .B(n773), .Z(n844) );
  NAND U937 ( .A(n292), .B(n636), .Z(n773) );
  IV U938 ( .A(n775), .Z(n849) );
  XNOR U939 ( .A(n780), .B(n781), .Z(n777) );
  NAND U940 ( .A(n382), .B(n506), .Z(n781) );
  XNOR U941 ( .A(n779), .B(n853), .Z(n780) );
  AND U942 ( .A(n573), .B(n337), .Z(n853) );
  XNOR U943 ( .A(n796), .B(n782), .Z(n843) );
  XNOR U944 ( .A(n860), .B(n793), .Z(n796) );
  XOR U945 ( .A(n861), .B(n788), .Z(n793) );
  NAND U946 ( .A(n220), .B(n792), .Z(n788) );
  NANDN U947 ( .B(n194), .A(n863), .Z(n862) );
  XNOR U948 ( .A(n794), .B(n795), .Z(n860) );
  XNOR U949 ( .A(n873), .B(n814), .Z(n804) );
  XNOR U950 ( .A(n801), .B(n802), .Z(n814) );
  NAND U951 ( .A(n320), .B(n613), .Z(n802) );
  XNOR U952 ( .A(n800), .B(n874), .Z(n801) );
  AND U953 ( .A(n548), .B(n361), .Z(n874) );
  XNOR U954 ( .A(n813), .B(n803), .Z(n873) );
  XNOR U955 ( .A(n808), .B(n882), .Z(n809) );
  AND U956 ( .A(n431), .B(n468), .Z(n882) );
  XOR U957 ( .A(n886), .B(n810), .Z(n881) );
  NAND U958 ( .A(n414), .B(n483), .Z(n810) );
  IV U959 ( .A(n812), .Z(n886) );
  XNOR U960 ( .A(n817), .B(n891), .Z(n820) );
  AND U961 ( .A(n681), .B(n288), .Z(n891) );
  XOR U962 ( .A(n895), .B(n821), .Z(n890) );
  NANDN U963 ( .B(n749), .A(n250), .Z(n821) );
  IV U964 ( .A(n823), .Z(n895) );
  XNOR U965 ( .A(n830), .B(n831), .Z(n825) );
  NANDN U966 ( .B(n195), .A(n899), .Z(n831) );
  ANDN U967 ( .A(n219), .B(n826), .Z(n900) );
  NAND U968 ( .A(n901), .B(n902), .Z(n829) );
  NANDN U969 ( .B(n903), .A(n904), .Z(n901) );
  XNOR U970 ( .A(n859), .B(n858), .Z(n766) );
  XNOR U971 ( .A(n905), .B(n869), .Z(n858) );
  XNOR U972 ( .A(n846), .B(n907), .Z(n847) );
  AND U973 ( .A(n707), .B(n292), .Z(n907) );
  XOR U974 ( .A(n911), .B(n848), .Z(n906) );
  NAND U975 ( .A(n337), .B(n636), .Z(n848) );
  IV U976 ( .A(n850), .Z(n911) );
  XNOR U977 ( .A(n855), .B(n856), .Z(n852) );
  NAND U978 ( .A(n431), .B(n506), .Z(n856) );
  XNOR U979 ( .A(n854), .B(n915), .Z(n855) );
  AND U980 ( .A(n573), .B(n382), .Z(n915) );
  XNOR U981 ( .A(n868), .B(n857), .Z(n905) );
  XOR U982 ( .A(n919), .B(n920), .Z(n857) );
  XNOR U983 ( .A(n921), .B(n872), .Z(n868) );
  NAND U984 ( .A(n255), .B(n792), .Z(n866) );
  XNOR U985 ( .A(n864), .B(n922), .Z(n865) );
  AND U986 ( .A(n863), .B(n220), .Z(n922) );
  XNOR U987 ( .A(n871), .B(n867), .Z(n921) );
  XOR U988 ( .A(n926), .B(n927), .Z(n867) );
  AND U989 ( .A(n928), .B(n929), .Z(n927) );
  XOR U990 ( .A(n930), .B(n931), .Z(n929) );
  XOR U991 ( .A(n926), .B(n932), .Z(n931) );
  XOR U992 ( .A(n913), .B(n933), .Z(n928) );
  XOR U993 ( .A(n926), .B(n914), .Z(n933) );
  NAND U994 ( .A(n506), .B(n483), .Z(n918) );
  XNOR U995 ( .A(n916), .B(n934), .Z(n917) );
  AND U996 ( .A(n573), .B(n431), .Z(n934) );
  XNOR U997 ( .A(n908), .B(n939), .Z(n909) );
  AND U998 ( .A(n707), .B(n337), .Z(n939) );
  XOR U999 ( .A(n940), .B(n941), .Z(n908) );
  ANDN U1000 ( .A(n942), .B(n943), .Z(n941) );
  XNOR U1001 ( .A(n944), .B(n940), .Z(n942) );
  XOR U1002 ( .A(n945), .B(n910), .Z(n938) );
  NAND U1003 ( .A(n382), .B(n636), .Z(n910) );
  IV U1004 ( .A(n912), .Z(n945) );
  XOR U1005 ( .A(n949), .B(n950), .Z(n926) );
  AND U1006 ( .A(n951), .B(n952), .Z(n950) );
  XOR U1007 ( .A(n953), .B(n954), .Z(n952) );
  XOR U1008 ( .A(n949), .B(n955), .Z(n954) );
  XOR U1009 ( .A(n947), .B(n956), .Z(n951) );
  XOR U1010 ( .A(n949), .B(n948), .Z(n956) );
  NAND U1011 ( .A(n506), .B(n548), .Z(n937) );
  XNOR U1012 ( .A(n935), .B(n957), .Z(n936) );
  AND U1013 ( .A(n483), .B(n573), .Z(n957) );
  XNOR U1014 ( .A(n940), .B(n962), .Z(n943) );
  AND U1015 ( .A(n707), .B(n382), .Z(n962) );
  XOR U1016 ( .A(n963), .B(n964), .Z(n940) );
  ANDN U1017 ( .A(n965), .B(n966), .Z(n964) );
  XNOR U1018 ( .A(n967), .B(n963), .Z(n965) );
  XOR U1019 ( .A(n968), .B(n944), .Z(n961) );
  NAND U1020 ( .A(n431), .B(n636), .Z(n944) );
  IV U1021 ( .A(n946), .Z(n968) );
  XOR U1022 ( .A(n972), .B(n973), .Z(n949) );
  AND U1023 ( .A(n974), .B(n975), .Z(n973) );
  XOR U1024 ( .A(n976), .B(n977), .Z(n975) );
  XOR U1025 ( .A(n972), .B(n978), .Z(n977) );
  XOR U1026 ( .A(n970), .B(n979), .Z(n974) );
  XOR U1027 ( .A(n972), .B(n971), .Z(n979) );
  NAND U1028 ( .A(n506), .B(n613), .Z(n960) );
  XNOR U1029 ( .A(n958), .B(n980), .Z(n959) );
  AND U1030 ( .A(n548), .B(n573), .Z(n980) );
  XNOR U1031 ( .A(n963), .B(n985), .Z(n966) );
  AND U1032 ( .A(n707), .B(n431), .Z(n985) );
  XOR U1033 ( .A(n986), .B(n987), .Z(n963) );
  ANDN U1034 ( .A(n988), .B(n989), .Z(n987) );
  XNOR U1035 ( .A(n990), .B(n986), .Z(n988) );
  XOR U1036 ( .A(n991), .B(n967), .Z(n984) );
  NAND U1037 ( .A(n636), .B(n483), .Z(n967) );
  IV U1038 ( .A(n969), .Z(n991) );
  XOR U1039 ( .A(n995), .B(n996), .Z(n972) );
  AND U1040 ( .A(n997), .B(n998), .Z(n996) );
  XOR U1041 ( .A(n999), .B(n1000), .Z(n998) );
  XOR U1042 ( .A(n995), .B(n1001), .Z(n1000) );
  XOR U1043 ( .A(n993), .B(n1002), .Z(n997) );
  XOR U1044 ( .A(n995), .B(n994), .Z(n1002) );
  XNOR U1045 ( .A(n1003), .B(n983), .Z(n994) );
  NAND U1046 ( .A(n506), .B(n681), .Z(n983) );
  IV U1047 ( .A(n982), .Z(n1003) );
  XNOR U1048 ( .A(n981), .B(n1004), .Z(n982) );
  AND U1049 ( .A(n613), .B(n573), .Z(n1004) );
  XOR U1050 ( .A(n1005), .B(n1006), .Z(n981) );
  ANDN U1051 ( .A(n1007), .B(n1008), .Z(n1006) );
  XNOR U1052 ( .A(n1009), .B(n1005), .Z(n1007) );
  XNOR U1053 ( .A(n1010), .B(n1011), .Z(n993) );
  IV U1054 ( .A(n989), .Z(n1011) );
  XNOR U1055 ( .A(n986), .B(n1012), .Z(n989) );
  AND U1056 ( .A(n483), .B(n707), .Z(n1012) );
  XOR U1057 ( .A(n1013), .B(n1014), .Z(n986) );
  ANDN U1058 ( .A(n1015), .B(n1016), .Z(n1014) );
  XNOR U1059 ( .A(n1017), .B(n1013), .Z(n1015) );
  XOR U1060 ( .A(n1018), .B(n990), .Z(n1010) );
  NAND U1061 ( .A(n636), .B(n548), .Z(n990) );
  IV U1062 ( .A(n992), .Z(n1018) );
  XOR U1063 ( .A(n1022), .B(n1023), .Z(n995) );
  AND U1064 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U1065 ( .A(n1026), .B(n1027), .Z(n1025) );
  XOR U1066 ( .A(n1022), .B(n1028), .Z(n1027) );
  XOR U1067 ( .A(n1020), .B(n1029), .Z(n1024) );
  XOR U1068 ( .A(n1022), .B(n1021), .Z(n1029) );
  XNOR U1069 ( .A(n1030), .B(n1009), .Z(n1021) );
  NANDN U1070 ( .B(n749), .A(n506), .Z(n1009) );
  IV U1071 ( .A(n1008), .Z(n1030) );
  XNOR U1072 ( .A(n1005), .B(n1031), .Z(n1008) );
  AND U1073 ( .A(n681), .B(n573), .Z(n1031) );
  XOR U1074 ( .A(n1032), .B(n1033), .Z(n1005) );
  ANDN U1075 ( .A(n1034), .B(n1035), .Z(n1033) );
  XNOR U1076 ( .A(n1036), .B(n1032), .Z(n1034) );
  XNOR U1077 ( .A(n1037), .B(n1038), .Z(n1020) );
  IV U1078 ( .A(n1016), .Z(n1038) );
  XNOR U1079 ( .A(n1013), .B(n1039), .Z(n1016) );
  AND U1080 ( .A(n548), .B(n707), .Z(n1039) );
  XOR U1081 ( .A(n1040), .B(n1041), .Z(n1013) );
  ANDN U1082 ( .A(n1042), .B(n1043), .Z(n1041) );
  XNOR U1083 ( .A(n1044), .B(n1040), .Z(n1042) );
  XOR U1084 ( .A(n1045), .B(n1017), .Z(n1037) );
  NAND U1085 ( .A(n636), .B(n613), .Z(n1017) );
  IV U1086 ( .A(n1019), .Z(n1045) );
  XOR U1087 ( .A(n1049), .B(n1050), .Z(n1022) );
  AND U1088 ( .A(n1051), .B(n1052), .Z(n1050) );
  XOR U1089 ( .A(n1053), .B(n1054), .Z(n1052) );
  XOR U1090 ( .A(n1049), .B(n1055), .Z(n1054) );
  XOR U1091 ( .A(n1047), .B(n1056), .Z(n1051) );
  XOR U1092 ( .A(n1049), .B(n1048), .Z(n1056) );
  XNOR U1093 ( .A(n1057), .B(n1036), .Z(n1048) );
  NANDN U1094 ( .B(n826), .A(n506), .Z(n1036) );
  IV U1095 ( .A(n1035), .Z(n1057) );
  XNOR U1096 ( .A(n1032), .B(n1058), .Z(n1035) );
  ANDN U1097 ( .A(n573), .B(n749), .Z(n1058) );
  XOR U1098 ( .A(n1059), .B(n1060), .Z(n1032) );
  ANDN U1099 ( .A(n1061), .B(n1062), .Z(n1060) );
  XNOR U1100 ( .A(n1063), .B(n1059), .Z(n1061) );
  XNOR U1101 ( .A(n1064), .B(n1065), .Z(n1047) );
  IV U1102 ( .A(n1043), .Z(n1065) );
  XNOR U1103 ( .A(n1040), .B(n1066), .Z(n1043) );
  AND U1104 ( .A(n613), .B(n707), .Z(n1066) );
  XOR U1105 ( .A(n1067), .B(n1068), .Z(n1040) );
  ANDN U1106 ( .A(n1069), .B(n1070), .Z(n1068) );
  XNOR U1107 ( .A(n1071), .B(n1067), .Z(n1069) );
  XOR U1108 ( .A(n1072), .B(n1044), .Z(n1064) );
  NAND U1109 ( .A(n636), .B(n681), .Z(n1044) );
  IV U1110 ( .A(n1046), .Z(n1072) );
  XOR U1111 ( .A(n1076), .B(n1077), .Z(n1049) );
  AND U1112 ( .A(n1078), .B(n1079), .Z(n1077) );
  XOR U1113 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR U1114 ( .A(n1076), .B(n1082), .Z(n1081) );
  XOR U1115 ( .A(n1074), .B(n1083), .Z(n1078) );
  XOR U1116 ( .A(n1076), .B(n1075), .Z(n1083) );
  XNOR U1117 ( .A(n1084), .B(n1063), .Z(n1075) );
  NAND U1118 ( .A(n506), .B(n899), .Z(n1063) );
  IV U1119 ( .A(n1062), .Z(n1084) );
  XNOR U1120 ( .A(n1059), .B(n1085), .Z(n1062) );
  ANDN U1121 ( .A(n573), .B(n826), .Z(n1085) );
  XOR U1122 ( .A(n1086), .B(n1087), .Z(n1059) );
  ANDN U1123 ( .A(n1088), .B(n1089), .Z(n1087) );
  XNOR U1124 ( .A(n1090), .B(n1086), .Z(n1088) );
  XNOR U1125 ( .A(n1091), .B(n1092), .Z(n1074) );
  IV U1126 ( .A(n1070), .Z(n1092) );
  XNOR U1127 ( .A(n1067), .B(n1093), .Z(n1070) );
  AND U1128 ( .A(n681), .B(n707), .Z(n1093) );
  XOR U1129 ( .A(n1094), .B(n1095), .Z(n1067) );
  ANDN U1130 ( .A(n1096), .B(n1097), .Z(n1095) );
  XNOR U1131 ( .A(n1098), .B(n1094), .Z(n1096) );
  XOR U1132 ( .A(n1099), .B(n1071), .Z(n1091) );
  NANDN U1133 ( .B(n749), .A(n636), .Z(n1071) );
  IV U1134 ( .A(n1073), .Z(n1099) );
  XOR U1135 ( .A(n1104), .B(n1105), .Z(n920) );
  XNOR U1136 ( .A(n1106), .B(n1103), .Z(n1104) );
  XNOR U1137 ( .A(n1094), .B(n1108), .Z(n1097) );
  ANDN U1138 ( .A(n707), .B(n749), .Z(n1108) );
  XOR U1139 ( .A(n1111), .B(n1109), .Z(n1110) );
  ANDN U1140 ( .A(n707), .B(n826), .Z(n1111) );
  AND U1141 ( .A(n899), .B(n636), .Z(n1112) );
  XOR U1142 ( .A(n1113), .B(n1114), .Z(n1109) );
  ANDN U1143 ( .A(n1115), .B(n1116), .Z(n1114) );
  XNOR U1144 ( .A(n1117), .B(n1113), .Z(n1115) );
  XOR U1145 ( .A(n1118), .B(n1098), .Z(n1107) );
  NANDN U1146 ( .B(n826), .A(n636), .Z(n1098) );
  IV U1147 ( .A(n1100), .Z(n1118) );
  NAND U1148 ( .A(n636), .B(n1119), .Z(n1117) );
  XNOR U1149 ( .A(n1113), .B(n1120), .Z(n1116) );
  AND U1150 ( .A(n899), .B(n707), .Z(n1120) );
  AND U1151 ( .A(n1121), .B(g_input[0]), .Z(n1113) );
  NANDN U1152 ( .B(n636), .A(n1122), .Z(n1121) );
  NAND U1153 ( .A(n1119), .B(n707), .Z(n1122) );
  XNOR U1154 ( .A(n1089), .B(n1090), .Z(n1102) );
  NAND U1155 ( .A(n506), .B(n1119), .Z(n1090) );
  XNOR U1156 ( .A(n1086), .B(n1125), .Z(n1089) );
  AND U1157 ( .A(n899), .B(n573), .Z(n1125) );
  AND U1158 ( .A(n1126), .B(g_input[0]), .Z(n1086) );
  NANDN U1159 ( .B(n506), .A(n1127), .Z(n1126) );
  NAND U1160 ( .A(n1119), .B(n573), .Z(n1127) );
  XOR U1161 ( .A(n1130), .B(n1131), .Z(n1103) );
  XOR U1162 ( .A(n1132), .B(n1133), .Z(n871) );
  AND U1163 ( .A(n1134), .B(n1135), .Z(n1133) );
  NANDN U1164 ( .B(n194), .A(n1136), .Z(n1135) );
  NANDN U1165 ( .B(n1137), .A(n1138), .Z(n194) );
  AND U1166 ( .A(n1139), .B(g_input[15]), .Z(n1138) );
  OR U1167 ( .A(n1140), .B(n1141), .Z(n1134) );
  IV U1168 ( .A(n870), .Z(n1132) );
  NAND U1169 ( .A(n292), .B(n792), .Z(n925) );
  XNOR U1170 ( .A(n923), .B(n1143), .Z(n924) );
  AND U1171 ( .A(n863), .B(n255), .Z(n1143) );
  XOR U1172 ( .A(n1151), .B(n1140), .Z(n1147) );
  NAND U1173 ( .A(n220), .B(n1136), .Z(n1140) );
  IV U1174 ( .A(n1142), .Z(n1151) );
  NAND U1175 ( .A(n337), .B(n792), .Z(n1146) );
  XNOR U1176 ( .A(n1144), .B(n1153), .Z(n1145) );
  AND U1177 ( .A(n863), .B(n292), .Z(n1153) );
  XNOR U1178 ( .A(n1148), .B(n1158), .Z(n1149) );
  AND U1179 ( .A(n220), .B(e_input[0]), .Z(n1158) );
  XNOR U1180 ( .A(n1139), .B(g_input[14]), .Z(n1137) );
  NOR U1181 ( .A(n1159), .B(n1160), .Z(n1139) );
  XOR U1182 ( .A(n1164), .B(n1150), .Z(n1157) );
  NAND U1183 ( .A(n255), .B(n1136), .Z(n1150) );
  IV U1184 ( .A(n1152), .Z(n1164) );
  NAND U1185 ( .A(n382), .B(n792), .Z(n1156) );
  XNOR U1186 ( .A(n1154), .B(n1166), .Z(n1155) );
  AND U1187 ( .A(n863), .B(n337), .Z(n1166) );
  XOR U1188 ( .A(n1167), .B(n1168), .Z(n1154) );
  ANDN U1189 ( .A(n1169), .B(n1170), .Z(n1168) );
  XNOR U1190 ( .A(n1171), .B(n1167), .Z(n1169) );
  XNOR U1191 ( .A(n1161), .B(n1173), .Z(n1162) );
  AND U1192 ( .A(n255), .B(e_input[0]), .Z(n1173) );
  XOR U1193 ( .A(n1159), .B(g_input[13]), .Z(n1160) );
  NANDN U1194 ( .B(n1174), .A(n1175), .Z(n1159) );
  XOR U1195 ( .A(n1179), .B(n1163), .Z(n1172) );
  NAND U1196 ( .A(n292), .B(n1136), .Z(n1163) );
  IV U1197 ( .A(n1165), .Z(n1179) );
  XNOR U1198 ( .A(n1181), .B(n1171), .Z(n999) );
  NAND U1199 ( .A(n431), .B(n792), .Z(n1171) );
  IV U1200 ( .A(n1170), .Z(n1181) );
  XNOR U1201 ( .A(n1167), .B(n1182), .Z(n1170) );
  AND U1202 ( .A(n863), .B(n382), .Z(n1182) );
  XOR U1203 ( .A(n1183), .B(n1184), .Z(n1167) );
  ANDN U1204 ( .A(n1185), .B(n1186), .Z(n1184) );
  XNOR U1205 ( .A(n1187), .B(n1183), .Z(n1185) );
  XNOR U1206 ( .A(n1188), .B(n1189), .Z(n1001) );
  IV U1207 ( .A(n1177), .Z(n1189) );
  XNOR U1208 ( .A(n1176), .B(n1190), .Z(n1177) );
  AND U1209 ( .A(n292), .B(e_input[0]), .Z(n1190) );
  XNOR U1210 ( .A(n1175), .B(g_input[12]), .Z(n1174) );
  NOR U1211 ( .A(n1191), .B(n1192), .Z(n1175) );
  XOR U1212 ( .A(n1193), .B(n1194), .Z(n1176) );
  ANDN U1213 ( .A(n1195), .B(n1196), .Z(n1194) );
  XNOR U1214 ( .A(n1197), .B(n1193), .Z(n1195) );
  XOR U1215 ( .A(n1198), .B(n1178), .Z(n1188) );
  NAND U1216 ( .A(n337), .B(n1136), .Z(n1178) );
  IV U1217 ( .A(n1180), .Z(n1198) );
  XNOR U1218 ( .A(n1200), .B(n1187), .Z(n1026) );
  NAND U1219 ( .A(n483), .B(n792), .Z(n1187) );
  IV U1220 ( .A(n1186), .Z(n1200) );
  XNOR U1221 ( .A(n1183), .B(n1201), .Z(n1186) );
  AND U1222 ( .A(n863), .B(n431), .Z(n1201) );
  XOR U1223 ( .A(n1202), .B(n1203), .Z(n1183) );
  ANDN U1224 ( .A(n1204), .B(n1205), .Z(n1203) );
  XNOR U1225 ( .A(n1206), .B(n1202), .Z(n1204) );
  XNOR U1226 ( .A(n1207), .B(n1208), .Z(n1028) );
  IV U1227 ( .A(n1196), .Z(n1208) );
  XNOR U1228 ( .A(n1193), .B(n1209), .Z(n1196) );
  AND U1229 ( .A(n337), .B(e_input[0]), .Z(n1209) );
  XOR U1230 ( .A(n1191), .B(g_input[11]), .Z(n1192) );
  NANDN U1231 ( .B(n1210), .A(n1211), .Z(n1191) );
  XOR U1232 ( .A(n1212), .B(n1213), .Z(n1193) );
  ANDN U1233 ( .A(n1214), .B(n1215), .Z(n1213) );
  XNOR U1234 ( .A(n1216), .B(n1212), .Z(n1214) );
  XOR U1235 ( .A(n1217), .B(n1197), .Z(n1207) );
  NAND U1236 ( .A(n382), .B(n1136), .Z(n1197) );
  IV U1237 ( .A(n1199), .Z(n1217) );
  XNOR U1238 ( .A(n1219), .B(n1206), .Z(n1053) );
  NAND U1239 ( .A(n548), .B(n792), .Z(n1206) );
  IV U1240 ( .A(n1205), .Z(n1219) );
  XNOR U1241 ( .A(n1202), .B(n1220), .Z(n1205) );
  AND U1242 ( .A(n863), .B(n483), .Z(n1220) );
  XOR U1243 ( .A(n1221), .B(n1222), .Z(n1202) );
  ANDN U1244 ( .A(n1223), .B(n1224), .Z(n1222) );
  XNOR U1245 ( .A(n1225), .B(n1221), .Z(n1223) );
  XNOR U1246 ( .A(n1226), .B(n1227), .Z(n1055) );
  IV U1247 ( .A(n1215), .Z(n1227) );
  XNOR U1248 ( .A(n1212), .B(n1228), .Z(n1215) );
  AND U1249 ( .A(n382), .B(e_input[0]), .Z(n1228) );
  XNOR U1250 ( .A(n1211), .B(g_input[10]), .Z(n1210) );
  NOR U1251 ( .A(n1229), .B(n1230), .Z(n1211) );
  XOR U1252 ( .A(n1231), .B(n1232), .Z(n1212) );
  ANDN U1253 ( .A(n1233), .B(n1234), .Z(n1232) );
  XNOR U1254 ( .A(n1235), .B(n1231), .Z(n1233) );
  XOR U1255 ( .A(n1236), .B(n1216), .Z(n1226) );
  NAND U1256 ( .A(n431), .B(n1136), .Z(n1216) );
  IV U1257 ( .A(n1218), .Z(n1236) );
  XNOR U1258 ( .A(n1238), .B(n1225), .Z(n1080) );
  NAND U1259 ( .A(n613), .B(n792), .Z(n1225) );
  IV U1260 ( .A(n1224), .Z(n1238) );
  XNOR U1261 ( .A(n1221), .B(n1239), .Z(n1224) );
  AND U1262 ( .A(n863), .B(n548), .Z(n1239) );
  XOR U1263 ( .A(n1240), .B(n1241), .Z(n1221) );
  ANDN U1264 ( .A(n1242), .B(n1243), .Z(n1241) );
  XNOR U1265 ( .A(n1244), .B(n1240), .Z(n1242) );
  XNOR U1266 ( .A(n1245), .B(n1246), .Z(n1082) );
  IV U1267 ( .A(n1234), .Z(n1246) );
  XNOR U1268 ( .A(n1231), .B(n1247), .Z(n1234) );
  AND U1269 ( .A(n431), .B(e_input[0]), .Z(n1247) );
  XOR U1270 ( .A(n1229), .B(g_input[9]), .Z(n1230) );
  NANDN U1271 ( .B(n1248), .A(n1249), .Z(n1229) );
  XOR U1272 ( .A(n1250), .B(n1251), .Z(n1231) );
  ANDN U1273 ( .A(n1252), .B(n1253), .Z(n1251) );
  XNOR U1274 ( .A(n1254), .B(n1250), .Z(n1252) );
  XOR U1275 ( .A(n1255), .B(n1235), .Z(n1245) );
  NAND U1276 ( .A(n483), .B(n1136), .Z(n1235) );
  IV U1277 ( .A(n1237), .Z(n1255) );
  NAND U1278 ( .A(n681), .B(n792), .Z(n1244) );
  XNOR U1279 ( .A(n1240), .B(n1257), .Z(n1243) );
  AND U1280 ( .A(n863), .B(n613), .Z(n1257) );
  XNOR U1281 ( .A(n1261), .B(n1258), .Z(n1260) );
  XNOR U1282 ( .A(n1250), .B(n1263), .Z(n1253) );
  AND U1283 ( .A(n483), .B(e_input[0]), .Z(n1263) );
  XNOR U1284 ( .A(n1267), .B(n1264), .Z(n1266) );
  XOR U1285 ( .A(n1268), .B(n1254), .Z(n1262) );
  NAND U1286 ( .A(n548), .B(n1136), .Z(n1254) );
  IV U1287 ( .A(n1256), .Z(n1268) );
  XNOR U1288 ( .A(n1269), .B(n1270), .Z(n1256) );
  AND U1289 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U1290 ( .A(n1265), .B(n1273), .Z(n1272) );
  XNOR U1291 ( .A(n1267), .B(n1269), .Z(n1273) );
  NAND U1292 ( .A(n613), .B(n1136), .Z(n1267) );
  XOR U1293 ( .A(n1264), .B(n1274), .Z(n1265) );
  AND U1294 ( .A(n548), .B(e_input[0]), .Z(n1274) );
  XNOR U1295 ( .A(n1278), .B(n1275), .Z(n1277) );
  XOR U1296 ( .A(n1259), .B(n1279), .Z(n1271) );
  XNOR U1297 ( .A(n1261), .B(n1269), .Z(n1279) );
  NANDN U1298 ( .B(n749), .A(n792), .Z(n1261) );
  XOR U1299 ( .A(n1258), .B(n1280), .Z(n1259) );
  AND U1300 ( .A(n863), .B(n681), .Z(n1280) );
  XOR U1301 ( .A(n1281), .B(n1282), .Z(n1258) );
  AND U1302 ( .A(n1283), .B(n1284), .Z(n1282) );
  XNOR U1303 ( .A(n1285), .B(n1281), .Z(n1284) );
  XOR U1304 ( .A(n1286), .B(n1287), .Z(n1269) );
  AND U1305 ( .A(n1288), .B(n1289), .Z(n1287) );
  XOR U1306 ( .A(n1276), .B(n1290), .Z(n1289) );
  XNOR U1307 ( .A(n1278), .B(n1286), .Z(n1290) );
  NAND U1308 ( .A(n681), .B(n1136), .Z(n1278) );
  XOR U1309 ( .A(n1275), .B(n1291), .Z(n1276) );
  AND U1310 ( .A(n613), .B(e_input[0]), .Z(n1291) );
  XNOR U1311 ( .A(n1295), .B(n1292), .Z(n1294) );
  XOR U1312 ( .A(n1283), .B(n1296), .Z(n1288) );
  XNOR U1313 ( .A(n1285), .B(n1286), .Z(n1296) );
  NANDN U1314 ( .B(n826), .A(n792), .Z(n1285) );
  XOR U1315 ( .A(n1281), .B(n1297), .Z(n1283) );
  ANDN U1316 ( .A(n863), .B(n749), .Z(n1297) );
  XOR U1317 ( .A(n1298), .B(n1299), .Z(n1281) );
  AND U1318 ( .A(n1300), .B(n1301), .Z(n1299) );
  XNOR U1319 ( .A(n1302), .B(n1298), .Z(n1301) );
  XOR U1320 ( .A(n1303), .B(n1304), .Z(n1286) );
  AND U1321 ( .A(n1305), .B(n1306), .Z(n1304) );
  XOR U1322 ( .A(n1293), .B(n1307), .Z(n1306) );
  XNOR U1323 ( .A(n1295), .B(n1303), .Z(n1307) );
  NANDN U1324 ( .B(n749), .A(n1136), .Z(n1295) );
  XOR U1325 ( .A(n1292), .B(n1308), .Z(n1293) );
  AND U1326 ( .A(n681), .B(e_input[0]), .Z(n1308) );
  XOR U1327 ( .A(n1300), .B(n1312), .Z(n1305) );
  XNOR U1328 ( .A(n1302), .B(n1303), .Z(n1312) );
  NAND U1329 ( .A(n792), .B(n899), .Z(n1302) );
  XOR U1330 ( .A(n1298), .B(n1313), .Z(n1300) );
  ANDN U1331 ( .A(n863), .B(n826), .Z(n1313) );
  NAND U1332 ( .A(n792), .B(n1119), .Z(n1316) );
  XNOR U1333 ( .A(n1314), .B(n1318), .Z(n1315) );
  AND U1334 ( .A(n899), .B(n863), .Z(n1318) );
  AND U1335 ( .A(n1319), .B(g_input[0]), .Z(n1314) );
  NANDN U1336 ( .B(n792), .A(n1320), .Z(n1319) );
  NAND U1337 ( .A(n1119), .B(n863), .Z(n1320) );
  XNOR U1338 ( .A(n1309), .B(n1324), .Z(n1310) );
  ANDN U1339 ( .A(e_input[0]), .B(n749), .Z(n1324) );
  XOR U1340 ( .A(n1327), .B(n1325), .Z(n1326) );
  ANDN U1341 ( .A(e_input[0]), .B(n826), .Z(n1327) );
  AND U1342 ( .A(n1136), .B(n899), .Z(n1328) );
  XOR U1343 ( .A(n1332), .B(n1311), .Z(n1323) );
  NANDN U1344 ( .B(n826), .A(n1136), .Z(n1311) );
  IV U1345 ( .A(n1317), .Z(n1332) );
  NAND U1346 ( .A(n1136), .B(n1119), .Z(n1331) );
  XNOR U1347 ( .A(n1329), .B(n1333), .Z(n1330) );
  AND U1348 ( .A(n899), .B(e_input[0]), .Z(n1333) );
  AND U1349 ( .A(n1334), .B(g_input[0]), .Z(n1329) );
  NANDN U1350 ( .B(n1136), .A(n1335), .Z(n1334) );
  NAND U1351 ( .A(n1119), .B(e_input[0]), .Z(n1335) );
  XNOR U1352 ( .A(n1337), .B(n889), .Z(n879) );
  XNOR U1353 ( .A(n876), .B(n877), .Z(n889) );
  NAND U1354 ( .A(n320), .B(n681), .Z(n877) );
  XNOR U1355 ( .A(n875), .B(n1338), .Z(n876) );
  AND U1356 ( .A(n613), .B(n361), .Z(n1338) );
  XNOR U1357 ( .A(n1342), .B(n1339), .Z(n1341) );
  XNOR U1358 ( .A(n888), .B(n878), .Z(n1337) );
  XOR U1359 ( .A(n1343), .B(n1344), .Z(n878) );
  XNOR U1360 ( .A(n883), .B(n1346), .Z(n884) );
  AND U1361 ( .A(n483), .B(n468), .Z(n1346) );
  XNOR U1362 ( .A(n1249), .B(g_input[8]), .Z(n1248) );
  NOR U1363 ( .A(n1347), .B(n1348), .Z(n1249) );
  XOR U1364 ( .A(n1349), .B(n1350), .Z(n883) );
  AND U1365 ( .A(n1351), .B(n1352), .Z(n1350) );
  XNOR U1366 ( .A(n1353), .B(n1349), .Z(n1352) );
  XOR U1367 ( .A(n1354), .B(n885), .Z(n1345) );
  NAND U1368 ( .A(n414), .B(n548), .Z(n885) );
  IV U1369 ( .A(n887), .Z(n1354) );
  XNOR U1370 ( .A(n1355), .B(n1356), .Z(n887) );
  AND U1371 ( .A(n1357), .B(n1358), .Z(n1356) );
  XOR U1372 ( .A(n1351), .B(n1359), .Z(n1358) );
  XNOR U1373 ( .A(n1353), .B(n1355), .Z(n1359) );
  NAND U1374 ( .A(n414), .B(n613), .Z(n1353) );
  XOR U1375 ( .A(n1349), .B(n1360), .Z(n1351) );
  AND U1376 ( .A(n548), .B(n468), .Z(n1360) );
  XOR U1377 ( .A(n1347), .B(g_input[7]), .Z(n1348) );
  NANDN U1378 ( .B(n1361), .A(n1362), .Z(n1347) );
  XOR U1379 ( .A(n1363), .B(n1364), .Z(n1349) );
  AND U1380 ( .A(n1365), .B(n1366), .Z(n1364) );
  XNOR U1381 ( .A(n1367), .B(n1363), .Z(n1366) );
  XOR U1382 ( .A(n1340), .B(n1368), .Z(n1357) );
  XNOR U1383 ( .A(n1342), .B(n1355), .Z(n1368) );
  NANDN U1384 ( .B(n749), .A(n320), .Z(n1342) );
  XOR U1385 ( .A(n1339), .B(n1369), .Z(n1340) );
  AND U1386 ( .A(n681), .B(n361), .Z(n1369) );
  XNOR U1387 ( .A(n1373), .B(n1370), .Z(n1372) );
  XOR U1388 ( .A(n1374), .B(n1375), .Z(n1355) );
  AND U1389 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR U1390 ( .A(n1365), .B(n1378), .Z(n1377) );
  XNOR U1391 ( .A(n1367), .B(n1374), .Z(n1378) );
  NAND U1392 ( .A(n414), .B(n681), .Z(n1367) );
  XOR U1393 ( .A(n1363), .B(n1379), .Z(n1365) );
  AND U1394 ( .A(n613), .B(n468), .Z(n1379) );
  XNOR U1395 ( .A(n1362), .B(g_input[6]), .Z(n1361) );
  NOR U1396 ( .A(n1380), .B(n1381), .Z(n1362) );
  XOR U1397 ( .A(n1382), .B(n1383), .Z(n1363) );
  AND U1398 ( .A(n1384), .B(n1385), .Z(n1383) );
  XNOR U1399 ( .A(n1386), .B(n1382), .Z(n1385) );
  XOR U1400 ( .A(n1371), .B(n1387), .Z(n1376) );
  XNOR U1401 ( .A(n1373), .B(n1374), .Z(n1387) );
  NANDN U1402 ( .B(n826), .A(n320), .Z(n1373) );
  XOR U1403 ( .A(n1370), .B(n1388), .Z(n1371) );
  ANDN U1404 ( .A(n361), .B(n749), .Z(n1388) );
  XNOR U1405 ( .A(n1392), .B(n1389), .Z(n1391) );
  XOR U1406 ( .A(n1393), .B(n1394), .Z(n1374) );
  AND U1407 ( .A(n1395), .B(n1396), .Z(n1394) );
  XOR U1408 ( .A(n1384), .B(n1397), .Z(n1396) );
  XNOR U1409 ( .A(n1386), .B(n1393), .Z(n1397) );
  NANDN U1410 ( .B(n749), .A(n414), .Z(n1386) );
  XOR U1411 ( .A(n1382), .B(n1398), .Z(n1384) );
  AND U1412 ( .A(n681), .B(n468), .Z(n1398) );
  XOR U1413 ( .A(n1380), .B(g_input[5]), .Z(n1381) );
  NANDN U1414 ( .B(n1399), .A(n1400), .Z(n1380) );
  XOR U1415 ( .A(n1401), .B(n1402), .Z(n1382) );
  ANDN U1416 ( .A(n1403), .B(n1404), .Z(n1402) );
  XNOR U1417 ( .A(n1405), .B(n1401), .Z(n1403) );
  XOR U1418 ( .A(n1390), .B(n1406), .Z(n1395) );
  XNOR U1419 ( .A(n1392), .B(n1393), .Z(n1406) );
  NAND U1420 ( .A(n320), .B(n899), .Z(n1392) );
  XOR U1421 ( .A(n1389), .B(n1407), .Z(n1390) );
  ANDN U1422 ( .A(n361), .B(n826), .Z(n1407) );
  XOR U1423 ( .A(n1408), .B(n1409), .Z(n1389) );
  ANDN U1424 ( .A(n1410), .B(n1411), .Z(n1409) );
  XNOR U1425 ( .A(n1412), .B(n1408), .Z(n1410) );
  NAND U1426 ( .A(n320), .B(n1119), .Z(n1412) );
  XNOR U1427 ( .A(n1408), .B(n1414), .Z(n1411) );
  AND U1428 ( .A(n899), .B(n361), .Z(n1414) );
  AND U1429 ( .A(n1415), .B(g_input[0]), .Z(n1408) );
  NANDN U1430 ( .B(n320), .A(n1416), .Z(n1415) );
  NAND U1431 ( .A(n1119), .B(n361), .Z(n1416) );
  XNOR U1432 ( .A(n1401), .B(n1420), .Z(n1404) );
  ANDN U1433 ( .A(n468), .B(n749), .Z(n1420) );
  XOR U1434 ( .A(n1421), .B(n1422), .Z(n1401) );
  AND U1435 ( .A(n1423), .B(n1424), .Z(n1422) );
  XOR U1436 ( .A(n1425), .B(n1421), .Z(n1424) );
  ANDN U1437 ( .A(n468), .B(n826), .Z(n1425) );
  XOR U1438 ( .A(n1426), .B(n1421), .Z(n1423) );
  AND U1439 ( .A(n899), .B(n414), .Z(n1426) );
  XOR U1440 ( .A(n1427), .B(n1428), .Z(n1421) );
  ANDN U1441 ( .A(n1429), .B(n1430), .Z(n1428) );
  XNOR U1442 ( .A(n1431), .B(n1427), .Z(n1429) );
  XOR U1443 ( .A(n1432), .B(n1405), .Z(n1419) );
  NANDN U1444 ( .B(n826), .A(n414), .Z(n1405) );
  IV U1445 ( .A(n1413), .Z(n1432) );
  XOR U1446 ( .A(n1433), .B(n1431), .Z(n1413) );
  NAND U1447 ( .A(n414), .B(n1119), .Z(n1431) );
  IV U1448 ( .A(n1430), .Z(n1433) );
  XNOR U1449 ( .A(n1427), .B(n1434), .Z(n1430) );
  AND U1450 ( .A(n899), .B(n468), .Z(n1434) );
  AND U1451 ( .A(n1435), .B(g_input[0]), .Z(n1427) );
  NANDN U1452 ( .B(n414), .A(n1436), .Z(n1435) );
  NAND U1453 ( .A(n1119), .B(n468), .Z(n1436) );
  XNOR U1454 ( .A(n892), .B(n1440), .Z(n893) );
  ANDN U1455 ( .A(n288), .B(n749), .Z(n1440) );
  XNOR U1456 ( .A(n1400), .B(g_input[4]), .Z(n1399) );
  NOR U1457 ( .A(n1441), .B(n1442), .Z(n1400) );
  XOR U1458 ( .A(n1443), .B(n1444), .Z(n892) );
  AND U1459 ( .A(n1445), .B(n1446), .Z(n1444) );
  XOR U1460 ( .A(n1447), .B(n1443), .Z(n1446) );
  ANDN U1461 ( .A(n288), .B(n826), .Z(n1447) );
  XOR U1462 ( .A(n1448), .B(n1443), .Z(n1445) );
  AND U1463 ( .A(n899), .B(n250), .Z(n1448) );
  XOR U1464 ( .A(n1449), .B(n1450), .Z(n1443) );
  ANDN U1465 ( .A(n1451), .B(n1452), .Z(n1450) );
  XNOR U1466 ( .A(n1453), .B(n1449), .Z(n1451) );
  XOR U1467 ( .A(n1454), .B(n894), .Z(n1439) );
  NANDN U1468 ( .B(n826), .A(n250), .Z(n894) );
  NANDN U1469 ( .B(n1455), .A(n1456), .Z(n1441) );
  IV U1470 ( .A(n896), .Z(n1454) );
  NAND U1471 ( .A(n250), .B(n1119), .Z(n1453) );
  XNOR U1472 ( .A(n1449), .B(n1457), .Z(n1452) );
  AND U1473 ( .A(n899), .B(n288), .Z(n1457) );
  AND U1474 ( .A(n1458), .B(g_input[0]), .Z(n1449) );
  NANDN U1475 ( .B(n250), .A(n1459), .Z(n1458) );
  NAND U1476 ( .A(n1119), .B(n288), .Z(n1459) );
  XNOR U1477 ( .A(n1460), .B(e_input[12]), .Z(n288) );
  NAND U1478 ( .A(n1461), .B(e_input[15]), .Z(n1460) );
  XOR U1479 ( .A(n1462), .B(e_input[12]), .Z(n1461) );
  XNOR U1480 ( .A(n903), .B(n904), .Z(n898) );
  NANDN U1481 ( .B(n195), .A(n1119), .Z(n904) );
  XNOR U1482 ( .A(n902), .B(n1464), .Z(n903) );
  AND U1483 ( .A(n899), .B(n219), .Z(n1464) );
  XNOR U1484 ( .A(n1456), .B(g_input[2]), .Z(n1455) );
  AND U1485 ( .A(n1466), .B(g_input[0]), .Z(n902) );
  NAND U1486 ( .A(n1467), .B(n195), .Z(n1466) );
  NANDN U1487 ( .B(n1468), .A(n1469), .Z(n195) );
  ANDN U1488 ( .A(e_input[15]), .B(n1470), .Z(n1469) );
  NAND U1489 ( .A(n1119), .B(n219), .Z(n1467) );
  XOR U1490 ( .A(n1470), .B(e_input[14]), .Z(n1468) );
  OR U1491 ( .A(n1463), .B(n1471), .Z(n1470) );
  XOR U1492 ( .A(n1471), .B(e_input[13]), .Z(n1463) );
  OR U1493 ( .A(n1462), .B(n1472), .Z(n1471) );
  XOR U1494 ( .A(n1472), .B(e_input[12]), .Z(n1462) );
  OR U1495 ( .A(n1418), .B(n1473), .Z(n1472) );
  XOR U1496 ( .A(n1473), .B(e_input[11]), .Z(n1418) );
  OR U1497 ( .A(n1417), .B(n1474), .Z(n1473) );
  XOR U1498 ( .A(n1474), .B(e_input[10]), .Z(n1417) );
  OR U1499 ( .A(n1438), .B(n1475), .Z(n1474) );
  XOR U1500 ( .A(n1475), .B(e_input[9]), .Z(n1438) );
  OR U1501 ( .A(n1437), .B(n1476), .Z(n1475) );
  XOR U1502 ( .A(n1476), .B(e_input[8]), .Z(n1437) );
  OR U1503 ( .A(n1129), .B(n1477), .Z(n1476) );
  XOR U1504 ( .A(n1477), .B(e_input[7]), .Z(n1129) );
  OR U1505 ( .A(n1128), .B(n1478), .Z(n1477) );
  XOR U1506 ( .A(n1478), .B(e_input[6]), .Z(n1128) );
  OR U1507 ( .A(n1124), .B(n1479), .Z(n1478) );
  XOR U1508 ( .A(n1479), .B(e_input[5]), .Z(n1124) );
  OR U1509 ( .A(n1123), .B(n1480), .Z(n1479) );
  XOR U1510 ( .A(n1480), .B(e_input[4]), .Z(n1123) );
  OR U1511 ( .A(n1322), .B(n1481), .Z(n1480) );
  XOR U1512 ( .A(n1481), .B(e_input[3]), .Z(n1322) );
  OR U1513 ( .A(n1321), .B(n1482), .Z(n1481) );
  XOR U1514 ( .A(n1482), .B(e_input[2]), .Z(n1321) );
  NANDN U1515 ( .B(e_input[0]), .A(n1336), .Z(n1482) );
  XNOR U1516 ( .A(e_input[0]), .B(e_input[1]), .Z(n1336) );
  XOR U1517 ( .A(g_input[0]), .B(g_input[1]), .Z(n1465) );
  NANDN U1518 ( .B(n838), .A(n110), .Z(n162) );
  IV U1519 ( .A(rst), .Z(n110) );
  NAND U1520 ( .A(n1483), .B(n1484), .Z(n838) );
  ANDN U1521 ( .A(n1485), .B(\_MxM/n[2] ), .Z(n1484) );
  NOR U1522 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n1485) );
  ANDN U1523 ( .A(n1486), .B(n104), .Z(n1483) );
  OR U1524 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n104) );
  NOR U1525 ( .A(\_MxM/n[0] ), .B(\_MxM/n[1] ), .Z(n1486) );
endmodule

