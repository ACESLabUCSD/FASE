
module MxM_W16_N100 ( clk, rst, A, X, Y );
  input [15:0] A;
  input [15:0] X;
  output [15:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229,
         \add_25/carry[6] , \add_25/carry[5] , \add_25/carry[4] ,
         \add_25/carry[3] , \add_25/carry[2] , n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715;
  wire   [15:0] Y0;
  wire   [6:0] n;

  DFF \n_reg[0]  ( .D(n229), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n228), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n227), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n226), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n225), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n224), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n223), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \Y0_reg[0]  ( .D(n222), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n221), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n220), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n219), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n218), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n217), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n216), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n215), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y0_reg[8]  ( .D(n214), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[8]) );
  DFF \Y0_reg[9]  ( .D(n213), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[9]) );
  DFF \Y0_reg[10]  ( .D(n212), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[10]) );
  DFF \Y0_reg[11]  ( .D(n211), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[11]) );
  DFF \Y0_reg[12]  ( .D(n210), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[12]) );
  DFF \Y0_reg[13]  ( .D(n209), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[13]) );
  DFF \Y0_reg[14]  ( .D(n208), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[14]) );
  DFF \Y0_reg[15]  ( .D(n207), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[15]) );
  DFF \Y_reg[15]  ( .D(n206), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[15]) );
  DFF \Y_reg[14]  ( .D(n205), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[14]) );
  DFF \Y_reg[13]  ( .D(n204), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[13]) );
  DFF \Y_reg[12]  ( .D(n203), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[12]) );
  DFF \Y_reg[11]  ( .D(n202), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[11]) );
  DFF \Y_reg[10]  ( .D(n201), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[10]) );
  DFF \Y_reg[9]  ( .D(n200), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[9]) );
  DFF \Y_reg[8]  ( .D(n199), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[8]) );
  DFF \Y_reg[7]  ( .D(n198), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n197), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n196), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n195), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n194), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n193), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n192), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n191), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  MUX U232 ( .IN0(n230), .IN1(n1543), .SEL(n1544), .F(n1527) );
  IV U233 ( .A(n1545), .Z(n230) );
  MUX U234 ( .IN0(n231), .IN1(n1210), .SEL(n1211), .F(n1187) );
  IV U235 ( .A(n1212), .Z(n231) );
  MUX U236 ( .IN0(n1618), .IN1(n1636), .SEL(n1620), .F(n1599) );
  XOR U237 ( .A(n1401), .B(n1391), .Z(n1207) );
  XOR U238 ( .A(n1213), .B(n1195), .Z(n1199) );
  MUX U239 ( .IN0(n232), .IN1(n960), .SEL(n961), .F(n890) );
  IV U240 ( .A(n962), .Z(n232) );
  MUX U241 ( .IN0(n233), .IN1(n1121), .SEL(n1122), .F(n1046) );
  IV U242 ( .A(n1123), .Z(n233) );
  MUX U243 ( .IN0(n234), .IN1(n1187), .SEL(n1188), .F(n1164) );
  IV U244 ( .A(n1189), .Z(n234) );
  MUX U245 ( .IN0(n235), .IN1(n1383), .SEL(n1384), .F(n1373) );
  IV U246 ( .A(n1385), .Z(n235) );
  XOR U247 ( .A(n1386), .B(n1378), .Z(n1184) );
  MUX U248 ( .IN0(n1338), .IN1(n1341), .SEL(n1339), .F(n1323) );
  MUX U249 ( .IN0(n236), .IN1(n685), .SEL(n686), .F(n634) );
  IV U250 ( .A(n687), .Z(n236) );
  MUX U251 ( .IN0(n237), .IN1(n1037), .SEL(n1038), .F(n960) );
  IV U252 ( .A(n1039), .Z(n237) );
  XNOR U253 ( .A(n1681), .B(n1682), .Z(n1125) );
  XOR U254 ( .A(n1188), .B(n1189), .Z(n1200) );
  MUX U255 ( .IN0(n238), .IN1(n1137), .SEL(n1138), .F(n1075) );
  IV U256 ( .A(n1139), .Z(n238) );
  XOR U257 ( .A(n1374), .B(n1375), .Z(n1182) );
  MUX U258 ( .IN0(n239), .IN1(n814), .SEL(n815), .F(n749) );
  IV U259 ( .A(n816), .Z(n239) );
  MUX U260 ( .IN0(X[8]), .IN1(n1666), .SEL(X[15]), .F(n697) );
  MUX U261 ( .IN0(n1379), .IN1(n240), .SEL(n1378), .F(n1370) );
  IV U262 ( .A(n1377), .Z(n240) );
  MUX U263 ( .IN0(X[13]), .IN1(n1692), .SEL(X[15]), .F(n479) );
  MUX U264 ( .IN0(n1554), .IN1(n1557), .SEL(n1555), .F(n1538) );
  MUX U265 ( .IN0(n241), .IN1(n1164), .SEL(n1165), .F(n1145) );
  IV U266 ( .A(n1166), .Z(n241) );
  MUX U267 ( .IN0(n242), .IN1(n1373), .SEL(n1374), .F(n1152) );
  IV U268 ( .A(n1375), .Z(n242) );
  XOR U269 ( .A(n1190), .B(n1172), .Z(n1176) );
  MUX U270 ( .IN0(X[9]), .IN1(n1667), .SEL(X[15]), .F(n643) );
  MUX U271 ( .IN0(n520), .IN1(n243), .SEL(n519), .F(n481) );
  IV U272 ( .A(n518), .Z(n243) );
  MUX U273 ( .IN0(X[11]), .IN1(n1647), .SEL(X[15]), .F(n549) );
  MUX U274 ( .IN0(n610), .IN1(n608), .SEL(n609), .F(n563) );
  MUX U275 ( .IN0(n244), .IN1(n403), .SEL(n402), .F(n411) );
  IV U276 ( .A(n414), .Z(n244) );
  MUX U277 ( .IN0(n245), .IN1(n1558), .SEL(n1559), .F(n1554) );
  IV U278 ( .A(n1560), .Z(n245) );
  XOR U279 ( .A(n1384), .B(n1385), .Z(n1205) );
  MUX U280 ( .IN0(n246), .IN1(n941), .SEL(n942), .F(n872) );
  IV U281 ( .A(n943), .Z(n246) );
  MUX U282 ( .IN0(n247), .IN1(n1000), .SEL(n1001), .F(n937) );
  IV U283 ( .A(n1002), .Z(n247) );
  MUX U284 ( .IN0(X[10]), .IN1(n1646), .SEL(X[15]), .F(n590) );
  MUX U285 ( .IN0(n700), .IN1(n248), .SEL(n699), .F(n645) );
  IV U286 ( .A(n698), .Z(n248) );
  MUX U287 ( .IN0(n776), .IN1(n774), .SEL(n775), .F(n709) );
  XNOR U288 ( .A(n1668), .B(n1122), .Z(n1126) );
  XOR U289 ( .A(n412), .B(n433), .Z(n431) );
  MUX U290 ( .IN0(n1599), .IN1(n1617), .SEL(n1601), .F(n1568) );
  MUX U291 ( .IN0(n1487), .IN1(n1509), .SEL(n1489), .F(n1469) );
  MUX U292 ( .IN0(n249), .IN1(n1145), .SEL(n1146), .F(n1083) );
  IV U293 ( .A(n1147), .Z(n249) );
  MUX U294 ( .IN0(n250), .IN1(n1390), .SEL(n1391), .F(n1377) );
  IV U295 ( .A(n1392), .Z(n250) );
  MUX U296 ( .IN0(n251), .IN1(n1112), .SEL(n1113), .F(n1037) );
  IV U297 ( .A(n1114), .Z(n251) );
  MUX U298 ( .IN0(A[11]), .IN1(n1421), .SEL(A[15]), .F(n566) );
  MUX U299 ( .IN0(n648), .IN1(n256), .SEL(n647), .F(n597) );
  MUX U300 ( .IN0(n909), .IN1(n907), .SEL(n908), .F(n839) );
  MUX U301 ( .IN0(n939), .IN1(n252), .SEL(n938), .F(n867) );
  IV U302 ( .A(n937), .Z(n252) );
  NAND U303 ( .A(n481), .B(n516), .Z(n515) );
  XOR U304 ( .A(n459), .B(n467), .Z(n465) );
  MUX U305 ( .IN0(n253), .IN1(n1405), .SEL(n1406), .F(n1390) );
  IV U306 ( .A(n1407), .Z(n253) );
  MUX U307 ( .IN0(n254), .IN1(n952), .SEL(n953), .F(n882) );
  IV U308 ( .A(n954), .Z(n254) );
  MUX U309 ( .IN0(n255), .IN1(n1008), .SEL(n1009), .F(n941) );
  IV U310 ( .A(n1010), .Z(n255) );
  MUX U311 ( .IN0(X[4]), .IN1(n1352), .SEL(X[15]), .F(n936) );
  XOR U312 ( .A(n1648), .B(n1633), .Z(n1573) );
  MUX U313 ( .IN0(n692), .IN1(n694), .SEL(n693), .F(n256) );
  IV U314 ( .A(n256), .Z(n646) );
  MUX U315 ( .IN0(n870), .IN1(n257), .SEL(n869), .F(n797) );
  IV U316 ( .A(n868), .Z(n257) );
  MUX U317 ( .IN0(n977), .IN1(n975), .SEL(n976), .F(n907) );
  MUX U318 ( .IN0(n1095), .IN1(n258), .SEL(n1094), .F(n1018) );
  IV U319 ( .A(n1093), .Z(n258) );
  XNOR U320 ( .A(n600), .B(n560), .Z(n564) );
  XOR U321 ( .A(n490), .B(n498), .Z(n496) );
  XOR U322 ( .A(n1165), .B(n1166), .Z(n1177) );
  MUX U323 ( .IN0(n1493), .IN1(n1503), .SEL(n1495), .F(n1479) );
  MUX U324 ( .IN0(n1568), .IN1(n1598), .SEL(n1570), .F(n1104) );
  XNOR U325 ( .A(n1345), .B(n1346), .Z(n1329) );
  MUX U326 ( .IN0(A[9]), .IN1(n1459), .SEL(A[15]), .F(n660) );
  MUX U327 ( .IN0(A[12]), .IN1(n1403), .SEL(A[15]), .F(n521) );
  XOR U328 ( .A(n569), .B(n612), .Z(n570) );
  MUX U329 ( .IN0(n964), .IN1(n966), .SEL(n965), .F(n896) );
  MUX U330 ( .IN0(n1006), .IN1(n1004), .SEL(n1005), .F(n931) );
  XOR U331 ( .A(n1094), .B(n1095), .Z(n1101) );
  XNOR U332 ( .A(n597), .B(n640), .Z(n598) );
  XNOR U333 ( .A(n701), .B(n654), .Z(n658) );
  MUX U334 ( .IN0(n259), .IN1(n885), .SEL(n886), .F(n817) );
  IV U335 ( .A(n887), .Z(n259) );
  MUX U336 ( .IN0(n744), .IN1(n746), .SEL(n745), .F(n260) );
  IV U337 ( .A(n260), .Z(n680) );
  XOR U338 ( .A(n527), .B(n535), .Z(n533) );
  MUX U339 ( .IN0(n1485), .IN1(n261), .SEL(n1335), .F(n1466) );
  IV U340 ( .A(n1334), .Z(n261) );
  MUX U341 ( .IN0(n1331), .IN1(n1329), .SEL(n1330), .F(n1302) );
  XOR U342 ( .A(n1376), .B(n1370), .Z(n1161) );
  MUX U343 ( .IN0(n262), .IN1(n1104), .SEL(n1105), .F(n1029) );
  IV U344 ( .A(n1106), .Z(n262) );
  MUX U345 ( .IN0(n263), .IN1(n1152), .SEL(n1153), .F(n1093) );
  IV U346 ( .A(n1154), .Z(n263) );
  XOR U347 ( .A(n1167), .B(n1138), .Z(n1142) );
  MUX U348 ( .IN0(n828), .IN1(n830), .SEL(n829), .F(n763) );
  MUX U349 ( .IN0(n1054), .IN1(n1052), .SEL(n1053), .F(n975) );
  XOR U350 ( .A(n1574), .B(n1113), .Z(n1117) );
  XNOR U351 ( .A(n649), .B(n605), .Z(n609) );
  MUX U352 ( .IN0(n264), .IN1(n688), .SEL(n689), .F(n637) );
  IV U353 ( .A(n690), .Z(n264) );
  MUX U354 ( .IN0(n265), .IN1(n803), .SEL(n804), .F(n743) );
  IV U355 ( .A(n805), .Z(n265) );
  NAND U356 ( .A(n867), .B(n935), .Z(n934) );
  MUX U357 ( .IN0(n809), .IN1(n811), .SEL(n810), .F(n744) );
  MUX U358 ( .IN0(n266), .IN1(n783), .SEL(n784), .F(n718) );
  IV U359 ( .A(Y0[5]), .Z(n266) );
  XOR U360 ( .A(n572), .B(n580), .Z(n578) );
  MUX U361 ( .IN0(n267), .IN1(n1538), .SEL(n1539), .F(n1521) );
  IV U362 ( .A(n1540), .Z(n267) );
  MUX U363 ( .IN0(A[1]), .IN1(n1694), .SEL(A[15]), .F(n1348) );
  MUX U364 ( .IN0(n268), .IN1(n749), .SEL(n750), .F(n685) );
  IV U365 ( .A(n751), .Z(n268) );
  MUX U366 ( .IN0(A[6]), .IN1(n1590), .SEL(A[15]), .F(n842) );
  MUX U367 ( .IN0(A[7]), .IN1(n1577), .SEL(A[15]), .F(n777) );
  MUX U368 ( .IN0(A[5]), .IN1(n1610), .SEL(A[15]), .F(n910) );
  MUX U369 ( .IN0(n269), .IN1(n1083), .SEL(n1084), .F(n1008) );
  IV U370 ( .A(n1085), .Z(n269) );
  XOR U371 ( .A(n1153), .B(n1154), .Z(n1159) );
  MUX U372 ( .IN0(n896), .IN1(n898), .SEL(n897), .F(n828) );
  XNOR U373 ( .A(n1135), .B(n1076), .Z(n1080) );
  XOR U374 ( .A(n487), .B(n522), .Z(n488) );
  MUX U375 ( .IN0(n270), .IN1(n552), .SEL(n553), .F(n505) );
  IV U376 ( .A(n554), .Z(n270) );
  NAND U377 ( .A(n645), .B(n696), .Z(n695) );
  MUX U378 ( .IN0(n799), .IN1(n797), .SEL(n798), .F(n741) );
  XNOR U379 ( .A(n831), .B(n771), .Z(n775) );
  MUX U380 ( .IN0(n271), .IN1(n1032), .SEL(n1033), .F(n955) );
  IV U381 ( .A(n1034), .Z(n271) );
  MUX U382 ( .IN0(n272), .IN1(n879), .SEL(n878), .F(n809) );
  IV U383 ( .A(n877), .Z(n272) );
  MUX U384 ( .IN0(n273), .IN1(n848), .SEL(n849), .F(n783) );
  IV U385 ( .A(Y0[4]), .Z(n273) );
  XOR U386 ( .A(n617), .B(n625), .Z(n623) );
  MUX U387 ( .IN0(n1302), .IN1(n274), .SEL(n1303), .F(n1275) );
  IV U388 ( .A(n1304), .Z(n274) );
  MUX U389 ( .IN0(n1394), .IN1(n275), .SEL(n1207), .F(n1381) );
  IV U390 ( .A(n1205), .Z(n275) );
  XNOR U391 ( .A(n1559), .B(n1560), .Z(n1546) );
  MUX U392 ( .IN0(n276), .IN1(n882), .SEL(n883), .F(n814) );
  IV U393 ( .A(n884), .Z(n276) );
  MUX U394 ( .IN0(A[3]), .IN1(n1671), .SEL(A[15]), .F(n277) );
  IV U395 ( .A(n277), .Z(n1055) );
  MUX U396 ( .IN0(A[4]), .IN1(n1628), .SEL(A[15]), .F(n278) );
  IV U397 ( .A(n278), .Z(n978) );
  MUX U398 ( .IN0(n1141), .IN1(n279), .SEL(n1142), .F(n1079) );
  IV U399 ( .A(n1143), .Z(n279) );
  XOR U400 ( .A(n1472), .B(n1473), .Z(n1334) );
  MUX U401 ( .IN0(n565), .IN1(n563), .SEL(n564), .F(n510) );
  MUX U402 ( .IN0(n280), .IN1(n872), .SEL(n873), .F(n803) );
  IV U403 ( .A(n874), .Z(n280) );
  XOR U404 ( .A(n780), .B(n843), .Z(n781) );
  MUX U405 ( .IN0(n1041), .IN1(n1043), .SEL(n1042), .F(n964) );
  MUX U406 ( .IN0(n1127), .IN1(n1125), .SEL(n1126), .F(n1052) );
  MUX U407 ( .IN0(n281), .IN1(n594), .SEL(n595), .F(n552) );
  IV U408 ( .A(n596), .Z(n281) );
  XOR U409 ( .A(n755), .B(n699), .Z(n693) );
  XNOR U410 ( .A(n766), .B(n706), .Z(n710) );
  MUX U411 ( .IN0(n282), .IN1(n817), .SEL(n818), .F(n752) );
  IV U412 ( .A(n819), .Z(n282) );
  XOR U413 ( .A(n930), .B(n868), .Z(n869) );
  MUX U414 ( .IN0(n1026), .IN1(n283), .SEL(n1025), .F(n947) );
  IV U415 ( .A(n1024), .Z(n283) );
  MUX U416 ( .IN0(n944), .IN1(n284), .SEL(n945), .F(n877) );
  IV U417 ( .A(n946), .Z(n284) );
  MUX U418 ( .IN0(n285), .IN1(n916), .SEL(n917), .F(n848) );
  IV U419 ( .A(Y0[3]), .Z(n285) );
  XOR U420 ( .A(n672), .B(n678), .Z(n667) );
  MUX U421 ( .IN0(n286), .IN1(n1332), .SEL(n1149), .F(n1305) );
  IV U422 ( .A(n1148), .Z(n286) );
  MUX U423 ( .IN0(n1248), .IN1(n287), .SEL(n1249), .F(n1221) );
  IV U424 ( .A(n1250), .Z(n287) );
  MUX U425 ( .IN0(X[1]), .IN1(n288), .SEL(X[15]), .F(n1365) );
  IV U426 ( .A(n1565), .Z(n288) );
  MUX U427 ( .IN0(X[6]), .IN1(n1357), .SEL(X[15]), .F(n802) );
  MUX U428 ( .IN0(X[3]), .IN1(n1551), .SEL(X[15]), .F(n1021) );
  MUX U429 ( .IN0(n1116), .IN1(n1118), .SEL(n1117), .F(n1041) );
  MUX U430 ( .IN0(X[14]), .IN1(n1697), .SEL(X[15]), .F(n448) );
  NAND U431 ( .A(n546), .B(n589), .Z(n588) );
  XOR U432 ( .A(n820), .B(n760), .Z(n764) );
  XNOR U433 ( .A(n899), .B(n836), .Z(n840) );
  MUX U434 ( .IN0(n289), .IN1(n955), .SEL(n956), .F(n885) );
  IV U435 ( .A(n957), .Z(n289) );
  XNOR U436 ( .A(n998), .B(n938), .Z(n932) );
  MUX U437 ( .IN0(n1011), .IN1(n290), .SEL(n1012), .F(n944) );
  IV U438 ( .A(n1013), .Z(n290) );
  MUX U439 ( .IN0(n291), .IN1(n490), .SEL(n491), .F(n459) );
  IV U440 ( .A(Y0[11]), .Z(n291) );
  XOR U441 ( .A(n718), .B(n726), .Z(n724) );
  MUX U442 ( .IN0(n1466), .IN1(n292), .SEL(n1311), .F(n1447) );
  IV U443 ( .A(n1309), .Z(n292) );
  MUX U444 ( .IN0(n1521), .IN1(n1537), .SEL(n1523), .F(n1504) );
  MUX U445 ( .IN0(n1198), .IN1(n293), .SEL(n1199), .F(n1175) );
  IV U446 ( .A(n1200), .Z(n293) );
  XOR U447 ( .A(n1146), .B(n1147), .Z(n1143) );
  XOR U448 ( .A(n1544), .B(n1545), .Z(n1359) );
  MUX U449 ( .IN0(n294), .IN1(n1029), .SEL(n1030), .F(n952) );
  IV U450 ( .A(n1031), .Z(n294) );
  MUX U451 ( .IN0(A[10]), .IN1(n1439), .SEL(A[15]), .F(n611) );
  XNOR U452 ( .A(n1336), .B(n1326), .Z(n1330) );
  XOR U453 ( .A(n663), .B(n713), .Z(n664) );
  MUX U454 ( .IN0(n711), .IN1(n709), .SEL(n710), .F(n657) );
  MUX U455 ( .IN0(n933), .IN1(n931), .SEL(n932), .F(n868) );
  MUX U456 ( .IN0(A[13]), .IN1(n1389), .SEL(A[15]), .F(n484) );
  MUX U457 ( .IN0(n295), .IN1(n752), .SEL(n753), .F(n688) );
  IV U458 ( .A(n754), .Z(n295) );
  XOR U459 ( .A(n888), .B(n825), .Z(n829) );
  XNOR U460 ( .A(n1044), .B(n972), .Z(n976) );
  MUX U461 ( .IN0(n296), .IN1(n1107), .SEL(n1108), .F(n1032) );
  IV U462 ( .A(n1109), .Z(n296) );
  MUX U463 ( .IN0(n297), .IN1(n1096), .SEL(n1097), .F(n1024) );
  IV U464 ( .A(n1098), .Z(n297) );
  MUX U465 ( .IN0(A[14]), .IN1(n1366), .SEL(A[15]), .F(n449) );
  MUX U466 ( .IN0(n507), .IN1(n298), .SEL(n506), .F(n475) );
  IV U467 ( .A(n505), .Z(n298) );
  XNOR U468 ( .A(n809), .B(n808), .Z(n861) );
  MUX U469 ( .IN0(Y0[13]), .IN1(n299), .SEL(n413), .F(n405) );
  IV U470 ( .A(n412), .Z(n299) );
  MUX U471 ( .IN0(n300), .IN1(n572), .SEL(n573), .F(n527) );
  IV U472 ( .A(Y0[9]), .Z(n300) );
  MUX U473 ( .IN0(n301), .IN1(n1061), .SEL(n1062), .F(n984) );
  IV U474 ( .A(Y0[1]), .Z(n301) );
  XOR U475 ( .A(n783), .B(n791), .Z(n789) );
  MUX U476 ( .IN0(n1447), .IN1(n302), .SEL(n1284), .F(n1428) );
  IV U477 ( .A(n1282), .Z(n302) );
  MUX U478 ( .IN0(n1221), .IN1(n303), .SEL(n1222), .F(n1198) );
  IV U479 ( .A(n1223), .Z(n303) );
  MUX U480 ( .IN0(n1504), .IN1(n1520), .SEL(n1506), .F(n1493) );
  MUX U481 ( .IN0(n1381), .IN1(n304), .SEL(n1184), .F(n1371) );
  IV U482 ( .A(n1182), .Z(n304) );
  MUX U483 ( .IN0(A[8]), .IN1(n1477), .SEL(A[15]), .F(n712) );
  MUX U484 ( .IN0(A[2]), .IN1(n1684), .SEL(A[15]), .F(n1128) );
  MUX U485 ( .IN0(n305), .IN1(n1075), .SEL(n1076), .F(n1000) );
  IV U486 ( .A(n1077), .Z(n305) );
  MUX U487 ( .IN0(n306), .IN1(n634), .SEL(n635), .F(n591) );
  IV U488 ( .A(n636), .Z(n306) );
  MUX U489 ( .IN0(n763), .IN1(n765), .SEL(n764), .F(n692) );
  MUX U490 ( .IN0(n841), .IN1(n839), .SEL(n840), .F(n774) );
  XOR U491 ( .A(n1058), .B(n1129), .Z(n1059) );
  MUX U492 ( .IN0(n1081), .IN1(n1079), .SEL(n1080), .F(n1004) );
  XNOR U493 ( .A(n510), .B(n511), .Z(n509) );
  MUX U494 ( .IN0(n307), .IN1(n637), .SEL(n638), .F(n594) );
  IV U495 ( .A(n639), .Z(n307) );
  XOR U496 ( .A(n804), .B(n805), .Z(n799) );
  XOR U497 ( .A(n1035), .B(n961), .Z(n965) );
  XNOR U498 ( .A(n1119), .B(n1049), .Z(n1053) );
  NAND U499 ( .A(n1018), .B(n1091), .Z(n1090) );
  XNOR U500 ( .A(n514), .B(n513), .Z(n507) );
  XNOR U501 ( .A(n909), .B(n908), .Z(n887) );
  MUX U502 ( .IN0(n949), .IN1(n947), .SEL(n948), .F(n308) );
  IV U503 ( .A(n308), .Z(n876) );
  MUX U504 ( .IN0(n1086), .IN1(n309), .SEL(n1087), .F(n1011) );
  IV U505 ( .A(n1088), .Z(n309) );
  MUX U506 ( .IN0(n680), .IN1(n310), .SEL(n681), .F(n631) );
  IV U507 ( .A(n682), .Z(n310) );
  MUX U508 ( .IN0(n311), .IN1(n459), .SEL(n460), .F(n412) );
  IV U509 ( .A(Y0[12]), .Z(n311) );
  MUX U510 ( .IN0(n312), .IN1(n617), .SEL(n618), .F(n572) );
  IV U511 ( .A(Y0[8]), .Z(n312) );
  XOR U512 ( .A(n848), .B(n856), .Z(n854) );
  MUX U513 ( .IN0(n1428), .IN1(n313), .SEL(n1257), .F(n1409) );
  IV U514 ( .A(n1255), .Z(n313) );
  MUX U515 ( .IN0(n314), .IN1(n1572), .SEL(n1573), .F(n1622) );
  IV U516 ( .A(n1642), .Z(n314) );
  NOR U517 ( .A(A[0]), .B(n1694), .Z(n1685) );
  XOR U518 ( .A(n1552), .B(n1539), .Z(n1360) );
  MUX U519 ( .IN0(n1371), .IN1(n315), .SEL(n1161), .F(n1099) );
  IV U520 ( .A(n1159), .Z(n315) );
  MUX U521 ( .IN0(n659), .IN1(n657), .SEL(n658), .F(n608) );
  XOR U522 ( .A(n913), .B(n979), .Z(n914) );
  MUX U523 ( .IN0(n593), .IN1(n316), .SEL(n592), .F(n546) );
  IV U524 ( .A(n591), .Z(n316) );
  MUX U525 ( .IN0(X[7]), .IN1(n1358), .SEL(X[15]), .F(n735) );
  XNOR U526 ( .A(n967), .B(n904), .Z(n908) );
  XOR U527 ( .A(n958), .B(n893), .Z(n897) );
  XNOR U528 ( .A(n1073), .B(n1001), .Z(n1005) );
  XNOR U529 ( .A(n1127), .B(n1126), .Z(n1109) );
  MUX U530 ( .IN0(n483), .IN1(n509), .SEL(n482), .F(n454) );
  XNOR U531 ( .A(n565), .B(n564), .Z(n554) );
  XNOR U532 ( .A(n776), .B(n775), .Z(n754) );
  XNOR U533 ( .A(n841), .B(n840), .Z(n819) );
  XNOR U534 ( .A(n947), .B(n1014), .Z(n948) );
  XNOR U535 ( .A(n690), .B(n689), .Z(n682) );
  XOR U536 ( .A(n796), .B(n737), .Z(n745) );
  XNOR U537 ( .A(n957), .B(n956), .Z(n946) );
  XNOR U538 ( .A(n1034), .B(n1033), .Z(n1013) );
  XNOR U539 ( .A(n473), .B(n472), .Z(n497) );
  MUX U540 ( .IN0(n317), .IN1(n666), .SEL(n667), .F(n617) );
  IV U541 ( .A(Y0[7]), .Z(n317) );
  MUX U542 ( .IN0(Y0[14]), .IN1(n405), .SEL(n406), .F(n395) );
  XOR U543 ( .A(n916), .B(n924), .Z(n922) );
  MUX U544 ( .IN0(n1275), .IN1(n318), .SEL(n1276), .F(n1248) );
  IV U545 ( .A(n1277), .Z(n318) );
  MUX U546 ( .IN0(n319), .IN1(n1359), .SEL(n1360), .F(n1532) );
  IV U547 ( .A(n1546), .Z(n319) );
  MUX U548 ( .IN0(n1409), .IN1(n320), .SEL(n1230), .F(n1394) );
  IV U549 ( .A(n1228), .Z(n320) );
  XOR U550 ( .A(n1670), .B(A[3]), .Z(n1671) );
  MUX U551 ( .IN0(n1175), .IN1(n321), .SEL(n1176), .F(n1141) );
  IV U552 ( .A(n1177), .Z(n321) );
  XOR U553 ( .A(n1640), .B(n1641), .Z(n1572) );
  XOR U554 ( .A(n1491), .B(n1482), .Z(n1335) );
  MUX U555 ( .IN0(X[5]), .IN1(n1353), .SEL(X[15]), .F(n865) );
  MUX U556 ( .IN0(X[2]), .IN1(n1550), .SEL(X[15]), .F(n1092) );
  XNOR U557 ( .A(n1331), .B(n1330), .Z(n1148) );
  XNOR U558 ( .A(n555), .B(n519), .Z(n513) );
  MUX U559 ( .IN0(n599), .IN1(n597), .SEL(n598), .F(n322) );
  IV U560 ( .A(n322), .Z(n551) );
  XOR U561 ( .A(n873), .B(n874), .Z(n870) );
  XOR U562 ( .A(n1110), .B(n1038), .Z(n1042) );
  MUX U563 ( .IN0(n1101), .IN1(n1361), .SEL(n1100), .F(n1023) );
  XNOR U564 ( .A(n1081), .B(n1080), .Z(n1098) );
  AND U565 ( .A(n443), .B(n420), .Z(n442) );
  XNOR U566 ( .A(n610), .B(n609), .Z(n596) );
  XNOR U567 ( .A(n659), .B(n658), .Z(n639) );
  XNOR U568 ( .A(n711), .B(n710), .Z(n690) );
  XNOR U569 ( .A(n933), .B(n932), .Z(n949) );
  XNOR U570 ( .A(n977), .B(n976), .Z(n957) );
  XNOR U571 ( .A(n1054), .B(n1053), .Z(n1034) );
  XNOR U572 ( .A(n1006), .B(n1005), .Z(n1026) );
  XNOR U573 ( .A(n1109), .B(n1108), .Z(n1088) );
  XNOR U574 ( .A(n474), .B(n475), .Z(n473) );
  XNOR U575 ( .A(n754), .B(n753), .Z(n746) );
  XNOR U576 ( .A(n819), .B(n818), .Z(n811) );
  XNOR U577 ( .A(n887), .B(n886), .Z(n879) );
  MUX U578 ( .IN0(n323), .IN1(n527), .SEL(n528), .F(n490) );
  IV U579 ( .A(Y0[10]), .Z(n323) );
  MUX U580 ( .IN0(n324), .IN1(n718), .SEL(n719), .F(n666) );
  IV U581 ( .A(Y0[6]), .Z(n324) );
  MUX U582 ( .IN0(n325), .IN1(n984), .SEL(n985), .F(n916) );
  IV U583 ( .A(Y0[2]), .Z(n325) );
  MUX U584 ( .IN0(Y0[15]), .IN1(n395), .SEL(n396), .F(n326) );
  IV U585 ( .A(n326), .Z(n392) );
  XOR U586 ( .A(n1062), .B(Y0[1]), .Z(n337) );
  ANDN U587 ( .A(n327), .B(n[0]), .Z(n229) );
  AND U588 ( .A(N8), .B(n327), .Z(n228) );
  AND U589 ( .A(N9), .B(n327), .Z(n227) );
  AND U590 ( .A(N10), .B(n327), .Z(n226) );
  AND U591 ( .A(N11), .B(n327), .Z(n225) );
  AND U592 ( .A(N12), .B(n327), .Z(n224) );
  AND U593 ( .A(n327), .B(n328), .Z(n223) );
  XOR U594 ( .A(n[6]), .B(\add_25/carry[6] ), .Z(n328) );
  ANDN U595 ( .A(n329), .B(rst), .Z(n327) );
  NAND U596 ( .A(n330), .B(n331), .Z(n329) );
  AND U597 ( .A(n[0]), .B(n332), .Z(n331) );
  NOR U598 ( .A(n333), .B(n[2]), .Z(n332) );
  AND U599 ( .A(n334), .B(n[6]), .Z(n330) );
  AND U600 ( .A(n[5]), .B(n[1]), .Z(n334) );
  NAND U601 ( .A(n335), .B(n336), .Z(n222) );
  OR U602 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U603 ( .B(n339), .A(Y0[0]), .Z(n335) );
  NAND U604 ( .A(n340), .B(n341), .Z(n221) );
  NANDN U605 ( .B(n338), .A(n342), .Z(n341) );
  NANDN U606 ( .B(n343), .A(rst), .Z(n340) );
  NAND U607 ( .A(n344), .B(n345), .Z(n220) );
  NANDN U608 ( .B(n338), .A(n346), .Z(n345) );
  NANDN U609 ( .B(n339), .A(Y0[2]), .Z(n344) );
  NAND U610 ( .A(n347), .B(n348), .Z(n219) );
  NANDN U611 ( .B(n338), .A(n349), .Z(n348) );
  NANDN U612 ( .B(n339), .A(Y0[3]), .Z(n347) );
  NAND U613 ( .A(n350), .B(n351), .Z(n218) );
  NANDN U614 ( .B(n338), .A(n352), .Z(n351) );
  NANDN U615 ( .B(n339), .A(Y0[4]), .Z(n350) );
  NAND U616 ( .A(n353), .B(n354), .Z(n217) );
  NANDN U617 ( .B(n338), .A(n355), .Z(n354) );
  NANDN U618 ( .B(n339), .A(Y0[5]), .Z(n353) );
  NAND U619 ( .A(n356), .B(n357), .Z(n216) );
  NANDN U620 ( .B(n338), .A(n358), .Z(n357) );
  NANDN U621 ( .B(n339), .A(Y0[6]), .Z(n356) );
  NAND U622 ( .A(n359), .B(n360), .Z(n215) );
  NANDN U623 ( .B(n338), .A(n361), .Z(n360) );
  NANDN U624 ( .B(n339), .A(Y0[7]), .Z(n359) );
  NAND U625 ( .A(n362), .B(n363), .Z(n214) );
  NANDN U626 ( .B(n338), .A(n364), .Z(n363) );
  NANDN U627 ( .B(n339), .A(Y0[8]), .Z(n362) );
  NAND U628 ( .A(n365), .B(n366), .Z(n213) );
  NANDN U629 ( .B(n338), .A(n367), .Z(n366) );
  NANDN U630 ( .B(n339), .A(Y0[9]), .Z(n365) );
  NAND U631 ( .A(n368), .B(n369), .Z(n212) );
  NANDN U632 ( .B(n338), .A(n370), .Z(n369) );
  NANDN U633 ( .B(n339), .A(Y0[10]), .Z(n368) );
  NAND U634 ( .A(n371), .B(n372), .Z(n211) );
  NANDN U635 ( .B(n338), .A(n373), .Z(n372) );
  NANDN U636 ( .B(n339), .A(Y0[11]), .Z(n371) );
  NAND U637 ( .A(n374), .B(n375), .Z(n210) );
  NANDN U638 ( .B(n338), .A(n376), .Z(n375) );
  NANDN U639 ( .B(n339), .A(Y0[12]), .Z(n374) );
  NAND U640 ( .A(n377), .B(n378), .Z(n209) );
  NANDN U641 ( .B(n338), .A(n379), .Z(n378) );
  NANDN U642 ( .B(n339), .A(Y0[13]), .Z(n377) );
  NAND U643 ( .A(n380), .B(n381), .Z(n208) );
  OR U644 ( .A(n382), .B(n338), .Z(n381) );
  NANDN U645 ( .B(n339), .A(Y0[14]), .Z(n380) );
  NAND U646 ( .A(n383), .B(n384), .Z(n207) );
  OR U647 ( .A(n338), .B(n385), .Z(n384) );
  NANDN U648 ( .B(n386), .A(n339), .Z(n338) );
  NANDN U649 ( .B(n339), .A(Y0[15]), .Z(n383) );
  NAND U650 ( .A(n387), .B(n388), .Z(n206) );
  NANDN U651 ( .B(n339), .A(Y[15]), .Z(n388) );
  AND U652 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U653 ( .B(n386), .A(Y[15]), .Z(n390) );
  OR U654 ( .A(n385), .B(n391), .Z(n389) );
  XOR U655 ( .A(n392), .B(n393), .Z(n385) );
  XNOR U656 ( .A(Y0[15]), .B(n394), .Z(n393) );
  NAND U657 ( .A(n397), .B(n398), .Z(n205) );
  NANDN U658 ( .B(n339), .A(Y[14]), .Z(n398) );
  AND U659 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U660 ( .B(n386), .A(Y[14]), .Z(n400) );
  OR U661 ( .A(n382), .B(n391), .Z(n399) );
  XOR U662 ( .A(n396), .B(Y0[15]), .Z(n382) );
  XOR U663 ( .A(n395), .B(n394), .Z(n396) );
  NAND U664 ( .A(n401), .B(n402), .Z(n394) );
  OR U665 ( .A(n403), .B(n404), .Z(n401) );
  NAND U666 ( .A(n407), .B(n408), .Z(n204) );
  NANDN U667 ( .B(n339), .A(Y[13]), .Z(n408) );
  AND U668 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U669 ( .B(n386), .A(Y[13]), .Z(n410) );
  NANDN U670 ( .B(n391), .A(n379), .Z(n409) );
  XNOR U671 ( .A(n406), .B(Y0[14]), .Z(n379) );
  XNOR U672 ( .A(n411), .B(n405), .Z(n406) );
  XNOR U673 ( .A(n404), .B(n414), .Z(n403) );
  OR U674 ( .A(n415), .B(n416), .Z(n404) );
  AND U675 ( .A(n417), .B(n418), .Z(n414) );
  OR U676 ( .A(n419), .B(n420), .Z(n418) );
  AND U677 ( .A(n421), .B(n422), .Z(n417) );
  OR U678 ( .A(n423), .B(n424), .Z(n422) );
  OR U679 ( .A(n425), .B(n426), .Z(n421) );
  NAND U680 ( .A(n427), .B(n428), .Z(n203) );
  NANDN U681 ( .B(n339), .A(Y[12]), .Z(n428) );
  AND U682 ( .A(n429), .B(n430), .Z(n427) );
  NANDN U683 ( .B(n386), .A(Y[12]), .Z(n430) );
  NANDN U684 ( .B(n391), .A(n376), .Z(n429) );
  XNOR U685 ( .A(n413), .B(Y0[13]), .Z(n376) );
  XNOR U686 ( .A(n431), .B(n432), .Z(n413) );
  AND U687 ( .A(n402), .B(n434), .Z(n433) );
  XOR U688 ( .A(n415), .B(n435), .Z(n434) );
  XOR U689 ( .A(n435), .B(n416), .Z(n415) );
  OR U690 ( .A(n436), .B(n437), .Z(n416) );
  IV U691 ( .A(n432), .Z(n435) );
  XNOR U692 ( .A(n426), .B(n425), .Z(n432) );
  OR U693 ( .A(n438), .B(n439), .Z(n425) );
  AND U694 ( .A(n440), .B(n441), .Z(n426) );
  XNOR U695 ( .A(n419), .B(n442), .Z(n441) );
  NAND U696 ( .A(n444), .B(n445), .Z(n420) );
  NANDN U697 ( .B(n446), .A(n447), .Z(n444) );
  NANDN U698 ( .B(n423), .A(n448), .Z(n443) );
  NANDN U699 ( .B(n424), .A(n449), .Z(n419) );
  AND U700 ( .A(n450), .B(n451), .Z(n440) );
  OR U701 ( .A(n452), .B(n453), .Z(n451) );
  XNOR U702 ( .A(n454), .B(n455), .Z(n450) );
  ANDN U703 ( .A(n456), .B(n457), .Z(n455) );
  XOR U704 ( .A(n454), .B(n458), .Z(n456) );
  NAND U705 ( .A(n461), .B(n462), .Z(n202) );
  NANDN U706 ( .B(n339), .A(Y[11]), .Z(n462) );
  AND U707 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U708 ( .B(n386), .A(Y[11]), .Z(n464) );
  NANDN U709 ( .B(n391), .A(n373), .Z(n463) );
  XNOR U710 ( .A(n460), .B(Y0[12]), .Z(n373) );
  XNOR U711 ( .A(n465), .B(n466), .Z(n460) );
  AND U712 ( .A(n402), .B(n468), .Z(n467) );
  XOR U713 ( .A(n436), .B(n469), .Z(n468) );
  XOR U714 ( .A(n469), .B(n437), .Z(n436) );
  OR U715 ( .A(n470), .B(n471), .Z(n437) );
  IV U716 ( .A(n466), .Z(n469) );
  XNOR U717 ( .A(n439), .B(n438), .Z(n466) );
  OR U718 ( .A(n472), .B(n473), .Z(n438) );
  XNOR U719 ( .A(n453), .B(n452), .Z(n439) );
  OR U720 ( .A(n474), .B(n475), .Z(n452) );
  XOR U721 ( .A(n458), .B(n457), .Z(n453) );
  XOR U722 ( .A(n454), .B(n476), .Z(n457) );
  AND U723 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U724 ( .B(n423), .A(n479), .Z(n478) );
  OR U725 ( .A(n480), .B(n481), .Z(n477) );
  XOR U726 ( .A(n446), .B(n447), .Z(n458) );
  NANDN U727 ( .B(n424), .A(n484), .Z(n447) );
  XNOR U728 ( .A(n445), .B(n485), .Z(n446) );
  AND U729 ( .A(n449), .B(n448), .Z(n485) );
  ANDN U730 ( .A(n486), .B(n487), .Z(n445) );
  NANDN U731 ( .B(n488), .A(n489), .Z(n486) );
  NAND U732 ( .A(n492), .B(n493), .Z(n201) );
  NANDN U733 ( .B(n339), .A(Y[10]), .Z(n493) );
  AND U734 ( .A(n494), .B(n495), .Z(n492) );
  NANDN U735 ( .B(n386), .A(Y[10]), .Z(n495) );
  NANDN U736 ( .B(n391), .A(n370), .Z(n494) );
  XNOR U737 ( .A(n491), .B(Y0[11]), .Z(n370) );
  XNOR U738 ( .A(n496), .B(n497), .Z(n491) );
  AND U739 ( .A(n402), .B(n499), .Z(n498) );
  XOR U740 ( .A(n470), .B(n500), .Z(n499) );
  XOR U741 ( .A(n500), .B(n471), .Z(n470) );
  OR U742 ( .A(n501), .B(n502), .Z(n471) );
  IV U743 ( .A(n497), .Z(n500) );
  OR U744 ( .A(n503), .B(n504), .Z(n472) );
  XOR U745 ( .A(n483), .B(n482), .Z(n474) );
  XNOR U746 ( .A(n508), .B(n509), .Z(n482) );
  ANDN U747 ( .A(n512), .B(n513), .Z(n511) );
  XOR U748 ( .A(n510), .B(n514), .Z(n512) );
  XNOR U749 ( .A(n515), .B(n480), .Z(n508) );
  NAND U750 ( .A(n479), .B(n449), .Z(n480) );
  NANDN U751 ( .B(n423), .A(n517), .Z(n516) );
  XOR U752 ( .A(n488), .B(n489), .Z(n483) );
  NANDN U753 ( .B(n424), .A(n521), .Z(n489) );
  AND U754 ( .A(n484), .B(n448), .Z(n522) );
  NAND U755 ( .A(n523), .B(n524), .Z(n487) );
  NANDN U756 ( .B(n525), .A(n526), .Z(n523) );
  NAND U757 ( .A(n529), .B(n530), .Z(n200) );
  NANDN U758 ( .B(n339), .A(Y[9]), .Z(n530) );
  AND U759 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U760 ( .B(n386), .A(Y[9]), .Z(n532) );
  NANDN U761 ( .B(n391), .A(n367), .Z(n531) );
  XNOR U762 ( .A(n528), .B(Y0[10]), .Z(n367) );
  XNOR U763 ( .A(n533), .B(n534), .Z(n528) );
  AND U764 ( .A(n402), .B(n536), .Z(n535) );
  XOR U765 ( .A(n501), .B(n537), .Z(n536) );
  XOR U766 ( .A(n537), .B(n502), .Z(n501) );
  OR U767 ( .A(n538), .B(n539), .Z(n502) );
  IV U768 ( .A(n534), .Z(n537) );
  XNOR U769 ( .A(n504), .B(n503), .Z(n534) );
  OR U770 ( .A(n540), .B(n541), .Z(n503) );
  XNOR U771 ( .A(n507), .B(n506), .Z(n504) );
  XOR U772 ( .A(n505), .B(n542), .Z(n506) );
  AND U773 ( .A(n543), .B(n544), .Z(n542) );
  OR U774 ( .A(n545), .B(n546), .Z(n544) );
  AND U775 ( .A(n547), .B(n548), .Z(n543) );
  NANDN U776 ( .B(n423), .A(n549), .Z(n548) );
  NAND U777 ( .A(n550), .B(n551), .Z(n547) );
  XNOR U778 ( .A(n518), .B(n556), .Z(n519) );
  AND U779 ( .A(n449), .B(n517), .Z(n556) );
  XOR U780 ( .A(n557), .B(n558), .Z(n518) );
  ANDN U781 ( .A(n559), .B(n560), .Z(n558) );
  XNOR U782 ( .A(n561), .B(n557), .Z(n559) );
  XOR U783 ( .A(n562), .B(n520), .Z(n555) );
  NAND U784 ( .A(n479), .B(n484), .Z(n520) );
  IV U785 ( .A(n510), .Z(n562) );
  XNOR U786 ( .A(n525), .B(n526), .Z(n514) );
  NANDN U787 ( .B(n424), .A(n566), .Z(n526) );
  XNOR U788 ( .A(n524), .B(n567), .Z(n525) );
  AND U789 ( .A(n521), .B(n448), .Z(n567) );
  ANDN U790 ( .A(n568), .B(n569), .Z(n524) );
  NANDN U791 ( .B(n570), .A(n571), .Z(n568) );
  NAND U792 ( .A(n574), .B(n575), .Z(n199) );
  NANDN U793 ( .B(n339), .A(Y[8]), .Z(n575) );
  AND U794 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U795 ( .B(n386), .A(Y[8]), .Z(n577) );
  NANDN U796 ( .B(n391), .A(n364), .Z(n576) );
  XNOR U797 ( .A(n573), .B(Y0[9]), .Z(n364) );
  XNOR U798 ( .A(n578), .B(n579), .Z(n573) );
  AND U799 ( .A(n402), .B(n581), .Z(n580) );
  XOR U800 ( .A(n538), .B(n582), .Z(n581) );
  XOR U801 ( .A(n582), .B(n539), .Z(n538) );
  OR U802 ( .A(n583), .B(n584), .Z(n539) );
  IV U803 ( .A(n579), .Z(n582) );
  XNOR U804 ( .A(n541), .B(n540), .Z(n579) );
  OR U805 ( .A(n585), .B(n586), .Z(n540) );
  XNOR U806 ( .A(n554), .B(n553), .Z(n541) );
  XOR U807 ( .A(n587), .B(n550), .Z(n553) );
  XNOR U808 ( .A(n588), .B(n545), .Z(n550) );
  NAND U809 ( .A(n549), .B(n449), .Z(n545) );
  NANDN U810 ( .B(n423), .A(n590), .Z(n589) );
  XNOR U811 ( .A(n551), .B(n552), .Z(n587) );
  XNOR U812 ( .A(n557), .B(n601), .Z(n560) );
  AND U813 ( .A(n484), .B(n517), .Z(n601) );
  XOR U814 ( .A(n602), .B(n603), .Z(n557) );
  ANDN U815 ( .A(n604), .B(n605), .Z(n603) );
  XNOR U816 ( .A(n606), .B(n602), .Z(n604) );
  XOR U817 ( .A(n607), .B(n561), .Z(n600) );
  NAND U818 ( .A(n479), .B(n521), .Z(n561) );
  IV U819 ( .A(n563), .Z(n607) );
  XNOR U820 ( .A(n570), .B(n571), .Z(n565) );
  NANDN U821 ( .B(n424), .A(n611), .Z(n571) );
  AND U822 ( .A(n566), .B(n448), .Z(n612) );
  NAND U823 ( .A(n613), .B(n614), .Z(n569) );
  NANDN U824 ( .B(n615), .A(n616), .Z(n613) );
  NAND U825 ( .A(n619), .B(n620), .Z(n198) );
  NANDN U826 ( .B(n339), .A(Y[7]), .Z(n620) );
  AND U827 ( .A(n621), .B(n622), .Z(n619) );
  NANDN U828 ( .B(n386), .A(Y[7]), .Z(n622) );
  NANDN U829 ( .B(n391), .A(n361), .Z(n621) );
  XNOR U830 ( .A(n618), .B(Y0[8]), .Z(n361) );
  XNOR U831 ( .A(n623), .B(n624), .Z(n618) );
  AND U832 ( .A(n402), .B(n626), .Z(n625) );
  XOR U833 ( .A(n583), .B(n627), .Z(n626) );
  XOR U834 ( .A(n627), .B(n584), .Z(n583) );
  OR U835 ( .A(n628), .B(n629), .Z(n584) );
  IV U836 ( .A(n624), .Z(n627) );
  XNOR U837 ( .A(n586), .B(n585), .Z(n624) );
  NANDN U838 ( .B(n630), .A(n631), .Z(n585) );
  XNOR U839 ( .A(n596), .B(n595), .Z(n586) );
  XOR U840 ( .A(n632), .B(n599), .Z(n595) );
  XNOR U841 ( .A(n592), .B(n593), .Z(n599) );
  NAND U842 ( .A(n549), .B(n484), .Z(n593) );
  XNOR U843 ( .A(n591), .B(n633), .Z(n592) );
  AND U844 ( .A(n449), .B(n590), .Z(n633) );
  XNOR U845 ( .A(n598), .B(n594), .Z(n632) );
  AND U846 ( .A(n641), .B(n642), .Z(n640) );
  NANDN U847 ( .B(n423), .A(n643), .Z(n642) );
  OR U848 ( .A(n644), .B(n645), .Z(n641) );
  XNOR U849 ( .A(n602), .B(n650), .Z(n605) );
  AND U850 ( .A(n521), .B(n517), .Z(n650) );
  XOR U851 ( .A(n651), .B(n652), .Z(n602) );
  ANDN U852 ( .A(n653), .B(n654), .Z(n652) );
  XNOR U853 ( .A(n655), .B(n651), .Z(n653) );
  XOR U854 ( .A(n656), .B(n606), .Z(n649) );
  NAND U855 ( .A(n479), .B(n566), .Z(n606) );
  IV U856 ( .A(n608), .Z(n656) );
  XNOR U857 ( .A(n615), .B(n616), .Z(n610) );
  NANDN U858 ( .B(n424), .A(n660), .Z(n616) );
  XNOR U859 ( .A(n614), .B(n661), .Z(n615) );
  AND U860 ( .A(n611), .B(n448), .Z(n661) );
  ANDN U861 ( .A(n662), .B(n663), .Z(n614) );
  NANDN U862 ( .B(n664), .A(n665), .Z(n662) );
  NAND U863 ( .A(n668), .B(n669), .Z(n197) );
  NANDN U864 ( .B(n339), .A(Y[6]), .Z(n669) );
  AND U865 ( .A(n670), .B(n671), .Z(n668) );
  NANDN U866 ( .B(n386), .A(Y[6]), .Z(n671) );
  NANDN U867 ( .B(n391), .A(n358), .Z(n670) );
  XNOR U868 ( .A(n667), .B(Y0[7]), .Z(n358) );
  XNOR U869 ( .A(n673), .B(n674), .Z(n672) );
  AND U870 ( .A(n402), .B(n675), .Z(n674) );
  XOR U871 ( .A(n628), .B(n678), .Z(n675) );
  XOR U872 ( .A(n678), .B(n629), .Z(n628) );
  OR U873 ( .A(n676), .B(n677), .Z(n629) );
  XNOR U874 ( .A(n630), .B(n631), .Z(n678) );
  XNOR U875 ( .A(n639), .B(n638), .Z(n630) );
  XOR U876 ( .A(n683), .B(n648), .Z(n638) );
  XNOR U877 ( .A(n635), .B(n636), .Z(n648) );
  NAND U878 ( .A(n549), .B(n521), .Z(n636) );
  XNOR U879 ( .A(n634), .B(n684), .Z(n635) );
  AND U880 ( .A(n484), .B(n590), .Z(n684) );
  XNOR U881 ( .A(n647), .B(n637), .Z(n683) );
  XNOR U882 ( .A(n691), .B(n646), .Z(n647) );
  XNOR U883 ( .A(n695), .B(n644), .Z(n691) );
  NAND U884 ( .A(n643), .B(n449), .Z(n644) );
  NANDN U885 ( .B(n423), .A(n697), .Z(n696) );
  XNOR U886 ( .A(n651), .B(n702), .Z(n654) );
  AND U887 ( .A(n566), .B(n517), .Z(n702) );
  XOR U888 ( .A(n703), .B(n704), .Z(n651) );
  ANDN U889 ( .A(n705), .B(n706), .Z(n704) );
  XNOR U890 ( .A(n707), .B(n703), .Z(n705) );
  XOR U891 ( .A(n708), .B(n655), .Z(n701) );
  NAND U892 ( .A(n479), .B(n611), .Z(n655) );
  IV U893 ( .A(n657), .Z(n708) );
  XNOR U894 ( .A(n664), .B(n665), .Z(n659) );
  NANDN U895 ( .B(n424), .A(n712), .Z(n665) );
  AND U896 ( .A(n660), .B(n448), .Z(n713) );
  NAND U897 ( .A(n714), .B(n715), .Z(n663) );
  NANDN U898 ( .B(n716), .A(n717), .Z(n714) );
  IV U899 ( .A(n666), .Z(n673) );
  NAND U900 ( .A(n720), .B(n721), .Z(n196) );
  NANDN U901 ( .B(n339), .A(Y[5]), .Z(n721) );
  AND U902 ( .A(n722), .B(n723), .Z(n720) );
  NANDN U903 ( .B(n386), .A(Y[5]), .Z(n723) );
  NANDN U904 ( .B(n391), .A(n355), .Z(n722) );
  XNOR U905 ( .A(n719), .B(Y0[6]), .Z(n355) );
  XNOR U906 ( .A(n724), .B(n725), .Z(n719) );
  AND U907 ( .A(n402), .B(n727), .Z(n726) );
  XOR U908 ( .A(n676), .B(n728), .Z(n727) );
  XOR U909 ( .A(n728), .B(n677), .Z(n676) );
  OR U910 ( .A(n729), .B(n730), .Z(n677) );
  IV U911 ( .A(n725), .Z(n728) );
  XOR U912 ( .A(n682), .B(n681), .Z(n725) );
  XNOR U913 ( .A(n680), .B(n731), .Z(n681) );
  AND U914 ( .A(n679), .B(n732), .Z(n731) );
  AND U915 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U916 ( .B(n423), .A(n735), .Z(n734) );
  OR U917 ( .A(n736), .B(n737), .Z(n733) );
  AND U918 ( .A(n738), .B(n739), .Z(n679) );
  NANDN U919 ( .B(n740), .A(n741), .Z(n739) );
  NANDN U920 ( .B(n742), .A(n743), .Z(n738) );
  XNOR U921 ( .A(n747), .B(n694), .Z(n689) );
  XNOR U922 ( .A(n686), .B(n687), .Z(n694) );
  NAND U923 ( .A(n549), .B(n566), .Z(n687) );
  XNOR U924 ( .A(n685), .B(n748), .Z(n686) );
  AND U925 ( .A(n521), .B(n590), .Z(n748) );
  XNOR U926 ( .A(n693), .B(n688), .Z(n747) );
  XNOR U927 ( .A(n698), .B(n756), .Z(n699) );
  AND U928 ( .A(n449), .B(n697), .Z(n756) );
  XOR U929 ( .A(n757), .B(n758), .Z(n698) );
  ANDN U930 ( .A(n759), .B(n760), .Z(n758) );
  XNOR U931 ( .A(n761), .B(n757), .Z(n759) );
  XOR U932 ( .A(n762), .B(n700), .Z(n755) );
  NAND U933 ( .A(n643), .B(n484), .Z(n700) );
  IV U934 ( .A(n692), .Z(n762) );
  XNOR U935 ( .A(n703), .B(n767), .Z(n706) );
  AND U936 ( .A(n611), .B(n517), .Z(n767) );
  XOR U937 ( .A(n768), .B(n769), .Z(n703) );
  ANDN U938 ( .A(n770), .B(n771), .Z(n769) );
  XNOR U939 ( .A(n772), .B(n768), .Z(n770) );
  XOR U940 ( .A(n773), .B(n707), .Z(n766) );
  NAND U941 ( .A(n479), .B(n660), .Z(n707) );
  IV U942 ( .A(n709), .Z(n773) );
  XNOR U943 ( .A(n716), .B(n717), .Z(n711) );
  NANDN U944 ( .B(n424), .A(n777), .Z(n717) );
  XNOR U945 ( .A(n715), .B(n778), .Z(n716) );
  AND U946 ( .A(n712), .B(n448), .Z(n778) );
  ANDN U947 ( .A(n779), .B(n780), .Z(n715) );
  NANDN U948 ( .B(n781), .A(n782), .Z(n779) );
  NAND U949 ( .A(n785), .B(n786), .Z(n195) );
  NANDN U950 ( .B(n339), .A(Y[4]), .Z(n786) );
  AND U951 ( .A(n787), .B(n788), .Z(n785) );
  NANDN U952 ( .B(n386), .A(Y[4]), .Z(n788) );
  NANDN U953 ( .B(n391), .A(n352), .Z(n787) );
  XNOR U954 ( .A(n784), .B(Y0[5]), .Z(n352) );
  XNOR U955 ( .A(n789), .B(n790), .Z(n784) );
  AND U956 ( .A(n402), .B(n792), .Z(n791) );
  XOR U957 ( .A(n729), .B(n793), .Z(n792) );
  XOR U958 ( .A(n793), .B(n730), .Z(n729) );
  OR U959 ( .A(n794), .B(n795), .Z(n730) );
  IV U960 ( .A(n790), .Z(n793) );
  XOR U961 ( .A(n746), .B(n745), .Z(n790) );
  XOR U962 ( .A(n740), .B(n741), .Z(n737) );
  XOR U963 ( .A(n800), .B(n742), .Z(n740) );
  NAND U964 ( .A(n449), .B(n735), .Z(n742) );
  NANDN U965 ( .B(n743), .A(n801), .Z(n800) );
  NANDN U966 ( .B(n423), .A(n802), .Z(n801) );
  XOR U967 ( .A(n806), .B(n736), .Z(n796) );
  OR U968 ( .A(n807), .B(n808), .Z(n736) );
  IV U969 ( .A(n744), .Z(n806) );
  XNOR U970 ( .A(n812), .B(n765), .Z(n753) );
  XNOR U971 ( .A(n750), .B(n751), .Z(n765) );
  NAND U972 ( .A(n549), .B(n611), .Z(n751) );
  XNOR U973 ( .A(n749), .B(n813), .Z(n750) );
  AND U974 ( .A(n566), .B(n590), .Z(n813) );
  XNOR U975 ( .A(n764), .B(n752), .Z(n812) );
  XNOR U976 ( .A(n757), .B(n821), .Z(n760) );
  AND U977 ( .A(n484), .B(n697), .Z(n821) );
  XOR U978 ( .A(n822), .B(n823), .Z(n757) );
  ANDN U979 ( .A(n824), .B(n825), .Z(n823) );
  XNOR U980 ( .A(n826), .B(n822), .Z(n824) );
  XOR U981 ( .A(n827), .B(n761), .Z(n820) );
  NAND U982 ( .A(n643), .B(n521), .Z(n761) );
  IV U983 ( .A(n763), .Z(n827) );
  XNOR U984 ( .A(n768), .B(n832), .Z(n771) );
  AND U985 ( .A(n660), .B(n517), .Z(n832) );
  XOR U986 ( .A(n833), .B(n834), .Z(n768) );
  ANDN U987 ( .A(n835), .B(n836), .Z(n834) );
  XNOR U988 ( .A(n837), .B(n833), .Z(n835) );
  XOR U989 ( .A(n838), .B(n772), .Z(n831) );
  NAND U990 ( .A(n479), .B(n712), .Z(n772) );
  IV U991 ( .A(n774), .Z(n838) );
  XNOR U992 ( .A(n781), .B(n782), .Z(n776) );
  NANDN U993 ( .B(n424), .A(n842), .Z(n782) );
  AND U994 ( .A(n777), .B(n448), .Z(n843) );
  NAND U995 ( .A(n844), .B(n845), .Z(n780) );
  NANDN U996 ( .B(n846), .A(n847), .Z(n844) );
  NAND U997 ( .A(n850), .B(n851), .Z(n194) );
  NANDN U998 ( .B(n339), .A(Y[3]), .Z(n851) );
  AND U999 ( .A(n852), .B(n853), .Z(n850) );
  NANDN U1000 ( .B(n386), .A(Y[3]), .Z(n853) );
  NANDN U1001 ( .B(n391), .A(n349), .Z(n852) );
  XNOR U1002 ( .A(n849), .B(Y0[4]), .Z(n349) );
  XNOR U1003 ( .A(n854), .B(n855), .Z(n849) );
  AND U1004 ( .A(n402), .B(n857), .Z(n856) );
  XOR U1005 ( .A(n794), .B(n858), .Z(n857) );
  XOR U1006 ( .A(n858), .B(n795), .Z(n794) );
  OR U1007 ( .A(n859), .B(n860), .Z(n795) );
  IV U1008 ( .A(n855), .Z(n858) );
  XOR U1009 ( .A(n811), .B(n810), .Z(n855) );
  XOR U1010 ( .A(n861), .B(n807), .Z(n810) );
  XOR U1011 ( .A(n799), .B(n798), .Z(n807) );
  XOR U1012 ( .A(n797), .B(n862), .Z(n798) );
  AND U1013 ( .A(n863), .B(n864), .Z(n862) );
  NANDN U1014 ( .B(n423), .A(n865), .Z(n864) );
  OR U1015 ( .A(n866), .B(n867), .Z(n863) );
  NAND U1016 ( .A(n484), .B(n735), .Z(n805) );
  XNOR U1017 ( .A(n803), .B(n871), .Z(n804) );
  AND U1018 ( .A(n802), .B(n449), .Z(n871) );
  NANDN U1019 ( .B(n875), .A(n876), .Z(n808) );
  XNOR U1020 ( .A(n880), .B(n830), .Z(n818) );
  XNOR U1021 ( .A(n815), .B(n816), .Z(n830) );
  NAND U1022 ( .A(n549), .B(n660), .Z(n816) );
  XNOR U1023 ( .A(n814), .B(n881), .Z(n815) );
  AND U1024 ( .A(n611), .B(n590), .Z(n881) );
  XNOR U1025 ( .A(n829), .B(n817), .Z(n880) );
  XNOR U1026 ( .A(n822), .B(n889), .Z(n825) );
  AND U1027 ( .A(n521), .B(n697), .Z(n889) );
  XOR U1028 ( .A(n890), .B(n891), .Z(n822) );
  ANDN U1029 ( .A(n892), .B(n893), .Z(n891) );
  XNOR U1030 ( .A(n894), .B(n890), .Z(n892) );
  XOR U1031 ( .A(n895), .B(n826), .Z(n888) );
  NAND U1032 ( .A(n643), .B(n566), .Z(n826) );
  IV U1033 ( .A(n828), .Z(n895) );
  XNOR U1034 ( .A(n833), .B(n900), .Z(n836) );
  AND U1035 ( .A(n712), .B(n517), .Z(n900) );
  XOR U1036 ( .A(n901), .B(n902), .Z(n833) );
  ANDN U1037 ( .A(n903), .B(n904), .Z(n902) );
  XNOR U1038 ( .A(n905), .B(n901), .Z(n903) );
  XOR U1039 ( .A(n906), .B(n837), .Z(n899) );
  NAND U1040 ( .A(n479), .B(n777), .Z(n837) );
  IV U1041 ( .A(n839), .Z(n906) );
  XNOR U1042 ( .A(n846), .B(n847), .Z(n841) );
  NANDN U1043 ( .B(n424), .A(n910), .Z(n847) );
  XNOR U1044 ( .A(n845), .B(n911), .Z(n846) );
  AND U1045 ( .A(n842), .B(n448), .Z(n911) );
  ANDN U1046 ( .A(n912), .B(n913), .Z(n845) );
  NANDN U1047 ( .B(n914), .A(n915), .Z(n912) );
  NAND U1048 ( .A(n918), .B(n919), .Z(n193) );
  NANDN U1049 ( .B(n339), .A(Y[2]), .Z(n919) );
  AND U1050 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1051 ( .B(n386), .A(Y[2]), .Z(n921) );
  NANDN U1052 ( .B(n391), .A(n346), .Z(n920) );
  XNOR U1053 ( .A(n917), .B(Y0[3]), .Z(n346) );
  XNOR U1054 ( .A(n922), .B(n923), .Z(n917) );
  AND U1055 ( .A(n402), .B(n925), .Z(n924) );
  XOR U1056 ( .A(n859), .B(n926), .Z(n925) );
  XOR U1057 ( .A(n926), .B(n860), .Z(n859) );
  OR U1058 ( .A(n927), .B(n928), .Z(n860) );
  IV U1059 ( .A(n923), .Z(n926) );
  XOR U1060 ( .A(n879), .B(n878), .Z(n923) );
  XOR U1061 ( .A(n929), .B(n875), .Z(n878) );
  XOR U1062 ( .A(n870), .B(n869), .Z(n875) );
  XNOR U1063 ( .A(n934), .B(n866), .Z(n930) );
  NAND U1064 ( .A(n449), .B(n865), .Z(n866) );
  NANDN U1065 ( .B(n423), .A(n936), .Z(n935) );
  NAND U1066 ( .A(n521), .B(n735), .Z(n874) );
  XNOR U1067 ( .A(n872), .B(n940), .Z(n873) );
  AND U1068 ( .A(n802), .B(n484), .Z(n940) );
  XNOR U1069 ( .A(n876), .B(n877), .Z(n929) );
  XNOR U1070 ( .A(n950), .B(n898), .Z(n886) );
  XNOR U1071 ( .A(n883), .B(n884), .Z(n898) );
  NAND U1072 ( .A(n549), .B(n712), .Z(n884) );
  XNOR U1073 ( .A(n882), .B(n951), .Z(n883) );
  AND U1074 ( .A(n660), .B(n590), .Z(n951) );
  XNOR U1075 ( .A(n897), .B(n885), .Z(n950) );
  XNOR U1076 ( .A(n890), .B(n959), .Z(n893) );
  AND U1077 ( .A(n566), .B(n697), .Z(n959) );
  XOR U1078 ( .A(n963), .B(n894), .Z(n958) );
  NAND U1079 ( .A(n643), .B(n611), .Z(n894) );
  IV U1080 ( .A(n896), .Z(n963) );
  XNOR U1081 ( .A(n901), .B(n968), .Z(n904) );
  AND U1082 ( .A(n777), .B(n517), .Z(n968) );
  XOR U1083 ( .A(n969), .B(n970), .Z(n901) );
  ANDN U1084 ( .A(n971), .B(n972), .Z(n970) );
  XNOR U1085 ( .A(n973), .B(n969), .Z(n971) );
  XOR U1086 ( .A(n974), .B(n905), .Z(n967) );
  NAND U1087 ( .A(n479), .B(n842), .Z(n905) );
  IV U1088 ( .A(n907), .Z(n974) );
  XNOR U1089 ( .A(n914), .B(n915), .Z(n909) );
  OR U1090 ( .A(n978), .B(n424), .Z(n915) );
  AND U1091 ( .A(n910), .B(n448), .Z(n979) );
  NAND U1092 ( .A(n980), .B(n981), .Z(n913) );
  NANDN U1093 ( .B(n982), .A(n983), .Z(n980) );
  NAND U1094 ( .A(n986), .B(n987), .Z(n192) );
  NANDN U1095 ( .B(n339), .A(Y[1]), .Z(n987) );
  AND U1096 ( .A(n988), .B(n989), .Z(n986) );
  NANDN U1097 ( .B(n386), .A(Y[1]), .Z(n989) );
  NANDN U1098 ( .B(n391), .A(n342), .Z(n988) );
  XNOR U1099 ( .A(n985), .B(Y0[2]), .Z(n342) );
  XNOR U1100 ( .A(n990), .B(n991), .Z(n985) );
  XOR U1101 ( .A(n984), .B(n992), .Z(n990) );
  AND U1102 ( .A(n402), .B(n993), .Z(n992) );
  XOR U1103 ( .A(n927), .B(n994), .Z(n993) );
  XOR U1104 ( .A(n994), .B(n928), .Z(n927) );
  NANDN U1105 ( .B(n995), .A(n996), .Z(n928) );
  IV U1106 ( .A(n991), .Z(n994) );
  XOR U1107 ( .A(n946), .B(n945), .Z(n991) );
  XNOR U1108 ( .A(n997), .B(n949), .Z(n945) );
  XNOR U1109 ( .A(n937), .B(n999), .Z(n938) );
  AND U1110 ( .A(n936), .B(n449), .Z(n999) );
  XOR U1111 ( .A(n1003), .B(n939), .Z(n998) );
  NAND U1112 ( .A(n484), .B(n865), .Z(n939) );
  IV U1113 ( .A(n931), .Z(n1003) );
  XNOR U1114 ( .A(n942), .B(n943), .Z(n933) );
  NAND U1115 ( .A(n566), .B(n735), .Z(n943) );
  XNOR U1116 ( .A(n941), .B(n1007), .Z(n942) );
  AND U1117 ( .A(n802), .B(n521), .Z(n1007) );
  XNOR U1118 ( .A(n948), .B(n944), .Z(n997) );
  AND U1119 ( .A(n1015), .B(n1016), .Z(n1014) );
  OR U1120 ( .A(n1017), .B(n1018), .Z(n1016) );
  AND U1121 ( .A(n1019), .B(n1020), .Z(n1015) );
  NANDN U1122 ( .B(n423), .A(n1021), .Z(n1020) );
  NANDN U1123 ( .B(n1022), .A(n1023), .Z(n1019) );
  XNOR U1124 ( .A(n1027), .B(n966), .Z(n956) );
  XNOR U1125 ( .A(n953), .B(n954), .Z(n966) );
  NAND U1126 ( .A(n549), .B(n777), .Z(n954) );
  XNOR U1127 ( .A(n952), .B(n1028), .Z(n953) );
  AND U1128 ( .A(n712), .B(n590), .Z(n1028) );
  XNOR U1129 ( .A(n965), .B(n955), .Z(n1027) );
  XNOR U1130 ( .A(n960), .B(n1036), .Z(n961) );
  AND U1131 ( .A(n611), .B(n697), .Z(n1036) );
  XOR U1132 ( .A(n1040), .B(n962), .Z(n1035) );
  NAND U1133 ( .A(n643), .B(n660), .Z(n962) );
  IV U1134 ( .A(n964), .Z(n1040) );
  XNOR U1135 ( .A(n969), .B(n1045), .Z(n972) );
  AND U1136 ( .A(n842), .B(n517), .Z(n1045) );
  XOR U1137 ( .A(n1046), .B(n1047), .Z(n969) );
  ANDN U1138 ( .A(n1048), .B(n1049), .Z(n1047) );
  XNOR U1139 ( .A(n1050), .B(n1046), .Z(n1048) );
  XOR U1140 ( .A(n1051), .B(n973), .Z(n1044) );
  NAND U1141 ( .A(n479), .B(n910), .Z(n973) );
  IV U1142 ( .A(n975), .Z(n1051) );
  XNOR U1143 ( .A(n982), .B(n983), .Z(n977) );
  OR U1144 ( .A(n1055), .B(n424), .Z(n983) );
  XNOR U1145 ( .A(n981), .B(n1056), .Z(n982) );
  ANDN U1146 ( .A(n448), .B(n978), .Z(n1056) );
  ANDN U1147 ( .A(n1057), .B(n1058), .Z(n981) );
  NANDN U1148 ( .B(n1059), .A(n1060), .Z(n1057) );
  NAND U1149 ( .A(n1063), .B(n1064), .Z(n191) );
  NANDN U1150 ( .B(n339), .A(Y[0]), .Z(n1064) );
  AND U1151 ( .A(n1065), .B(n1066), .Z(n1063) );
  NANDN U1152 ( .B(n386), .A(Y[0]), .Z(n1066) );
  IV U1153 ( .A(n1067), .Z(n386) );
  OR U1154 ( .A(n391), .B(n337), .Z(n1065) );
  IV U1155 ( .A(Y0[1]), .Z(n343) );
  XOR U1156 ( .A(n1068), .B(n1069), .Z(n1062) );
  XNOR U1157 ( .A(n1070), .B(n1061), .Z(n1068) );
  NAND U1158 ( .A(Y0[0]), .B(n995), .Z(n1061) );
  NAND U1159 ( .A(n1071), .B(n402), .Z(n1070) );
  XOR U1160 ( .A(A[15]), .B(X[15]), .Z(n402) );
  XNOR U1161 ( .A(n996), .B(n1069), .Z(n1071) );
  XNOR U1162 ( .A(n995), .B(n1069), .Z(n996) );
  XNOR U1163 ( .A(n1013), .B(n1012), .Z(n1069) );
  XNOR U1164 ( .A(n1072), .B(n1026), .Z(n1012) );
  XNOR U1165 ( .A(n1000), .B(n1074), .Z(n1001) );
  AND U1166 ( .A(n936), .B(n484), .Z(n1074) );
  XOR U1167 ( .A(n1078), .B(n1002), .Z(n1073) );
  NAND U1168 ( .A(n521), .B(n865), .Z(n1002) );
  IV U1169 ( .A(n1004), .Z(n1078) );
  XNOR U1170 ( .A(n1009), .B(n1010), .Z(n1006) );
  NAND U1171 ( .A(n611), .B(n735), .Z(n1010) );
  XNOR U1172 ( .A(n1008), .B(n1082), .Z(n1009) );
  AND U1173 ( .A(n802), .B(n566), .Z(n1082) );
  XNOR U1174 ( .A(n1025), .B(n1011), .Z(n1072) );
  XNOR U1175 ( .A(n1089), .B(n1022), .Z(n1025) );
  XOR U1176 ( .A(n1090), .B(n1017), .Z(n1022) );
  NAND U1177 ( .A(n449), .B(n1021), .Z(n1017) );
  NANDN U1178 ( .B(n423), .A(n1092), .Z(n1091) );
  XNOR U1179 ( .A(n1023), .B(n1024), .Z(n1089) );
  XNOR U1180 ( .A(n1102), .B(n1043), .Z(n1033) );
  XNOR U1181 ( .A(n1030), .B(n1031), .Z(n1043) );
  NAND U1182 ( .A(n549), .B(n842), .Z(n1031) );
  XNOR U1183 ( .A(n1029), .B(n1103), .Z(n1030) );
  AND U1184 ( .A(n777), .B(n590), .Z(n1103) );
  XNOR U1185 ( .A(n1042), .B(n1032), .Z(n1102) );
  XNOR U1186 ( .A(n1037), .B(n1111), .Z(n1038) );
  AND U1187 ( .A(n660), .B(n697), .Z(n1111) );
  XOR U1188 ( .A(n1115), .B(n1039), .Z(n1110) );
  NAND U1189 ( .A(n643), .B(n712), .Z(n1039) );
  IV U1190 ( .A(n1041), .Z(n1115) );
  XNOR U1191 ( .A(n1046), .B(n1120), .Z(n1049) );
  AND U1192 ( .A(n910), .B(n517), .Z(n1120) );
  XOR U1193 ( .A(n1124), .B(n1050), .Z(n1119) );
  NANDN U1194 ( .B(n978), .A(n479), .Z(n1050) );
  IV U1195 ( .A(n1052), .Z(n1124) );
  XNOR U1196 ( .A(n1059), .B(n1060), .Z(n1054) );
  NANDN U1197 ( .B(n424), .A(n1128), .Z(n1060) );
  ANDN U1198 ( .A(n448), .B(n1055), .Z(n1129) );
  NAND U1199 ( .A(n1130), .B(n1131), .Z(n1058) );
  NANDN U1200 ( .B(n1132), .A(n1133), .Z(n1130) );
  XNOR U1201 ( .A(n1088), .B(n1087), .Z(n995) );
  XNOR U1202 ( .A(n1134), .B(n1098), .Z(n1087) );
  XNOR U1203 ( .A(n1075), .B(n1136), .Z(n1076) );
  AND U1204 ( .A(n936), .B(n521), .Z(n1136) );
  XOR U1205 ( .A(n1140), .B(n1077), .Z(n1135) );
  NAND U1206 ( .A(n566), .B(n865), .Z(n1077) );
  IV U1207 ( .A(n1079), .Z(n1140) );
  XNOR U1208 ( .A(n1084), .B(n1085), .Z(n1081) );
  NAND U1209 ( .A(n660), .B(n735), .Z(n1085) );
  XNOR U1210 ( .A(n1083), .B(n1144), .Z(n1084) );
  AND U1211 ( .A(n802), .B(n611), .Z(n1144) );
  XNOR U1212 ( .A(n1097), .B(n1086), .Z(n1134) );
  XOR U1213 ( .A(n1148), .B(n1149), .Z(n1086) );
  XNOR U1214 ( .A(n1150), .B(n1101), .Z(n1097) );
  NAND U1215 ( .A(n484), .B(n1021), .Z(n1095) );
  XNOR U1216 ( .A(n1093), .B(n1151), .Z(n1094) );
  AND U1217 ( .A(n1092), .B(n449), .Z(n1151) );
  XNOR U1218 ( .A(n1100), .B(n1096), .Z(n1150) );
  XOR U1219 ( .A(n1155), .B(n1156), .Z(n1096) );
  AND U1220 ( .A(n1157), .B(n1158), .Z(n1156) );
  XOR U1221 ( .A(n1159), .B(n1160), .Z(n1158) );
  XOR U1222 ( .A(n1155), .B(n1161), .Z(n1160) );
  XOR U1223 ( .A(n1142), .B(n1162), .Z(n1157) );
  XOR U1224 ( .A(n1155), .B(n1143), .Z(n1162) );
  NAND U1225 ( .A(n735), .B(n712), .Z(n1147) );
  XNOR U1226 ( .A(n1145), .B(n1163), .Z(n1146) );
  AND U1227 ( .A(n802), .B(n660), .Z(n1163) );
  XNOR U1228 ( .A(n1137), .B(n1168), .Z(n1138) );
  AND U1229 ( .A(n936), .B(n566), .Z(n1168) );
  XOR U1230 ( .A(n1169), .B(n1170), .Z(n1137) );
  ANDN U1231 ( .A(n1171), .B(n1172), .Z(n1170) );
  XNOR U1232 ( .A(n1173), .B(n1169), .Z(n1171) );
  XOR U1233 ( .A(n1174), .B(n1139), .Z(n1167) );
  NAND U1234 ( .A(n611), .B(n865), .Z(n1139) );
  IV U1235 ( .A(n1141), .Z(n1174) );
  XOR U1236 ( .A(n1178), .B(n1179), .Z(n1155) );
  AND U1237 ( .A(n1180), .B(n1181), .Z(n1179) );
  XOR U1238 ( .A(n1182), .B(n1183), .Z(n1181) );
  XOR U1239 ( .A(n1178), .B(n1184), .Z(n1183) );
  XOR U1240 ( .A(n1176), .B(n1185), .Z(n1180) );
  XOR U1241 ( .A(n1178), .B(n1177), .Z(n1185) );
  NAND U1242 ( .A(n735), .B(n777), .Z(n1166) );
  XNOR U1243 ( .A(n1164), .B(n1186), .Z(n1165) );
  AND U1244 ( .A(n712), .B(n802), .Z(n1186) );
  XNOR U1245 ( .A(n1169), .B(n1191), .Z(n1172) );
  AND U1246 ( .A(n936), .B(n611), .Z(n1191) );
  XOR U1247 ( .A(n1192), .B(n1193), .Z(n1169) );
  ANDN U1248 ( .A(n1194), .B(n1195), .Z(n1193) );
  XNOR U1249 ( .A(n1196), .B(n1192), .Z(n1194) );
  XOR U1250 ( .A(n1197), .B(n1173), .Z(n1190) );
  NAND U1251 ( .A(n660), .B(n865), .Z(n1173) );
  IV U1252 ( .A(n1175), .Z(n1197) );
  XOR U1253 ( .A(n1201), .B(n1202), .Z(n1178) );
  AND U1254 ( .A(n1203), .B(n1204), .Z(n1202) );
  XOR U1255 ( .A(n1205), .B(n1206), .Z(n1204) );
  XOR U1256 ( .A(n1201), .B(n1207), .Z(n1206) );
  XOR U1257 ( .A(n1199), .B(n1208), .Z(n1203) );
  XOR U1258 ( .A(n1201), .B(n1200), .Z(n1208) );
  NAND U1259 ( .A(n735), .B(n842), .Z(n1189) );
  XNOR U1260 ( .A(n1187), .B(n1209), .Z(n1188) );
  AND U1261 ( .A(n777), .B(n802), .Z(n1209) );
  XNOR U1262 ( .A(n1192), .B(n1214), .Z(n1195) );
  AND U1263 ( .A(n936), .B(n660), .Z(n1214) );
  XOR U1264 ( .A(n1215), .B(n1216), .Z(n1192) );
  ANDN U1265 ( .A(n1217), .B(n1218), .Z(n1216) );
  XNOR U1266 ( .A(n1219), .B(n1215), .Z(n1217) );
  XOR U1267 ( .A(n1220), .B(n1196), .Z(n1213) );
  NAND U1268 ( .A(n865), .B(n712), .Z(n1196) );
  IV U1269 ( .A(n1198), .Z(n1220) );
  XOR U1270 ( .A(n1224), .B(n1225), .Z(n1201) );
  AND U1271 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U1272 ( .A(n1228), .B(n1229), .Z(n1227) );
  XOR U1273 ( .A(n1224), .B(n1230), .Z(n1229) );
  XOR U1274 ( .A(n1222), .B(n1231), .Z(n1226) );
  XOR U1275 ( .A(n1224), .B(n1223), .Z(n1231) );
  XNOR U1276 ( .A(n1232), .B(n1212), .Z(n1223) );
  NAND U1277 ( .A(n735), .B(n910), .Z(n1212) );
  IV U1278 ( .A(n1211), .Z(n1232) );
  XNOR U1279 ( .A(n1210), .B(n1233), .Z(n1211) );
  AND U1280 ( .A(n842), .B(n802), .Z(n1233) );
  XOR U1281 ( .A(n1234), .B(n1235), .Z(n1210) );
  ANDN U1282 ( .A(n1236), .B(n1237), .Z(n1235) );
  XNOR U1283 ( .A(n1238), .B(n1234), .Z(n1236) );
  XNOR U1284 ( .A(n1239), .B(n1240), .Z(n1222) );
  IV U1285 ( .A(n1218), .Z(n1240) );
  XNOR U1286 ( .A(n1215), .B(n1241), .Z(n1218) );
  AND U1287 ( .A(n712), .B(n936), .Z(n1241) );
  XOR U1288 ( .A(n1242), .B(n1243), .Z(n1215) );
  ANDN U1289 ( .A(n1244), .B(n1245), .Z(n1243) );
  XNOR U1290 ( .A(n1246), .B(n1242), .Z(n1244) );
  XOR U1291 ( .A(n1247), .B(n1219), .Z(n1239) );
  NAND U1292 ( .A(n865), .B(n777), .Z(n1219) );
  IV U1293 ( .A(n1221), .Z(n1247) );
  XOR U1294 ( .A(n1251), .B(n1252), .Z(n1224) );
  AND U1295 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U1296 ( .A(n1255), .B(n1256), .Z(n1254) );
  XOR U1297 ( .A(n1251), .B(n1257), .Z(n1256) );
  XOR U1298 ( .A(n1249), .B(n1258), .Z(n1253) );
  XOR U1299 ( .A(n1251), .B(n1250), .Z(n1258) );
  XNOR U1300 ( .A(n1259), .B(n1238), .Z(n1250) );
  NANDN U1301 ( .B(n978), .A(n735), .Z(n1238) );
  IV U1302 ( .A(n1237), .Z(n1259) );
  XNOR U1303 ( .A(n1234), .B(n1260), .Z(n1237) );
  AND U1304 ( .A(n910), .B(n802), .Z(n1260) );
  XOR U1305 ( .A(n1261), .B(n1262), .Z(n1234) );
  ANDN U1306 ( .A(n1263), .B(n1264), .Z(n1262) );
  XNOR U1307 ( .A(n1265), .B(n1261), .Z(n1263) );
  XNOR U1308 ( .A(n1266), .B(n1267), .Z(n1249) );
  IV U1309 ( .A(n1245), .Z(n1267) );
  XNOR U1310 ( .A(n1242), .B(n1268), .Z(n1245) );
  AND U1311 ( .A(n777), .B(n936), .Z(n1268) );
  XOR U1312 ( .A(n1269), .B(n1270), .Z(n1242) );
  ANDN U1313 ( .A(n1271), .B(n1272), .Z(n1270) );
  XNOR U1314 ( .A(n1273), .B(n1269), .Z(n1271) );
  XOR U1315 ( .A(n1274), .B(n1246), .Z(n1266) );
  NAND U1316 ( .A(n865), .B(n842), .Z(n1246) );
  IV U1317 ( .A(n1248), .Z(n1274) );
  XOR U1318 ( .A(n1278), .B(n1279), .Z(n1251) );
  AND U1319 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U1320 ( .A(n1282), .B(n1283), .Z(n1281) );
  XOR U1321 ( .A(n1278), .B(n1284), .Z(n1283) );
  XOR U1322 ( .A(n1276), .B(n1285), .Z(n1280) );
  XOR U1323 ( .A(n1278), .B(n1277), .Z(n1285) );
  XNOR U1324 ( .A(n1286), .B(n1265), .Z(n1277) );
  NANDN U1325 ( .B(n1055), .A(n735), .Z(n1265) );
  IV U1326 ( .A(n1264), .Z(n1286) );
  XNOR U1327 ( .A(n1261), .B(n1287), .Z(n1264) );
  ANDN U1328 ( .A(n802), .B(n978), .Z(n1287) );
  XOR U1329 ( .A(n1288), .B(n1289), .Z(n1261) );
  ANDN U1330 ( .A(n1290), .B(n1291), .Z(n1289) );
  XNOR U1331 ( .A(n1292), .B(n1288), .Z(n1290) );
  XNOR U1332 ( .A(n1293), .B(n1294), .Z(n1276) );
  IV U1333 ( .A(n1272), .Z(n1294) );
  XNOR U1334 ( .A(n1269), .B(n1295), .Z(n1272) );
  AND U1335 ( .A(n842), .B(n936), .Z(n1295) );
  XOR U1336 ( .A(n1296), .B(n1297), .Z(n1269) );
  ANDN U1337 ( .A(n1298), .B(n1299), .Z(n1297) );
  XNOR U1338 ( .A(n1300), .B(n1296), .Z(n1298) );
  XOR U1339 ( .A(n1301), .B(n1273), .Z(n1293) );
  NAND U1340 ( .A(n865), .B(n910), .Z(n1273) );
  IV U1341 ( .A(n1275), .Z(n1301) );
  XOR U1342 ( .A(n1305), .B(n1306), .Z(n1278) );
  AND U1343 ( .A(n1307), .B(n1308), .Z(n1306) );
  XOR U1344 ( .A(n1309), .B(n1310), .Z(n1308) );
  XOR U1345 ( .A(n1305), .B(n1311), .Z(n1310) );
  XOR U1346 ( .A(n1303), .B(n1312), .Z(n1307) );
  XOR U1347 ( .A(n1305), .B(n1304), .Z(n1312) );
  XNOR U1348 ( .A(n1313), .B(n1292), .Z(n1304) );
  NAND U1349 ( .A(n735), .B(n1128), .Z(n1292) );
  IV U1350 ( .A(n1291), .Z(n1313) );
  XNOR U1351 ( .A(n1288), .B(n1314), .Z(n1291) );
  ANDN U1352 ( .A(n802), .B(n1055), .Z(n1314) );
  XOR U1353 ( .A(n1315), .B(n1316), .Z(n1288) );
  ANDN U1354 ( .A(n1317), .B(n1318), .Z(n1316) );
  XNOR U1355 ( .A(n1319), .B(n1315), .Z(n1317) );
  XNOR U1356 ( .A(n1320), .B(n1321), .Z(n1303) );
  IV U1357 ( .A(n1299), .Z(n1321) );
  XNOR U1358 ( .A(n1296), .B(n1322), .Z(n1299) );
  AND U1359 ( .A(n910), .B(n936), .Z(n1322) );
  XOR U1360 ( .A(n1323), .B(n1324), .Z(n1296) );
  ANDN U1361 ( .A(n1325), .B(n1326), .Z(n1324) );
  XNOR U1362 ( .A(n1327), .B(n1323), .Z(n1325) );
  XOR U1363 ( .A(n1328), .B(n1300), .Z(n1320) );
  NANDN U1364 ( .B(n978), .A(n865), .Z(n1300) );
  IV U1365 ( .A(n1302), .Z(n1328) );
  XOR U1366 ( .A(n1333), .B(n1334), .Z(n1149) );
  XNOR U1367 ( .A(n1335), .B(n1332), .Z(n1333) );
  XNOR U1368 ( .A(n1323), .B(n1337), .Z(n1326) );
  ANDN U1369 ( .A(n936), .B(n978), .Z(n1337) );
  XOR U1370 ( .A(n1340), .B(n1338), .Z(n1339) );
  ANDN U1371 ( .A(n936), .B(n1055), .Z(n1340) );
  AND U1372 ( .A(n1128), .B(n865), .Z(n1341) );
  XOR U1373 ( .A(n1342), .B(n1343), .Z(n1338) );
  ANDN U1374 ( .A(n1344), .B(n1345), .Z(n1343) );
  XNOR U1375 ( .A(n1346), .B(n1342), .Z(n1344) );
  XOR U1376 ( .A(n1347), .B(n1327), .Z(n1336) );
  NANDN U1377 ( .B(n1055), .A(n865), .Z(n1327) );
  IV U1378 ( .A(n1329), .Z(n1347) );
  NAND U1379 ( .A(n865), .B(n1348), .Z(n1346) );
  XNOR U1380 ( .A(n1342), .B(n1349), .Z(n1345) );
  AND U1381 ( .A(n1128), .B(n936), .Z(n1349) );
  AND U1382 ( .A(n1350), .B(A[0]), .Z(n1342) );
  NANDN U1383 ( .B(n865), .A(n1351), .Z(n1350) );
  NAND U1384 ( .A(n1348), .B(n936), .Z(n1351) );
  XNOR U1385 ( .A(n1318), .B(n1319), .Z(n1331) );
  NAND U1386 ( .A(n735), .B(n1348), .Z(n1319) );
  XNOR U1387 ( .A(n1315), .B(n1354), .Z(n1318) );
  AND U1388 ( .A(n1128), .B(n802), .Z(n1354) );
  AND U1389 ( .A(n1355), .B(A[0]), .Z(n1315) );
  NANDN U1390 ( .B(n735), .A(n1356), .Z(n1355) );
  NAND U1391 ( .A(n1348), .B(n802), .Z(n1356) );
  XOR U1392 ( .A(n1359), .B(n1360), .Z(n1332) );
  XOR U1393 ( .A(n1361), .B(n1362), .Z(n1100) );
  AND U1394 ( .A(n1363), .B(n1364), .Z(n1362) );
  NANDN U1395 ( .B(n423), .A(n1365), .Z(n1364) );
  NANDN U1396 ( .B(n1366), .A(n1367), .Z(n423) );
  AND U1397 ( .A(n1368), .B(A[15]), .Z(n1367) );
  OR U1398 ( .A(n1369), .B(n1370), .Z(n1363) );
  IV U1399 ( .A(n1099), .Z(n1361) );
  NAND U1400 ( .A(n521), .B(n1021), .Z(n1154) );
  XNOR U1401 ( .A(n1152), .B(n1372), .Z(n1153) );
  AND U1402 ( .A(n1092), .B(n484), .Z(n1372) );
  XOR U1403 ( .A(n1380), .B(n1369), .Z(n1376) );
  NAND U1404 ( .A(n449), .B(n1365), .Z(n1369) );
  IV U1405 ( .A(n1371), .Z(n1380) );
  NAND U1406 ( .A(n566), .B(n1021), .Z(n1375) );
  XNOR U1407 ( .A(n1373), .B(n1382), .Z(n1374) );
  AND U1408 ( .A(n1092), .B(n521), .Z(n1382) );
  XNOR U1409 ( .A(n1377), .B(n1387), .Z(n1378) );
  AND U1410 ( .A(n449), .B(X[0]), .Z(n1387) );
  XNOR U1411 ( .A(n1368), .B(A[14]), .Z(n1366) );
  NOR U1412 ( .A(n1388), .B(n1389), .Z(n1368) );
  XOR U1413 ( .A(n1393), .B(n1379), .Z(n1386) );
  NAND U1414 ( .A(n484), .B(n1365), .Z(n1379) );
  IV U1415 ( .A(n1381), .Z(n1393) );
  NAND U1416 ( .A(n611), .B(n1021), .Z(n1385) );
  XNOR U1417 ( .A(n1383), .B(n1395), .Z(n1384) );
  AND U1418 ( .A(n1092), .B(n566), .Z(n1395) );
  XOR U1419 ( .A(n1396), .B(n1397), .Z(n1383) );
  ANDN U1420 ( .A(n1398), .B(n1399), .Z(n1397) );
  XNOR U1421 ( .A(n1400), .B(n1396), .Z(n1398) );
  XNOR U1422 ( .A(n1390), .B(n1402), .Z(n1391) );
  AND U1423 ( .A(n484), .B(X[0]), .Z(n1402) );
  XOR U1424 ( .A(n1388), .B(A[13]), .Z(n1389) );
  NANDN U1425 ( .B(n1403), .A(n1404), .Z(n1388) );
  XOR U1426 ( .A(n1408), .B(n1392), .Z(n1401) );
  NAND U1427 ( .A(n521), .B(n1365), .Z(n1392) );
  IV U1428 ( .A(n1394), .Z(n1408) );
  XNOR U1429 ( .A(n1410), .B(n1400), .Z(n1228) );
  NAND U1430 ( .A(n660), .B(n1021), .Z(n1400) );
  IV U1431 ( .A(n1399), .Z(n1410) );
  XNOR U1432 ( .A(n1396), .B(n1411), .Z(n1399) );
  AND U1433 ( .A(n1092), .B(n611), .Z(n1411) );
  XOR U1434 ( .A(n1412), .B(n1413), .Z(n1396) );
  ANDN U1435 ( .A(n1414), .B(n1415), .Z(n1413) );
  XNOR U1436 ( .A(n1416), .B(n1412), .Z(n1414) );
  XNOR U1437 ( .A(n1417), .B(n1418), .Z(n1230) );
  IV U1438 ( .A(n1406), .Z(n1418) );
  XNOR U1439 ( .A(n1405), .B(n1419), .Z(n1406) );
  AND U1440 ( .A(n521), .B(X[0]), .Z(n1419) );
  XNOR U1441 ( .A(n1404), .B(A[12]), .Z(n1403) );
  NOR U1442 ( .A(n1420), .B(n1421), .Z(n1404) );
  XOR U1443 ( .A(n1422), .B(n1423), .Z(n1405) );
  ANDN U1444 ( .A(n1424), .B(n1425), .Z(n1423) );
  XNOR U1445 ( .A(n1426), .B(n1422), .Z(n1424) );
  XOR U1446 ( .A(n1427), .B(n1407), .Z(n1417) );
  NAND U1447 ( .A(n566), .B(n1365), .Z(n1407) );
  IV U1448 ( .A(n1409), .Z(n1427) );
  XNOR U1449 ( .A(n1429), .B(n1416), .Z(n1255) );
  NAND U1450 ( .A(n712), .B(n1021), .Z(n1416) );
  IV U1451 ( .A(n1415), .Z(n1429) );
  XNOR U1452 ( .A(n1412), .B(n1430), .Z(n1415) );
  AND U1453 ( .A(n1092), .B(n660), .Z(n1430) );
  XOR U1454 ( .A(n1431), .B(n1432), .Z(n1412) );
  ANDN U1455 ( .A(n1433), .B(n1434), .Z(n1432) );
  XNOR U1456 ( .A(n1435), .B(n1431), .Z(n1433) );
  XNOR U1457 ( .A(n1436), .B(n1437), .Z(n1257) );
  IV U1458 ( .A(n1425), .Z(n1437) );
  XNOR U1459 ( .A(n1422), .B(n1438), .Z(n1425) );
  AND U1460 ( .A(n566), .B(X[0]), .Z(n1438) );
  XOR U1461 ( .A(n1420), .B(A[11]), .Z(n1421) );
  NANDN U1462 ( .B(n1439), .A(n1440), .Z(n1420) );
  XOR U1463 ( .A(n1441), .B(n1442), .Z(n1422) );
  ANDN U1464 ( .A(n1443), .B(n1444), .Z(n1442) );
  XNOR U1465 ( .A(n1445), .B(n1441), .Z(n1443) );
  XOR U1466 ( .A(n1446), .B(n1426), .Z(n1436) );
  NAND U1467 ( .A(n611), .B(n1365), .Z(n1426) );
  IV U1468 ( .A(n1428), .Z(n1446) );
  XNOR U1469 ( .A(n1448), .B(n1435), .Z(n1282) );
  NAND U1470 ( .A(n777), .B(n1021), .Z(n1435) );
  IV U1471 ( .A(n1434), .Z(n1448) );
  XNOR U1472 ( .A(n1431), .B(n1449), .Z(n1434) );
  AND U1473 ( .A(n1092), .B(n712), .Z(n1449) );
  XOR U1474 ( .A(n1450), .B(n1451), .Z(n1431) );
  ANDN U1475 ( .A(n1452), .B(n1453), .Z(n1451) );
  XNOR U1476 ( .A(n1454), .B(n1450), .Z(n1452) );
  XNOR U1477 ( .A(n1455), .B(n1456), .Z(n1284) );
  IV U1478 ( .A(n1444), .Z(n1456) );
  XNOR U1479 ( .A(n1441), .B(n1457), .Z(n1444) );
  AND U1480 ( .A(n611), .B(X[0]), .Z(n1457) );
  XNOR U1481 ( .A(n1440), .B(A[10]), .Z(n1439) );
  NOR U1482 ( .A(n1458), .B(n1459), .Z(n1440) );
  XOR U1483 ( .A(n1460), .B(n1461), .Z(n1441) );
  ANDN U1484 ( .A(n1462), .B(n1463), .Z(n1461) );
  XNOR U1485 ( .A(n1464), .B(n1460), .Z(n1462) );
  XOR U1486 ( .A(n1465), .B(n1445), .Z(n1455) );
  NAND U1487 ( .A(n660), .B(n1365), .Z(n1445) );
  IV U1488 ( .A(n1447), .Z(n1465) );
  XNOR U1489 ( .A(n1467), .B(n1454), .Z(n1309) );
  NAND U1490 ( .A(n842), .B(n1021), .Z(n1454) );
  IV U1491 ( .A(n1453), .Z(n1467) );
  XNOR U1492 ( .A(n1450), .B(n1468), .Z(n1453) );
  AND U1493 ( .A(n1092), .B(n777), .Z(n1468) );
  XOR U1494 ( .A(n1469), .B(n1470), .Z(n1450) );
  ANDN U1495 ( .A(n1471), .B(n1472), .Z(n1470) );
  XNOR U1496 ( .A(n1473), .B(n1469), .Z(n1471) );
  XNOR U1497 ( .A(n1474), .B(n1475), .Z(n1311) );
  IV U1498 ( .A(n1463), .Z(n1475) );
  XNOR U1499 ( .A(n1460), .B(n1476), .Z(n1463) );
  AND U1500 ( .A(n660), .B(X[0]), .Z(n1476) );
  XOR U1501 ( .A(n1458), .B(A[9]), .Z(n1459) );
  NANDN U1502 ( .B(n1477), .A(n1478), .Z(n1458) );
  XOR U1503 ( .A(n1479), .B(n1480), .Z(n1460) );
  ANDN U1504 ( .A(n1481), .B(n1482), .Z(n1480) );
  XNOR U1505 ( .A(n1483), .B(n1479), .Z(n1481) );
  XOR U1506 ( .A(n1484), .B(n1464), .Z(n1474) );
  NAND U1507 ( .A(n712), .B(n1365), .Z(n1464) );
  IV U1508 ( .A(n1466), .Z(n1484) );
  NAND U1509 ( .A(n910), .B(n1021), .Z(n1473) );
  XNOR U1510 ( .A(n1469), .B(n1486), .Z(n1472) );
  AND U1511 ( .A(n1092), .B(n842), .Z(n1486) );
  XNOR U1512 ( .A(n1490), .B(n1487), .Z(n1489) );
  XNOR U1513 ( .A(n1479), .B(n1492), .Z(n1482) );
  AND U1514 ( .A(n712), .B(X[0]), .Z(n1492) );
  XNOR U1515 ( .A(n1496), .B(n1493), .Z(n1495) );
  XOR U1516 ( .A(n1497), .B(n1483), .Z(n1491) );
  NAND U1517 ( .A(n777), .B(n1365), .Z(n1483) );
  IV U1518 ( .A(n1485), .Z(n1497) );
  XNOR U1519 ( .A(n1498), .B(n1499), .Z(n1485) );
  AND U1520 ( .A(n1500), .B(n1501), .Z(n1499) );
  XOR U1521 ( .A(n1494), .B(n1502), .Z(n1501) );
  XNOR U1522 ( .A(n1496), .B(n1498), .Z(n1502) );
  NAND U1523 ( .A(n842), .B(n1365), .Z(n1496) );
  XOR U1524 ( .A(n1493), .B(n1503), .Z(n1494) );
  AND U1525 ( .A(n777), .B(X[0]), .Z(n1503) );
  XNOR U1526 ( .A(n1507), .B(n1504), .Z(n1506) );
  XOR U1527 ( .A(n1488), .B(n1508), .Z(n1500) );
  XNOR U1528 ( .A(n1490), .B(n1498), .Z(n1508) );
  NANDN U1529 ( .B(n978), .A(n1021), .Z(n1490) );
  XOR U1530 ( .A(n1487), .B(n1509), .Z(n1488) );
  AND U1531 ( .A(n1092), .B(n910), .Z(n1509) );
  XOR U1532 ( .A(n1510), .B(n1511), .Z(n1487) );
  AND U1533 ( .A(n1512), .B(n1513), .Z(n1511) );
  XNOR U1534 ( .A(n1514), .B(n1510), .Z(n1513) );
  XOR U1535 ( .A(n1515), .B(n1516), .Z(n1498) );
  AND U1536 ( .A(n1517), .B(n1518), .Z(n1516) );
  XOR U1537 ( .A(n1505), .B(n1519), .Z(n1518) );
  XNOR U1538 ( .A(n1507), .B(n1515), .Z(n1519) );
  NAND U1539 ( .A(n910), .B(n1365), .Z(n1507) );
  XOR U1540 ( .A(n1504), .B(n1520), .Z(n1505) );
  AND U1541 ( .A(n842), .B(X[0]), .Z(n1520) );
  XNOR U1542 ( .A(n1524), .B(n1521), .Z(n1523) );
  XOR U1543 ( .A(n1512), .B(n1525), .Z(n1517) );
  XNOR U1544 ( .A(n1514), .B(n1515), .Z(n1525) );
  NANDN U1545 ( .B(n1055), .A(n1021), .Z(n1514) );
  XOR U1546 ( .A(n1510), .B(n1526), .Z(n1512) );
  ANDN U1547 ( .A(n1092), .B(n978), .Z(n1526) );
  XOR U1548 ( .A(n1527), .B(n1528), .Z(n1510) );
  AND U1549 ( .A(n1529), .B(n1530), .Z(n1528) );
  XNOR U1550 ( .A(n1531), .B(n1527), .Z(n1530) );
  XOR U1551 ( .A(n1532), .B(n1533), .Z(n1515) );
  AND U1552 ( .A(n1534), .B(n1535), .Z(n1533) );
  XOR U1553 ( .A(n1522), .B(n1536), .Z(n1535) );
  XNOR U1554 ( .A(n1524), .B(n1532), .Z(n1536) );
  NANDN U1555 ( .B(n978), .A(n1365), .Z(n1524) );
  XOR U1556 ( .A(n1521), .B(n1537), .Z(n1522) );
  AND U1557 ( .A(n910), .B(X[0]), .Z(n1537) );
  XOR U1558 ( .A(n1529), .B(n1541), .Z(n1534) );
  XNOR U1559 ( .A(n1531), .B(n1532), .Z(n1541) );
  NAND U1560 ( .A(n1021), .B(n1128), .Z(n1531) );
  XOR U1561 ( .A(n1527), .B(n1542), .Z(n1529) );
  ANDN U1562 ( .A(n1092), .B(n1055), .Z(n1542) );
  NAND U1563 ( .A(n1021), .B(n1348), .Z(n1545) );
  XNOR U1564 ( .A(n1543), .B(n1547), .Z(n1544) );
  AND U1565 ( .A(n1128), .B(n1092), .Z(n1547) );
  AND U1566 ( .A(n1548), .B(A[0]), .Z(n1543) );
  NANDN U1567 ( .B(n1021), .A(n1549), .Z(n1548) );
  NAND U1568 ( .A(n1348), .B(n1092), .Z(n1549) );
  XNOR U1569 ( .A(n1538), .B(n1553), .Z(n1539) );
  ANDN U1570 ( .A(X[0]), .B(n978), .Z(n1553) );
  XOR U1571 ( .A(n1556), .B(n1554), .Z(n1555) );
  ANDN U1572 ( .A(X[0]), .B(n1055), .Z(n1556) );
  AND U1573 ( .A(n1365), .B(n1128), .Z(n1557) );
  XOR U1574 ( .A(n1561), .B(n1540), .Z(n1552) );
  NANDN U1575 ( .B(n1055), .A(n1365), .Z(n1540) );
  IV U1576 ( .A(n1546), .Z(n1561) );
  NAND U1577 ( .A(n1365), .B(n1348), .Z(n1560) );
  XNOR U1578 ( .A(n1558), .B(n1562), .Z(n1559) );
  AND U1579 ( .A(n1128), .B(X[0]), .Z(n1562) );
  AND U1580 ( .A(n1563), .B(A[0]), .Z(n1558) );
  NANDN U1581 ( .B(n1365), .A(n1564), .Z(n1563) );
  NAND U1582 ( .A(n1348), .B(X[0]), .Z(n1564) );
  XNOR U1583 ( .A(n1566), .B(n1118), .Z(n1108) );
  XNOR U1584 ( .A(n1105), .B(n1106), .Z(n1118) );
  NAND U1585 ( .A(n549), .B(n910), .Z(n1106) );
  XNOR U1586 ( .A(n1104), .B(n1567), .Z(n1105) );
  AND U1587 ( .A(n842), .B(n590), .Z(n1567) );
  XNOR U1588 ( .A(n1571), .B(n1568), .Z(n1570) );
  XNOR U1589 ( .A(n1117), .B(n1107), .Z(n1566) );
  XOR U1590 ( .A(n1572), .B(n1573), .Z(n1107) );
  XNOR U1591 ( .A(n1112), .B(n1575), .Z(n1113) );
  AND U1592 ( .A(n712), .B(n697), .Z(n1575) );
  XNOR U1593 ( .A(n1478), .B(A[8]), .Z(n1477) );
  NOR U1594 ( .A(n1576), .B(n1577), .Z(n1478) );
  XOR U1595 ( .A(n1578), .B(n1579), .Z(n1112) );
  AND U1596 ( .A(n1580), .B(n1581), .Z(n1579) );
  XNOR U1597 ( .A(n1582), .B(n1578), .Z(n1581) );
  XOR U1598 ( .A(n1583), .B(n1114), .Z(n1574) );
  NAND U1599 ( .A(n643), .B(n777), .Z(n1114) );
  IV U1600 ( .A(n1116), .Z(n1583) );
  XNOR U1601 ( .A(n1584), .B(n1585), .Z(n1116) );
  AND U1602 ( .A(n1586), .B(n1587), .Z(n1585) );
  XOR U1603 ( .A(n1580), .B(n1588), .Z(n1587) );
  XNOR U1604 ( .A(n1582), .B(n1584), .Z(n1588) );
  NAND U1605 ( .A(n643), .B(n842), .Z(n1582) );
  XOR U1606 ( .A(n1578), .B(n1589), .Z(n1580) );
  AND U1607 ( .A(n777), .B(n697), .Z(n1589) );
  XOR U1608 ( .A(n1576), .B(A[7]), .Z(n1577) );
  NANDN U1609 ( .B(n1590), .A(n1591), .Z(n1576) );
  XOR U1610 ( .A(n1592), .B(n1593), .Z(n1578) );
  AND U1611 ( .A(n1594), .B(n1595), .Z(n1593) );
  XNOR U1612 ( .A(n1596), .B(n1592), .Z(n1595) );
  XOR U1613 ( .A(n1569), .B(n1597), .Z(n1586) );
  XNOR U1614 ( .A(n1571), .B(n1584), .Z(n1597) );
  NANDN U1615 ( .B(n978), .A(n549), .Z(n1571) );
  XOR U1616 ( .A(n1568), .B(n1598), .Z(n1569) );
  AND U1617 ( .A(n910), .B(n590), .Z(n1598) );
  XNOR U1618 ( .A(n1602), .B(n1599), .Z(n1601) );
  XOR U1619 ( .A(n1603), .B(n1604), .Z(n1584) );
  AND U1620 ( .A(n1605), .B(n1606), .Z(n1604) );
  XOR U1621 ( .A(n1594), .B(n1607), .Z(n1606) );
  XNOR U1622 ( .A(n1596), .B(n1603), .Z(n1607) );
  NAND U1623 ( .A(n643), .B(n910), .Z(n1596) );
  XOR U1624 ( .A(n1592), .B(n1608), .Z(n1594) );
  AND U1625 ( .A(n842), .B(n697), .Z(n1608) );
  XNOR U1626 ( .A(n1591), .B(A[6]), .Z(n1590) );
  NOR U1627 ( .A(n1609), .B(n1610), .Z(n1591) );
  XOR U1628 ( .A(n1611), .B(n1612), .Z(n1592) );
  AND U1629 ( .A(n1613), .B(n1614), .Z(n1612) );
  XNOR U1630 ( .A(n1615), .B(n1611), .Z(n1614) );
  XOR U1631 ( .A(n1600), .B(n1616), .Z(n1605) );
  XNOR U1632 ( .A(n1602), .B(n1603), .Z(n1616) );
  NANDN U1633 ( .B(n1055), .A(n549), .Z(n1602) );
  XOR U1634 ( .A(n1599), .B(n1617), .Z(n1600) );
  ANDN U1635 ( .A(n590), .B(n978), .Z(n1617) );
  XNOR U1636 ( .A(n1621), .B(n1618), .Z(n1620) );
  XOR U1637 ( .A(n1622), .B(n1623), .Z(n1603) );
  AND U1638 ( .A(n1624), .B(n1625), .Z(n1623) );
  XOR U1639 ( .A(n1613), .B(n1626), .Z(n1625) );
  XNOR U1640 ( .A(n1615), .B(n1622), .Z(n1626) );
  NANDN U1641 ( .B(n978), .A(n643), .Z(n1615) );
  XOR U1642 ( .A(n1611), .B(n1627), .Z(n1613) );
  AND U1643 ( .A(n910), .B(n697), .Z(n1627) );
  XOR U1644 ( .A(n1609), .B(A[5]), .Z(n1610) );
  NANDN U1645 ( .B(n1628), .A(n1629), .Z(n1609) );
  XOR U1646 ( .A(n1630), .B(n1631), .Z(n1611) );
  ANDN U1647 ( .A(n1632), .B(n1633), .Z(n1631) );
  XNOR U1648 ( .A(n1634), .B(n1630), .Z(n1632) );
  XOR U1649 ( .A(n1619), .B(n1635), .Z(n1624) );
  XNOR U1650 ( .A(n1621), .B(n1622), .Z(n1635) );
  NAND U1651 ( .A(n549), .B(n1128), .Z(n1621) );
  XOR U1652 ( .A(n1618), .B(n1636), .Z(n1619) );
  ANDN U1653 ( .A(n590), .B(n1055), .Z(n1636) );
  XOR U1654 ( .A(n1637), .B(n1638), .Z(n1618) );
  ANDN U1655 ( .A(n1639), .B(n1640), .Z(n1638) );
  XNOR U1656 ( .A(n1641), .B(n1637), .Z(n1639) );
  NAND U1657 ( .A(n549), .B(n1348), .Z(n1641) );
  XNOR U1658 ( .A(n1637), .B(n1643), .Z(n1640) );
  AND U1659 ( .A(n1128), .B(n590), .Z(n1643) );
  AND U1660 ( .A(n1644), .B(A[0]), .Z(n1637) );
  NANDN U1661 ( .B(n549), .A(n1645), .Z(n1644) );
  NAND U1662 ( .A(n1348), .B(n590), .Z(n1645) );
  XNOR U1663 ( .A(n1630), .B(n1649), .Z(n1633) );
  ANDN U1664 ( .A(n697), .B(n978), .Z(n1649) );
  XOR U1665 ( .A(n1650), .B(n1651), .Z(n1630) );
  AND U1666 ( .A(n1652), .B(n1653), .Z(n1651) );
  XOR U1667 ( .A(n1654), .B(n1650), .Z(n1653) );
  ANDN U1668 ( .A(n697), .B(n1055), .Z(n1654) );
  XOR U1669 ( .A(n1655), .B(n1650), .Z(n1652) );
  AND U1670 ( .A(n1128), .B(n643), .Z(n1655) );
  XOR U1671 ( .A(n1656), .B(n1657), .Z(n1650) );
  ANDN U1672 ( .A(n1658), .B(n1659), .Z(n1657) );
  XNOR U1673 ( .A(n1660), .B(n1656), .Z(n1658) );
  XOR U1674 ( .A(n1661), .B(n1634), .Z(n1648) );
  NANDN U1675 ( .B(n1055), .A(n643), .Z(n1634) );
  IV U1676 ( .A(n1642), .Z(n1661) );
  XOR U1677 ( .A(n1662), .B(n1660), .Z(n1642) );
  NAND U1678 ( .A(n643), .B(n1348), .Z(n1660) );
  IV U1679 ( .A(n1659), .Z(n1662) );
  XNOR U1680 ( .A(n1656), .B(n1663), .Z(n1659) );
  AND U1681 ( .A(n1128), .B(n697), .Z(n1663) );
  AND U1682 ( .A(n1664), .B(A[0]), .Z(n1656) );
  NANDN U1683 ( .B(n643), .A(n1665), .Z(n1664) );
  NAND U1684 ( .A(n1348), .B(n697), .Z(n1665) );
  XNOR U1685 ( .A(n1121), .B(n1669), .Z(n1122) );
  ANDN U1686 ( .A(n517), .B(n978), .Z(n1669) );
  XNOR U1687 ( .A(n1629), .B(A[4]), .Z(n1628) );
  NOR U1688 ( .A(n1670), .B(n1671), .Z(n1629) );
  XOR U1689 ( .A(n1672), .B(n1673), .Z(n1121) );
  AND U1690 ( .A(n1674), .B(n1675), .Z(n1673) );
  XOR U1691 ( .A(n1676), .B(n1672), .Z(n1675) );
  ANDN U1692 ( .A(n517), .B(n1055), .Z(n1676) );
  XOR U1693 ( .A(n1677), .B(n1672), .Z(n1674) );
  AND U1694 ( .A(n1128), .B(n479), .Z(n1677) );
  XOR U1695 ( .A(n1678), .B(n1679), .Z(n1672) );
  ANDN U1696 ( .A(n1680), .B(n1681), .Z(n1679) );
  XNOR U1697 ( .A(n1682), .B(n1678), .Z(n1680) );
  XOR U1698 ( .A(n1683), .B(n1123), .Z(n1668) );
  NANDN U1699 ( .B(n1055), .A(n479), .Z(n1123) );
  NANDN U1700 ( .B(n1684), .A(n1685), .Z(n1670) );
  IV U1701 ( .A(n1125), .Z(n1683) );
  NAND U1702 ( .A(n479), .B(n1348), .Z(n1682) );
  XNOR U1703 ( .A(n1678), .B(n1686), .Z(n1681) );
  AND U1704 ( .A(n1128), .B(n517), .Z(n1686) );
  AND U1705 ( .A(n1687), .B(A[0]), .Z(n1678) );
  NANDN U1706 ( .B(n479), .A(n1688), .Z(n1687) );
  NAND U1707 ( .A(n1348), .B(n517), .Z(n1688) );
  XNOR U1708 ( .A(n1689), .B(X[12]), .Z(n517) );
  NAND U1709 ( .A(n1690), .B(X[15]), .Z(n1689) );
  XOR U1710 ( .A(n1691), .B(X[12]), .Z(n1690) );
  XNOR U1711 ( .A(n1132), .B(n1133), .Z(n1127) );
  NANDN U1712 ( .B(n424), .A(n1348), .Z(n1133) );
  XNOR U1713 ( .A(n1131), .B(n1693), .Z(n1132) );
  AND U1714 ( .A(n1128), .B(n448), .Z(n1693) );
  XNOR U1715 ( .A(n1685), .B(A[2]), .Z(n1684) );
  AND U1716 ( .A(n1695), .B(A[0]), .Z(n1131) );
  NAND U1717 ( .A(n1696), .B(n424), .Z(n1695) );
  NANDN U1718 ( .B(n1697), .A(n1698), .Z(n424) );
  ANDN U1719 ( .A(X[15]), .B(n1699), .Z(n1698) );
  NAND U1720 ( .A(n1348), .B(n448), .Z(n1696) );
  XOR U1721 ( .A(n1699), .B(X[14]), .Z(n1697) );
  OR U1722 ( .A(n1692), .B(n1700), .Z(n1699) );
  XOR U1723 ( .A(n1700), .B(X[13]), .Z(n1692) );
  OR U1724 ( .A(n1691), .B(n1701), .Z(n1700) );
  XOR U1725 ( .A(n1701), .B(X[12]), .Z(n1691) );
  OR U1726 ( .A(n1647), .B(n1702), .Z(n1701) );
  XOR U1727 ( .A(n1702), .B(X[11]), .Z(n1647) );
  OR U1728 ( .A(n1646), .B(n1703), .Z(n1702) );
  XOR U1729 ( .A(n1703), .B(X[10]), .Z(n1646) );
  OR U1730 ( .A(n1667), .B(n1704), .Z(n1703) );
  XOR U1731 ( .A(n1704), .B(X[9]), .Z(n1667) );
  OR U1732 ( .A(n1666), .B(n1705), .Z(n1704) );
  XOR U1733 ( .A(n1705), .B(X[8]), .Z(n1666) );
  OR U1734 ( .A(n1358), .B(n1706), .Z(n1705) );
  XOR U1735 ( .A(n1706), .B(X[7]), .Z(n1358) );
  OR U1736 ( .A(n1357), .B(n1707), .Z(n1706) );
  XOR U1737 ( .A(n1707), .B(X[6]), .Z(n1357) );
  OR U1738 ( .A(n1353), .B(n1708), .Z(n1707) );
  XOR U1739 ( .A(n1708), .B(X[5]), .Z(n1353) );
  OR U1740 ( .A(n1352), .B(n1709), .Z(n1708) );
  XOR U1741 ( .A(n1709), .B(X[4]), .Z(n1352) );
  OR U1742 ( .A(n1551), .B(n1710), .Z(n1709) );
  XOR U1743 ( .A(n1710), .B(X[3]), .Z(n1551) );
  OR U1744 ( .A(n1550), .B(n1711), .Z(n1710) );
  XOR U1745 ( .A(n1711), .B(X[2]), .Z(n1550) );
  NANDN U1746 ( .B(X[0]), .A(n1565), .Z(n1711) );
  XNOR U1747 ( .A(X[0]), .B(X[1]), .Z(n1565) );
  XOR U1748 ( .A(A[0]), .B(A[1]), .Z(n1694) );
  NANDN U1749 ( .B(n1067), .A(n339), .Z(n391) );
  IV U1750 ( .A(rst), .Z(n339) );
  NAND U1751 ( .A(n1712), .B(n1713), .Z(n1067) );
  ANDN U1752 ( .A(n1714), .B(n[2]), .Z(n1713) );
  NOR U1753 ( .A(n[6]), .B(n[5]), .Z(n1714) );
  ANDN U1754 ( .A(n1715), .B(n333), .Z(n1712) );
  OR U1755 ( .A(n[4]), .B(n[3]), .Z(n333) );
  NOR U1756 ( .A(n[0]), .B(n[1]), .Z(n1715) );
endmodule

