
module MxM_TG_W16_N100 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MxM/n91 , \_MxM/n88 , \_MxM/n85 , \_MxM/n82 , \_MxM/n79 ,
         \_MxM/n76 , \_MxM/n73 , \_MxM/n70 , \_MxM/n67 , \_MxM/n64 ,
         \_MxM/n61 , \_MxM/n58 , \_MxM/n55 , \_MxM/n52 , \_MxM/n49 ,
         \_MxM/n46 , \_MxM/N17 , \_MxM/N16 , \_MxM/N15 , \_MxM/N14 ,
         \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N9 , \_MxM/N8 , \_MxM/N7 ,
         \_MxM/N6 , \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] ,
         \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/Y1[0] ,
         \_MxM/Y1[1] , \_MxM/Y1[2] , \_MxM/Y1[3] , \_MxM/Y1[4] , \_MxM/Y1[5] ,
         \_MxM/Y1[6] , \_MxM/Y1[7] , \_MxM/Y1[8] , \_MxM/Y1[9] , \_MxM/Y1[10] ,
         \_MxM/Y1[11] , \_MxM/Y1[12] , \_MxM/Y1[13] , \_MxM/Y1[14] ,
         \_MxM/Y1[15] , \_MxM/Y0[15] , \_MxM/Y0[14] , \_MxM/Y0[13] ,
         \_MxM/Y0[12] , \_MxM/Y0[11] , \_MxM/Y0[10] , \_MxM/Y0[9] ,
         \_MxM/Y0[8] , \_MxM/Y0[7] , \_MxM/Y0[6] , \_MxM/Y0[5] , \_MxM/Y0[4] ,
         \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] , \_MxM/Y0[0] ,
         \_MxM/add_43/carry[6] , \_MxM/add_43/carry[5] ,
         \_MxM/add_43/carry[4] , \_MxM/add_43/carry[3] ,
         \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374;

  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n46 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/Y1[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n49 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/Y1[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n52 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/Y1[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n55 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/Y1[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n58 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/Y1[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n61 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/Y1[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n64 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/Y1[9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n67 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/Y1[8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n70 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n73 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n76 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n79 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n82 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n85 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n88 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n91 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N14 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N13 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N12 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N11 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  MUX U1 ( .IN0(n1), .IN1(n1296), .SEL(n1297), .F(n1277) );
  IV U2 ( .A(n1298), .Z(n1) );
  MUX U3 ( .IN0(n2), .IN1(n841), .SEL(n842), .F(n820) );
  IV U4 ( .A(n843), .Z(n2) );
  XOR U5 ( .A(n1061), .B(n1051), .Z(n861) );
  MUX U6 ( .IN0(n995), .IN1(n998), .SEL(n996), .F(n980) );
  XOR U7 ( .A(n1033), .B(n1034), .Z(n836) );
  MUX U8 ( .IN0(n3), .IN1(n556), .SEL(n557), .F(n495) );
  IV U9 ( .A(n558), .Z(n3) );
  MUX U10 ( .IN0(e_input[12]), .IN1(n1348), .SEL(e_input[15]), .F(n223) );
  MUX U11 ( .IN0(n1277), .IN1(n1295), .SEL(n1279), .F(n1257) );
  XOR U12 ( .A(n1043), .B(n1044), .Z(n859) );
  MUX U13 ( .IN0(n4), .IN1(n801), .SEL(n802), .F(n734) );
  IV U14 ( .A(n803), .Z(n4) );
  XOR U15 ( .A(n844), .B(n826), .Z(n830) );
  MUX U16 ( .IN0(n1038), .IN1(n5), .SEL(n1037), .F(n1027) );
  IV U17 ( .A(n1036), .Z(n5) );
  MUX U18 ( .IN0(e_input[8]), .IN1(n1324), .SEL(e_input[15]), .F(n382) );
  XNOR U19 ( .A(n1326), .B(n776), .Z(n780) );
  MUX U20 ( .IN0(n6), .IN1(n1082), .SEL(n1083), .F(n1065) );
  IV U21 ( .A(n1084), .Z(n6) );
  MUX U22 ( .IN0(n1226), .IN1(n1256), .SEL(n1228), .F(n754) );
  XOR U23 ( .A(n802), .B(n803), .Z(n799) );
  MUX U24 ( .IN0(n7), .IN1(n1032), .SEL(n1033), .F(n808) );
  IV U25 ( .A(n1034), .Z(n7) );
  MUX U26 ( .IN0(n8), .IN1(n437), .SEL(n438), .F(n383) );
  IV U27 ( .A(n439), .Z(n8) );
  MUX U28 ( .IN0(n598), .IN1(n9), .SEL(n597), .F(n533) );
  IV U29 ( .A(n596), .Z(n9) );
  MUX U30 ( .IN0(e_input[13]), .IN1(n1349), .SEL(e_input[15]), .F(n188) );
  MUX U31 ( .IN0(n10), .IN1(n1042), .SEL(n1043), .F(n1032) );
  IV U32 ( .A(n1044), .Z(n10) );
  MUX U33 ( .IN0(n11), .IN1(n1050), .SEL(n1051), .F(n1036) );
  IV U34 ( .A(n1052), .Z(n11) );
  MUX U35 ( .IN0(n12), .IN1(n734), .SEL(n735), .F(n664) );
  IV U36 ( .A(n736), .Z(n12) );
  MUX U37 ( .IN0(n13), .IN1(n726), .SEL(n727), .F(n656) );
  IV U38 ( .A(n728), .Z(n13) );
  MUX U39 ( .IN0(n14), .IN1(n548), .SEL(n549), .F(n487) );
  IV U40 ( .A(n550), .Z(n14) );
  MUX U41 ( .IN0(e_input[9]), .IN1(n1325), .SEL(e_input[15]), .F(n335) );
  MUX U42 ( .IN0(n573), .IN1(n571), .SEL(n572), .F(n510) );
  MUX U43 ( .IN0(n226), .IN1(n15), .SEL(n225), .F(n190) );
  IV U44 ( .A(n224), .Z(n15) );
  MUX U45 ( .IN0(n16), .IN1(n1194), .SEL(n1195), .F(n1177) );
  IV U46 ( .A(n1196), .Z(n16) );
  XOR U47 ( .A(n821), .B(n822), .Z(n831) );
  MUX U48 ( .IN0(n17), .IN1(n754), .SEL(n755), .F(n685) );
  IV U49 ( .A(n756), .Z(n17) );
  MUX U50 ( .IN0(n18), .IN1(n693), .SEL(n694), .F(n619) );
  IV U51 ( .A(n695), .Z(n18) );
  MUX U52 ( .IN0(n19), .IN1(n656), .SEL(n657), .F(n596) );
  IV U53 ( .A(n658), .Z(n19) );
  MUX U54 ( .IN0(g_input[11]), .IN1(n1081), .SEL(g_input[15]), .F(n267) );
  XOR U55 ( .A(n745), .B(n746), .Z(n751) );
  MUX U56 ( .IN0(n499), .IN1(n501), .SEL(n500), .F(n441) );
  MUX U57 ( .IN0(n536), .IN1(n20), .SEL(n535), .F(n470) );
  IV U58 ( .A(n534), .Z(n20) );
  XNOR U59 ( .A(n771), .B(n705), .Z(n709) );
  XOR U60 ( .A(n842), .B(n843), .Z(n854) );
  MUX U61 ( .IN0(g_input[1]), .IN1(n1351), .SEL(g_input[15]), .F(n1005) );
  XOR U62 ( .A(n1035), .B(n1027), .Z(n817) );
  MUX U63 ( .IN0(g_input[2]), .IN1(n1342), .SEL(g_input[15]), .F(n782) );
  MUX U64 ( .IN0(n21), .IN1(n611), .SEL(n612), .F(n548) );
  IV U65 ( .A(n613), .Z(n21) );
  MUX U66 ( .IN0(n22), .IN1(n495), .SEL(n496), .F(n437) );
  IV U67 ( .A(n497), .Z(n22) );
  MUX U68 ( .IN0(g_input[10]), .IN1(n1097), .SEL(g_input[15]), .F(n307) );
  MUX U69 ( .IN0(n746), .IN1(n23), .SEL(n745), .F(n674) );
  IV U70 ( .A(n744), .Z(n23) );
  MUX U71 ( .IN0(n454), .IN1(n452), .SEL(n453), .F(n394) );
  MUX U72 ( .IN0(n377), .IN1(n379), .SEL(n378), .F(n24) );
  IV U73 ( .A(n24), .Z(n338) );
  XNOR U74 ( .A(n724), .B(n657), .Z(n661) );
  XNOR U75 ( .A(n700), .B(n633), .Z(n637) );
  MUX U76 ( .IN0(n1212), .IN1(n1215), .SEL(n1213), .F(n1194) );
  XOR U77 ( .A(n1297), .B(n1298), .Z(n1230) );
  XOR U78 ( .A(n809), .B(n810), .Z(n815) );
  MUX U79 ( .IN0(n25), .IN1(n664), .SEL(n665), .F(n600) );
  IV U80 ( .A(n666), .Z(n25) );
  MUX U81 ( .IN0(g_input[9]), .IN1(n1117), .SEL(g_input[15]), .F(n350) );
  XNOR U82 ( .A(n789), .B(n727), .Z(n731) );
  MUX U83 ( .IN0(n441), .IN1(n443), .SEL(n442), .F(n377) );
  MUX U84 ( .IN0(n396), .IN1(n394), .SEL(n395), .F(n347) );
  MUX U85 ( .IN0(n385), .IN1(n26), .SEL(n384), .F(n337) );
  IV U86 ( .A(n383), .Z(n26) );
  XNOR U87 ( .A(n628), .B(n568), .Z(n572) );
  NAND U88 ( .A(n533), .B(n594), .Z(n593) );
  MUX U89 ( .IN0(n27), .IN1(n989), .SEL(n805), .F(n962) );
  IV U90 ( .A(n804), .Z(n27) );
  MUX U91 ( .IN0(n1160), .IN1(n1176), .SEL(n1162), .F(n1149) );
  MUX U92 ( .IN0(n28), .IN1(n808), .SEL(n809), .F(n744) );
  IV U93 ( .A(n810), .Z(n28) );
  MUX U94 ( .IN0(n29), .IN1(n600), .SEL(n601), .F(n538) );
  IV U95 ( .A(n602), .Z(n29) );
  XOR U96 ( .A(n714), .B(n783), .Z(n715) );
  MUX U97 ( .IN0(n349), .IN1(n347), .SEL(n348), .F(n304) );
  MUX U98 ( .IN0(e_input[10]), .IN1(n1303), .SEL(e_input[15]), .F(n286) );
  XOR U99 ( .A(n589), .B(n534), .Z(n535) );
  XNOR U100 ( .A(n563), .B(n507), .Z(n511) );
  XOR U101 ( .A(n435), .B(n384), .Z(n378) );
  MUX U102 ( .IN0(n424), .IN1(n426), .SEL(n425), .F(n30) );
  IV U103 ( .A(n30), .Z(n365) );
  XOR U104 ( .A(n580), .B(n583), .Z(n581) );
  MUX U105 ( .IN0(n932), .IN1(n31), .SEL(n933), .F(n905) );
  IV U106 ( .A(n934), .Z(n31) );
  MUX U107 ( .IN0(n32), .IN1(n1065), .SEL(n1066), .F(n1050) );
  IV U108 ( .A(n1067), .Z(n32) );
  XOR U109 ( .A(n1128), .B(n1129), .Z(n991) );
  MUX U110 ( .IN0(n625), .IN1(n627), .SEL(n626), .F(n560) );
  XOR U111 ( .A(n458), .B(n514), .Z(n459) );
  MUX U112 ( .IN0(e_input[6]), .IN1(n1014), .SEL(e_input[15]), .F(n475) );
  MUX U113 ( .IN0(n33), .IN1(n326), .SEL(n327), .F(n287) );
  IV U114 ( .A(n328), .Z(n33) );
  XNOR U115 ( .A(n654), .B(n597), .Z(n591) );
  MUX U116 ( .IN0(n34), .IN1(n551), .SEL(n552), .F(n490) );
  IV U117 ( .A(n553), .Z(n34) );
  XNOR U118 ( .A(n502), .B(n449), .Z(n453) );
  NAND U119 ( .A(n337), .B(n381), .Z(n380) );
  XOR U120 ( .A(n519), .B(n522), .Z(n520) );
  MUX U121 ( .IN0(n35), .IN1(n1118), .SEL(n1119), .F(n1099) );
  IV U122 ( .A(n1120), .Z(n35) );
  MUX U123 ( .IN0(n36), .IN1(n1016), .SEL(n1017), .F(n1188) );
  IV U124 ( .A(n1204), .Z(n36) );
  MUX U125 ( .IN0(n1143), .IN1(n1165), .SEL(n1145), .F(n1125) );
  XOR U126 ( .A(n823), .B(n794), .Z(n798) );
  MUX U127 ( .IN0(g_input[3]), .IN1(n1329), .SEL(g_input[15]), .F(n37) );
  IV U128 ( .A(n37), .Z(n711) );
  MUX U129 ( .IN0(n38), .IN1(n685), .SEL(n686), .F(n611) );
  IV U130 ( .A(n687), .Z(n38) );
  MUX U131 ( .IN0(n781), .IN1(n779), .SEL(n780), .F(n708) );
  XOR U132 ( .A(n577), .B(n640), .Z(n578) );
  MUX U133 ( .IN0(n560), .IN1(n562), .SEL(n561), .F(n499) );
  MUX U134 ( .IN0(n266), .IN1(n264), .SEL(n265), .F(n216) );
  MUX U135 ( .IN0(g_input[12]), .IN1(n1063), .SEL(g_input[15]), .F(n227) );
  XOR U136 ( .A(n477), .B(n478), .Z(n472) );
  MUX U137 ( .IN0(n39), .IN1(n432), .SEL(n433), .F(n373) );
  IV U138 ( .A(n434), .Z(n39) );
  XNOR U139 ( .A(n444), .B(n391), .Z(n395) );
  XNOR U140 ( .A(n293), .B(n332), .Z(n294) );
  MUX U141 ( .IN0(n667), .IN1(n40), .SEL(n668), .F(n603) );
  IV U142 ( .A(n669), .Z(n40) );
  MUX U143 ( .IN0(n41), .IN1(n313), .SEL(n107), .F(n273) );
  IV U144 ( .A(\_MxM/Y0[8] ), .Z(n41) );
  XOR U145 ( .A(n461), .B(n464), .Z(n462) );
  MUX U146 ( .IN0(n1086), .IN1(n42), .SEL(n914), .F(n1069) );
  IV U147 ( .A(n912), .Z(n42) );
  MUX U148 ( .IN0(e_input[1]), .IN1(n43), .SEL(e_input[15]), .F(n1022) );
  IV U149 ( .A(n1223), .Z(n43) );
  MUX U150 ( .IN0(n829), .IN1(n44), .SEL(n830), .F(n797) );
  IV U151 ( .A(n831), .Z(n44) );
  XNOR U152 ( .A(n1002), .B(n1003), .Z(n986) );
  MUX U153 ( .IN0(n768), .IN1(n770), .SEL(n769), .F(n697) );
  MUX U154 ( .IN0(e_input[2]), .IN1(n1208), .SEL(e_input[15]), .F(n743) );
  MUX U155 ( .IN0(n512), .IN1(n510), .SEL(n511), .F(n452) );
  XOR U156 ( .A(n353), .B(n398), .Z(n354) );
  MUX U157 ( .IN0(n45), .IN1(n747), .SEL(n748), .F(n680) );
  IV U158 ( .A(n749), .Z(n45) );
  MUX U159 ( .IN0(n46), .IN1(n688), .SEL(n689), .F(n614) );
  IV U160 ( .A(n690), .Z(n46) );
  XOR U161 ( .A(n554), .B(n496), .Z(n500) );
  MUX U162 ( .IN0(n47), .IN1(n476), .SEL(n477), .F(n423) );
  IV U163 ( .A(n478), .Z(n47) );
  MUX U164 ( .IN0(n48), .IN1(n373), .SEL(n374), .F(n329) );
  IV U165 ( .A(n375), .Z(n48) );
  NAND U166 ( .A(n247), .B(n285), .Z(n284) );
  XNOR U167 ( .A(n296), .B(n261), .Z(n265) );
  MUX U168 ( .IN0(n49), .IN1(n545), .SEL(n544), .F(n482) );
  IV U169 ( .A(n543), .Z(n49) );
  MUX U170 ( .IN0(n50), .IN1(n199), .SEL(n200), .F(n169) );
  IV U171 ( .A(\_MxM/Y0[11] ), .Z(n50) );
  XOR U172 ( .A(n403), .B(n406), .Z(n404) );
  MUX U173 ( .IN0(n959), .IN1(n51), .SEL(n960), .F(n932) );
  IV U174 ( .A(n961), .Z(n51) );
  MUX U175 ( .IN0(n1122), .IN1(n52), .SEL(n968), .F(n1105) );
  IV U176 ( .A(n966), .Z(n52) );
  MUX U177 ( .IN0(n852), .IN1(n53), .SEL(n853), .F(n829) );
  IV U178 ( .A(n854), .Z(n53) );
  MUX U179 ( .IN0(n1054), .IN1(n54), .SEL(n861), .F(n1040) );
  IV U180 ( .A(n859), .Z(n54) );
  XOR U181 ( .A(n1210), .B(n1195), .Z(n1017) );
  MUX U182 ( .IN0(e_input[4]), .IN1(n1009), .SEL(e_input[15]), .F(n595) );
  XOR U183 ( .A(n1232), .B(n765), .Z(n769) );
  MUX U184 ( .IN0(n662), .IN1(n660), .SEL(n661), .F(n590) );
  MUX U185 ( .IN0(n55), .IN1(n538), .SEL(n539), .F(n476) );
  IV U186 ( .A(n540), .Z(n55) );
  MUX U187 ( .IN0(e_input[11]), .IN1(n1304), .SEL(e_input[15]), .F(n250) );
  MUX U188 ( .IN0(n56), .IN1(n614), .SEL(n615), .F(n551) );
  IV U189 ( .A(n616), .Z(n56) );
  XNOR U190 ( .A(n256), .B(n225), .Z(n219) );
  MUX U191 ( .IN0(n57), .IN1(n253), .SEL(n254), .F(n211) );
  IV U192 ( .A(n255), .Z(n57) );
  MUX U193 ( .IN0(e_input[14]), .IN1(n1354), .SEL(e_input[15]), .F(n158) );
  XNOR U194 ( .A(n606), .B(n670), .Z(n607) );
  MUX U195 ( .IN0(n482), .IN1(n484), .SEL(n483), .F(n424) );
  MUX U196 ( .IN0(n58), .IN1(n645), .SEL(n113), .F(n580) );
  IV U197 ( .A(\_MxM/Y0[2] ), .Z(n58) );
  XNOR U198 ( .A(n169), .B(n170), .Z(n127) );
  XOR U199 ( .A(n357), .B(n363), .Z(n108) );
  MUX U200 ( .IN0(n1105), .IN1(n59), .SEL(n941), .F(n1086) );
  IV U201 ( .A(n939), .Z(n59) );
  MUX U202 ( .IN0(n60), .IN1(n1216), .SEL(n1217), .F(n1212) );
  IV U203 ( .A(n1218), .Z(n60) );
  MUX U204 ( .IN0(n1040), .IN1(n61), .SEL(n838), .F(n1028) );
  IV U205 ( .A(n836), .Z(n61) );
  MUX U206 ( .IN0(n797), .IN1(n62), .SEL(n798), .F(n730) );
  IV U207 ( .A(n799), .Z(n62) );
  XNOR U208 ( .A(n993), .B(n983), .Z(n987) );
  MUX U209 ( .IN0(g_input[5]), .IN1(n1269), .SEL(g_input[15]), .F(n574) );
  MUX U210 ( .IN0(n710), .IN1(n708), .SEL(n709), .F(n636) );
  MUX U211 ( .IN0(n340), .IN1(n63), .SEL(n339), .F(n293) );
  IV U212 ( .A(n338), .Z(n63) );
  XOR U213 ( .A(n270), .B(n308), .Z(n271) );
  MUX U214 ( .IN0(n64), .IN1(n757), .SEL(n758), .F(n688) );
  IV U215 ( .A(n759), .Z(n64) );
  NAND U216 ( .A(n674), .B(n742), .Z(n741) );
  XOR U217 ( .A(n691), .B(n622), .Z(n626) );
  XOR U218 ( .A(n539), .B(n540), .Z(n536) );
  MUX U219 ( .IN0(n65), .IN1(n490), .SEL(n491), .F(n432) );
  IV U220 ( .A(n492), .Z(n65) );
  XNOR U221 ( .A(n386), .B(n344), .Z(n348) );
  MUX U222 ( .IN0(n66), .IN1(n290), .SEL(n291), .F(n253) );
  IV U223 ( .A(n292), .Z(n66) );
  MUX U224 ( .IN0(n289), .IN1(n67), .SEL(n288), .F(n247) );
  IV U225 ( .A(n287), .Z(n67) );
  XNOR U226 ( .A(n216), .B(n217), .Z(n215) );
  XNOR U227 ( .A(n592), .B(n591), .Z(n608) );
  XNOR U228 ( .A(n220), .B(n219), .Z(n213) );
  XOR U229 ( .A(n469), .B(n417), .Z(n425) );
  MUX U230 ( .IN0(n68), .IN1(n519), .SEL(n111), .F(n461) );
  IV U231 ( .A(\_MxM/Y0[4] ), .Z(n68) );
  MUX U232 ( .IN0(\_MxM/Y0[13] ), .IN1(n127), .SEL(n126), .F(n123) );
  XOR U233 ( .A(n273), .B(n276), .Z(n274) );
  XOR U234 ( .A(n1147), .B(n1138), .Z(n992) );
  MUX U235 ( .IN0(n69), .IN1(n429), .SEL(n430), .F(n370) );
  IV U236 ( .A(n431), .Z(n69) );
  MUX U237 ( .IN0(e_input[3]), .IN1(n1209), .SEL(e_input[15]), .F(n677) );
  MUX U238 ( .IN0(n638), .IN1(n636), .SEL(n637), .F(n571) );
  MUX U239 ( .IN0(e_input[5]), .IN1(n1010), .SEL(e_input[15]), .F(n531) );
  MUX U240 ( .IN0(n306), .IN1(n304), .SEL(n305), .F(n264) );
  XOR U241 ( .A(n760), .B(n694), .Z(n698) );
  XNOR U242 ( .A(n781), .B(n780), .Z(n759) );
  MUX U243 ( .IN0(n682), .IN1(n70), .SEL(n681), .F(n606) );
  IV U244 ( .A(n680), .Z(n70) );
  MUX U245 ( .IN0(e_input[7]), .IN1(n1015), .SEL(e_input[15]), .F(n415) );
  MUX U246 ( .IN0(n295), .IN1(n293), .SEL(n294), .F(n71) );
  IV U247 ( .A(n71), .Z(n252) );
  NAND U248 ( .A(n190), .B(n222), .Z(n221) );
  XOR U249 ( .A(n196), .B(n228), .Z(n197) );
  MUX U250 ( .IN0(n603), .IN1(n72), .SEL(n604), .F(n543) );
  IV U251 ( .A(n605), .Z(n72) );
  XNOR U252 ( .A(n396), .B(n395), .Z(n375) );
  MUX U253 ( .IN0(n213), .IN1(n73), .SEL(n212), .F(n184) );
  IV U254 ( .A(n211), .Z(n73) );
  XNOR U255 ( .A(n492), .B(n491), .Z(n484) );
  MUX U256 ( .IN0(n74), .IN1(n461), .SEL(n110), .F(n403) );
  IV U257 ( .A(\_MxM/Y0[5] ), .Z(n74) );
  MUX U258 ( .IN0(n75), .IN1(n273), .SEL(n106), .F(n233) );
  IV U259 ( .A(\_MxM/Y0[9] ), .Z(n75) );
  MUX U260 ( .IN0(n76), .IN1(n121), .SEL(n120), .F(n125) );
  IV U261 ( .A(n128), .Z(n76) );
  MUX U262 ( .IN0(n905), .IN1(n77), .SEL(n906), .F(n878) );
  IV U263 ( .A(n907), .Z(n77) );
  MUX U264 ( .IN0(n1184), .IN1(n1198), .SEL(n1186), .F(n1166) );
  XNOR U265 ( .A(n1217), .B(n1218), .Z(n1204) );
  XOR U266 ( .A(n1328), .B(g_input[3]), .Z(n1329) );
  MUX U267 ( .IN0(g_input[6]), .IN1(n1248), .SEL(g_input[15]), .F(n513) );
  MUX U268 ( .IN0(n78), .IN1(n487), .SEL(n488), .F(n429) );
  IV U269 ( .A(n489), .Z(n78) );
  MUX U270 ( .IN0(g_input[7]), .IN1(n1235), .SEL(g_input[15]), .F(n455) );
  MUX U271 ( .IN0(g_input[8]), .IN1(n1133), .SEL(g_input[15]), .F(n397) );
  XNOR U272 ( .A(n1028), .B(n1029), .Z(n1018) );
  XNOR U273 ( .A(n988), .B(n987), .Z(n804) );
  MUX U274 ( .IN0(n592), .IN1(n590), .SEL(n591), .F(n534) );
  XNOR U275 ( .A(n732), .B(n731), .Z(n749) );
  XOR U276 ( .A(n617), .B(n557), .Z(n561) );
  MUX U277 ( .IN0(n79), .IN1(n329), .SEL(n330), .F(n290) );
  IV U278 ( .A(n331), .Z(n79) );
  XNOR U279 ( .A(n341), .B(n301), .Z(n305) );
  MUX U280 ( .IN0(g_input[13]), .IN1(n1049), .SEL(g_input[15]), .F(n193) );
  XNOR U281 ( .A(n662), .B(n661), .Z(n682) );
  XNOR U282 ( .A(n759), .B(n758), .Z(n739) );
  XNOR U283 ( .A(n638), .B(n637), .Z(n616) );
  XNOR U284 ( .A(n573), .B(n572), .Z(n553) );
  AND U285 ( .A(n153), .B(n134), .Z(n152) );
  XNOR U286 ( .A(n690), .B(n689), .Z(n669) );
  XNOR U287 ( .A(n482), .B(n481), .Z(n527) );
  MUX U288 ( .IN0(n80), .IN1(n580), .SEL(n112), .F(n519) );
  IV U289 ( .A(\_MxM/Y0[3] ), .Z(n80) );
  XNOR U290 ( .A(n434), .B(n433), .Z(n426) );
  XNOR U291 ( .A(n375), .B(n374), .Z(n367) );
  MUX U292 ( .IN0(n81), .IN1(n356), .SEL(n108), .F(n313) );
  IV U293 ( .A(\_MxM/Y0[7] ), .Z(n81) );
  XNOR U294 ( .A(n183), .B(n184), .Z(n182) );
  XOR U295 ( .A(n233), .B(n236), .Z(n234) );
  MUX U296 ( .IN0(\_MxM/Y0[14] ), .IN1(n123), .SEL(n124), .F(n117) );
  MUX U297 ( .IN0(n988), .IN1(n986), .SEL(n987), .F(n959) );
  MUX U298 ( .IN0(n1141), .IN1(n82), .SEL(n992), .F(n1122) );
  IV U299 ( .A(n991), .Z(n82) );
  MUX U300 ( .IN0(n83), .IN1(n1230), .SEL(n1231), .F(n1281) );
  IV U301 ( .A(n1299), .Z(n83) );
  MUX U302 ( .IN0(n878), .IN1(n84), .SEL(n879), .F(n852) );
  IV U303 ( .A(n880), .Z(n84) );
  NOR U304 ( .A(g_input[0]), .B(n1351), .Z(n1343) );
  MUX U305 ( .IN0(n1069), .IN1(n85), .SEL(n887), .F(n1054) );
  IV U306 ( .A(n885), .Z(n85) );
  MUX U307 ( .IN0(n86), .IN1(n820), .SEL(n821), .F(n801) );
  IV U308 ( .A(n822), .Z(n86) );
  MUX U309 ( .IN0(n87), .IN1(n825), .SEL(n826), .F(n791) );
  IV U310 ( .A(n827), .Z(n87) );
  MUX U311 ( .IN0(n1149), .IN1(n1159), .SEL(n1151), .F(n1135) );
  XOR U312 ( .A(n1202), .B(n1203), .Z(n1016) );
  MUX U313 ( .IN0(g_input[4]), .IN1(n1287), .SEL(g_input[15]), .F(n88) );
  IV U314 ( .A(n88), .Z(n639) );
  MUX U315 ( .IN0(n89), .IN1(n343), .SEL(n344), .F(n298) );
  IV U316 ( .A(n345), .Z(n89) );
  MUX U317 ( .IN0(n90), .IN1(n370), .SEL(n371), .F(n326) );
  IV U318 ( .A(n372), .Z(n90) );
  MUX U319 ( .IN0(n732), .IN1(n730), .SEL(n731), .F(n660) );
  MUX U320 ( .IN0(n697), .IN1(n699), .SEL(n698), .F(n625) );
  MUX U321 ( .IN0(n751), .IN1(n1018), .SEL(n750), .F(n679) );
  XOR U322 ( .A(n493), .B(n438), .Z(n442) );
  MUX U323 ( .IN0(n472), .IN1(n470), .SEL(n471), .F(n421) );
  XNOR U324 ( .A(n710), .B(n709), .Z(n690) );
  MUX U325 ( .IN0(n737), .IN1(n91), .SEL(n738), .F(n667) );
  IV U326 ( .A(n739), .Z(n91) );
  MUX U327 ( .IN0(n608), .IN1(n606), .SEL(n607), .F(n92) );
  IV U328 ( .A(n92), .Z(n542) );
  XNOR U329 ( .A(n512), .B(n511), .Z(n492) );
  XNOR U330 ( .A(n454), .B(n453), .Z(n434) );
  XNOR U331 ( .A(n349), .B(n348), .Z(n331) );
  XNOR U332 ( .A(n306), .B(n305), .Z(n292) );
  XNOR U333 ( .A(n266), .B(n265), .Z(n255) );
  MUX U334 ( .IN0(n192), .IN1(n215), .SEL(n191), .F(n164) );
  MUX U335 ( .IN0(g_input[14]), .IN1(n1023), .SEL(g_input[15]), .F(n159) );
  XNOR U336 ( .A(n616), .B(n615), .Z(n605) );
  XNOR U337 ( .A(n553), .B(n552), .Z(n545) );
  MUX U338 ( .IN0(n365), .IN1(n93), .SEL(n366), .F(n323) );
  IV U339 ( .A(n367), .Z(n93) );
  MUX U340 ( .IN0(n94), .IN1(n403), .SEL(n109), .F(n356) );
  IV U341 ( .A(\_MxM/Y0[6] ), .Z(n94) );
  MUX U342 ( .IN0(n95), .IN1(n233), .SEL(n105), .F(n199) );
  IV U343 ( .A(\_MxM/Y0[10] ), .Z(n95) );
  MUX U344 ( .IN0(n96), .IN1(n717), .SEL(n718), .F(n645) );
  IV U345 ( .A(\_MxM/Y0[1] ), .Z(n96) );
  XNOR U346 ( .A(n182), .B(n181), .Z(n203) );
  MUX U347 ( .IN0(\_MxM/Y0[15] ), .IN1(n117), .SEL(n118), .F(n97) );
  IV U348 ( .A(n97), .Z(n114) );
  MUX U349 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n98), .F(\_MxM/n91 ) );
  MUX U350 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n98), .F(\_MxM/n88 ) );
  MUX U351 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n98), .F(\_MxM/n85 ) );
  MUX U352 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n98), .F(\_MxM/n82 ) );
  MUX U353 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n98), .F(\_MxM/n79 ) );
  MUX U354 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n98), .F(\_MxM/n76 ) );
  MUX U355 ( .IN0(\_MxM/Y1[6] ), .IN1(o[6]), .SEL(n98), .F(\_MxM/n73 ) );
  MUX U356 ( .IN0(\_MxM/Y1[7] ), .IN1(o[7]), .SEL(n98), .F(\_MxM/n70 ) );
  MUX U357 ( .IN0(\_MxM/Y1[8] ), .IN1(o[8]), .SEL(n98), .F(\_MxM/n67 ) );
  MUX U358 ( .IN0(\_MxM/Y1[9] ), .IN1(o[9]), .SEL(n98), .F(\_MxM/n64 ) );
  MUX U359 ( .IN0(\_MxM/Y1[10] ), .IN1(o[10]), .SEL(n98), .F(\_MxM/n61 ) );
  MUX U360 ( .IN0(\_MxM/Y1[11] ), .IN1(o[11]), .SEL(n98), .F(\_MxM/n58 ) );
  MUX U361 ( .IN0(\_MxM/Y1[12] ), .IN1(o[12]), .SEL(n98), .F(\_MxM/n55 ) );
  MUX U362 ( .IN0(\_MxM/Y1[13] ), .IN1(o[13]), .SEL(n98), .F(\_MxM/n52 ) );
  IV U363 ( .A(n99), .Z(n98) );
  MUX U364 ( .IN0(o[14]), .IN1(\_MxM/Y1[14] ), .SEL(n99), .F(\_MxM/n49 ) );
  MUX U365 ( .IN0(o[15]), .IN1(\_MxM/Y1[15] ), .SEL(n99), .F(\_MxM/n46 ) );
  AND U366 ( .A(n100), .B(n101), .Z(n99) );
  ANDN U367 ( .A(n102), .B(\_MxM/n[2] ), .Z(n101) );
  NOR U368 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n102) );
  ANDN U369 ( .A(n103), .B(n104), .Z(n100) );
  ANDN U370 ( .A(\_MxM/N11 ), .B(\_MxM/n[1] ), .Z(n103) );
  XNOR U371 ( .A(n105), .B(\_MxM/Y0[10] ), .Z(\_MxM/Y1[9] ) );
  XNOR U372 ( .A(n106), .B(\_MxM/Y0[9] ), .Z(\_MxM/Y1[8] ) );
  XNOR U373 ( .A(n107), .B(\_MxM/Y0[8] ), .Z(\_MxM/Y1[7] ) );
  XNOR U374 ( .A(n108), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XNOR U375 ( .A(n109), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XNOR U376 ( .A(n110), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U377 ( .A(n111), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U378 ( .A(n112), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U379 ( .A(n113), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U380 ( .A(n114), .B(n115), .Z(\_MxM/Y1[15] ) );
  XNOR U381 ( .A(\_MxM/Y0[15] ), .B(n116), .Z(n115) );
  XNOR U382 ( .A(n118), .B(\_MxM/Y0[15] ), .Z(\_MxM/Y1[14] ) );
  XOR U383 ( .A(n117), .B(n116), .Z(n118) );
  NAND U384 ( .A(n119), .B(n120), .Z(n116) );
  OR U385 ( .A(n121), .B(n122), .Z(n119) );
  XNOR U386 ( .A(n124), .B(\_MxM/Y0[14] ), .Z(\_MxM/Y1[13] ) );
  XNOR U387 ( .A(n125), .B(n123), .Z(n124) );
  XNOR U388 ( .A(n122), .B(n128), .Z(n121) );
  OR U389 ( .A(n129), .B(n130), .Z(n122) );
  AND U390 ( .A(n131), .B(n132), .Z(n128) );
  OR U391 ( .A(n133), .B(n134), .Z(n132) );
  AND U392 ( .A(n135), .B(n136), .Z(n131) );
  OR U393 ( .A(n137), .B(n138), .Z(n136) );
  OR U394 ( .A(n139), .B(n140), .Z(n135) );
  XNOR U395 ( .A(n126), .B(\_MxM/Y0[13] ), .Z(\_MxM/Y1[12] ) );
  XNOR U396 ( .A(n141), .B(n142), .Z(n126) );
  XNOR U397 ( .A(n127), .B(n143), .Z(n141) );
  AND U398 ( .A(n120), .B(n144), .Z(n143) );
  XOR U399 ( .A(n129), .B(n145), .Z(n144) );
  XOR U400 ( .A(n145), .B(n130), .Z(n129) );
  OR U401 ( .A(n146), .B(n147), .Z(n130) );
  IV U402 ( .A(n142), .Z(n145) );
  XNOR U403 ( .A(n140), .B(n139), .Z(n142) );
  OR U404 ( .A(n148), .B(n149), .Z(n139) );
  AND U405 ( .A(n150), .B(n151), .Z(n140) );
  XNOR U406 ( .A(n133), .B(n152), .Z(n151) );
  NAND U407 ( .A(n154), .B(n155), .Z(n134) );
  NANDN U408 ( .B(n156), .A(n157), .Z(n154) );
  NANDN U409 ( .B(n137), .A(n158), .Z(n153) );
  NANDN U410 ( .B(n138), .A(n159), .Z(n133) );
  AND U411 ( .A(n160), .B(n161), .Z(n150) );
  OR U412 ( .A(n162), .B(n163), .Z(n161) );
  XNOR U413 ( .A(n164), .B(n165), .Z(n160) );
  ANDN U414 ( .A(n166), .B(n167), .Z(n165) );
  XOR U415 ( .A(n164), .B(n168), .Z(n166) );
  ANDN U416 ( .A(n171), .B(n172), .Z(n170) );
  XOR U417 ( .A(\_MxM/Y0[12] ), .B(n173), .Z(n171) );
  XNOR U418 ( .A(n172), .B(\_MxM/Y0[12] ), .Z(\_MxM/Y1[11] ) );
  XNOR U419 ( .A(n174), .B(n175), .Z(n172) );
  XNOR U420 ( .A(n173), .B(n176), .Z(n174) );
  AND U421 ( .A(n120), .B(n177), .Z(n176) );
  XOR U422 ( .A(n146), .B(n178), .Z(n177) );
  XOR U423 ( .A(n178), .B(n147), .Z(n146) );
  OR U424 ( .A(n179), .B(n180), .Z(n147) );
  IV U425 ( .A(n175), .Z(n178) );
  XNOR U426 ( .A(n149), .B(n148), .Z(n175) );
  OR U427 ( .A(n181), .B(n182), .Z(n148) );
  XNOR U428 ( .A(n163), .B(n162), .Z(n149) );
  OR U429 ( .A(n183), .B(n184), .Z(n162) );
  XOR U430 ( .A(n168), .B(n167), .Z(n163) );
  XOR U431 ( .A(n164), .B(n185), .Z(n167) );
  AND U432 ( .A(n186), .B(n187), .Z(n185) );
  NANDN U433 ( .B(n137), .A(n188), .Z(n187) );
  OR U434 ( .A(n189), .B(n190), .Z(n186) );
  XOR U435 ( .A(n156), .B(n157), .Z(n168) );
  NANDN U436 ( .B(n138), .A(n193), .Z(n157) );
  XNOR U437 ( .A(n155), .B(n194), .Z(n156) );
  AND U438 ( .A(n159), .B(n158), .Z(n194) );
  ANDN U439 ( .A(n195), .B(n196), .Z(n155) );
  NANDN U440 ( .B(n197), .A(n198), .Z(n195) );
  IV U441 ( .A(n169), .Z(n173) );
  XNOR U442 ( .A(n200), .B(\_MxM/Y0[11] ), .Z(\_MxM/Y1[10] ) );
  XNOR U443 ( .A(n202), .B(n203), .Z(n200) );
  XNOR U444 ( .A(n201), .B(n204), .Z(n202) );
  AND U445 ( .A(n120), .B(n205), .Z(n204) );
  XOR U446 ( .A(n179), .B(n206), .Z(n205) );
  XOR U447 ( .A(n206), .B(n180), .Z(n179) );
  OR U448 ( .A(n207), .B(n208), .Z(n180) );
  IV U449 ( .A(n203), .Z(n206) );
  OR U450 ( .A(n209), .B(n210), .Z(n181) );
  XOR U451 ( .A(n192), .B(n191), .Z(n183) );
  XNOR U452 ( .A(n214), .B(n215), .Z(n191) );
  ANDN U453 ( .A(n218), .B(n219), .Z(n217) );
  XOR U454 ( .A(n216), .B(n220), .Z(n218) );
  XNOR U455 ( .A(n221), .B(n189), .Z(n214) );
  NAND U456 ( .A(n188), .B(n159), .Z(n189) );
  NANDN U457 ( .B(n137), .A(n223), .Z(n222) );
  XOR U458 ( .A(n197), .B(n198), .Z(n192) );
  NANDN U459 ( .B(n138), .A(n227), .Z(n198) );
  AND U460 ( .A(n193), .B(n158), .Z(n228) );
  NAND U461 ( .A(n229), .B(n230), .Z(n196) );
  NANDN U462 ( .B(n231), .A(n232), .Z(n229) );
  IV U463 ( .A(n199), .Z(n201) );
  XNOR U464 ( .A(n234), .B(n235), .Z(n105) );
  AND U465 ( .A(n120), .B(n237), .Z(n236) );
  XOR U466 ( .A(n207), .B(n238), .Z(n237) );
  XOR U467 ( .A(n238), .B(n208), .Z(n207) );
  OR U468 ( .A(n239), .B(n240), .Z(n208) );
  IV U469 ( .A(n235), .Z(n238) );
  XNOR U470 ( .A(n210), .B(n209), .Z(n235) );
  OR U471 ( .A(n241), .B(n242), .Z(n209) );
  XNOR U472 ( .A(n213), .B(n212), .Z(n210) );
  XOR U473 ( .A(n211), .B(n243), .Z(n212) );
  AND U474 ( .A(n244), .B(n245), .Z(n243) );
  OR U475 ( .A(n246), .B(n247), .Z(n245) );
  AND U476 ( .A(n248), .B(n249), .Z(n244) );
  NANDN U477 ( .B(n137), .A(n250), .Z(n249) );
  NAND U478 ( .A(n251), .B(n252), .Z(n248) );
  XNOR U479 ( .A(n224), .B(n257), .Z(n225) );
  AND U480 ( .A(n159), .B(n223), .Z(n257) );
  XOR U481 ( .A(n258), .B(n259), .Z(n224) );
  ANDN U482 ( .A(n260), .B(n261), .Z(n259) );
  XNOR U483 ( .A(n262), .B(n258), .Z(n260) );
  XOR U484 ( .A(n263), .B(n226), .Z(n256) );
  NAND U485 ( .A(n188), .B(n193), .Z(n226) );
  IV U486 ( .A(n216), .Z(n263) );
  XNOR U487 ( .A(n231), .B(n232), .Z(n220) );
  NANDN U488 ( .B(n138), .A(n267), .Z(n232) );
  XNOR U489 ( .A(n230), .B(n268), .Z(n231) );
  AND U490 ( .A(n227), .B(n158), .Z(n268) );
  ANDN U491 ( .A(n269), .B(n270), .Z(n230) );
  NANDN U492 ( .B(n271), .A(n272), .Z(n269) );
  XNOR U493 ( .A(n274), .B(n275), .Z(n106) );
  AND U494 ( .A(n120), .B(n277), .Z(n276) );
  XOR U495 ( .A(n239), .B(n278), .Z(n277) );
  XOR U496 ( .A(n278), .B(n240), .Z(n239) );
  OR U497 ( .A(n279), .B(n280), .Z(n240) );
  IV U498 ( .A(n275), .Z(n278) );
  XNOR U499 ( .A(n242), .B(n241), .Z(n275) );
  OR U500 ( .A(n281), .B(n282), .Z(n241) );
  XNOR U501 ( .A(n255), .B(n254), .Z(n242) );
  XOR U502 ( .A(n283), .B(n251), .Z(n254) );
  XNOR U503 ( .A(n284), .B(n246), .Z(n251) );
  NAND U504 ( .A(n250), .B(n159), .Z(n246) );
  NANDN U505 ( .B(n137), .A(n286), .Z(n285) );
  XNOR U506 ( .A(n252), .B(n253), .Z(n283) );
  XNOR U507 ( .A(n258), .B(n297), .Z(n261) );
  AND U508 ( .A(n193), .B(n223), .Z(n297) );
  XOR U509 ( .A(n298), .B(n299), .Z(n258) );
  ANDN U510 ( .A(n300), .B(n301), .Z(n299) );
  XNOR U511 ( .A(n302), .B(n298), .Z(n300) );
  XOR U512 ( .A(n303), .B(n262), .Z(n296) );
  NAND U513 ( .A(n188), .B(n227), .Z(n262) );
  IV U514 ( .A(n264), .Z(n303) );
  XNOR U515 ( .A(n271), .B(n272), .Z(n266) );
  NANDN U516 ( .B(n138), .A(n307), .Z(n272) );
  AND U517 ( .A(n267), .B(n158), .Z(n308) );
  NAND U518 ( .A(n309), .B(n310), .Z(n270) );
  NANDN U519 ( .B(n311), .A(n312), .Z(n309) );
  XNOR U520 ( .A(n314), .B(n315), .Z(n107) );
  XNOR U521 ( .A(n316), .B(n317), .Z(n314) );
  AND U522 ( .A(n120), .B(n318), .Z(n317) );
  XOR U523 ( .A(n279), .B(n319), .Z(n318) );
  XOR U524 ( .A(n319), .B(n280), .Z(n279) );
  OR U525 ( .A(n320), .B(n321), .Z(n280) );
  IV U526 ( .A(n315), .Z(n319) );
  XNOR U527 ( .A(n282), .B(n281), .Z(n315) );
  NANDN U528 ( .B(n322), .A(n323), .Z(n281) );
  XNOR U529 ( .A(n292), .B(n291), .Z(n282) );
  XOR U530 ( .A(n324), .B(n295), .Z(n291) );
  XNOR U531 ( .A(n288), .B(n289), .Z(n295) );
  NAND U532 ( .A(n250), .B(n193), .Z(n289) );
  XNOR U533 ( .A(n287), .B(n325), .Z(n288) );
  AND U534 ( .A(n159), .B(n286), .Z(n325) );
  XNOR U535 ( .A(n294), .B(n290), .Z(n324) );
  AND U536 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U537 ( .B(n137), .A(n335), .Z(n334) );
  OR U538 ( .A(n336), .B(n337), .Z(n333) );
  XNOR U539 ( .A(n298), .B(n342), .Z(n301) );
  AND U540 ( .A(n227), .B(n223), .Z(n342) );
  XOR U541 ( .A(n346), .B(n302), .Z(n341) );
  NAND U542 ( .A(n188), .B(n267), .Z(n302) );
  IV U543 ( .A(n304), .Z(n346) );
  XNOR U544 ( .A(n311), .B(n312), .Z(n306) );
  NANDN U545 ( .B(n138), .A(n350), .Z(n312) );
  XNOR U546 ( .A(n310), .B(n351), .Z(n311) );
  AND U547 ( .A(n307), .B(n158), .Z(n351) );
  ANDN U548 ( .A(n352), .B(n353), .Z(n310) );
  NANDN U549 ( .B(n354), .A(n355), .Z(n352) );
  IV U550 ( .A(n313), .Z(n316) );
  XNOR U551 ( .A(n358), .B(n359), .Z(n357) );
  AND U552 ( .A(n120), .B(n360), .Z(n359) );
  XOR U553 ( .A(n320), .B(n363), .Z(n360) );
  XOR U554 ( .A(n363), .B(n321), .Z(n320) );
  OR U555 ( .A(n361), .B(n362), .Z(n321) );
  XNOR U556 ( .A(n322), .B(n323), .Z(n363) );
  XNOR U557 ( .A(n331), .B(n330), .Z(n322) );
  XOR U558 ( .A(n368), .B(n340), .Z(n330) );
  XNOR U559 ( .A(n327), .B(n328), .Z(n340) );
  NAND U560 ( .A(n250), .B(n227), .Z(n328) );
  XNOR U561 ( .A(n326), .B(n369), .Z(n327) );
  AND U562 ( .A(n193), .B(n286), .Z(n369) );
  XNOR U563 ( .A(n339), .B(n329), .Z(n368) );
  XNOR U564 ( .A(n376), .B(n338), .Z(n339) );
  XNOR U565 ( .A(n380), .B(n336), .Z(n376) );
  NAND U566 ( .A(n335), .B(n159), .Z(n336) );
  NANDN U567 ( .B(n137), .A(n382), .Z(n381) );
  XNOR U568 ( .A(n343), .B(n387), .Z(n344) );
  AND U569 ( .A(n267), .B(n223), .Z(n387) );
  XOR U570 ( .A(n388), .B(n389), .Z(n343) );
  ANDN U571 ( .A(n390), .B(n391), .Z(n389) );
  XNOR U572 ( .A(n392), .B(n388), .Z(n390) );
  XOR U573 ( .A(n393), .B(n345), .Z(n386) );
  NAND U574 ( .A(n188), .B(n307), .Z(n345) );
  IV U575 ( .A(n347), .Z(n393) );
  XNOR U576 ( .A(n354), .B(n355), .Z(n349) );
  NANDN U577 ( .B(n138), .A(n397), .Z(n355) );
  AND U578 ( .A(n350), .B(n158), .Z(n398) );
  NAND U579 ( .A(n399), .B(n400), .Z(n353) );
  NANDN U580 ( .B(n401), .A(n402), .Z(n399) );
  IV U581 ( .A(n356), .Z(n358) );
  XNOR U582 ( .A(n404), .B(n405), .Z(n109) );
  AND U583 ( .A(n120), .B(n407), .Z(n406) );
  XOR U584 ( .A(n361), .B(n408), .Z(n407) );
  XOR U585 ( .A(n408), .B(n362), .Z(n361) );
  OR U586 ( .A(n409), .B(n410), .Z(n362) );
  IV U587 ( .A(n405), .Z(n408) );
  XOR U588 ( .A(n367), .B(n366), .Z(n405) );
  XNOR U589 ( .A(n365), .B(n411), .Z(n366) );
  AND U590 ( .A(n364), .B(n412), .Z(n411) );
  AND U591 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U592 ( .B(n137), .A(n415), .Z(n414) );
  OR U593 ( .A(n416), .B(n417), .Z(n413) );
  AND U594 ( .A(n418), .B(n419), .Z(n364) );
  NANDN U595 ( .B(n420), .A(n421), .Z(n419) );
  NANDN U596 ( .B(n422), .A(n423), .Z(n418) );
  XNOR U597 ( .A(n427), .B(n379), .Z(n374) );
  XNOR U598 ( .A(n371), .B(n372), .Z(n379) );
  NAND U599 ( .A(n250), .B(n267), .Z(n372) );
  XNOR U600 ( .A(n370), .B(n428), .Z(n371) );
  AND U601 ( .A(n227), .B(n286), .Z(n428) );
  XNOR U602 ( .A(n378), .B(n373), .Z(n427) );
  XNOR U603 ( .A(n383), .B(n436), .Z(n384) );
  AND U604 ( .A(n159), .B(n382), .Z(n436) );
  XOR U605 ( .A(n440), .B(n385), .Z(n435) );
  NAND U606 ( .A(n335), .B(n193), .Z(n385) );
  IV U607 ( .A(n377), .Z(n440) );
  XNOR U608 ( .A(n388), .B(n445), .Z(n391) );
  AND U609 ( .A(n307), .B(n223), .Z(n445) );
  XOR U610 ( .A(n446), .B(n447), .Z(n388) );
  ANDN U611 ( .A(n448), .B(n449), .Z(n447) );
  XNOR U612 ( .A(n450), .B(n446), .Z(n448) );
  XOR U613 ( .A(n451), .B(n392), .Z(n444) );
  NAND U614 ( .A(n188), .B(n350), .Z(n392) );
  IV U615 ( .A(n394), .Z(n451) );
  XNOR U616 ( .A(n401), .B(n402), .Z(n396) );
  NANDN U617 ( .B(n138), .A(n455), .Z(n402) );
  XNOR U618 ( .A(n400), .B(n456), .Z(n401) );
  AND U619 ( .A(n397), .B(n158), .Z(n456) );
  ANDN U620 ( .A(n457), .B(n458), .Z(n400) );
  NANDN U621 ( .B(n459), .A(n460), .Z(n457) );
  XNOR U622 ( .A(n462), .B(n463), .Z(n110) );
  AND U623 ( .A(n120), .B(n465), .Z(n464) );
  XOR U624 ( .A(n409), .B(n466), .Z(n465) );
  XOR U625 ( .A(n466), .B(n410), .Z(n409) );
  OR U626 ( .A(n467), .B(n468), .Z(n410) );
  IV U627 ( .A(n463), .Z(n466) );
  XOR U628 ( .A(n426), .B(n425), .Z(n463) );
  XOR U629 ( .A(n420), .B(n421), .Z(n417) );
  XOR U630 ( .A(n473), .B(n422), .Z(n420) );
  NAND U631 ( .A(n159), .B(n415), .Z(n422) );
  NANDN U632 ( .B(n423), .A(n474), .Z(n473) );
  NANDN U633 ( .B(n137), .A(n475), .Z(n474) );
  XOR U634 ( .A(n479), .B(n416), .Z(n469) );
  OR U635 ( .A(n480), .B(n481), .Z(n416) );
  IV U636 ( .A(n424), .Z(n479) );
  XNOR U637 ( .A(n485), .B(n443), .Z(n433) );
  XNOR U638 ( .A(n430), .B(n431), .Z(n443) );
  NAND U639 ( .A(n250), .B(n307), .Z(n431) );
  XNOR U640 ( .A(n429), .B(n486), .Z(n430) );
  AND U641 ( .A(n267), .B(n286), .Z(n486) );
  XNOR U642 ( .A(n442), .B(n432), .Z(n485) );
  XNOR U643 ( .A(n437), .B(n494), .Z(n438) );
  AND U644 ( .A(n193), .B(n382), .Z(n494) );
  XOR U645 ( .A(n498), .B(n439), .Z(n493) );
  NAND U646 ( .A(n335), .B(n227), .Z(n439) );
  IV U647 ( .A(n441), .Z(n498) );
  XNOR U648 ( .A(n446), .B(n503), .Z(n449) );
  AND U649 ( .A(n350), .B(n223), .Z(n503) );
  XOR U650 ( .A(n504), .B(n505), .Z(n446) );
  ANDN U651 ( .A(n506), .B(n507), .Z(n505) );
  XNOR U652 ( .A(n508), .B(n504), .Z(n506) );
  XOR U653 ( .A(n509), .B(n450), .Z(n502) );
  NAND U654 ( .A(n188), .B(n397), .Z(n450) );
  IV U655 ( .A(n452), .Z(n509) );
  XNOR U656 ( .A(n459), .B(n460), .Z(n454) );
  NANDN U657 ( .B(n138), .A(n513), .Z(n460) );
  AND U658 ( .A(n455), .B(n158), .Z(n514) );
  NAND U659 ( .A(n515), .B(n516), .Z(n458) );
  NANDN U660 ( .B(n517), .A(n518), .Z(n515) );
  XNOR U661 ( .A(n520), .B(n521), .Z(n111) );
  AND U662 ( .A(n120), .B(n523), .Z(n522) );
  XOR U663 ( .A(n467), .B(n524), .Z(n523) );
  XOR U664 ( .A(n524), .B(n468), .Z(n467) );
  OR U665 ( .A(n525), .B(n526), .Z(n468) );
  IV U666 ( .A(n521), .Z(n524) );
  XOR U667 ( .A(n484), .B(n483), .Z(n521) );
  XOR U668 ( .A(n527), .B(n480), .Z(n483) );
  XOR U669 ( .A(n472), .B(n471), .Z(n480) );
  XOR U670 ( .A(n470), .B(n528), .Z(n471) );
  AND U671 ( .A(n529), .B(n530), .Z(n528) );
  NANDN U672 ( .B(n137), .A(n531), .Z(n530) );
  OR U673 ( .A(n532), .B(n533), .Z(n529) );
  NAND U674 ( .A(n193), .B(n415), .Z(n478) );
  XNOR U675 ( .A(n476), .B(n537), .Z(n477) );
  AND U676 ( .A(n475), .B(n159), .Z(n537) );
  NANDN U677 ( .B(n541), .A(n542), .Z(n481) );
  XNOR U678 ( .A(n546), .B(n501), .Z(n491) );
  XNOR U679 ( .A(n488), .B(n489), .Z(n501) );
  NAND U680 ( .A(n250), .B(n350), .Z(n489) );
  XNOR U681 ( .A(n487), .B(n547), .Z(n488) );
  AND U682 ( .A(n307), .B(n286), .Z(n547) );
  XNOR U683 ( .A(n500), .B(n490), .Z(n546) );
  XNOR U684 ( .A(n495), .B(n555), .Z(n496) );
  AND U685 ( .A(n227), .B(n382), .Z(n555) );
  XOR U686 ( .A(n559), .B(n497), .Z(n554) );
  NAND U687 ( .A(n335), .B(n267), .Z(n497) );
  IV U688 ( .A(n499), .Z(n559) );
  XNOR U689 ( .A(n504), .B(n564), .Z(n507) );
  AND U690 ( .A(n397), .B(n223), .Z(n564) );
  XOR U691 ( .A(n565), .B(n566), .Z(n504) );
  ANDN U692 ( .A(n567), .B(n568), .Z(n566) );
  XNOR U693 ( .A(n569), .B(n565), .Z(n567) );
  XOR U694 ( .A(n570), .B(n508), .Z(n563) );
  NAND U695 ( .A(n188), .B(n455), .Z(n508) );
  IV U696 ( .A(n510), .Z(n570) );
  XNOR U697 ( .A(n517), .B(n518), .Z(n512) );
  NANDN U698 ( .B(n138), .A(n574), .Z(n518) );
  XNOR U699 ( .A(n516), .B(n575), .Z(n517) );
  AND U700 ( .A(n513), .B(n158), .Z(n575) );
  ANDN U701 ( .A(n576), .B(n577), .Z(n516) );
  NANDN U702 ( .B(n578), .A(n579), .Z(n576) );
  XNOR U703 ( .A(n581), .B(n582), .Z(n112) );
  AND U704 ( .A(n120), .B(n584), .Z(n583) );
  XOR U705 ( .A(n525), .B(n585), .Z(n584) );
  XOR U706 ( .A(n585), .B(n526), .Z(n525) );
  OR U707 ( .A(n586), .B(n587), .Z(n526) );
  IV U708 ( .A(n582), .Z(n585) );
  XOR U709 ( .A(n545), .B(n544), .Z(n582) );
  XOR U710 ( .A(n588), .B(n541), .Z(n544) );
  XOR U711 ( .A(n536), .B(n535), .Z(n541) );
  XNOR U712 ( .A(n593), .B(n532), .Z(n589) );
  NAND U713 ( .A(n159), .B(n531), .Z(n532) );
  NANDN U714 ( .B(n137), .A(n595), .Z(n594) );
  NAND U715 ( .A(n227), .B(n415), .Z(n540) );
  XNOR U716 ( .A(n538), .B(n599), .Z(n539) );
  AND U717 ( .A(n475), .B(n193), .Z(n599) );
  XNOR U718 ( .A(n542), .B(n543), .Z(n588) );
  XNOR U719 ( .A(n609), .B(n562), .Z(n552) );
  XNOR U720 ( .A(n549), .B(n550), .Z(n562) );
  NAND U721 ( .A(n250), .B(n397), .Z(n550) );
  XNOR U722 ( .A(n548), .B(n610), .Z(n549) );
  AND U723 ( .A(n350), .B(n286), .Z(n610) );
  XNOR U724 ( .A(n561), .B(n551), .Z(n609) );
  XNOR U725 ( .A(n556), .B(n618), .Z(n557) );
  AND U726 ( .A(n267), .B(n382), .Z(n618) );
  XOR U727 ( .A(n619), .B(n620), .Z(n556) );
  ANDN U728 ( .A(n621), .B(n622), .Z(n620) );
  XNOR U729 ( .A(n623), .B(n619), .Z(n621) );
  XOR U730 ( .A(n624), .B(n558), .Z(n617) );
  NAND U731 ( .A(n335), .B(n307), .Z(n558) );
  IV U732 ( .A(n560), .Z(n624) );
  XNOR U733 ( .A(n565), .B(n629), .Z(n568) );
  AND U734 ( .A(n455), .B(n223), .Z(n629) );
  XOR U735 ( .A(n630), .B(n631), .Z(n565) );
  ANDN U736 ( .A(n632), .B(n633), .Z(n631) );
  XNOR U737 ( .A(n634), .B(n630), .Z(n632) );
  XOR U738 ( .A(n635), .B(n569), .Z(n628) );
  NAND U739 ( .A(n188), .B(n513), .Z(n569) );
  IV U740 ( .A(n571), .Z(n635) );
  XNOR U741 ( .A(n578), .B(n579), .Z(n573) );
  OR U742 ( .A(n639), .B(n138), .Z(n579) );
  AND U743 ( .A(n574), .B(n158), .Z(n640) );
  NAND U744 ( .A(n641), .B(n642), .Z(n577) );
  NANDN U745 ( .B(n643), .A(n644), .Z(n641) );
  XNOR U746 ( .A(n646), .B(n647), .Z(n113) );
  XOR U747 ( .A(n645), .B(n648), .Z(n646) );
  AND U748 ( .A(n120), .B(n649), .Z(n648) );
  XOR U749 ( .A(n586), .B(n650), .Z(n649) );
  XOR U750 ( .A(n650), .B(n587), .Z(n586) );
  NANDN U751 ( .B(n651), .A(n652), .Z(n587) );
  IV U752 ( .A(n647), .Z(n650) );
  XOR U753 ( .A(n605), .B(n604), .Z(n647) );
  XNOR U754 ( .A(n653), .B(n608), .Z(n604) );
  XNOR U755 ( .A(n596), .B(n655), .Z(n597) );
  AND U756 ( .A(n595), .B(n159), .Z(n655) );
  XOR U757 ( .A(n659), .B(n598), .Z(n654) );
  NAND U758 ( .A(n193), .B(n531), .Z(n598) );
  IV U759 ( .A(n590), .Z(n659) );
  XNOR U760 ( .A(n601), .B(n602), .Z(n592) );
  NAND U761 ( .A(n267), .B(n415), .Z(n602) );
  XNOR U762 ( .A(n600), .B(n663), .Z(n601) );
  AND U763 ( .A(n475), .B(n227), .Z(n663) );
  XNOR U764 ( .A(n607), .B(n603), .Z(n653) );
  AND U765 ( .A(n671), .B(n672), .Z(n670) );
  OR U766 ( .A(n673), .B(n674), .Z(n672) );
  AND U767 ( .A(n675), .B(n676), .Z(n671) );
  NANDN U768 ( .B(n137), .A(n677), .Z(n676) );
  NANDN U769 ( .B(n678), .A(n679), .Z(n675) );
  XNOR U770 ( .A(n683), .B(n627), .Z(n615) );
  XNOR U771 ( .A(n612), .B(n613), .Z(n627) );
  NAND U772 ( .A(n250), .B(n455), .Z(n613) );
  XNOR U773 ( .A(n611), .B(n684), .Z(n612) );
  AND U774 ( .A(n397), .B(n286), .Z(n684) );
  XNOR U775 ( .A(n626), .B(n614), .Z(n683) );
  XNOR U776 ( .A(n619), .B(n692), .Z(n622) );
  AND U777 ( .A(n307), .B(n382), .Z(n692) );
  XOR U778 ( .A(n696), .B(n623), .Z(n691) );
  NAND U779 ( .A(n335), .B(n350), .Z(n623) );
  IV U780 ( .A(n625), .Z(n696) );
  XNOR U781 ( .A(n630), .B(n701), .Z(n633) );
  AND U782 ( .A(n513), .B(n223), .Z(n701) );
  XOR U783 ( .A(n702), .B(n703), .Z(n630) );
  ANDN U784 ( .A(n704), .B(n705), .Z(n703) );
  XNOR U785 ( .A(n706), .B(n702), .Z(n704) );
  XOR U786 ( .A(n707), .B(n634), .Z(n700) );
  NAND U787 ( .A(n188), .B(n574), .Z(n634) );
  IV U788 ( .A(n636), .Z(n707) );
  XNOR U789 ( .A(n643), .B(n644), .Z(n638) );
  OR U790 ( .A(n711), .B(n138), .Z(n644) );
  XNOR U791 ( .A(n642), .B(n712), .Z(n643) );
  ANDN U792 ( .A(n158), .B(n639), .Z(n712) );
  ANDN U793 ( .A(n713), .B(n714), .Z(n642) );
  NANDN U794 ( .B(n715), .A(n716), .Z(n713) );
  XNOR U795 ( .A(n718), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U796 ( .A(n719), .B(n720), .Z(n718) );
  XNOR U797 ( .A(n721), .B(n717), .Z(n719) );
  NAND U798 ( .A(\_MxM/Y0[0] ), .B(n651), .Z(n717) );
  NAND U799 ( .A(n722), .B(n120), .Z(n721) );
  XOR U800 ( .A(e_input[15]), .B(g_input[15]), .Z(n120) );
  XNOR U801 ( .A(n652), .B(n720), .Z(n722) );
  XNOR U802 ( .A(n651), .B(n720), .Z(n652) );
  XNOR U803 ( .A(n669), .B(n668), .Z(n720) );
  XNOR U804 ( .A(n723), .B(n682), .Z(n668) );
  XNOR U805 ( .A(n656), .B(n725), .Z(n657) );
  AND U806 ( .A(n595), .B(n193), .Z(n725) );
  XOR U807 ( .A(n729), .B(n658), .Z(n724) );
  NAND U808 ( .A(n227), .B(n531), .Z(n658) );
  IV U809 ( .A(n660), .Z(n729) );
  XNOR U810 ( .A(n665), .B(n666), .Z(n662) );
  NAND U811 ( .A(n307), .B(n415), .Z(n666) );
  XNOR U812 ( .A(n664), .B(n733), .Z(n665) );
  AND U813 ( .A(n475), .B(n267), .Z(n733) );
  XNOR U814 ( .A(n681), .B(n667), .Z(n723) );
  XNOR U815 ( .A(n740), .B(n678), .Z(n681) );
  XOR U816 ( .A(n741), .B(n673), .Z(n678) );
  NAND U817 ( .A(n159), .B(n677), .Z(n673) );
  NANDN U818 ( .B(n137), .A(n743), .Z(n742) );
  XNOR U819 ( .A(n679), .B(n680), .Z(n740) );
  XNOR U820 ( .A(n752), .B(n699), .Z(n689) );
  XNOR U821 ( .A(n686), .B(n687), .Z(n699) );
  NAND U822 ( .A(n250), .B(n513), .Z(n687) );
  XNOR U823 ( .A(n685), .B(n753), .Z(n686) );
  AND U824 ( .A(n455), .B(n286), .Z(n753) );
  XNOR U825 ( .A(n698), .B(n688), .Z(n752) );
  XNOR U826 ( .A(n693), .B(n761), .Z(n694) );
  AND U827 ( .A(n350), .B(n382), .Z(n761) );
  XOR U828 ( .A(n762), .B(n763), .Z(n693) );
  ANDN U829 ( .A(n764), .B(n765), .Z(n763) );
  XNOR U830 ( .A(n766), .B(n762), .Z(n764) );
  XOR U831 ( .A(n767), .B(n695), .Z(n760) );
  NAND U832 ( .A(n335), .B(n397), .Z(n695) );
  IV U833 ( .A(n697), .Z(n767) );
  XNOR U834 ( .A(n702), .B(n772), .Z(n705) );
  AND U835 ( .A(n574), .B(n223), .Z(n772) );
  XOR U836 ( .A(n773), .B(n774), .Z(n702) );
  ANDN U837 ( .A(n775), .B(n776), .Z(n774) );
  XNOR U838 ( .A(n777), .B(n773), .Z(n775) );
  XOR U839 ( .A(n778), .B(n706), .Z(n771) );
  NANDN U840 ( .B(n639), .A(n188), .Z(n706) );
  IV U841 ( .A(n708), .Z(n778) );
  XNOR U842 ( .A(n715), .B(n716), .Z(n710) );
  NANDN U843 ( .B(n138), .A(n782), .Z(n716) );
  ANDN U844 ( .A(n158), .B(n711), .Z(n783) );
  NAND U845 ( .A(n784), .B(n785), .Z(n714) );
  NANDN U846 ( .B(n786), .A(n787), .Z(n784) );
  XNOR U847 ( .A(n739), .B(n738), .Z(n651) );
  XNOR U848 ( .A(n788), .B(n749), .Z(n738) );
  XNOR U849 ( .A(n726), .B(n790), .Z(n727) );
  AND U850 ( .A(n595), .B(n227), .Z(n790) );
  XOR U851 ( .A(n791), .B(n792), .Z(n726) );
  ANDN U852 ( .A(n793), .B(n794), .Z(n792) );
  XNOR U853 ( .A(n795), .B(n791), .Z(n793) );
  XOR U854 ( .A(n796), .B(n728), .Z(n789) );
  NAND U855 ( .A(n267), .B(n531), .Z(n728) );
  IV U856 ( .A(n730), .Z(n796) );
  XNOR U857 ( .A(n735), .B(n736), .Z(n732) );
  NAND U858 ( .A(n350), .B(n415), .Z(n736) );
  XNOR U859 ( .A(n734), .B(n800), .Z(n735) );
  AND U860 ( .A(n475), .B(n307), .Z(n800) );
  XNOR U861 ( .A(n748), .B(n737), .Z(n788) );
  XOR U862 ( .A(n804), .B(n805), .Z(n737) );
  XNOR U863 ( .A(n806), .B(n751), .Z(n748) );
  NAND U864 ( .A(n193), .B(n677), .Z(n746) );
  XNOR U865 ( .A(n744), .B(n807), .Z(n745) );
  AND U866 ( .A(n743), .B(n159), .Z(n807) );
  XNOR U867 ( .A(n750), .B(n747), .Z(n806) );
  XOR U868 ( .A(n811), .B(n812), .Z(n747) );
  AND U869 ( .A(n813), .B(n814), .Z(n812) );
  XOR U870 ( .A(n815), .B(n816), .Z(n814) );
  XOR U871 ( .A(n811), .B(n817), .Z(n816) );
  XOR U872 ( .A(n798), .B(n818), .Z(n813) );
  XOR U873 ( .A(n811), .B(n799), .Z(n818) );
  NAND U874 ( .A(n415), .B(n397), .Z(n803) );
  XNOR U875 ( .A(n801), .B(n819), .Z(n802) );
  AND U876 ( .A(n475), .B(n350), .Z(n819) );
  XNOR U877 ( .A(n791), .B(n824), .Z(n794) );
  AND U878 ( .A(n595), .B(n267), .Z(n824) );
  XOR U879 ( .A(n828), .B(n795), .Z(n823) );
  NAND U880 ( .A(n307), .B(n531), .Z(n795) );
  IV U881 ( .A(n797), .Z(n828) );
  XOR U882 ( .A(n832), .B(n833), .Z(n811) );
  AND U883 ( .A(n834), .B(n835), .Z(n833) );
  XOR U884 ( .A(n836), .B(n837), .Z(n835) );
  XOR U885 ( .A(n832), .B(n838), .Z(n837) );
  XOR U886 ( .A(n830), .B(n839), .Z(n834) );
  XOR U887 ( .A(n832), .B(n831), .Z(n839) );
  NAND U888 ( .A(n415), .B(n455), .Z(n822) );
  XNOR U889 ( .A(n820), .B(n840), .Z(n821) );
  AND U890 ( .A(n397), .B(n475), .Z(n840) );
  XNOR U891 ( .A(n825), .B(n845), .Z(n826) );
  AND U892 ( .A(n595), .B(n307), .Z(n845) );
  XOR U893 ( .A(n846), .B(n847), .Z(n825) );
  ANDN U894 ( .A(n848), .B(n849), .Z(n847) );
  XNOR U895 ( .A(n850), .B(n846), .Z(n848) );
  XOR U896 ( .A(n851), .B(n827), .Z(n844) );
  NAND U897 ( .A(n350), .B(n531), .Z(n827) );
  IV U898 ( .A(n829), .Z(n851) );
  XOR U899 ( .A(n855), .B(n856), .Z(n832) );
  AND U900 ( .A(n857), .B(n858), .Z(n856) );
  XOR U901 ( .A(n859), .B(n860), .Z(n858) );
  XOR U902 ( .A(n855), .B(n861), .Z(n860) );
  XOR U903 ( .A(n853), .B(n862), .Z(n857) );
  XOR U904 ( .A(n855), .B(n854), .Z(n862) );
  NAND U905 ( .A(n415), .B(n513), .Z(n843) );
  XNOR U906 ( .A(n841), .B(n863), .Z(n842) );
  AND U907 ( .A(n455), .B(n475), .Z(n863) );
  XOR U908 ( .A(n864), .B(n865), .Z(n841) );
  ANDN U909 ( .A(n866), .B(n867), .Z(n865) );
  XNOR U910 ( .A(n868), .B(n864), .Z(n866) );
  XNOR U911 ( .A(n869), .B(n870), .Z(n853) );
  IV U912 ( .A(n849), .Z(n870) );
  XNOR U913 ( .A(n846), .B(n871), .Z(n849) );
  AND U914 ( .A(n595), .B(n350), .Z(n871) );
  XOR U915 ( .A(n872), .B(n873), .Z(n846) );
  ANDN U916 ( .A(n874), .B(n875), .Z(n873) );
  XNOR U917 ( .A(n876), .B(n872), .Z(n874) );
  XOR U918 ( .A(n877), .B(n850), .Z(n869) );
  NAND U919 ( .A(n531), .B(n397), .Z(n850) );
  IV U920 ( .A(n852), .Z(n877) );
  XOR U921 ( .A(n881), .B(n882), .Z(n855) );
  AND U922 ( .A(n883), .B(n884), .Z(n882) );
  XOR U923 ( .A(n885), .B(n886), .Z(n884) );
  XOR U924 ( .A(n881), .B(n887), .Z(n886) );
  XOR U925 ( .A(n879), .B(n888), .Z(n883) );
  XOR U926 ( .A(n881), .B(n880), .Z(n888) );
  XNOR U927 ( .A(n889), .B(n868), .Z(n880) );
  NAND U928 ( .A(n415), .B(n574), .Z(n868) );
  IV U929 ( .A(n867), .Z(n889) );
  XNOR U930 ( .A(n864), .B(n890), .Z(n867) );
  AND U931 ( .A(n513), .B(n475), .Z(n890) );
  XOR U932 ( .A(n891), .B(n892), .Z(n864) );
  ANDN U933 ( .A(n893), .B(n894), .Z(n892) );
  XNOR U934 ( .A(n895), .B(n891), .Z(n893) );
  XNOR U935 ( .A(n896), .B(n897), .Z(n879) );
  IV U936 ( .A(n875), .Z(n897) );
  XNOR U937 ( .A(n872), .B(n898), .Z(n875) );
  AND U938 ( .A(n397), .B(n595), .Z(n898) );
  XOR U939 ( .A(n899), .B(n900), .Z(n872) );
  ANDN U940 ( .A(n901), .B(n902), .Z(n900) );
  XNOR U941 ( .A(n903), .B(n899), .Z(n901) );
  XOR U942 ( .A(n904), .B(n876), .Z(n896) );
  NAND U943 ( .A(n531), .B(n455), .Z(n876) );
  IV U944 ( .A(n878), .Z(n904) );
  XOR U945 ( .A(n908), .B(n909), .Z(n881) );
  AND U946 ( .A(n910), .B(n911), .Z(n909) );
  XOR U947 ( .A(n912), .B(n913), .Z(n911) );
  XOR U948 ( .A(n908), .B(n914), .Z(n913) );
  XOR U949 ( .A(n906), .B(n915), .Z(n910) );
  XOR U950 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U951 ( .A(n916), .B(n895), .Z(n907) );
  NANDN U952 ( .B(n639), .A(n415), .Z(n895) );
  IV U953 ( .A(n894), .Z(n916) );
  XNOR U954 ( .A(n891), .B(n917), .Z(n894) );
  AND U955 ( .A(n574), .B(n475), .Z(n917) );
  XOR U956 ( .A(n918), .B(n919), .Z(n891) );
  ANDN U957 ( .A(n920), .B(n921), .Z(n919) );
  XNOR U958 ( .A(n922), .B(n918), .Z(n920) );
  XNOR U959 ( .A(n923), .B(n924), .Z(n906) );
  IV U960 ( .A(n902), .Z(n924) );
  XNOR U961 ( .A(n899), .B(n925), .Z(n902) );
  AND U962 ( .A(n455), .B(n595), .Z(n925) );
  XOR U963 ( .A(n926), .B(n927), .Z(n899) );
  ANDN U964 ( .A(n928), .B(n929), .Z(n927) );
  XNOR U965 ( .A(n930), .B(n926), .Z(n928) );
  XOR U966 ( .A(n931), .B(n903), .Z(n923) );
  NAND U967 ( .A(n531), .B(n513), .Z(n903) );
  IV U968 ( .A(n905), .Z(n931) );
  XOR U969 ( .A(n935), .B(n936), .Z(n908) );
  AND U970 ( .A(n937), .B(n938), .Z(n936) );
  XOR U971 ( .A(n939), .B(n940), .Z(n938) );
  XOR U972 ( .A(n935), .B(n941), .Z(n940) );
  XOR U973 ( .A(n933), .B(n942), .Z(n937) );
  XOR U974 ( .A(n935), .B(n934), .Z(n942) );
  XNOR U975 ( .A(n943), .B(n922), .Z(n934) );
  NANDN U976 ( .B(n711), .A(n415), .Z(n922) );
  IV U977 ( .A(n921), .Z(n943) );
  XNOR U978 ( .A(n918), .B(n944), .Z(n921) );
  ANDN U979 ( .A(n475), .B(n639), .Z(n944) );
  XOR U980 ( .A(n945), .B(n946), .Z(n918) );
  ANDN U981 ( .A(n947), .B(n948), .Z(n946) );
  XNOR U982 ( .A(n949), .B(n945), .Z(n947) );
  XNOR U983 ( .A(n950), .B(n951), .Z(n933) );
  IV U984 ( .A(n929), .Z(n951) );
  XNOR U985 ( .A(n926), .B(n952), .Z(n929) );
  AND U986 ( .A(n513), .B(n595), .Z(n952) );
  XOR U987 ( .A(n953), .B(n954), .Z(n926) );
  ANDN U988 ( .A(n955), .B(n956), .Z(n954) );
  XNOR U989 ( .A(n957), .B(n953), .Z(n955) );
  XOR U990 ( .A(n958), .B(n930), .Z(n950) );
  NAND U991 ( .A(n531), .B(n574), .Z(n930) );
  IV U992 ( .A(n932), .Z(n958) );
  XOR U993 ( .A(n962), .B(n963), .Z(n935) );
  AND U994 ( .A(n964), .B(n965), .Z(n963) );
  XOR U995 ( .A(n966), .B(n967), .Z(n965) );
  XOR U996 ( .A(n962), .B(n968), .Z(n967) );
  XOR U997 ( .A(n960), .B(n969), .Z(n964) );
  XOR U998 ( .A(n962), .B(n961), .Z(n969) );
  XNOR U999 ( .A(n970), .B(n949), .Z(n961) );
  NAND U1000 ( .A(n415), .B(n782), .Z(n949) );
  IV U1001 ( .A(n948), .Z(n970) );
  XNOR U1002 ( .A(n945), .B(n971), .Z(n948) );
  ANDN U1003 ( .A(n475), .B(n711), .Z(n971) );
  XOR U1004 ( .A(n972), .B(n973), .Z(n945) );
  ANDN U1005 ( .A(n974), .B(n975), .Z(n973) );
  XNOR U1006 ( .A(n976), .B(n972), .Z(n974) );
  XNOR U1007 ( .A(n977), .B(n978), .Z(n960) );
  IV U1008 ( .A(n956), .Z(n978) );
  XNOR U1009 ( .A(n953), .B(n979), .Z(n956) );
  AND U1010 ( .A(n574), .B(n595), .Z(n979) );
  XOR U1011 ( .A(n980), .B(n981), .Z(n953) );
  ANDN U1012 ( .A(n982), .B(n983), .Z(n981) );
  XNOR U1013 ( .A(n984), .B(n980), .Z(n982) );
  XOR U1014 ( .A(n985), .B(n957), .Z(n977) );
  NANDN U1015 ( .B(n639), .A(n531), .Z(n957) );
  IV U1016 ( .A(n959), .Z(n985) );
  XOR U1017 ( .A(n990), .B(n991), .Z(n805) );
  XNOR U1018 ( .A(n992), .B(n989), .Z(n990) );
  XNOR U1019 ( .A(n980), .B(n994), .Z(n983) );
  ANDN U1020 ( .A(n595), .B(n639), .Z(n994) );
  XOR U1021 ( .A(n997), .B(n995), .Z(n996) );
  ANDN U1022 ( .A(n595), .B(n711), .Z(n997) );
  AND U1023 ( .A(n782), .B(n531), .Z(n998) );
  XOR U1024 ( .A(n999), .B(n1000), .Z(n995) );
  ANDN U1025 ( .A(n1001), .B(n1002), .Z(n1000) );
  XNOR U1026 ( .A(n1003), .B(n999), .Z(n1001) );
  XOR U1027 ( .A(n1004), .B(n984), .Z(n993) );
  NANDN U1028 ( .B(n711), .A(n531), .Z(n984) );
  IV U1029 ( .A(n986), .Z(n1004) );
  NAND U1030 ( .A(n531), .B(n1005), .Z(n1003) );
  XNOR U1031 ( .A(n999), .B(n1006), .Z(n1002) );
  AND U1032 ( .A(n782), .B(n595), .Z(n1006) );
  AND U1033 ( .A(n1007), .B(g_input[0]), .Z(n999) );
  NANDN U1034 ( .B(n531), .A(n1008), .Z(n1007) );
  NAND U1035 ( .A(n1005), .B(n595), .Z(n1008) );
  XNOR U1036 ( .A(n975), .B(n976), .Z(n988) );
  NAND U1037 ( .A(n415), .B(n1005), .Z(n976) );
  XNOR U1038 ( .A(n972), .B(n1011), .Z(n975) );
  AND U1039 ( .A(n782), .B(n475), .Z(n1011) );
  AND U1040 ( .A(n1012), .B(g_input[0]), .Z(n972) );
  NANDN U1041 ( .B(n415), .A(n1013), .Z(n1012) );
  NAND U1042 ( .A(n1005), .B(n475), .Z(n1013) );
  XOR U1043 ( .A(n1016), .B(n1017), .Z(n989) );
  XOR U1044 ( .A(n1018), .B(n1019), .Z(n750) );
  AND U1045 ( .A(n1020), .B(n1021), .Z(n1019) );
  NANDN U1046 ( .B(n137), .A(n1022), .Z(n1021) );
  NANDN U1047 ( .B(n1023), .A(n1024), .Z(n137) );
  AND U1048 ( .A(n1025), .B(g_input[15]), .Z(n1024) );
  OR U1049 ( .A(n1026), .B(n1027), .Z(n1020) );
  AND U1050 ( .A(n817), .B(n1030), .Z(n1029) );
  XNOR U1051 ( .A(n1028), .B(n815), .Z(n1030) );
  NAND U1052 ( .A(n227), .B(n677), .Z(n810) );
  XNOR U1053 ( .A(n808), .B(n1031), .Z(n809) );
  AND U1054 ( .A(n743), .B(n193), .Z(n1031) );
  XOR U1055 ( .A(n1039), .B(n1026), .Z(n1035) );
  NAND U1056 ( .A(n159), .B(n1022), .Z(n1026) );
  IV U1057 ( .A(n1028), .Z(n1039) );
  NAND U1058 ( .A(n267), .B(n677), .Z(n1034) );
  XNOR U1059 ( .A(n1032), .B(n1041), .Z(n1033) );
  AND U1060 ( .A(n743), .B(n227), .Z(n1041) );
  XNOR U1061 ( .A(n1045), .B(n1046), .Z(n838) );
  IV U1062 ( .A(n1037), .Z(n1046) );
  XNOR U1063 ( .A(n1036), .B(n1047), .Z(n1037) );
  AND U1064 ( .A(n159), .B(e_input[0]), .Z(n1047) );
  XNOR U1065 ( .A(n1025), .B(g_input[14]), .Z(n1023) );
  NOR U1066 ( .A(n1048), .B(n1049), .Z(n1025) );
  XOR U1067 ( .A(n1053), .B(n1038), .Z(n1045) );
  NAND U1068 ( .A(n193), .B(n1022), .Z(n1038) );
  IV U1069 ( .A(n1040), .Z(n1053) );
  NAND U1070 ( .A(n307), .B(n677), .Z(n1044) );
  XNOR U1071 ( .A(n1042), .B(n1055), .Z(n1043) );
  AND U1072 ( .A(n743), .B(n267), .Z(n1055) );
  XOR U1073 ( .A(n1056), .B(n1057), .Z(n1042) );
  ANDN U1074 ( .A(n1058), .B(n1059), .Z(n1057) );
  XNOR U1075 ( .A(n1060), .B(n1056), .Z(n1058) );
  XNOR U1076 ( .A(n1050), .B(n1062), .Z(n1051) );
  AND U1077 ( .A(n193), .B(e_input[0]), .Z(n1062) );
  XOR U1078 ( .A(n1048), .B(g_input[13]), .Z(n1049) );
  NANDN U1079 ( .B(n1063), .A(n1064), .Z(n1048) );
  XOR U1080 ( .A(n1068), .B(n1052), .Z(n1061) );
  NAND U1081 ( .A(n227), .B(n1022), .Z(n1052) );
  IV U1082 ( .A(n1054), .Z(n1068) );
  XNOR U1083 ( .A(n1070), .B(n1060), .Z(n885) );
  NAND U1084 ( .A(n350), .B(n677), .Z(n1060) );
  IV U1085 ( .A(n1059), .Z(n1070) );
  XNOR U1086 ( .A(n1056), .B(n1071), .Z(n1059) );
  AND U1087 ( .A(n743), .B(n307), .Z(n1071) );
  XOR U1088 ( .A(n1072), .B(n1073), .Z(n1056) );
  ANDN U1089 ( .A(n1074), .B(n1075), .Z(n1073) );
  XNOR U1090 ( .A(n1076), .B(n1072), .Z(n1074) );
  XNOR U1091 ( .A(n1077), .B(n1078), .Z(n887) );
  IV U1092 ( .A(n1066), .Z(n1078) );
  XNOR U1093 ( .A(n1065), .B(n1079), .Z(n1066) );
  AND U1094 ( .A(n227), .B(e_input[0]), .Z(n1079) );
  XNOR U1095 ( .A(n1064), .B(g_input[12]), .Z(n1063) );
  NOR U1096 ( .A(n1080), .B(n1081), .Z(n1064) );
  XOR U1097 ( .A(n1085), .B(n1067), .Z(n1077) );
  NAND U1098 ( .A(n267), .B(n1022), .Z(n1067) );
  IV U1099 ( .A(n1069), .Z(n1085) );
  XNOR U1100 ( .A(n1087), .B(n1076), .Z(n912) );
  NAND U1101 ( .A(n397), .B(n677), .Z(n1076) );
  IV U1102 ( .A(n1075), .Z(n1087) );
  XNOR U1103 ( .A(n1072), .B(n1088), .Z(n1075) );
  AND U1104 ( .A(n743), .B(n350), .Z(n1088) );
  XOR U1105 ( .A(n1089), .B(n1090), .Z(n1072) );
  ANDN U1106 ( .A(n1091), .B(n1092), .Z(n1090) );
  XNOR U1107 ( .A(n1093), .B(n1089), .Z(n1091) );
  XNOR U1108 ( .A(n1094), .B(n1095), .Z(n914) );
  IV U1109 ( .A(n1083), .Z(n1095) );
  XNOR U1110 ( .A(n1082), .B(n1096), .Z(n1083) );
  AND U1111 ( .A(n267), .B(e_input[0]), .Z(n1096) );
  XOR U1112 ( .A(n1080), .B(g_input[11]), .Z(n1081) );
  NANDN U1113 ( .B(n1097), .A(n1098), .Z(n1080) );
  XOR U1114 ( .A(n1099), .B(n1100), .Z(n1082) );
  ANDN U1115 ( .A(n1101), .B(n1102), .Z(n1100) );
  XNOR U1116 ( .A(n1103), .B(n1099), .Z(n1101) );
  XOR U1117 ( .A(n1104), .B(n1084), .Z(n1094) );
  NAND U1118 ( .A(n307), .B(n1022), .Z(n1084) );
  IV U1119 ( .A(n1086), .Z(n1104) );
  XNOR U1120 ( .A(n1106), .B(n1093), .Z(n939) );
  NAND U1121 ( .A(n455), .B(n677), .Z(n1093) );
  IV U1122 ( .A(n1092), .Z(n1106) );
  XNOR U1123 ( .A(n1089), .B(n1107), .Z(n1092) );
  AND U1124 ( .A(n743), .B(n397), .Z(n1107) );
  XOR U1125 ( .A(n1108), .B(n1109), .Z(n1089) );
  ANDN U1126 ( .A(n1110), .B(n1111), .Z(n1109) );
  XNOR U1127 ( .A(n1112), .B(n1108), .Z(n1110) );
  XNOR U1128 ( .A(n1113), .B(n1114), .Z(n941) );
  IV U1129 ( .A(n1102), .Z(n1114) );
  XNOR U1130 ( .A(n1099), .B(n1115), .Z(n1102) );
  AND U1131 ( .A(n307), .B(e_input[0]), .Z(n1115) );
  XNOR U1132 ( .A(n1098), .B(g_input[10]), .Z(n1097) );
  NOR U1133 ( .A(n1116), .B(n1117), .Z(n1098) );
  XOR U1134 ( .A(n1121), .B(n1103), .Z(n1113) );
  NAND U1135 ( .A(n350), .B(n1022), .Z(n1103) );
  IV U1136 ( .A(n1105), .Z(n1121) );
  XNOR U1137 ( .A(n1123), .B(n1112), .Z(n966) );
  NAND U1138 ( .A(n513), .B(n677), .Z(n1112) );
  IV U1139 ( .A(n1111), .Z(n1123) );
  XNOR U1140 ( .A(n1108), .B(n1124), .Z(n1111) );
  AND U1141 ( .A(n743), .B(n455), .Z(n1124) );
  XOR U1142 ( .A(n1125), .B(n1126), .Z(n1108) );
  ANDN U1143 ( .A(n1127), .B(n1128), .Z(n1126) );
  XNOR U1144 ( .A(n1129), .B(n1125), .Z(n1127) );
  XNOR U1145 ( .A(n1130), .B(n1131), .Z(n968) );
  IV U1146 ( .A(n1119), .Z(n1131) );
  XNOR U1147 ( .A(n1118), .B(n1132), .Z(n1119) );
  AND U1148 ( .A(n350), .B(e_input[0]), .Z(n1132) );
  XOR U1149 ( .A(n1116), .B(g_input[9]), .Z(n1117) );
  NANDN U1150 ( .B(n1133), .A(n1134), .Z(n1116) );
  XOR U1151 ( .A(n1135), .B(n1136), .Z(n1118) );
  ANDN U1152 ( .A(n1137), .B(n1138), .Z(n1136) );
  XNOR U1153 ( .A(n1139), .B(n1135), .Z(n1137) );
  XOR U1154 ( .A(n1140), .B(n1120), .Z(n1130) );
  NAND U1155 ( .A(n397), .B(n1022), .Z(n1120) );
  IV U1156 ( .A(n1122), .Z(n1140) );
  NAND U1157 ( .A(n574), .B(n677), .Z(n1129) );
  XNOR U1158 ( .A(n1125), .B(n1142), .Z(n1128) );
  AND U1159 ( .A(n743), .B(n513), .Z(n1142) );
  XNOR U1160 ( .A(n1146), .B(n1143), .Z(n1145) );
  XNOR U1161 ( .A(n1135), .B(n1148), .Z(n1138) );
  AND U1162 ( .A(n397), .B(e_input[0]), .Z(n1148) );
  XNOR U1163 ( .A(n1152), .B(n1149), .Z(n1151) );
  XOR U1164 ( .A(n1153), .B(n1139), .Z(n1147) );
  NAND U1165 ( .A(n455), .B(n1022), .Z(n1139) );
  IV U1166 ( .A(n1141), .Z(n1153) );
  XNOR U1167 ( .A(n1154), .B(n1155), .Z(n1141) );
  AND U1168 ( .A(n1156), .B(n1157), .Z(n1155) );
  XOR U1169 ( .A(n1150), .B(n1158), .Z(n1157) );
  XNOR U1170 ( .A(n1152), .B(n1154), .Z(n1158) );
  NAND U1171 ( .A(n513), .B(n1022), .Z(n1152) );
  XOR U1172 ( .A(n1149), .B(n1159), .Z(n1150) );
  AND U1173 ( .A(n455), .B(e_input[0]), .Z(n1159) );
  XNOR U1174 ( .A(n1163), .B(n1160), .Z(n1162) );
  XOR U1175 ( .A(n1144), .B(n1164), .Z(n1156) );
  XNOR U1176 ( .A(n1146), .B(n1154), .Z(n1164) );
  NANDN U1177 ( .B(n639), .A(n677), .Z(n1146) );
  XOR U1178 ( .A(n1143), .B(n1165), .Z(n1144) );
  AND U1179 ( .A(n743), .B(n574), .Z(n1165) );
  XOR U1180 ( .A(n1166), .B(n1167), .Z(n1143) );
  AND U1181 ( .A(n1168), .B(n1169), .Z(n1167) );
  XNOR U1182 ( .A(n1170), .B(n1166), .Z(n1169) );
  XOR U1183 ( .A(n1171), .B(n1172), .Z(n1154) );
  AND U1184 ( .A(n1173), .B(n1174), .Z(n1172) );
  XOR U1185 ( .A(n1161), .B(n1175), .Z(n1174) );
  XNOR U1186 ( .A(n1163), .B(n1171), .Z(n1175) );
  NAND U1187 ( .A(n574), .B(n1022), .Z(n1163) );
  XOR U1188 ( .A(n1160), .B(n1176), .Z(n1161) );
  AND U1189 ( .A(n513), .B(e_input[0]), .Z(n1176) );
  XOR U1190 ( .A(n1177), .B(n1178), .Z(n1160) );
  AND U1191 ( .A(n1179), .B(n1180), .Z(n1178) );
  XNOR U1192 ( .A(n1181), .B(n1177), .Z(n1180) );
  XOR U1193 ( .A(n1168), .B(n1182), .Z(n1173) );
  XNOR U1194 ( .A(n1170), .B(n1171), .Z(n1182) );
  NANDN U1195 ( .B(n711), .A(n677), .Z(n1170) );
  XOR U1196 ( .A(n1166), .B(n1183), .Z(n1168) );
  ANDN U1197 ( .A(n743), .B(n639), .Z(n1183) );
  XNOR U1198 ( .A(n1187), .B(n1184), .Z(n1186) );
  XOR U1199 ( .A(n1188), .B(n1189), .Z(n1171) );
  AND U1200 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U1201 ( .A(n1179), .B(n1192), .Z(n1191) );
  XNOR U1202 ( .A(n1181), .B(n1188), .Z(n1192) );
  NANDN U1203 ( .B(n639), .A(n1022), .Z(n1181) );
  XOR U1204 ( .A(n1177), .B(n1193), .Z(n1179) );
  AND U1205 ( .A(n574), .B(e_input[0]), .Z(n1193) );
  XOR U1206 ( .A(n1185), .B(n1197), .Z(n1190) );
  XNOR U1207 ( .A(n1187), .B(n1188), .Z(n1197) );
  NAND U1208 ( .A(n677), .B(n782), .Z(n1187) );
  XOR U1209 ( .A(n1184), .B(n1198), .Z(n1185) );
  ANDN U1210 ( .A(n743), .B(n711), .Z(n1198) );
  XOR U1211 ( .A(n1199), .B(n1200), .Z(n1184) );
  ANDN U1212 ( .A(n1201), .B(n1202), .Z(n1200) );
  XNOR U1213 ( .A(n1203), .B(n1199), .Z(n1201) );
  NAND U1214 ( .A(n677), .B(n1005), .Z(n1203) );
  XNOR U1215 ( .A(n1199), .B(n1205), .Z(n1202) );
  AND U1216 ( .A(n782), .B(n743), .Z(n1205) );
  AND U1217 ( .A(n1206), .B(g_input[0]), .Z(n1199) );
  NANDN U1218 ( .B(n677), .A(n1207), .Z(n1206) );
  NAND U1219 ( .A(n1005), .B(n743), .Z(n1207) );
  XNOR U1220 ( .A(n1194), .B(n1211), .Z(n1195) );
  ANDN U1221 ( .A(e_input[0]), .B(n639), .Z(n1211) );
  XOR U1222 ( .A(n1214), .B(n1212), .Z(n1213) );
  ANDN U1223 ( .A(e_input[0]), .B(n711), .Z(n1214) );
  AND U1224 ( .A(n1022), .B(n782), .Z(n1215) );
  XOR U1225 ( .A(n1219), .B(n1196), .Z(n1210) );
  NANDN U1226 ( .B(n711), .A(n1022), .Z(n1196) );
  IV U1227 ( .A(n1204), .Z(n1219) );
  NAND U1228 ( .A(n1022), .B(n1005), .Z(n1218) );
  XNOR U1229 ( .A(n1216), .B(n1220), .Z(n1217) );
  AND U1230 ( .A(n782), .B(e_input[0]), .Z(n1220) );
  AND U1231 ( .A(n1221), .B(g_input[0]), .Z(n1216) );
  NANDN U1232 ( .B(n1022), .A(n1222), .Z(n1221) );
  NAND U1233 ( .A(n1005), .B(e_input[0]), .Z(n1222) );
  XNOR U1234 ( .A(n1224), .B(n770), .Z(n758) );
  XNOR U1235 ( .A(n755), .B(n756), .Z(n770) );
  NAND U1236 ( .A(n250), .B(n574), .Z(n756) );
  XNOR U1237 ( .A(n754), .B(n1225), .Z(n755) );
  AND U1238 ( .A(n513), .B(n286), .Z(n1225) );
  XNOR U1239 ( .A(n1229), .B(n1226), .Z(n1228) );
  XNOR U1240 ( .A(n769), .B(n757), .Z(n1224) );
  XOR U1241 ( .A(n1230), .B(n1231), .Z(n757) );
  XNOR U1242 ( .A(n762), .B(n1233), .Z(n765) );
  AND U1243 ( .A(n397), .B(n382), .Z(n1233) );
  XNOR U1244 ( .A(n1134), .B(g_input[8]), .Z(n1133) );
  NOR U1245 ( .A(n1234), .B(n1235), .Z(n1134) );
  XOR U1246 ( .A(n1236), .B(n1237), .Z(n762) );
  AND U1247 ( .A(n1238), .B(n1239), .Z(n1237) );
  XNOR U1248 ( .A(n1240), .B(n1236), .Z(n1239) );
  XOR U1249 ( .A(n1241), .B(n766), .Z(n1232) );
  NAND U1250 ( .A(n335), .B(n455), .Z(n766) );
  IV U1251 ( .A(n768), .Z(n1241) );
  XNOR U1252 ( .A(n1242), .B(n1243), .Z(n768) );
  AND U1253 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U1254 ( .A(n1238), .B(n1246), .Z(n1245) );
  XNOR U1255 ( .A(n1240), .B(n1242), .Z(n1246) );
  NAND U1256 ( .A(n335), .B(n513), .Z(n1240) );
  XOR U1257 ( .A(n1236), .B(n1247), .Z(n1238) );
  AND U1258 ( .A(n455), .B(n382), .Z(n1247) );
  XOR U1259 ( .A(n1234), .B(g_input[7]), .Z(n1235) );
  NANDN U1260 ( .B(n1248), .A(n1249), .Z(n1234) );
  XOR U1261 ( .A(n1250), .B(n1251), .Z(n1236) );
  AND U1262 ( .A(n1252), .B(n1253), .Z(n1251) );
  XNOR U1263 ( .A(n1254), .B(n1250), .Z(n1253) );
  XOR U1264 ( .A(n1227), .B(n1255), .Z(n1244) );
  XNOR U1265 ( .A(n1229), .B(n1242), .Z(n1255) );
  NANDN U1266 ( .B(n639), .A(n250), .Z(n1229) );
  XOR U1267 ( .A(n1226), .B(n1256), .Z(n1227) );
  AND U1268 ( .A(n574), .B(n286), .Z(n1256) );
  XOR U1269 ( .A(n1257), .B(n1258), .Z(n1226) );
  AND U1270 ( .A(n1259), .B(n1260), .Z(n1258) );
  XNOR U1271 ( .A(n1261), .B(n1257), .Z(n1260) );
  XOR U1272 ( .A(n1262), .B(n1263), .Z(n1242) );
  AND U1273 ( .A(n1264), .B(n1265), .Z(n1263) );
  XOR U1274 ( .A(n1252), .B(n1266), .Z(n1265) );
  XNOR U1275 ( .A(n1254), .B(n1262), .Z(n1266) );
  NAND U1276 ( .A(n335), .B(n574), .Z(n1254) );
  XOR U1277 ( .A(n1250), .B(n1267), .Z(n1252) );
  AND U1278 ( .A(n513), .B(n382), .Z(n1267) );
  XNOR U1279 ( .A(n1249), .B(g_input[6]), .Z(n1248) );
  NOR U1280 ( .A(n1268), .B(n1269), .Z(n1249) );
  XOR U1281 ( .A(n1270), .B(n1271), .Z(n1250) );
  AND U1282 ( .A(n1272), .B(n1273), .Z(n1271) );
  XNOR U1283 ( .A(n1274), .B(n1270), .Z(n1273) );
  XOR U1284 ( .A(n1259), .B(n1275), .Z(n1264) );
  XNOR U1285 ( .A(n1261), .B(n1262), .Z(n1275) );
  NANDN U1286 ( .B(n711), .A(n250), .Z(n1261) );
  XOR U1287 ( .A(n1257), .B(n1276), .Z(n1259) );
  ANDN U1288 ( .A(n286), .B(n639), .Z(n1276) );
  XNOR U1289 ( .A(n1280), .B(n1277), .Z(n1279) );
  XOR U1290 ( .A(n1281), .B(n1282), .Z(n1262) );
  AND U1291 ( .A(n1283), .B(n1284), .Z(n1282) );
  XOR U1292 ( .A(n1272), .B(n1285), .Z(n1284) );
  XNOR U1293 ( .A(n1274), .B(n1281), .Z(n1285) );
  NANDN U1294 ( .B(n639), .A(n335), .Z(n1274) );
  XOR U1295 ( .A(n1270), .B(n1286), .Z(n1272) );
  AND U1296 ( .A(n574), .B(n382), .Z(n1286) );
  XOR U1297 ( .A(n1268), .B(g_input[5]), .Z(n1269) );
  NANDN U1298 ( .B(n1287), .A(n1288), .Z(n1268) );
  XOR U1299 ( .A(n1289), .B(n1290), .Z(n1270) );
  ANDN U1300 ( .A(n1291), .B(n1292), .Z(n1290) );
  XNOR U1301 ( .A(n1293), .B(n1289), .Z(n1291) );
  XOR U1302 ( .A(n1278), .B(n1294), .Z(n1283) );
  XNOR U1303 ( .A(n1280), .B(n1281), .Z(n1294) );
  NAND U1304 ( .A(n250), .B(n782), .Z(n1280) );
  XOR U1305 ( .A(n1277), .B(n1295), .Z(n1278) );
  ANDN U1306 ( .A(n286), .B(n711), .Z(n1295) );
  NAND U1307 ( .A(n250), .B(n1005), .Z(n1298) );
  XNOR U1308 ( .A(n1296), .B(n1300), .Z(n1297) );
  AND U1309 ( .A(n782), .B(n286), .Z(n1300) );
  AND U1310 ( .A(n1301), .B(g_input[0]), .Z(n1296) );
  NANDN U1311 ( .B(n250), .A(n1302), .Z(n1301) );
  NAND U1312 ( .A(n1005), .B(n286), .Z(n1302) );
  XNOR U1313 ( .A(n1305), .B(n1306), .Z(n1231) );
  IV U1314 ( .A(n1292), .Z(n1306) );
  XNOR U1315 ( .A(n1289), .B(n1307), .Z(n1292) );
  ANDN U1316 ( .A(n382), .B(n639), .Z(n1307) );
  XOR U1317 ( .A(n1308), .B(n1309), .Z(n1289) );
  AND U1318 ( .A(n1310), .B(n1311), .Z(n1309) );
  XOR U1319 ( .A(n1312), .B(n1308), .Z(n1311) );
  ANDN U1320 ( .A(n382), .B(n711), .Z(n1312) );
  XOR U1321 ( .A(n1313), .B(n1308), .Z(n1310) );
  AND U1322 ( .A(n782), .B(n335), .Z(n1313) );
  XOR U1323 ( .A(n1314), .B(n1315), .Z(n1308) );
  ANDN U1324 ( .A(n1316), .B(n1317), .Z(n1315) );
  XNOR U1325 ( .A(n1318), .B(n1314), .Z(n1316) );
  XOR U1326 ( .A(n1319), .B(n1293), .Z(n1305) );
  NANDN U1327 ( .B(n711), .A(n335), .Z(n1293) );
  IV U1328 ( .A(n1299), .Z(n1319) );
  XOR U1329 ( .A(n1320), .B(n1318), .Z(n1299) );
  NAND U1330 ( .A(n335), .B(n1005), .Z(n1318) );
  IV U1331 ( .A(n1317), .Z(n1320) );
  XNOR U1332 ( .A(n1314), .B(n1321), .Z(n1317) );
  AND U1333 ( .A(n782), .B(n382), .Z(n1321) );
  AND U1334 ( .A(n1322), .B(g_input[0]), .Z(n1314) );
  NANDN U1335 ( .B(n335), .A(n1323), .Z(n1322) );
  NAND U1336 ( .A(n1005), .B(n382), .Z(n1323) );
  XNOR U1337 ( .A(n773), .B(n1327), .Z(n776) );
  ANDN U1338 ( .A(n223), .B(n639), .Z(n1327) );
  XNOR U1339 ( .A(n1288), .B(g_input[4]), .Z(n1287) );
  NOR U1340 ( .A(n1328), .B(n1329), .Z(n1288) );
  XOR U1341 ( .A(n1330), .B(n1331), .Z(n773) );
  AND U1342 ( .A(n1332), .B(n1333), .Z(n1331) );
  XOR U1343 ( .A(n1334), .B(n1330), .Z(n1333) );
  ANDN U1344 ( .A(n223), .B(n711), .Z(n1334) );
  XOR U1345 ( .A(n1335), .B(n1330), .Z(n1332) );
  AND U1346 ( .A(n782), .B(n188), .Z(n1335) );
  XOR U1347 ( .A(n1336), .B(n1337), .Z(n1330) );
  ANDN U1348 ( .A(n1338), .B(n1339), .Z(n1337) );
  XNOR U1349 ( .A(n1340), .B(n1336), .Z(n1338) );
  XOR U1350 ( .A(n1341), .B(n777), .Z(n1326) );
  NANDN U1351 ( .B(n711), .A(n188), .Z(n777) );
  NANDN U1352 ( .B(n1342), .A(n1343), .Z(n1328) );
  IV U1353 ( .A(n779), .Z(n1341) );
  XOR U1354 ( .A(n1344), .B(n1340), .Z(n779) );
  NAND U1355 ( .A(n188), .B(n1005), .Z(n1340) );
  IV U1356 ( .A(n1339), .Z(n1344) );
  XNOR U1357 ( .A(n1336), .B(n1345), .Z(n1339) );
  AND U1358 ( .A(n782), .B(n223), .Z(n1345) );
  AND U1359 ( .A(n1346), .B(g_input[0]), .Z(n1336) );
  NANDN U1360 ( .B(n188), .A(n1347), .Z(n1346) );
  NAND U1361 ( .A(n1005), .B(n223), .Z(n1347) );
  XNOR U1362 ( .A(n786), .B(n787), .Z(n781) );
  NANDN U1363 ( .B(n138), .A(n1005), .Z(n787) );
  XNOR U1364 ( .A(n785), .B(n1350), .Z(n786) );
  AND U1365 ( .A(n782), .B(n158), .Z(n1350) );
  XNOR U1366 ( .A(n1343), .B(g_input[2]), .Z(n1342) );
  AND U1367 ( .A(n1352), .B(g_input[0]), .Z(n785) );
  NAND U1368 ( .A(n1353), .B(n138), .Z(n1352) );
  NANDN U1369 ( .B(n1354), .A(n1355), .Z(n138) );
  ANDN U1370 ( .A(e_input[15]), .B(n1356), .Z(n1355) );
  NAND U1371 ( .A(n1005), .B(n158), .Z(n1353) );
  XOR U1372 ( .A(n1356), .B(e_input[14]), .Z(n1354) );
  OR U1373 ( .A(n1349), .B(n1357), .Z(n1356) );
  XOR U1374 ( .A(n1357), .B(e_input[13]), .Z(n1349) );
  OR U1375 ( .A(n1348), .B(n1358), .Z(n1357) );
  XOR U1376 ( .A(n1358), .B(e_input[12]), .Z(n1348) );
  OR U1377 ( .A(n1304), .B(n1359), .Z(n1358) );
  XOR U1378 ( .A(n1359), .B(e_input[11]), .Z(n1304) );
  OR U1379 ( .A(n1303), .B(n1360), .Z(n1359) );
  XOR U1380 ( .A(n1360), .B(e_input[10]), .Z(n1303) );
  OR U1381 ( .A(n1325), .B(n1361), .Z(n1360) );
  XOR U1382 ( .A(n1361), .B(e_input[9]), .Z(n1325) );
  OR U1383 ( .A(n1324), .B(n1362), .Z(n1361) );
  XOR U1384 ( .A(n1362), .B(e_input[8]), .Z(n1324) );
  OR U1385 ( .A(n1015), .B(n1363), .Z(n1362) );
  XOR U1386 ( .A(n1363), .B(e_input[7]), .Z(n1015) );
  OR U1387 ( .A(n1014), .B(n1364), .Z(n1363) );
  XOR U1388 ( .A(n1364), .B(e_input[6]), .Z(n1014) );
  OR U1389 ( .A(n1010), .B(n1365), .Z(n1364) );
  XOR U1390 ( .A(n1365), .B(e_input[5]), .Z(n1010) );
  OR U1391 ( .A(n1009), .B(n1366), .Z(n1365) );
  XOR U1392 ( .A(n1366), .B(e_input[4]), .Z(n1009) );
  OR U1393 ( .A(n1209), .B(n1367), .Z(n1366) );
  XOR U1394 ( .A(n1367), .B(e_input[3]), .Z(n1209) );
  OR U1395 ( .A(n1208), .B(n1368), .Z(n1367) );
  XOR U1396 ( .A(n1368), .B(e_input[2]), .Z(n1208) );
  NANDN U1397 ( .B(e_input[0]), .A(n1223), .Z(n1368) );
  XNOR U1398 ( .A(e_input[0]), .B(e_input[1]), .Z(n1223) );
  XOR U1399 ( .A(g_input[0]), .B(g_input[1]), .Z(n1351) );
  AND U1400 ( .A(n1369), .B(n1370), .Z(\_MxM/N17 ) );
  XOR U1401 ( .A(\_MxM/n[6] ), .B(\_MxM/add_43/carry[6] ), .Z(n1370) );
  AND U1402 ( .A(\_MxM/N9 ), .B(n1369), .Z(\_MxM/N16 ) );
  AND U1403 ( .A(\_MxM/N8 ), .B(n1369), .Z(\_MxM/N15 ) );
  AND U1404 ( .A(\_MxM/N7 ), .B(n1369), .Z(\_MxM/N14 ) );
  AND U1405 ( .A(\_MxM/N6 ), .B(n1369), .Z(\_MxM/N13 ) );
  AND U1406 ( .A(\_MxM/N5 ), .B(n1369), .Z(\_MxM/N12 ) );
  NAND U1407 ( .A(n1371), .B(n1372), .Z(n1369) );
  ANDN U1408 ( .A(n1373), .B(n104), .Z(n1372) );
  OR U1409 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n104) );
  NOR U1410 ( .A(\_MxM/N11 ), .B(\_MxM/n[2] ), .Z(n1373) );
  AND U1411 ( .A(\_MxM/n[6] ), .B(n1374), .Z(n1371) );
  AND U1412 ( .A(\_MxM/n[5] ), .B(\_MxM/n[1] ), .Z(n1374) );
  IV U1413 ( .A(\_MxM/n[0] ), .Z(\_MxM/N11 ) );
endmodule

