
module MAC_TG_N32 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MAC/_MULT/X__[0] , \_MAC/_MULT/A__[0] , n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236;
  wire   [31:0] o_reg;
  assign \_MAC/_MULT/X__[0]  = e_input[0];
  assign \_MAC/_MULT/A__[0]  = g_input[0];

  DFF \o_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[0])
         );
  DFF \o_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[1])
         );
  DFF \o_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[2])
         );
  DFF \o_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[3])
         );
  DFF \o_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[4])
         );
  DFF \o_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[5])
         );
  DFF \o_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[6])
         );
  DFF \o_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[7])
         );
  DFF \o_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[8])
         );
  DFF \o_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[9])
         );
  DFF \o_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[10]) );
  DFF \o_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[11]) );
  DFF \o_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[12]) );
  DFF \o_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[13]) );
  DFF \o_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[14]) );
  DFF \o_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[15]) );
  DFF \o_reg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[16]) );
  DFF \o_reg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[17]) );
  DFF \o_reg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[18]) );
  DFF \o_reg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[19]) );
  DFF \o_reg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[20]) );
  DFF \o_reg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[21]) );
  DFF \o_reg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[22]) );
  DFF \o_reg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[23]) );
  DFF \o_reg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[24]) );
  DFF \o_reg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[25]) );
  DFF \o_reg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[26]) );
  DFF \o_reg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[27]) );
  DFF \o_reg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[28]) );
  DFF \o_reg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[29]) );
  DFF \o_reg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[30]) );
  DFF \o_reg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[31]) );
  MUX U35 ( .IN0(n3766), .IN1(n3764), .SEL(n3765), .F(n3726) );
  MUX U36 ( .IN0(n4135), .IN1(n4133), .SEL(n4134), .F(n4116) );
  MUX U37 ( .IN0(n4538), .IN1(n33), .SEL(n4143), .F(n4525) );
  IV U38 ( .A(n4142), .Z(n33) );
  MUX U39 ( .IN0(n5013), .IN1(n34), .SEL(n4891), .F(n5000) );
  IV U40 ( .A(n4890), .Z(n34) );
  MUX U41 ( .IN0(n35), .IN1(n1982), .SEL(n1983), .F(n1881) );
  IV U42 ( .A(n1984), .Z(n35) );
  MUX U43 ( .IN0(n36), .IN1(n2943), .SEL(n2944), .F(n2819) );
  IV U44 ( .A(n2945), .Z(n36) );
  MUX U45 ( .IN0(n874), .IN1(n872), .SEL(n873), .F(n835) );
  MUX U46 ( .IN0(n903), .IN1(n905), .SEL(n904), .F(n863) );
  MUX U47 ( .IN0(n1411), .IN1(n1409), .SEL(n1410), .F(n1335) );
  MUX U48 ( .IN0(n1541), .IN1(n1543), .SEL(n1542), .F(n37) );
  IV U49 ( .A(n37), .Z(n1460) );
  MUX U50 ( .IN0(n1855), .IN1(n1853), .SEL(n1854), .F(n1756) );
  MUX U51 ( .IN0(n2316), .IN1(n2314), .SEL(n2315), .F(n2202) );
  MUX U52 ( .IN0(n2391), .IN1(n2389), .SEL(n2390), .F(n2273) );
  MUX U53 ( .IN0(n2693), .IN1(n38), .SEL(n2692), .F(n2561) );
  IV U54 ( .A(n2691), .Z(n38) );
  MUX U55 ( .IN0(n2712), .IN1(n2710), .SEL(n2711), .F(n2582) );
  MUX U56 ( .IN0(n3029), .IN1(n3027), .SEL(n3028), .F(n2889) );
  MUX U57 ( .IN0(n1097), .IN1(n1095), .SEL(n1096), .F(n1035) );
  MUX U58 ( .IN0(n1311), .IN1(n39), .SEL(n1310), .F(n1235) );
  IV U59 ( .A(n1309), .Z(n39) );
  MUX U60 ( .IN0(n1977), .IN1(n40), .SEL(n1978), .F(n1871) );
  IV U61 ( .A(n1979), .Z(n40) );
  MUX U62 ( .IN0(n41), .IN1(n2614), .SEL(n2615), .F(n2492) );
  IV U63 ( .A(n2616), .Z(n41) );
  XNOR U64 ( .A(n736), .B(n735), .Z(n733) );
  MUX U65 ( .IN0(n42), .IN1(n1168), .SEL(n1169), .F(n1106) );
  IV U66 ( .A(n1170), .Z(n42) );
  MUX U67 ( .IN0(n43), .IN1(n1529), .SEL(n1530), .F(n1443) );
  IV U68 ( .A(n1531), .Z(n43) );
  MUX U69 ( .IN0(n2327), .IN1(n2325), .SEL(n2326), .F(n2212) );
  OR U70 ( .A(n752), .B(n753), .Z(n730) );
  AND U71 ( .A(n843), .B(n844), .Z(n802) );
  MUX U72 ( .IN0(n934), .IN1(n44), .SEL(n933), .F(n890) );
  IV U73 ( .A(n932), .Z(n44) );
  MUX U74 ( .IN0(n1694), .IN1(n45), .SEL(n1695), .F(n1605) );
  IV U75 ( .A(n1696), .Z(n45) );
  MUX U76 ( .IN0(n2098), .IN1(n46), .SEL(n2099), .F(n1993) );
  IV U77 ( .A(n2100), .Z(n46) );
  OR U78 ( .A(n810), .B(n811), .Z(n779) );
  XNOR U79 ( .A(n3720), .B(n3685), .Z(n3689) );
  XNOR U80 ( .A(n4127), .B(n4113), .Z(n4117) );
  XOR U81 ( .A(n3741), .B(n3706), .Z(n3710) );
  MUX U82 ( .IN0(n4525), .IN1(n47), .SEL(n4126), .F(n4512) );
  IV U83 ( .A(n4125), .Z(n47) );
  XOR U84 ( .A(n4489), .B(n4490), .Z(n4091) );
  XOR U85 ( .A(n4476), .B(n4477), .Z(n4074) );
  MUX U86 ( .IN0(n3538), .IN1(n3536), .SEL(n3537), .F(n3498) );
  XNOR U87 ( .A(n4059), .B(n4045), .Z(n4049) );
  MUX U88 ( .IN0(n48), .IN1(n4626), .SEL(n4627), .F(n4615) );
  IV U89 ( .A(n4628), .Z(n48) );
  XOR U90 ( .A(n5005), .B(n4997), .Z(n4873) );
  MUX U91 ( .IN0(n4299), .IN1(n49), .SEL(n4300), .F(n4278) );
  IV U92 ( .A(n4301), .Z(n49) );
  MUX U93 ( .IN0(n4608), .IN1(n50), .SEL(n4266), .F(n4597) );
  IV U94 ( .A(n4264), .Z(n50) );
  MUX U95 ( .IN0(n51), .IN1(n4232), .SEL(n4233), .F(n4211) );
  IV U96 ( .A(n4234), .Z(n51) );
  MUX U97 ( .IN0(n4822), .IN1(n52), .SEL(n4823), .F(n4801) );
  IV U98 ( .A(n4824), .Z(n52) );
  XNOR U99 ( .A(n3974), .B(n3960), .Z(n3964) );
  XOR U100 ( .A(n4953), .B(n4945), .Z(n4789) );
  MUX U101 ( .IN0(n3272), .IN1(n3270), .SEL(n3271), .F(n3232) );
  XOR U102 ( .A(n4374), .B(n4363), .Z(n3922) );
  MUX U103 ( .IN0(n3911), .IN1(n3909), .SEL(n3910), .F(n3211) );
  MUX U104 ( .IN0(n53), .IN1(n919), .SEL(n920), .F(n877) );
  IV U105 ( .A(n921), .Z(n53) );
  MUX U106 ( .IN0(n54), .IN1(n910), .SEL(n911), .F(n868) );
  IV U107 ( .A(n912), .Z(n54) );
  MUX U108 ( .IN0(n55), .IN1(n1475), .SEL(n1476), .F(n1396) );
  IV U109 ( .A(n1477), .Z(n55) );
  MUX U110 ( .IN0(n56), .IN1(n1619), .SEL(n1620), .F(n1526) );
  IV U111 ( .A(n1621), .Z(n56) );
  MUX U112 ( .IN0(n57), .IN1(n1611), .SEL(n1612), .F(n1518) );
  IV U113 ( .A(n1613), .Z(n57) );
  MUX U114 ( .IN0(n58), .IN1(n2095), .SEL(n2096), .F(n1990) );
  IV U115 ( .A(n2097), .Z(n58) );
  MUX U116 ( .IN0(n59), .IN1(n2269), .SEL(n2270), .F(n2156) );
  IV U117 ( .A(n2271), .Z(n59) );
  MUX U118 ( .IN0(n60), .IN1(n2416), .SEL(n2417), .F(n2305) );
  IV U119 ( .A(n2418), .Z(n60) );
  MUX U120 ( .IN0(n61), .IN1(n2756), .SEL(n2757), .F(n2628) );
  IV U121 ( .A(n2758), .Z(n61) );
  XOR U122 ( .A(n3900), .B(n3901), .Z(n3917) );
  MUX U123 ( .IN0(n1007), .IN1(n1009), .SEL(n1008), .F(n949) );
  MUX U124 ( .IN0(n1018), .IN1(n1016), .SEL(n1017), .F(n958) );
  MUX U125 ( .IN0(n1256), .IN1(n1258), .SEL(n1257), .F(n1188) );
  MUX U126 ( .IN0(n1575), .IN1(n1573), .SEL(n1574), .F(n1488) );
  MUX U127 ( .IN0(n1639), .IN1(n1641), .SEL(n1640), .F(n1541) );
  MUX U128 ( .IN0(n1656), .IN1(n1658), .SEL(n1657), .F(n1564) );
  MUX U129 ( .IN0(n1805), .IN1(n1803), .SEL(n1804), .F(n1706) );
  MUX U130 ( .IN0(n1877), .IN1(n1875), .SEL(n1876), .F(n1784) );
  MUX U131 ( .IN0(n2057), .IN1(n2055), .SEL(n2056), .F(n1950) );
  MUX U132 ( .IN0(n2195), .IN1(n99), .SEL(n2194), .F(n2082) );
  MUX U133 ( .IN0(n2341), .IN1(n2339), .SEL(n2340), .F(n2223) );
  MUX U134 ( .IN0(n2431), .IN1(n2429), .SEL(n2430), .F(n2314) );
  MUX U135 ( .IN0(n2512), .IN1(n2510), .SEL(n2511), .F(n2389) );
  MUX U136 ( .IN0(n2792), .IN1(n2794), .SEL(n2793), .F(n2665) );
  MUX U137 ( .IN0(n2815), .IN1(n2813), .SEL(n2814), .F(n2691) );
  MUX U138 ( .IN0(n2841), .IN1(n2839), .SEL(n2840), .F(n2710) );
  MUX U139 ( .IN0(n2932), .IN1(n2930), .SEL(n2931), .F(n2801) );
  MUX U140 ( .IN0(n837), .IN1(n835), .SEL(n836), .F(n794) );
  MUX U141 ( .IN0(n62), .IN1(n898), .SEL(n899), .F(n860) );
  IV U142 ( .A(n900), .Z(n62) );
  MUX U143 ( .IN0(n63), .IN1(n1116), .SEL(n1117), .F(n1056) );
  IV U144 ( .A(n1118), .Z(n63) );
  MUX U145 ( .IN0(n64), .IN1(n1380), .SEL(n1381), .F(n1309) );
  IV U146 ( .A(n1382), .Z(n64) );
  MUX U147 ( .IN0(n65), .IN1(n1391), .SEL(n1392), .F(n1317) );
  IV U148 ( .A(n1393), .Z(n65) );
  MUX U149 ( .IN0(n2079), .IN1(n66), .SEL(n2080), .F(n1977) );
  IV U150 ( .A(n2081), .Z(n66) );
  MUX U151 ( .IN0(n67), .IN1(n2871), .SEL(n2872), .F(n2742) );
  IV U152 ( .A(n2873), .Z(n67) );
  MUX U153 ( .IN0(n68), .IN1(n989), .SEL(n990), .F(n932) );
  IV U154 ( .A(n991), .Z(n68) );
  OR U155 ( .A(n1109), .B(n1110), .Z(n1049) );
  MUX U156 ( .IN0(n69), .IN1(n1230), .SEL(n1231), .F(n1168) );
  IV U157 ( .A(n1232), .Z(n69) );
  MUX U158 ( .IN0(n70), .IN1(n1907), .SEL(n1908), .F(n1810) );
  IV U159 ( .A(n1909), .Z(n70) );
  MUX U160 ( .IN0(n2452), .IN1(n2450), .SEL(n2451), .F(n2325) );
  OR U161 ( .A(n732), .B(n733), .Z(n712) );
  OR U162 ( .A(n781), .B(n782), .Z(n752) );
  AND U163 ( .A(n880), .B(n881), .Z(n843) );
  AND U164 ( .A(n1142), .B(n1143), .Z(n1082) );
  MUX U165 ( .IN0(n71), .IN1(n1607), .SEL(n1606), .F(n1512) );
  IV U166 ( .A(n1605), .Z(n71) );
  NANDN U167 ( .B(n1794), .A(n1795), .Z(n1697) );
  MUX U168 ( .IN0(n2209), .IN1(n72), .SEL(n2210), .F(n2098) );
  IV U169 ( .A(n2211), .Z(n72) );
  OR U170 ( .A(n851), .B(n852), .Z(n810) );
  OR U171 ( .A(n1090), .B(n1091), .Z(n1032) );
  MUX U172 ( .IN0(n73), .IN1(n773), .SEL(n774), .F(n744) );
  IV U173 ( .A(o_reg[28]), .Z(n73) );
  MUX U174 ( .IN0(n74), .IN1(n4540), .SEL(n4541), .F(n4527) );
  IV U175 ( .A(n4542), .Z(n74) );
  XOR U176 ( .A(n4530), .B(n4522), .Z(n4126) );
  MUX U177 ( .IN0(n75), .IN1(n3667), .SEL(n3668), .F(n3629) );
  IV U178 ( .A(n3669), .Z(n75) );
  MUX U179 ( .IN0(n3652), .IN1(n3650), .SEL(n3651), .F(n3612) );
  XNOR U180 ( .A(n4110), .B(n4096), .Z(n4100) );
  XOR U181 ( .A(n4491), .B(n4483), .Z(n4075) );
  XOR U182 ( .A(n4463), .B(n4464), .Z(n4057) );
  MUX U183 ( .IN0(n3557), .IN1(n3559), .SEL(n3558), .F(n3519) );
  XOR U184 ( .A(n4450), .B(n4451), .Z(n4040) );
  MUX U185 ( .IN0(n3500), .IN1(n3498), .SEL(n3499), .F(n3460) );
  XNOR U186 ( .A(n4042), .B(n4028), .Z(n4032) );
  MUX U187 ( .IN0(n4641), .IN1(n76), .SEL(n4326), .F(n4630) );
  IV U188 ( .A(n4325), .Z(n76) );
  MUX U189 ( .IN0(n4322), .IN1(n4320), .SEL(n4321), .F(n4299) );
  MUX U190 ( .IN0(n4887), .IN1(n4885), .SEL(n4886), .F(n4864) );
  MUX U191 ( .IN0(n77), .IN1(n4615), .SEL(n4616), .F(n4604) );
  IV U192 ( .A(n4617), .Z(n77) );
  MUX U193 ( .IN0(n5000), .IN1(n78), .SEL(n4873), .F(n4987) );
  IV U194 ( .A(n4871), .Z(n78) );
  XOR U195 ( .A(n4426), .B(n4418), .Z(n3990) );
  XNOR U196 ( .A(n3991), .B(n3977), .Z(n3981) );
  XOR U197 ( .A(n4398), .B(n4399), .Z(n3972) );
  MUX U198 ( .IN0(n3348), .IN1(n3346), .SEL(n3347), .F(n3308) );
  MUX U199 ( .IN0(n4597), .IN1(n79), .SEL(n4245), .F(n4586) );
  IV U200 ( .A(n4243), .Z(n79) );
  MUX U201 ( .IN0(n4236), .IN1(n80), .SEL(n4237), .F(n4215) );
  IV U202 ( .A(n4238), .Z(n80) );
  XOR U203 ( .A(n4385), .B(n4386), .Z(n3955) );
  MUX U204 ( .IN0(n3329), .IN1(n3331), .SEL(n3330), .F(n3291) );
  MUX U205 ( .IN0(n4780), .IN1(n81), .SEL(n4781), .F(n4759) );
  IV U206 ( .A(n4782), .Z(n81) );
  MUX U207 ( .IN0(n3931), .IN1(n3929), .SEL(n3930), .F(n3909) );
  XOR U208 ( .A(n4367), .B(n4368), .Z(n3921) );
  XOR U209 ( .A(n4927), .B(n4919), .Z(n4747) );
  XOR U210 ( .A(n4732), .B(n4733), .Z(n4729) );
  MUX U211 ( .IN0(n82), .IN1(n3182), .SEL(n3183), .F(n3053) );
  IV U212 ( .A(n3184), .Z(n82) );
  MUX U213 ( .IN0(n83), .IN1(n3207), .SEL(n3208), .F(n3079) );
  IV U214 ( .A(n3209), .Z(n83) );
  MUX U215 ( .IN0(n84), .IN1(n1121), .SEL(n1122), .F(n1061) );
  IV U216 ( .A(n1123), .Z(n84) );
  MUX U217 ( .IN0(n85), .IN1(n1130), .SEL(n1131), .F(n1070) );
  IV U218 ( .A(n1132), .Z(n85) );
  MUX U219 ( .IN0(n86), .IN1(n1484), .SEL(n1485), .F(n1405) );
  IV U220 ( .A(n1486), .Z(n86) );
  MUX U221 ( .IN0(n87), .IN1(n1849), .SEL(n1850), .F(n1752) );
  IV U222 ( .A(n1851), .Z(n87) );
  MUX U223 ( .IN0(n88), .IN1(n1799), .SEL(n1800), .F(n1702) );
  IV U224 ( .A(n1801), .Z(n88) );
  MUX U225 ( .IN0(n89), .IN1(n1920), .SEL(n1921), .F(n1823) );
  IV U226 ( .A(n1922), .Z(n89) );
  MUX U227 ( .IN0(n90), .IN1(n1937), .SEL(n1938), .F(n1840) );
  IV U228 ( .A(n1939), .Z(n90) );
  MUX U229 ( .IN0(n91), .IN1(n2219), .SEL(n2220), .F(n2106) );
  IV U230 ( .A(n2221), .Z(n91) );
  MUX U231 ( .IN0(n92), .IN1(n2310), .SEL(n2311), .F(n2198) );
  IV U232 ( .A(n2312), .Z(n92) );
  MUX U233 ( .IN0(n93), .IN1(n2359), .SEL(n2360), .F(n2243) );
  IV U234 ( .A(n2361), .Z(n93) );
  MUX U235 ( .IN0(n94), .IN1(n2376), .SEL(n2377), .F(n2260) );
  IV U236 ( .A(n2378), .Z(n94) );
  MUX U237 ( .IN0(n95), .IN1(n2661), .SEL(n2662), .F(n2537) );
  IV U238 ( .A(n2663), .Z(n95) );
  MUX U239 ( .IN0(n96), .IN1(n2797), .SEL(n2798), .F(n2670) );
  IV U240 ( .A(n2799), .Z(n96) );
  MUX U241 ( .IN0(n97), .IN1(n2859), .SEL(n2860), .F(n2730) );
  IV U242 ( .A(n2861), .Z(n97) );
  MUX U243 ( .IN0(n98), .IN1(n2876), .SEL(n2877), .F(n2747) );
  IV U244 ( .A(n2878), .Z(n98) );
  MUX U245 ( .IN0(n960), .IN1(n958), .SEL(n959), .F(n914) );
  MUX U246 ( .IN0(n949), .IN1(n951), .SEL(n950), .F(n903) );
  MUX U247 ( .IN0(n1267), .IN1(n1265), .SEL(n1266), .F(n1197) );
  MUX U248 ( .IN0(n1225), .IN1(n1223), .SEL(n1224), .F(n1159) );
  MUX U249 ( .IN0(n1479), .IN1(n1481), .SEL(n1480), .F(n1400) );
  MUX U250 ( .IN0(n1524), .IN1(n1522), .SEL(n1523), .F(n1436) );
  MUX U251 ( .IN0(n1667), .IN1(n1665), .SEL(n1666), .F(n1573) );
  MUX U252 ( .IN0(n1730), .IN1(n1732), .SEL(n1731), .F(n1639) );
  MUX U253 ( .IN0(n1988), .IN1(n1986), .SEL(n1987), .F(n1875) );
  MUX U254 ( .IN0(n2007), .IN1(n2005), .SEL(n2006), .F(n1900) );
  MUX U255 ( .IN0(n2275), .IN1(n2273), .SEL(n2274), .F(n2160) );
  MUX U256 ( .IN0(n2299), .IN1(n2301), .SEL(n2300), .F(n99) );
  IV U257 ( .A(n99), .Z(n2193) );
  MUX U258 ( .IN0(n2462), .IN1(n2460), .SEL(n2461), .F(n2339) );
  MUX U259 ( .IN0(n2552), .IN1(n2550), .SEL(n2551), .F(n2429) );
  MUX U260 ( .IN0(n2762), .IN1(n2760), .SEL(n2761), .F(n2632) );
  MUX U261 ( .IN0(n2949), .IN1(n2947), .SEL(n2948), .F(n2813) );
  MUX U262 ( .IN0(n3068), .IN1(n3066), .SEL(n3067), .F(n2930) );
  XOR U263 ( .A(n429), .B(n4349), .Z(n3103) );
  MUX U264 ( .IN0(n827), .IN1(n100), .SEL(n826), .F(n783) );
  IV U265 ( .A(n825), .Z(n100) );
  MUX U266 ( .IN0(n101), .IN1(n1056), .SEL(n1057), .F(n997) );
  IV U267 ( .A(n1058), .Z(n101) );
  OR U268 ( .A(n1302), .B(n1303), .Z(n1240) );
  MUX U269 ( .IN0(n102), .IN1(n1738), .SEL(n1739), .F(n1647) );
  IV U270 ( .A(n1740), .Z(n102) );
  MUX U271 ( .IN0(n2184), .IN1(n103), .SEL(n2185), .F(n2079) );
  IV U272 ( .A(n2186), .Z(n103) );
  MUX U273 ( .IN0(n2725), .IN1(n104), .SEL(n2726), .F(n2597) );
  IV U274 ( .A(n2727), .Z(n104) );
  MUX U275 ( .IN0(n105), .IN1(n2783), .SEL(n2784), .F(n2656) );
  IV U276 ( .A(n2785), .Z(n105) );
  MUX U277 ( .IN0(n106), .IN1(n3009), .SEL(n3010), .F(n2871) );
  IV U278 ( .A(n3011), .Z(n106) );
  XNOR U279 ( .A(n788), .B(n763), .Z(n761) );
  NOR U280 ( .A(n1049), .B(n1050), .Z(n980) );
  MUX U281 ( .IN0(n107), .IN1(n1106), .SEL(n1107), .F(n1044) );
  IV U282 ( .A(n1108), .Z(n107) );
  MUX U283 ( .IN0(n108), .IN1(n1370), .SEL(n1371), .F(n1298) );
  IV U284 ( .A(n1372), .Z(n108) );
  MUX U285 ( .IN0(n2574), .IN1(n2572), .SEL(n2573), .F(n2450) );
  AND U286 ( .A(n922), .B(n923), .Z(n880) );
  ANDN U287 ( .A(n1344), .B(n1345), .Z(n1274) );
  MUX U288 ( .IN0(n1512), .IN1(n1514), .SEL(n1513), .F(n1426) );
  MUX U289 ( .IN0(n1888), .IN1(n109), .SEL(n1889), .F(n1791) );
  IV U290 ( .A(n1890), .Z(n109) );
  ANDN U291 ( .A(n1959), .B(n1960), .Z(n1862) );
  MUX U292 ( .IN0(n2321), .IN1(n110), .SEL(n2322), .F(n2209) );
  IV U293 ( .A(n2323), .Z(n110) );
  ANDN U294 ( .A(n711), .B(n710), .Z(n709) );
  OR U295 ( .A(n750), .B(n751), .Z(n728) );
  OR U296 ( .A(n888), .B(n889), .Z(n851) );
  OR U297 ( .A(n1213), .B(n1214), .Z(n1151) );
  NAND U298 ( .A(n699), .B(n700), .Z(n698) );
  MUX U299 ( .IN0(n111), .IN1(n804), .SEL(n805), .F(n773) );
  IV U300 ( .A(o_reg[27]), .Z(n111) );
  MUX U301 ( .IN0(n112), .IN1(n968), .SEL(n969), .F(n924) );
  IV U302 ( .A(o_reg[23]), .Z(n112) );
  MUX U303 ( .IN0(n113), .IN1(n4146), .SEL(n4147), .F(n4129) );
  IV U304 ( .A(n4148), .Z(n113) );
  MUX U305 ( .IN0(n114), .IN1(n3773), .SEL(n3774), .F(n3735) );
  IV U306 ( .A(n3775), .Z(n114) );
  MUX U307 ( .IN0(n115), .IN1(n3781), .SEL(n3782), .F(n3743) );
  IV U308 ( .A(n3783), .Z(n115) );
  XOR U309 ( .A(n4543), .B(n4535), .Z(n4143) );
  MUX U310 ( .IN0(n116), .IN1(n4527), .SEL(n4528), .F(n4514) );
  IV U311 ( .A(n4529), .Z(n116) );
  MUX U312 ( .IN0(n117), .IN1(n3776), .SEL(n3777), .F(n3738) );
  IV U313 ( .A(n3778), .Z(n117) );
  MUX U314 ( .IN0(n3690), .IN1(n3688), .SEL(n3689), .F(n3650) );
  MUX U315 ( .IN0(n3709), .IN1(n3711), .SEL(n3710), .F(n3671) );
  MUX U316 ( .IN0(n118), .IN1(n3608), .SEL(n3609), .F(n3570) );
  IV U317 ( .A(n3610), .Z(n118) );
  MUX U318 ( .IN0(n119), .IN1(n3629), .SEL(n3630), .F(n3591) );
  IV U319 ( .A(n3631), .Z(n119) );
  XOR U320 ( .A(n4504), .B(n4496), .Z(n4092) );
  XNOR U321 ( .A(n4093), .B(n4079), .Z(n4083) );
  XOR U322 ( .A(n4465), .B(n4457), .Z(n4041) );
  MUX U323 ( .IN0(n120), .IN1(n5009), .SEL(n5010), .F(n4996) );
  IV U324 ( .A(n5011), .Z(n120) );
  XOR U325 ( .A(n3551), .B(n3516), .Z(n3520) );
  MUX U326 ( .IN0(n121), .IN1(n4621), .SEL(n4622), .F(n4610) );
  IV U327 ( .A(n4623), .Z(n121) );
  XOR U328 ( .A(n4437), .B(n4438), .Z(n4023) );
  MUX U329 ( .IN0(n122), .IN1(n3426), .SEL(n3427), .F(n3388) );
  IV U330 ( .A(n3428), .Z(n122) );
  XNOR U331 ( .A(n4025), .B(n4011), .Z(n4015) );
  XNOR U332 ( .A(n3454), .B(n3419), .Z(n3423) );
  XOR U333 ( .A(n4624), .B(n4616), .Z(n4287) );
  XOR U334 ( .A(n4879), .B(n4861), .Z(n4865) );
  XOR U335 ( .A(n4293), .B(n4275), .Z(n4279) );
  MUX U336 ( .IN0(n4987), .IN1(n123), .SEL(n4852), .F(n4974) );
  IV U337 ( .A(n4850), .Z(n123) );
  XOR U338 ( .A(n3437), .B(n3402), .Z(n3406) );
  XOR U339 ( .A(n4413), .B(n4405), .Z(n3973) );
  MUX U340 ( .IN0(n124), .IN1(n5154), .SEL(n5155), .F(n5136) );
  IV U341 ( .A(n5156), .Z(n124) );
  MUX U342 ( .IN0(n4801), .IN1(n125), .SEL(n4802), .F(n4780) );
  IV U343 ( .A(n4803), .Z(n125) );
  MUX U344 ( .IN0(n3310), .IN1(n3308), .SEL(n3309), .F(n3270) );
  MUX U345 ( .IN0(n3948), .IN1(n3946), .SEL(n3947), .F(n3929) );
  MUX U346 ( .IN0(n4586), .IN1(n126), .SEL(n4224), .F(n4575) );
  IV U347 ( .A(n4222), .Z(n126) );
  MUX U348 ( .IN0(n4215), .IN1(n127), .SEL(n4216), .F(n4194) );
  IV U349 ( .A(n4217), .Z(n127) );
  XOR U350 ( .A(n4940), .B(n4932), .Z(n4768) );
  XOR U351 ( .A(n4751), .B(n4752), .Z(n4761) );
  MUX U352 ( .IN0(n128), .IN1(n4755), .SEL(n4756), .F(n4723) );
  IV U353 ( .A(n4757), .Z(n128) );
  MUX U354 ( .IN0(n129), .IN1(n3228), .SEL(n3229), .F(n3191) );
  IV U355 ( .A(n3230), .Z(n129) );
  MUX U356 ( .IN0(n130), .IN1(n4738), .SEL(n4739), .F(n3124) );
  IV U357 ( .A(n4740), .Z(n130) );
  MUX U358 ( .IN0(n3253), .IN1(n3255), .SEL(n3254), .F(n3186) );
  MUX U359 ( .IN0(n131), .IN1(n954), .SEL(n955), .F(n910) );
  IV U360 ( .A(n956), .Z(n131) );
  MUX U361 ( .IN0(n132), .IN1(n1184), .SEL(n1185), .F(n1121) );
  IV U362 ( .A(n1186), .Z(n132) );
  MUX U363 ( .IN0(n133), .IN1(n1357), .SEL(n1358), .F(n1287) );
  IV U364 ( .A(n1359), .Z(n133) );
  MUX U365 ( .IN0(n134), .IN1(n1661), .SEL(n1662), .F(n1569) );
  IV U366 ( .A(n1663), .Z(n134) );
  MUX U367 ( .IN0(n135), .IN1(n1823), .SEL(n1824), .F(n1726) );
  IV U368 ( .A(n1825), .Z(n135) );
  MUX U369 ( .IN0(n136), .IN1(n2235), .SEL(n2236), .F(n2122) );
  IV U370 ( .A(n2237), .Z(n136) );
  MUX U371 ( .IN0(n137), .IN1(n2243), .SEL(n2244), .F(n2130) );
  IV U372 ( .A(n2245), .Z(n137) );
  MUX U373 ( .IN0(n138), .IN1(n2456), .SEL(n2457), .F(n2335) );
  IV U374 ( .A(n2458), .Z(n138) );
  MUX U375 ( .IN0(n139), .IN1(n2670), .SEL(n2671), .F(n2546) );
  IV U376 ( .A(n2672), .Z(n139) );
  MUX U377 ( .IN0(n140), .IN1(n2722), .SEL(n2723), .F(n2594) );
  IV U378 ( .A(n2724), .Z(n140) );
  MUX U379 ( .IN0(n141), .IN1(n2730), .SEL(n2731), .F(n2602) );
  IV U380 ( .A(n2732), .Z(n141) );
  MUX U381 ( .IN0(n142), .IN1(n2917), .SEL(n2918), .F(n2788) );
  IV U382 ( .A(n2919), .Z(n142) );
  MUX U383 ( .IN0(n143), .IN1(n3921), .SEL(n3922), .F(n4355) );
  IV U384 ( .A(n4369), .Z(n143) );
  MUX U385 ( .IN0(n1076), .IN1(n1074), .SEL(n1075), .F(n1016) );
  MUX U386 ( .IN0(n1065), .IN1(n1067), .SEL(n1066), .F(n1007) );
  MUX U387 ( .IN0(n1337), .IN1(n1335), .SEL(n1336), .F(n1265) );
  MUX U388 ( .IN0(n1400), .IN1(n1402), .SEL(n1401), .F(n1326) );
  MUX U389 ( .IN0(n1708), .IN1(n1706), .SEL(n1707), .F(n1615) );
  MUX U390 ( .IN0(n1844), .IN1(n1846), .SEL(n1845), .F(n1747) );
  MUX U391 ( .IN0(n2029), .IN1(n2031), .SEL(n2030), .F(n1924) );
  MUX U392 ( .IN0(n2093), .IN1(n2091), .SEL(n2092), .F(n1986) );
  MUX U393 ( .IN0(n2112), .IN1(n2110), .SEL(n2111), .F(n2005) );
  MUX U394 ( .IN0(n2264), .IN1(n2266), .SEL(n2265), .F(n2151) );
  MUX U395 ( .IN0(n2420), .IN1(n2422), .SEL(n2421), .F(n2299) );
  MUX U396 ( .IN0(n2484), .IN1(n2486), .SEL(n2485), .F(n2363) );
  MUX U397 ( .IN0(n2569), .IN1(n144), .SEL(n2568), .F(n2446) );
  IV U398 ( .A(n2567), .Z(n144) );
  MUX U399 ( .IN0(n2751), .IN1(n2753), .SEL(n2752), .F(n2623) );
  MUX U400 ( .IN0(n2803), .IN1(n2801), .SEL(n2802), .F(n2674) );
  MUX U401 ( .IN0(n2891), .IN1(n2889), .SEL(n2890), .F(n2760) );
  MUX U402 ( .IN0(n3001), .IN1(n3003), .SEL(n3002), .F(n2863) );
  MUX U403 ( .IN0(n2979), .IN1(n2977), .SEL(n2978), .F(n2839) );
  MUX U404 ( .IN0(n3085), .IN1(n3083), .SEL(n3084), .F(n2947) );
  XOR U405 ( .A(n3098), .B(n3099), .Z(n3104) );
  MUX U406 ( .IN0(n145), .IN1(n840), .SEL(n841), .F(n799) );
  IV U407 ( .A(n842), .Z(n145) );
  AND U408 ( .A(n822), .B(n818), .Z(n821) );
  XNOR U409 ( .A(n828), .B(n790), .Z(n795) );
  MUX U410 ( .IN0(n146), .IN1(n860), .SEL(n861), .F(n825) );
  IV U411 ( .A(n862), .Z(n146) );
  OR U412 ( .A(n1099), .B(n1100), .Z(n1093) );
  MUX U413 ( .IN0(n147), .IN1(n1179), .SEL(n1180), .F(n1116) );
  IV U414 ( .A(n1181), .Z(n147) );
  MUX U415 ( .IN0(n148), .IN1(n1383), .SEL(n1384), .F(n1302) );
  IV U416 ( .A(n1385), .Z(n148) );
  MUX U417 ( .IN0(n149), .IN1(n1451), .SEL(n1452), .F(n1380) );
  IV U418 ( .A(n1453), .Z(n149) );
  MUX U419 ( .IN0(n150), .IN1(n1470), .SEL(n1471), .F(n1391) );
  IV U420 ( .A(n1472), .Z(n150) );
  MUX U421 ( .IN0(n1818), .IN1(n151), .SEL(n1819), .F(n1721) );
  IV U422 ( .A(n1820), .Z(n151) );
  XNOR U423 ( .A(n1944), .B(n1850), .Z(n1854) );
  MUX U424 ( .IN0(n152), .IN1(n2037), .SEL(n2038), .F(n1932) );
  IV U425 ( .A(n2039), .Z(n152) );
  XNOR U426 ( .A(n2267), .B(n2157), .Z(n2163) );
  MUX U427 ( .IN0(n153), .IN1(n2295), .SEL(n2296), .F(n2184) );
  IV U428 ( .A(n2297), .Z(n153) );
  MUX U429 ( .IN0(n2354), .IN1(n154), .SEL(n2355), .F(n2238) );
  IV U430 ( .A(n2356), .Z(n154) );
  MUX U431 ( .IN0(n155), .IN1(n2492), .SEL(n2493), .F(n2371) );
  IV U432 ( .A(n2494), .Z(n155) );
  MUX U433 ( .IN0(n156), .IN1(n2912), .SEL(n2913), .F(n2783) );
  IV U434 ( .A(n2914), .Z(n156) );
  MUX U435 ( .IN0(n157), .IN1(n3144), .SEL(n3145), .F(n3009) );
  IV U436 ( .A(n3146), .Z(n157) );
  MUX U437 ( .IN0(n1171), .IN1(n1173), .SEL(n1172), .F(n1109) );
  MUX U438 ( .IN0(n1687), .IN1(n1685), .SEL(n1686), .F(n1602) );
  MUX U439 ( .IN0(n158), .IN1(n2230), .SEL(n2231), .F(n2117) );
  IV U440 ( .A(n2232), .Z(n158) );
  MUX U441 ( .IN0(n2702), .IN1(n159), .SEL(n2701), .F(n2572) );
  IV U442 ( .A(n2700), .Z(n159) );
  MUX U443 ( .IN0(n160), .IN1(n2717), .SEL(n2718), .F(n2589) );
  IV U444 ( .A(n2719), .Z(n160) );
  XNOR U445 ( .A(n717), .B(n716), .Z(n713) );
  OR U446 ( .A(n890), .B(n891), .Z(n853) );
  AND U447 ( .A(n1024), .B(n1025), .Z(n966) );
  ANDN U448 ( .A(n1582), .B(n1583), .Z(n1497) );
  NANDN U449 ( .B(n1697), .A(n1698), .Z(n1591) );
  MUX U450 ( .IN0(n1791), .IN1(n161), .SEL(n1792), .F(n1694) );
  IV U451 ( .A(n1793), .Z(n161) );
  NANDN U452 ( .B(n2101), .A(n2102), .Z(n1996) );
  ANDN U453 ( .A(n2171), .B(n2172), .Z(n2064) );
  MUX U454 ( .IN0(n2436), .IN1(n162), .SEL(n2437), .F(n2321) );
  IV U455 ( .A(n2438), .Z(n162) );
  OR U456 ( .A(n730), .B(n731), .Z(n710) );
  OR U457 ( .A(n779), .B(n780), .Z(n750) );
  OR U458 ( .A(n930), .B(n931), .Z(n888) );
  OR U459 ( .A(n1151), .B(n1152), .Z(n1090) );
  MUX U460 ( .IN0(n1428), .IN1(n1426), .SEL(n1427), .F(n1352) );
  MUX U461 ( .IN0(n163), .IN1(n691), .SEL(n692), .F(n689) );
  IV U462 ( .A(o_reg[30]), .Z(n163) );
  MUX U463 ( .IN0(n164), .IN1(n845), .SEL(n846), .F(n804) );
  IV U464 ( .A(o_reg[26]), .Z(n164) );
  MUX U465 ( .IN0(n165), .IN1(n1084), .SEL(n1085), .F(n1026) );
  IV U466 ( .A(o_reg[21]), .Z(n165) );
  MUX U467 ( .IN0(n1346), .IN1(n166), .SEL(n1347), .F(n1276) );
  IV U468 ( .A(o_reg[17]), .Z(n166) );
  MUX U469 ( .IN0(n1676), .IN1(n167), .SEL(n1677), .F(n1584) );
  IV U470 ( .A(o_reg[13]), .Z(n167) );
  MUX U471 ( .IN0(n2066), .IN1(n168), .SEL(n680), .F(n1961) );
  IV U472 ( .A(o_reg[9]), .Z(n168) );
  MUX U473 ( .IN0(n2521), .IN1(n169), .SEL(n684), .F(n2400) );
  IV U474 ( .A(o_reg[5]), .Z(n169) );
  MUX U475 ( .IN0(n170), .IN1(n3768), .SEL(n3769), .F(n3730) );
  IV U476 ( .A(n3770), .Z(n170) );
  MUX U477 ( .IN0(n3785), .IN1(n3787), .SEL(n3786), .F(n3747) );
  XNOR U478 ( .A(n4144), .B(n4130), .Z(n4134) );
  XOR U479 ( .A(n4515), .B(n4516), .Z(n4125) );
  MUX U480 ( .IN0(n171), .IN1(n4534), .SEL(n4535), .F(n4521) );
  IV U481 ( .A(n4536), .Z(n171) );
  MUX U482 ( .IN0(n3738), .IN1(n172), .SEL(n3739), .F(n3700) );
  IV U483 ( .A(n3740), .Z(n172) );
  XOR U484 ( .A(n4502), .B(n4503), .Z(n4108) );
  MUX U485 ( .IN0(n3614), .IN1(n3612), .SEL(n3613), .F(n3574) );
  XOR U486 ( .A(n3665), .B(n3630), .Z(n3634) );
  MUX U487 ( .IN0(n4084), .IN1(n4082), .SEL(n4083), .F(n4065) );
  MUX U488 ( .IN0(n173), .IN1(n3532), .SEL(n3533), .F(n3494) );
  IV U489 ( .A(n3534), .Z(n173) );
  XOR U490 ( .A(n4478), .B(n4470), .Z(n4058) );
  MUX U491 ( .IN0(n174), .IN1(n4316), .SEL(n4317), .F(n4295) );
  IV U492 ( .A(n4318), .Z(n174) );
  MUX U493 ( .IN0(n175), .IN1(n5002), .SEL(n5003), .F(n4989) );
  IV U494 ( .A(n5004), .Z(n175) );
  MUX U495 ( .IN0(n176), .IN1(n4881), .SEL(n4882), .F(n4860) );
  IV U496 ( .A(n4883), .Z(n176) );
  MUX U497 ( .IN0(n3519), .IN1(n3521), .SEL(n3520), .F(n3481) );
  MUX U498 ( .IN0(n177), .IN1(n3477), .SEL(n3478), .F(n3439) );
  IV U499 ( .A(n3479), .Z(n177) );
  MUX U500 ( .IN0(n178), .IN1(n4996), .SEL(n4997), .F(n4983) );
  IV U501 ( .A(n4998), .Z(n178) );
  MUX U502 ( .IN0(n3462), .IN1(n3460), .SEL(n3461), .F(n3422) );
  MUX U503 ( .IN0(n4016), .IN1(n4014), .SEL(n4015), .F(n3997) );
  MUX U504 ( .IN0(n4630), .IN1(n179), .SEL(n4308), .F(n4619) );
  IV U505 ( .A(n4306), .Z(n179) );
  MUX U506 ( .IN0(n180), .IN1(n4610), .SEL(n4611), .F(n4599) );
  IV U507 ( .A(n4612), .Z(n180) );
  XOR U508 ( .A(n4439), .B(n4431), .Z(n4007) );
  MUX U509 ( .IN0(n181), .IN1(n4423), .SEL(n4424), .F(n4410) );
  IV U510 ( .A(n4425), .Z(n181) );
  MUX U511 ( .IN0(n182), .IN1(n4888), .SEL(n4735), .F(n4867) );
  IV U512 ( .A(n4734), .Z(n182) );
  MUX U513 ( .IN0(n4864), .IN1(n183), .SEL(n4865), .F(n4843) );
  IV U514 ( .A(n4866), .Z(n183) );
  MUX U515 ( .IN0(n184), .IN1(n3380), .SEL(n3381), .F(n3342) );
  IV U516 ( .A(n3382), .Z(n184) );
  MUX U517 ( .IN0(n185), .IN1(n3984), .SEL(n3985), .F(n3967) );
  IV U518 ( .A(n3986), .Z(n185) );
  MUX U519 ( .IN0(n186), .IN1(n4697), .SEL(n4698), .F(n4682) );
  IV U520 ( .A(n4699), .Z(n186) );
  MUX U521 ( .IN0(n187), .IN1(n4692), .SEL(n4693), .F(n4676) );
  IV U522 ( .A(n4694), .Z(n187) );
  MUX U523 ( .IN0(n188), .IN1(n4604), .SEL(n4605), .F(n4593) );
  IV U524 ( .A(n4606), .Z(n188) );
  MUX U525 ( .IN0(n4278), .IN1(n189), .SEL(n4279), .F(n4257) );
  IV U526 ( .A(n4280), .Z(n189) );
  MUX U527 ( .IN0(n190), .IN1(n5069), .SEL(n5070), .F(n5054) );
  IV U528 ( .A(n5071), .Z(n190) );
  MUX U529 ( .IN0(n191), .IN1(n5064), .SEL(n5065), .F(n5048) );
  IV U530 ( .A(n5066), .Z(n191) );
  MUX U531 ( .IN0(n192), .IN1(n4813), .SEL(n4814), .F(n4792) );
  IV U532 ( .A(n4815), .Z(n192) );
  MUX U533 ( .IN0(n193), .IN1(n3845), .SEL(n3846), .F(n3829) );
  IV U534 ( .A(n3847), .Z(n193) );
  XOR U535 ( .A(n4228), .B(n4229), .Z(n4238) );
  XOR U536 ( .A(n4966), .B(n4958), .Z(n4810) );
  MUX U537 ( .IN0(n194), .IN1(n4797), .SEL(n4798), .F(n4776) );
  IV U538 ( .A(n4799), .Z(n194) );
  XOR U539 ( .A(n3399), .B(n3364), .Z(n3368) );
  XOR U540 ( .A(n4207), .B(n4208), .Z(n4217) );
  XOR U541 ( .A(n4400), .B(n4392), .Z(n3956) );
  MUX U542 ( .IN0(n195), .IN1(n5174), .SEL(n5175), .F(n5170) );
  IV U543 ( .A(n5176), .Z(n195) );
  MUX U544 ( .IN0(n196), .IN1(n4937), .SEL(n4938), .F(n4924) );
  IV U545 ( .A(n4939), .Z(n196) );
  XNOR U546 ( .A(n3957), .B(n3943), .Z(n3947) );
  MUX U547 ( .IN0(n197), .IN1(n3287), .SEL(n3288), .F(n3249) );
  IV U548 ( .A(n3289), .Z(n197) );
  XNOR U549 ( .A(n3302), .B(n3267), .Z(n3271) );
  XOR U550 ( .A(n4580), .B(n4572), .Z(n4203) );
  XOR U551 ( .A(n4186), .B(n4187), .Z(n4196) );
  MUX U552 ( .IN0(n198), .IN1(n4190), .SEL(n4191), .F(n4165) );
  IV U553 ( .A(n4192), .Z(n198) );
  MUX U554 ( .IN0(n199), .IN1(n963), .SEL(n964), .F(n919) );
  IV U555 ( .A(n965), .Z(n199) );
  MUX U556 ( .IN0(n200), .IN1(n1003), .SEL(n1004), .F(n944) );
  IV U557 ( .A(n1005), .Z(n200) );
  MUX U558 ( .IN0(n201), .IN1(n1012), .SEL(n1013), .F(n954) );
  IV U559 ( .A(n1014), .Z(n201) );
  MUX U560 ( .IN0(n202), .IN1(n1244), .SEL(n1245), .F(n1176) );
  IV U561 ( .A(n1246), .Z(n202) );
  MUX U562 ( .IN0(n203), .IN1(n1261), .SEL(n1262), .F(n1193) );
  IV U563 ( .A(n1263), .Z(n203) );
  MUX U564 ( .IN0(n204), .IN1(n1295), .SEL(n1296), .F(n1227) );
  IV U565 ( .A(n1297), .Z(n204) );
  MUX U566 ( .IN0(n205), .IN1(n1287), .SEL(n1288), .F(n1219) );
  IV U567 ( .A(n1289), .Z(n205) );
  MUX U568 ( .IN0(n206), .IN1(n1396), .SEL(n1397), .F(n1322) );
  IV U569 ( .A(n1398), .Z(n206) );
  MUX U570 ( .IN0(n207), .IN1(n1635), .SEL(n1636), .F(n1547) );
  IV U571 ( .A(n1637), .Z(n207) );
  MUX U572 ( .IN0(n208), .IN1(n1743), .SEL(n1744), .F(n1652) );
  IV U573 ( .A(n1745), .Z(n208) );
  MUX U574 ( .IN0(n209), .IN1(n1807), .SEL(n1808), .F(n1710) );
  IV U575 ( .A(n1809), .Z(n209) );
  MUX U576 ( .IN0(n210), .IN1(n1990), .SEL(n1991), .F(n1885) );
  IV U577 ( .A(n1992), .Z(n210) );
  MUX U578 ( .IN0(n211), .IN1(n2001), .SEL(n2002), .F(n1896) );
  IV U579 ( .A(n2003), .Z(n211) );
  MUX U580 ( .IN0(n212), .IN1(n2147), .SEL(n2148), .F(n2042) );
  IV U581 ( .A(n2149), .Z(n212) );
  MUX U582 ( .IN0(n213), .IN1(n2464), .SEL(n2465), .F(n2343) );
  IV U583 ( .A(n2466), .Z(n213) );
  MUX U584 ( .IN0(n214), .IN1(n2619), .SEL(n2620), .F(n2497) );
  IV U585 ( .A(n2621), .Z(n214) );
  MUX U586 ( .IN0(n215), .IN1(n2973), .SEL(n2974), .F(n2835) );
  IV U587 ( .A(n2975), .Z(n215) );
  MUX U588 ( .IN0(n216), .IN1(n3149), .SEL(n3150), .F(n3014) );
  IV U589 ( .A(n3151), .Z(n216) );
  MUX U590 ( .IN0(n217), .IN1(n3079), .SEL(n3080), .F(n2943) );
  IV U591 ( .A(n3081), .Z(n217) );
  NAND U592 ( .A(n4354), .B(n4358), .Z(n4357) );
  MUX U593 ( .IN0(n4922), .IN1(n218), .SEL(n4747), .F(n3136) );
  IV U594 ( .A(n4745), .Z(n218) );
  MUX U595 ( .IN0(n4727), .IN1(n219), .SEL(n4728), .F(n3112) );
  IV U596 ( .A(n4729), .Z(n219) );
  MUX U597 ( .IN0(n3213), .IN1(n3211), .SEL(n3212), .F(n3083) );
  MUX U598 ( .IN0(n1125), .IN1(n1127), .SEL(n1126), .F(n1065) );
  MUX U599 ( .IN0(n1136), .IN1(n1134), .SEL(n1135), .F(n1074) );
  MUX U600 ( .IN0(n1438), .IN1(n1436), .SEL(n1437), .F(n1361) );
  MUX U601 ( .IN0(n1490), .IN1(n1488), .SEL(n1489), .F(n1409) );
  MUX U602 ( .IN0(n1564), .IN1(n1566), .SEL(n1565), .F(n1479) );
  MUX U603 ( .IN0(n1827), .IN1(n1829), .SEL(n1828), .F(n1730) );
  MUX U604 ( .IN0(n1883), .IN1(n220), .SEL(n1882), .F(n1783) );
  IV U605 ( .A(n1881), .Z(n220) );
  MUX U606 ( .IN0(n1941), .IN1(n1943), .SEL(n1942), .F(n1844) );
  MUX U607 ( .IN0(n2204), .IN1(n2202), .SEL(n2203), .F(n2091) );
  MUX U608 ( .IN0(n2225), .IN1(n2223), .SEL(n2224), .F(n2110) );
  MUX U609 ( .IN0(n2247), .IN1(n2249), .SEL(n2248), .F(n2134) );
  MUX U610 ( .IN0(n2380), .IN1(n2382), .SEL(n2381), .F(n2264) );
  MUX U611 ( .IN0(n2541), .IN1(n2543), .SEL(n2542), .F(n2420) );
  MUX U612 ( .IN0(n2676), .IN1(n2674), .SEL(n2675), .F(n2550) );
  MUX U613 ( .IN0(n2734), .IN1(n2736), .SEL(n2735), .F(n2606) );
  MUX U614 ( .IN0(n2880), .IN1(n2882), .SEL(n2881), .F(n2751) );
  MUX U615 ( .IN0(n3057), .IN1(n3059), .SEL(n3058), .F(n2921) );
  XNOR U616 ( .A(n3189), .B(n3063), .Z(n3067) );
  XNOR U617 ( .A(n1095), .B(n1100), .Z(n1154) );
  MUX U618 ( .IN0(n221), .IN1(n1317), .SEL(n1318), .F(n1247) );
  IV U619 ( .A(n1319), .Z(n221) );
  MUX U620 ( .IN0(n1537), .IN1(n222), .SEL(n1538), .F(n1451) );
  IV U621 ( .A(n1539), .Z(n222) );
  MUX U622 ( .IN0(n223), .IN1(n1647), .SEL(n1648), .F(n1555) );
  IV U623 ( .A(n1649), .Z(n223) );
  XNOR U624 ( .A(n1847), .B(n1753), .Z(n1759) );
  XNOR U625 ( .A(n1797), .B(n1703), .Z(n1707) );
  MUX U626 ( .IN0(n2020), .IN1(n224), .SEL(n2021), .F(n1915) );
  IV U627 ( .A(n2022), .Z(n224) );
  MUX U628 ( .IN0(n225), .IN1(n2142), .SEL(n2143), .F(n2037) );
  IV U629 ( .A(n2144), .Z(n225) );
  XNOR U630 ( .A(n2383), .B(n2270), .Z(n2274) );
  MUX U631 ( .IN0(n2475), .IN1(n226), .SEL(n2476), .F(n2354) );
  IV U632 ( .A(n2477), .Z(n226) );
  MUX U633 ( .IN0(n2563), .IN1(n2561), .SEL(n2562), .F(n2449) );
  MUX U634 ( .IN0(n227), .IN1(n2742), .SEL(n2743), .F(n2614) );
  IV U635 ( .A(n2744), .Z(n227) );
  XNOR U636 ( .A(n2754), .B(n2629), .Z(n2633) );
  XNOR U637 ( .A(n2704), .B(n2579), .Z(n2583) );
  MUX U638 ( .IN0(n2992), .IN1(n228), .SEL(n2993), .F(n2854) );
  IV U639 ( .A(n2994), .Z(n228) );
  MUX U640 ( .IN0(n2969), .IN1(n229), .SEL(n2968), .F(n2829) );
  IV U641 ( .A(n2967), .Z(n229) );
  XNOR U642 ( .A(n3156), .B(n3024), .Z(n3028) );
  MUX U643 ( .IN0(n796), .IN1(n794), .SEL(n795), .F(n760) );
  MUX U644 ( .IN0(n791), .IN1(n230), .SEL(n790), .F(n763) );
  IV U645 ( .A(n789), .Z(n230) );
  XOR U646 ( .A(n783), .B(n823), .Z(n816) );
  MUX U647 ( .IN0(n231), .IN1(n1041), .SEL(n1042), .F(n986) );
  IV U648 ( .A(n1043), .Z(n231) );
  NANDN U649 ( .B(n1240), .A(n1241), .Z(n1233) );
  MUX U650 ( .IN0(n232), .IN1(n1443), .SEL(n1444), .F(n1370) );
  IV U651 ( .A(n1445), .Z(n232) );
  MUX U652 ( .IN0(n233), .IN1(n1810), .SEL(n1811), .F(n1713) );
  IV U653 ( .A(n1812), .Z(n233) );
  MUX U654 ( .IN0(n1871), .IN1(n234), .SEL(n1872), .F(n1777) );
  IV U655 ( .A(n1873), .Z(n234) );
  MUX U656 ( .IN0(n235), .IN1(n2346), .SEL(n2347), .F(n2230) );
  IV U657 ( .A(n2348), .Z(n235) );
  MUX U658 ( .IN0(n236), .IN1(n2826), .SEL(n2827), .F(n2700) );
  IV U659 ( .A(n2828), .Z(n236) );
  MUX U660 ( .IN0(n237), .IN1(n2846), .SEL(n2847), .F(n2717) );
  IV U661 ( .A(n2848), .Z(n237) );
  AND U662 ( .A(n771), .B(n772), .Z(n742) );
  AND U663 ( .A(n966), .B(n967), .Z(n922) );
  XNOR U664 ( .A(n999), .B(n998), .Z(n991) );
  AND U665 ( .A(n1205), .B(n1206), .Z(n1142) );
  ANDN U666 ( .A(n1497), .B(n1498), .Z(n1418) );
  MUX U667 ( .IN0(n1993), .IN1(n238), .SEL(n1994), .F(n1888) );
  IV U668 ( .A(n1995), .Z(n238) );
  MUX U669 ( .IN0(n2212), .IN1(n2324), .SEL(n2214), .F(n2101) );
  ANDN U670 ( .A(n2282), .B(n2283), .Z(n2171) );
  MUX U671 ( .IN0(n2557), .IN1(n239), .SEL(n2558), .F(n2436) );
  IV U672 ( .A(n2559), .Z(n239) );
  ANDN U673 ( .A(n713), .B(n712), .Z(n708) );
  XNOR U674 ( .A(n815), .B(n812), .Z(n811) );
  OR U675 ( .A(n1032), .B(n1033), .Z(n974) );
  OR U676 ( .A(n1282), .B(n1283), .Z(n1213) );
  XNOR U677 ( .A(n1512), .B(n1511), .Z(n1590) );
  OR U678 ( .A(n728), .B(n729), .Z(n701) );
  MUX U679 ( .IN0(n240), .IN1(n744), .SEL(n745), .F(n691) );
  IV U680 ( .A(o_reg[29]), .Z(n240) );
  MUX U681 ( .IN0(n241), .IN1(n882), .SEL(n883), .F(n845) );
  IV U682 ( .A(o_reg[25]), .Z(n241) );
  MUX U683 ( .IN0(n242), .IN1(n1144), .SEL(n1145), .F(n1084) );
  IV U684 ( .A(o_reg[20]), .Z(n242) );
  MUX U685 ( .IN0(n1420), .IN1(n243), .SEL(n1421), .F(n1346) );
  IV U686 ( .A(o_reg[16]), .Z(n243) );
  MUX U687 ( .IN0(n1769), .IN1(n244), .SEL(n1770), .F(n1676) );
  IV U688 ( .A(o_reg[12]), .Z(n244) );
  MUX U689 ( .IN0(n2173), .IN1(n245), .SEL(n681), .F(n2066) );
  IV U690 ( .A(o_reg[8]), .Z(n245) );
  MUX U691 ( .IN0(n246), .IN1(n2643), .SEL(n685), .F(n2521) );
  IV U692 ( .A(o_reg[4]), .Z(n246) );
  MUX U693 ( .IN0(n247), .IN1(n3760), .SEL(n3761), .F(n3722) );
  IV U694 ( .A(n3762), .Z(n247) );
  MUX U695 ( .IN0(n248), .IN1(n3730), .SEL(n3731), .F(n3692) );
  IV U696 ( .A(n3732), .Z(n248) );
  MUX U697 ( .IN0(n249), .IN1(n4137), .SEL(n4138), .F(n4120) );
  IV U698 ( .A(n4139), .Z(n249) );
  MUX U699 ( .IN0(n250), .IN1(n4129), .SEL(n4130), .F(n4112) );
  IV U700 ( .A(n4131), .Z(n250) );
  MUX U701 ( .IN0(n251), .IN1(n3735), .SEL(n3736), .F(n3697) );
  IV U702 ( .A(n3737), .Z(n251) );
  MUX U703 ( .IN0(n252), .IN1(n3743), .SEL(n3744), .F(n3705) );
  IV U704 ( .A(n3745), .Z(n252) );
  MUX U705 ( .IN0(n253), .IN1(n4547), .SEL(n4548), .F(n4534) );
  IV U706 ( .A(n4549), .Z(n253) );
  MUX U707 ( .IN0(n254), .IN1(n4514), .SEL(n4515), .F(n4501) );
  IV U708 ( .A(n4516), .Z(n254) );
  MUX U709 ( .IN0(n255), .IN1(n4140), .SEL(n3756), .F(n4123) );
  IV U710 ( .A(n3754), .Z(n255) );
  MUX U711 ( .IN0(n256), .IN1(n3788), .SEL(n3203), .F(n3750) );
  IV U712 ( .A(n3202), .Z(n256) );
  XNOR U713 ( .A(n3682), .B(n3647), .Z(n3651) );
  XOR U714 ( .A(n4517), .B(n4509), .Z(n4109) );
  MUX U715 ( .IN0(n4101), .IN1(n4099), .SEL(n4100), .F(n4082) );
  MUX U716 ( .IN0(n3671), .IN1(n3673), .SEL(n3672), .F(n3633) );
  MUX U717 ( .IN0(n257), .IN1(n3578), .SEL(n3579), .F(n3540) );
  IV U718 ( .A(n3580), .Z(n257) );
  MUX U719 ( .IN0(n258), .IN1(n4069), .SEL(n4070), .F(n4052) );
  IV U720 ( .A(n4071), .Z(n258) );
  MUX U721 ( .IN0(n259), .IN1(n4061), .SEL(n4062), .F(n4044) );
  IV U722 ( .A(n4063), .Z(n259) );
  MUX U723 ( .IN0(n260), .IN1(n3583), .SEL(n3584), .F(n3545) );
  IV U724 ( .A(n3585), .Z(n260) );
  MUX U725 ( .IN0(n3624), .IN1(n261), .SEL(n3625), .F(n3586) );
  IV U726 ( .A(n3626), .Z(n261) );
  XNOR U727 ( .A(n3568), .B(n3533), .Z(n3537) );
  MUX U728 ( .IN0(n262), .IN1(n4072), .SEL(n3604), .F(n4055) );
  IV U729 ( .A(n3602), .Z(n262) );
  MUX U730 ( .IN0(n263), .IN1(n3515), .SEL(n3516), .F(n3477) );
  IV U731 ( .A(n3517), .Z(n263) );
  MUX U732 ( .IN0(n264), .IN1(n4632), .SEL(n4633), .F(n4621) );
  IV U733 ( .A(n4634), .Z(n264) );
  MUX U734 ( .IN0(n265), .IN1(n4449), .SEL(n4450), .F(n4436) );
  IV U735 ( .A(n4451), .Z(n265) );
  MUX U736 ( .IN0(n266), .IN1(n3456), .SEL(n3457), .F(n3418) );
  IV U737 ( .A(n3458), .Z(n266) );
  MUX U738 ( .IN0(n267), .IN1(n4469), .SEL(n4470), .F(n4456) );
  IV U739 ( .A(n4471), .Z(n267) );
  MUX U740 ( .IN0(n4033), .IN1(n4031), .SEL(n4032), .F(n4014) );
  MUX U741 ( .IN0(n268), .IN1(n4989), .SEL(n4990), .F(n4976) );
  IV U742 ( .A(n4991), .Z(n268) );
  XOR U743 ( .A(n4856), .B(n4857), .Z(n4866) );
  MUX U744 ( .IN0(n269), .IN1(n4001), .SEL(n4002), .F(n3984) );
  IV U745 ( .A(n4003), .Z(n269) );
  MUX U746 ( .IN0(n270), .IN1(n3993), .SEL(n3994), .F(n3976) );
  IV U747 ( .A(n3995), .Z(n270) );
  XOR U748 ( .A(n4314), .B(n4296), .Z(n4300) );
  XOR U749 ( .A(n4270), .B(n4271), .Z(n4280) );
  MUX U750 ( .IN0(n4447), .IN1(n271), .SEL(n4024), .F(n4434) );
  IV U751 ( .A(n4023), .Z(n271) );
  XOR U752 ( .A(n4835), .B(n4836), .Z(n4845) );
  MUX U753 ( .IN0(n272), .IN1(n4839), .SEL(n4840), .F(n4818) );
  IV U754 ( .A(n4841), .Z(n272) );
  MUX U755 ( .IN0(n3424), .IN1(n3422), .SEL(n3423), .F(n3384) );
  MUX U756 ( .IN0(n3472), .IN1(n273), .SEL(n3473), .F(n3434) );
  IV U757 ( .A(n3474), .Z(n273) );
  XOR U758 ( .A(n4613), .B(n4605), .Z(n4266) );
  XOR U759 ( .A(n4249), .B(n4250), .Z(n4259) );
  MUX U760 ( .IN0(n274), .IN1(n4253), .SEL(n4254), .F(n4232) );
  IV U761 ( .A(n4255), .Z(n274) );
  XOR U762 ( .A(n4979), .B(n4971), .Z(n4831) );
  XOR U763 ( .A(n4814), .B(n4815), .Z(n4824) );
  MUX U764 ( .IN0(n275), .IN1(n4004), .SEL(n3452), .F(n3987) );
  IV U765 ( .A(n3450), .Z(n275) );
  MUX U766 ( .IN0(n3405), .IN1(n3407), .SEL(n3406), .F(n3367) );
  MUX U767 ( .IN0(n276), .IN1(n3363), .SEL(n3364), .F(n3325) );
  IV U768 ( .A(n3365), .Z(n276) );
  MUX U769 ( .IN0(n277), .IN1(n4347), .SEL(n4348), .F(n4686) );
  IV U770 ( .A(n4700), .Z(n277) );
  MUX U771 ( .IN0(n4676), .IN1(n4691), .SEL(n4678), .F(n4660) );
  MUX U772 ( .IN0(n278), .IN1(n4588), .SEL(n4589), .F(n4577) );
  IV U773 ( .A(n4590), .Z(n278) );
  MUX U774 ( .IN0(n279), .IN1(n4397), .SEL(n4398), .F(n4384) );
  IV U775 ( .A(n4399), .Z(n279) );
  MUX U776 ( .IN0(n280), .IN1(n4912), .SEL(n4913), .F(n5058) );
  IV U777 ( .A(n5072), .Z(n280) );
  MUX U778 ( .IN0(n5048), .IN1(n5063), .SEL(n5050), .F(n5032) );
  MUX U779 ( .IN0(n281), .IN1(n3304), .SEL(n3305), .F(n3266) );
  IV U780 ( .A(n3306), .Z(n281) );
  MUX U781 ( .IN0(n3965), .IN1(n3963), .SEL(n3964), .F(n3946) );
  MUX U782 ( .IN0(n282), .IN1(n3798), .SEL(n3799), .F(n3839) );
  IV U783 ( .A(n3853), .Z(n282) );
  MUX U784 ( .IN0(n3829), .IN1(n3844), .SEL(n3831), .F(n3813) );
  MUX U785 ( .IN0(n283), .IN1(n5099), .SEL(n5100), .F(n5146) );
  IV U786 ( .A(n5162), .Z(n283) );
  MUX U787 ( .IN0(n284), .IN1(n4404), .SEL(n4405), .F(n4391) );
  IV U788 ( .A(n4406), .Z(n284) );
  MUX U789 ( .IN0(n285), .IN1(n3925), .SEL(n3926), .F(n3905) );
  IV U790 ( .A(n3927), .Z(n285) );
  MUX U791 ( .IN0(n286), .IN1(n3279), .SEL(n3280), .F(n3241) );
  IV U792 ( .A(n3281), .Z(n286) );
  MUX U793 ( .IN0(n4395), .IN1(n287), .SEL(n3956), .F(n4382) );
  IV U794 ( .A(n3955), .Z(n287) );
  MUX U795 ( .IN0(n288), .IN1(n5191), .SEL(n5192), .F(n5187) );
  IV U796 ( .A(n5193), .Z(n288) );
  MUX U797 ( .IN0(n289), .IN1(n3236), .SEL(n3237), .F(n3199) );
  IV U798 ( .A(n3238), .Z(n289) );
  MUX U799 ( .IN0(n290), .IN1(n3913), .SEL(n3914), .F(n3215) );
  IV U800 ( .A(n3915), .Z(n290) );
  MUX U801 ( .IN0(n3320), .IN1(n291), .SEL(n3321), .F(n3282) );
  IV U802 ( .A(n3322), .Z(n291) );
  MUX U803 ( .IN0(n4575), .IN1(n292), .SEL(n4203), .F(n4564) );
  IV U804 ( .A(n4201), .Z(n292) );
  XOR U805 ( .A(n4209), .B(n4191), .Z(n4195) );
  XOR U806 ( .A(n4174), .B(n4175), .Z(n4171) );
  MUX U807 ( .IN0(n5095), .IN1(n5123), .SEL(n5097), .F(n3141) );
  MUX U808 ( .IN0(n4935), .IN1(n293), .SEL(n4768), .F(n4922) );
  IV U809 ( .A(n4766), .Z(n293) );
  MUX U810 ( .IN0(n4759), .IN1(n294), .SEL(n4760), .F(n4727) );
  IV U811 ( .A(n4761), .Z(n294) );
  MUX U812 ( .IN0(n295), .IN1(n4723), .SEL(n4724), .F(n3108) );
  IV U813 ( .A(n4725), .Z(n295) );
  MUX U814 ( .IN0(n296), .IN1(n3936), .SEL(n3300), .F(n3919) );
  IV U815 ( .A(n3298), .Z(n296) );
  XOR U816 ( .A(n3285), .B(n3250), .Z(n3254) );
  XNOR U817 ( .A(n3226), .B(n3192), .Z(n3196) );
  MUX U818 ( .IN0(n297), .IN1(n1021), .SEL(n1022), .F(n963) );
  IV U819 ( .A(n1023), .Z(n297) );
  MUX U820 ( .IN0(n298), .IN1(n1070), .SEL(n1071), .F(n1012) );
  IV U821 ( .A(n1072), .Z(n298) );
  MUX U822 ( .IN0(n299), .IN1(n1061), .SEL(n1062), .F(n1003) );
  IV U823 ( .A(n1063), .Z(n299) );
  MUX U824 ( .IN0(n300), .IN1(n1322), .SEL(n1323), .F(n1252) );
  IV U825 ( .A(n1324), .Z(n300) );
  MUX U826 ( .IN0(n301), .IN1(n1405), .SEL(n1406), .F(n1331) );
  IV U827 ( .A(n1407), .Z(n301) );
  MUX U828 ( .IN0(n302), .IN1(n1518), .SEL(n1519), .F(n1432) );
  IV U829 ( .A(n1520), .Z(n302) );
  MUX U830 ( .IN0(n303), .IN1(n1726), .SEL(n1727), .F(n1635) );
  IV U831 ( .A(n1728), .Z(n303) );
  MUX U832 ( .IN0(n304), .IN1(n1832), .SEL(n1833), .F(n1735) );
  IV U833 ( .A(n1834), .Z(n304) );
  MUX U834 ( .IN0(n305), .IN1(n1840), .SEL(n1841), .F(n1743) );
  IV U835 ( .A(n1842), .Z(n305) );
  MUX U836 ( .IN0(n306), .IN1(n2009), .SEL(n2010), .F(n1904) );
  IV U837 ( .A(n2011), .Z(n306) );
  MUX U838 ( .IN0(n307), .IN1(n2130), .SEL(n2131), .F(n2025) );
  IV U839 ( .A(n2132), .Z(n307) );
  MUX U840 ( .IN0(n308), .IN1(n2252), .SEL(n2253), .F(n2139) );
  IV U841 ( .A(n2254), .Z(n308) );
  MUX U842 ( .IN0(n309), .IN1(n2260), .SEL(n2261), .F(n2147) );
  IV U843 ( .A(n2262), .Z(n309) );
  MUX U844 ( .IN0(n310), .IN1(n2425), .SEL(n2426), .F(n2310) );
  IV U845 ( .A(n2427), .Z(n310) );
  MUX U846 ( .IN0(n311), .IN1(n2602), .SEL(n2603), .F(n2480) );
  IV U847 ( .A(n2604), .Z(n311) );
  MUX U848 ( .IN0(n312), .IN1(n2653), .SEL(n2654), .F(n2529) );
  IV U849 ( .A(n2655), .Z(n312) );
  MUX U850 ( .IN0(n313), .IN1(n2678), .SEL(n2679), .F(n2554) );
  IV U851 ( .A(n2680), .Z(n313) );
  MUX U852 ( .IN0(n314), .IN1(n2739), .SEL(n2740), .F(n2611) );
  IV U853 ( .A(n2741), .Z(n314) );
  MUX U854 ( .IN0(n315), .IN1(n2747), .SEL(n2748), .F(n2619) );
  IV U855 ( .A(n2749), .Z(n315) );
  MUX U856 ( .IN0(n316), .IN1(n2714), .SEL(n2715), .F(n2586) );
  IV U857 ( .A(n2716), .Z(n316) );
  MUX U858 ( .IN0(n317), .IN1(n2788), .SEL(n2789), .F(n2661) );
  IV U859 ( .A(n2790), .Z(n317) );
  MUX U860 ( .IN0(n318), .IN1(n2823), .SEL(n2824), .F(n2695) );
  IV U861 ( .A(n2825), .Z(n318) );
  MUX U862 ( .IN0(n319), .IN1(n3132), .SEL(n3133), .F(n2997) );
  IV U863 ( .A(n3134), .Z(n319) );
  MUX U864 ( .IN0(n916), .IN1(n914), .SEL(n915), .F(n872) );
  MUX U865 ( .IN0(n320), .IN1(n1165), .SEL(n1166), .F(n1103) );
  IV U866 ( .A(n1167), .Z(n320) );
  MUX U867 ( .IN0(n1199), .IN1(n1197), .SEL(n1198), .F(n1134) );
  MUX U868 ( .IN0(n1188), .IN1(n1190), .SEL(n1189), .F(n1125) );
  MUX U869 ( .IN0(n1293), .IN1(n1291), .SEL(n1292), .F(n1223) );
  MUX U870 ( .IN0(n1379), .IN1(n321), .SEL(n1378), .F(n1308) );
  IV U871 ( .A(n1377), .Z(n321) );
  MUX U872 ( .IN0(n322), .IN1(n1885), .SEL(n1886), .F(n1788) );
  IV U873 ( .A(n1887), .Z(n322) );
  MUX U874 ( .IN0(n1617), .IN1(n1615), .SEL(n1616), .F(n1522) );
  MUX U875 ( .IN0(n1924), .IN1(n1926), .SEL(n1925), .F(n1827) );
  MUX U876 ( .IN0(n2046), .IN1(n2048), .SEL(n2047), .F(n1941) );
  MUX U877 ( .IN0(n2307), .IN1(n323), .SEL(n2306), .F(n2192) );
  IV U878 ( .A(n2305), .Z(n323) );
  MUX U879 ( .IN0(n2363), .IN1(n2365), .SEL(n2364), .F(n2247) );
  MUX U880 ( .IN0(n2501), .IN1(n2503), .SEL(n2502), .F(n2380) );
  MUX U881 ( .IN0(n2863), .IN1(n2865), .SEL(n2864), .F(n2734) );
  MUX U882 ( .IN0(n3018), .IN1(n3020), .SEL(n3019), .F(n2880) );
  MUX U883 ( .IN0(n2921), .IN1(n2923), .SEL(n2922), .F(n2792) );
  XNOR U884 ( .A(n3205), .B(n3080), .Z(n3084) );
  MUX U885 ( .IN0(n863), .IN1(n865), .SEL(n864), .F(n324) );
  IV U886 ( .A(n324), .Z(n818) );
  MUX U887 ( .IN0(n325), .IN1(n940), .SEL(n941), .F(n898) );
  IV U888 ( .A(n942), .Z(n325) );
  MUX U889 ( .IN0(n326), .IN1(n1247), .SEL(n1248), .F(n1179) );
  IV U890 ( .A(n1249), .Z(n326) );
  XNOR U891 ( .A(n1383), .B(n1454), .Z(n1384) );
  XOR U892 ( .A(n1558), .B(n1476), .Z(n1480) );
  XNOR U893 ( .A(n1659), .B(n1570), .Z(n1574) );
  MUX U894 ( .IN0(n1721), .IN1(n327), .SEL(n1722), .F(n1630) );
  IV U895 ( .A(n1723), .Z(n327) );
  MUX U896 ( .IN0(n328), .IN1(n1835), .SEL(n1836), .F(n1738) );
  IV U897 ( .A(n1837), .Z(n328) );
  NAND U898 ( .A(n1783), .B(n1879), .Z(n1878) );
  XNOR U899 ( .A(n2049), .B(n1947), .Z(n1951) );
  XNOR U900 ( .A(n1999), .B(n1897), .Z(n1901) );
  MUX U901 ( .IN0(n2125), .IN1(n329), .SEL(n2126), .F(n2020) );
  IV U902 ( .A(n2127), .Z(n329) );
  XNOR U903 ( .A(n2196), .B(n2088), .Z(n2092) );
  MUX U904 ( .IN0(n330), .IN1(n2255), .SEL(n2256), .F(n2142) );
  IV U905 ( .A(n2257), .Z(n330) );
  XNOR U906 ( .A(n2333), .B(n2220), .Z(n2224) );
  MUX U907 ( .IN0(n331), .IN1(n2411), .SEL(n2412), .F(n2295) );
  IV U908 ( .A(n2413), .Z(n331) );
  XNOR U909 ( .A(n2504), .B(n2386), .Z(n2390) );
  MUX U910 ( .IN0(n2597), .IN1(n332), .SEL(n2598), .F(n2475) );
  IV U911 ( .A(n2599), .Z(n332) );
  XNOR U912 ( .A(n2795), .B(n2671), .Z(n2675) );
  NAND U913 ( .A(n2690), .B(n2817), .Z(n2816) );
  XNOR U914 ( .A(n2833), .B(n2707), .Z(n2711) );
  XNOR U915 ( .A(n2883), .B(n2757), .Z(n2761) );
  MUX U916 ( .IN0(n3127), .IN1(n333), .SEL(n3128), .F(n2992) );
  IV U917 ( .A(n3129), .Z(n333) );
  MUX U918 ( .IN0(n334), .IN1(n3048), .SEL(n3049), .F(n2912) );
  IV U919 ( .A(n3050), .Z(n334) );
  MUX U920 ( .IN0(n3104), .IN1(n429), .SEL(n3103), .F(n2966) );
  XNOR U921 ( .A(n3164), .B(n3163), .Z(n3146) );
  MUX U922 ( .IN0(n335), .IN1(n1298), .SEL(n1299), .F(n1230) );
  IV U923 ( .A(n1300), .Z(n335) );
  MUX U924 ( .IN0(n336), .IN1(n1622), .SEL(n1623), .F(n1529) );
  IV U925 ( .A(n1624), .Z(n336) );
  MUX U926 ( .IN0(n337), .IN1(n2012), .SEL(n2013), .F(n1907) );
  IV U927 ( .A(n2014), .Z(n337) );
  MUX U928 ( .IN0(n338), .IN1(n2467), .SEL(n2468), .F(n2346) );
  IV U929 ( .A(n2469), .Z(n338) );
  MUX U930 ( .IN0(n2831), .IN1(n2829), .SEL(n2830), .F(n339) );
  IV U931 ( .A(n339), .Z(n2699) );
  MUX U932 ( .IN0(n340), .IN1(n2984), .SEL(n2985), .F(n2846) );
  IV U933 ( .A(n2986), .Z(n340) );
  OR U934 ( .A(n763), .B(n764), .Z(n758) );
  MUX U935 ( .IN0(n341), .IN1(n768), .SEL(n769), .F(n739) );
  IV U936 ( .A(n770), .Z(n341) );
  XOR U937 ( .A(n1049), .B(n1044), .Z(n1092) );
  ANDN U938 ( .A(n1418), .B(n1419), .Z(n1344) );
  ANDN U939 ( .A(n1767), .B(n1768), .Z(n1674) );
  XOR U940 ( .A(n2324), .B(n2212), .Z(n2213) );
  ANDN U941 ( .A(n2398), .B(n2399), .Z(n2282) );
  MUX U942 ( .IN0(n2681), .IN1(n342), .SEL(n2682), .F(n2557) );
  IV U943 ( .A(n2683), .Z(n342) );
  AND U944 ( .A(n742), .B(n743), .Z(n699) );
  XNOR U945 ( .A(n711), .B(n710), .Z(n702) );
  XNOR U946 ( .A(n753), .B(n752), .Z(n751) );
  XNOR U947 ( .A(n854), .B(n853), .Z(n852) );
  XNOR U948 ( .A(n1108), .B(n1107), .Z(n1091) );
  OR U949 ( .A(n1352), .B(n1353), .Z(n1282) );
  XOR U950 ( .A(n1591), .B(n1605), .Z(n1682) );
  XOR U951 ( .A(n1891), .B(n1888), .Z(n1966) );
  MUX U952 ( .IN0(n343), .IN1(n924), .SEL(n925), .F(n882) );
  IV U953 ( .A(o_reg[24]), .Z(n343) );
  XNOR U954 ( .A(n931), .B(n930), .Z(n971) );
  MUX U955 ( .IN0(n344), .IN1(n1207), .SEL(n1208), .F(n1144) );
  IV U956 ( .A(o_reg[19]), .Z(n344) );
  MUX U957 ( .IN0(n1499), .IN1(n345), .SEL(n1500), .F(n1420) );
  IV U958 ( .A(o_reg[15]), .Z(n345) );
  MUX U959 ( .IN0(n1864), .IN1(n346), .SEL(n1865), .F(n1769) );
  IV U960 ( .A(o_reg[11]), .Z(n346) );
  MUX U961 ( .IN0(n2284), .IN1(n347), .SEL(n682), .F(n2173) );
  IV U962 ( .A(o_reg[7]), .Z(n347) );
  MUX U963 ( .IN0(n348), .IN1(n2769), .SEL(n723), .F(n2643) );
  IV U964 ( .A(o_reg[3]), .Z(n348) );
  MUX U965 ( .IN0(o_reg[31]), .IN1(n349), .SEL(n690), .F(n686) );
  IV U966 ( .A(n689), .Z(n349) );
  MUX U967 ( .IN0(n350), .IN1(n4156), .SEL(n4157), .F(n4137) );
  IV U968 ( .A(n4158), .Z(n350) );
  MUX U969 ( .IN0(n3728), .IN1(n3726), .SEL(n3727), .F(n3688) );
  MUX U970 ( .IN0(n351), .IN1(n4159), .SEL(n3791), .F(n4140) );
  IV U971 ( .A(n3790), .Z(n351) );
  MUX U972 ( .IN0(n3747), .IN1(n3749), .SEL(n3748), .F(n3709) );
  MUX U973 ( .IN0(n352), .IN1(n3654), .SEL(n3655), .F(n3616) );
  IV U974 ( .A(n3656), .Z(n352) );
  MUX U975 ( .IN0(n353), .IN1(n3646), .SEL(n3647), .F(n3608) );
  IV U976 ( .A(n3648), .Z(n353) );
  MUX U977 ( .IN0(n4118), .IN1(n4116), .SEL(n4117), .F(n4099) );
  MUX U978 ( .IN0(n354), .IN1(n4521), .SEL(n4522), .F(n4508) );
  IV U979 ( .A(n4523), .Z(n354) );
  MUX U980 ( .IN0(n355), .IN1(n4086), .SEL(n4087), .F(n4069) );
  IV U981 ( .A(n4088), .Z(n355) );
  MUX U982 ( .IN0(n356), .IN1(n4078), .SEL(n4079), .F(n4061) );
  IV U983 ( .A(n4080), .Z(n356) );
  MUX U984 ( .IN0(n4512), .IN1(n357), .SEL(n4109), .F(n4499) );
  IV U985 ( .A(n4108), .Z(n357) );
  MUX U986 ( .IN0(n3662), .IN1(n358), .SEL(n3663), .F(n3624) );
  IV U987 ( .A(n3664), .Z(n358) );
  MUX U988 ( .IN0(n359), .IN1(n4475), .SEL(n4476), .F(n4462) );
  IV U989 ( .A(n4477), .Z(n359) );
  MUX U990 ( .IN0(n3576), .IN1(n3574), .SEL(n3575), .F(n3536) );
  MUX U991 ( .IN0(n360), .IN1(n4089), .SEL(n3642), .F(n4072) );
  IV U992 ( .A(n3640), .Z(n360) );
  XOR U993 ( .A(n3627), .B(n3592), .Z(n3596) );
  MUX U994 ( .IN0(n361), .IN1(n3545), .SEL(n3546), .F(n3507) );
  IV U995 ( .A(n3547), .Z(n361) );
  MUX U996 ( .IN0(n362), .IN1(n3502), .SEL(n3503), .F(n3464) );
  IV U997 ( .A(n3504), .Z(n362) );
  MUX U998 ( .IN0(n363), .IN1(n3494), .SEL(n3495), .F(n3456) );
  IV U999 ( .A(n3496), .Z(n363) );
  MUX U1000 ( .IN0(n4050), .IN1(n4048), .SEL(n4049), .F(n4031) );
  MUX U1001 ( .IN0(n364), .IN1(n4311), .SEL(n4312), .F(n4290) );
  IV U1002 ( .A(n4313), .Z(n364) );
  MUX U1003 ( .IN0(n365), .IN1(n4637), .SEL(n4638), .F(n4626) );
  IV U1004 ( .A(n4639), .Z(n365) );
  MUX U1005 ( .IN0(n366), .IN1(n4018), .SEL(n4019), .F(n4001) );
  IV U1006 ( .A(n4020), .Z(n366) );
  MUX U1007 ( .IN0(n367), .IN1(n4010), .SEL(n4011), .F(n3993) );
  IV U1008 ( .A(n4012), .Z(n367) );
  MUX U1009 ( .IN0(n4460), .IN1(n368), .SEL(n4041), .F(n4447) );
  IV U1010 ( .A(n4040), .Z(n368) );
  MUX U1011 ( .IN0(n369), .IN1(n4456), .SEL(n4457), .F(n4443) );
  IV U1012 ( .A(n4458), .Z(n369) );
  MUX U1013 ( .IN0(n3481), .IN1(n3483), .SEL(n3482), .F(n3443) );
  MUX U1014 ( .IN0(n370), .IN1(n3439), .SEL(n3440), .F(n3401) );
  IV U1015 ( .A(n3441), .Z(n370) );
  MUX U1016 ( .IN0(n3510), .IN1(n371), .SEL(n3511), .F(n3472) );
  IV U1017 ( .A(n3512), .Z(n371) );
  MUX U1018 ( .IN0(n372), .IN1(n4323), .SEL(n3896), .F(n4302) );
  IV U1019 ( .A(n3895), .Z(n372) );
  XOR U1020 ( .A(n4992), .B(n4984), .Z(n4852) );
  MUX U1021 ( .IN0(n373), .IN1(n4021), .SEL(n3490), .F(n4004) );
  IV U1022 ( .A(n3488), .Z(n373) );
  MUX U1023 ( .IN0(n374), .IN1(n3393), .SEL(n3394), .F(n3355) );
  IV U1024 ( .A(n3395), .Z(n374) );
  XNOR U1025 ( .A(n3416), .B(n3381), .Z(n3385) );
  MUX U1026 ( .IN0(n4619), .IN1(n375), .SEL(n4287), .F(n4608) );
  IV U1027 ( .A(n4285), .Z(n375) );
  MUX U1028 ( .IN0(n4843), .IN1(n376), .SEL(n4844), .F(n4822) );
  IV U1029 ( .A(n4845), .Z(n376) );
  MUX U1030 ( .IN0(n377), .IN1(n4818), .SEL(n4819), .F(n4797) );
  IV U1031 ( .A(n4820), .Z(n377) );
  MUX U1032 ( .IN0(n378), .IN1(n3350), .SEL(n3351), .F(n3312) );
  IV U1033 ( .A(n3352), .Z(n378) );
  MUX U1034 ( .IN0(n3982), .IN1(n3980), .SEL(n3981), .F(n3963) );
  MUX U1035 ( .IN0(n379), .IN1(n3850), .SEL(n3851), .F(n3835) );
  IV U1036 ( .A(n3852), .Z(n379) );
  MUX U1037 ( .IN0(n380), .IN1(n4227), .SEL(n4228), .F(n4206) );
  IV U1038 ( .A(n4229), .Z(n380) );
  MUX U1039 ( .IN0(n4682), .IN1(n4696), .SEL(n4684), .F(n4666) );
  MUX U1040 ( .IN0(n381), .IN1(n4712), .SEL(n4713), .F(n4708) );
  IV U1041 ( .A(n4714), .Z(n381) );
  MUX U1042 ( .IN0(n382), .IN1(n4593), .SEL(n4594), .F(n4582) );
  IV U1043 ( .A(n4595), .Z(n382) );
  XOR U1044 ( .A(n4272), .B(n4254), .Z(n4258) );
  MUX U1045 ( .IN0(n5054), .IN1(n5068), .SEL(n5056), .F(n5038) );
  MUX U1046 ( .IN0(n383), .IN1(n5084), .SEL(n5085), .F(n5080) );
  IV U1047 ( .A(n5086), .Z(n383) );
  XOR U1048 ( .A(n4964), .B(n4965), .Z(n4829) );
  MUX U1049 ( .IN0(n384), .IN1(n4957), .SEL(n4958), .F(n4944) );
  IV U1050 ( .A(n4959), .Z(n384) );
  MUX U1051 ( .IN0(n385), .IN1(n4792), .SEL(n4793), .F(n4771) );
  IV U1052 ( .A(n4794), .Z(n385) );
  MUX U1053 ( .IN0(n386), .IN1(n3942), .SEL(n3943), .F(n3925) );
  IV U1054 ( .A(n3944), .Z(n386) );
  MUX U1055 ( .IN0(n387), .IN1(n3866), .SEL(n3867), .F(n3862) );
  IV U1056 ( .A(n3868), .Z(n387) );
  MUX U1057 ( .IN0(n388), .IN1(n4333), .SEL(n4334), .F(n4329) );
  IV U1058 ( .A(n4335), .Z(n388) );
  XOR U1059 ( .A(n4589), .B(n4590), .Z(n4243) );
  MUX U1060 ( .IN0(n4408), .IN1(n389), .SEL(n3973), .F(n4395) );
  IV U1061 ( .A(n3972), .Z(n389) );
  MUX U1062 ( .IN0(n390), .IN1(n4384), .SEL(n4385), .F(n4371) );
  IV U1063 ( .A(n4386), .Z(n390) );
  MUX U1064 ( .IN0(n5142), .IN1(n5158), .SEL(n5144), .F(n5124) );
  MUX U1065 ( .IN0(n5136), .IN1(n5151), .SEL(n5138), .F(n5118) );
  MUX U1066 ( .IN0(n391), .IN1(n4898), .SEL(n4899), .F(n4894) );
  IV U1067 ( .A(n4900), .Z(n391) );
  XOR U1068 ( .A(n4951), .B(n4952), .Z(n4808) );
  MUX U1069 ( .IN0(n392), .IN1(n3933), .SEL(n3934), .F(n3913) );
  IV U1070 ( .A(n3935), .Z(n392) );
  MUX U1071 ( .IN0(n3358), .IN1(n393), .SEL(n3359), .F(n3320) );
  IV U1072 ( .A(n3360), .Z(n393) );
  MUX U1073 ( .IN0(n394), .IN1(n4566), .SEL(n4567), .F(n4555) );
  IV U1074 ( .A(n4568), .Z(n394) );
  XOR U1075 ( .A(n4938), .B(n4939), .Z(n4787) );
  MUX U1076 ( .IN0(n395), .IN1(n4391), .SEL(n4392), .F(n4378) );
  IV U1077 ( .A(n4393), .Z(n395) );
  MUX U1078 ( .IN0(n396), .IN1(n3953), .SEL(n3338), .F(n3936) );
  IV U1079 ( .A(n3336), .Z(n396) );
  XOR U1080 ( .A(n3323), .B(n3288), .Z(n3292) );
  XNOR U1081 ( .A(n3272), .B(n3271), .Z(n3284) );
  MUX U1082 ( .IN0(n3877), .IN1(n3880), .SEL(n3878), .F(n3760) );
  MUX U1083 ( .IN0(n397), .IN1(n4165), .SEL(n4166), .F(n4146) );
  IV U1084 ( .A(n4167), .Z(n397) );
  XOR U1085 ( .A(n4569), .B(n4561), .Z(n4182) );
  MUX U1086 ( .IN0(n4194), .IN1(n398), .SEL(n4195), .F(n4169) );
  IV U1087 ( .A(n4196), .Z(n398) );
  MUX U1088 ( .IN0(n5187), .IN1(n5190), .SEL(n5188), .F(n3158) );
  XOR U1089 ( .A(n4774), .B(n4756), .Z(n4760) );
  MUX U1090 ( .IN0(n399), .IN1(n3191), .SEL(n3192), .F(n3062) );
  IV U1091 ( .A(n3193), .Z(n399) );
  MUX U1092 ( .IN0(n400), .IN1(n3174), .SEL(n3175), .F(n3045) );
  IV U1093 ( .A(n3176), .Z(n400) );
  XNOR U1094 ( .A(n3234), .B(n3233), .Z(n3246) );
  MUX U1095 ( .IN0(n401), .IN1(n994), .SEL(n995), .F(n937) );
  IV U1096 ( .A(n996), .Z(n401) );
  MUX U1097 ( .IN0(n402), .IN1(n1079), .SEL(n1080), .F(n1021) );
  IV U1098 ( .A(n1081), .Z(n402) );
  MUX U1099 ( .IN0(n403), .IN1(n1193), .SEL(n1194), .F(n1130) );
  IV U1100 ( .A(n1195), .Z(n403) );
  MUX U1101 ( .IN0(n404), .IN1(n1367), .SEL(n1368), .F(n1295) );
  IV U1102 ( .A(n1369), .Z(n404) );
  MUX U1103 ( .IN0(n405), .IN1(n1448), .SEL(n1449), .F(n1377) );
  IV U1104 ( .A(n1450), .Z(n405) );
  MUX U1105 ( .IN0(n406), .IN1(n1432), .SEL(n1433), .F(n1357) );
  IV U1106 ( .A(n1434), .Z(n406) );
  MUX U1107 ( .IN0(n407), .IN1(n1467), .SEL(n1468), .F(n1388) );
  IV U1108 ( .A(n1469), .Z(n407) );
  MUX U1109 ( .IN0(n408), .IN1(n1652), .SEL(n1653), .F(n1560) );
  IV U1110 ( .A(n1654), .Z(n408) );
  MUX U1111 ( .IN0(n409), .IN1(n1710), .SEL(n1711), .F(n1619) );
  IV U1112 ( .A(n1712), .Z(n409) );
  MUX U1113 ( .IN0(n410), .IN1(n1815), .SEL(n1816), .F(n1718) );
  IV U1114 ( .A(n1817), .Z(n410) );
  MUX U1115 ( .IN0(n411), .IN1(n2042), .SEL(n2043), .F(n1937) );
  IV U1116 ( .A(n2044), .Z(n411) );
  MUX U1117 ( .IN0(n412), .IN1(n2025), .SEL(n2026), .F(n1920) );
  IV U1118 ( .A(n2027), .Z(n412) );
  MUX U1119 ( .IN0(n413), .IN1(n2114), .SEL(n2115), .F(n2009) );
  IV U1120 ( .A(n2116), .Z(n413) );
  MUX U1121 ( .IN0(n414), .IN1(n2206), .SEL(n2207), .F(n2095) );
  IV U1122 ( .A(n2208), .Z(n414) );
  MUX U1123 ( .IN0(n415), .IN1(n2198), .SEL(n2199), .F(n2087) );
  IV U1124 ( .A(n2200), .Z(n415) );
  MUX U1125 ( .IN0(n416), .IN1(n2292), .SEL(n2293), .F(n2181) );
  IV U1126 ( .A(n2294), .Z(n416) );
  MUX U1127 ( .IN0(n417), .IN1(n2497), .SEL(n2498), .F(n2376) );
  IV U1128 ( .A(n2499), .Z(n417) );
  MUX U1129 ( .IN0(n418), .IN1(n2480), .SEL(n2481), .F(n2359) );
  IV U1130 ( .A(n2482), .Z(n418) );
  MUX U1131 ( .IN0(n419), .IN1(n2537), .SEL(n2538), .F(n2416) );
  IV U1132 ( .A(n2539), .Z(n419) );
  MUX U1133 ( .IN0(n420), .IN1(n2586), .SEL(n2587), .F(n2464) );
  IV U1134 ( .A(n2588), .Z(n420) );
  MUX U1135 ( .IN0(n421), .IN1(n2706), .SEL(n2707), .F(n2578) );
  IV U1136 ( .A(n2708), .Z(n421) );
  MUX U1137 ( .IN0(n422), .IN1(n2805), .SEL(n2806), .F(n2678) );
  IV U1138 ( .A(n2807), .Z(n422) );
  MUX U1139 ( .IN0(n423), .IN1(n2997), .SEL(n2998), .F(n2859) );
  IV U1140 ( .A(n2999), .Z(n423) );
  MUX U1141 ( .IN0(n424), .IN1(n3014), .SEL(n3015), .F(n2876) );
  IV U1142 ( .A(n3016), .Z(n424) );
  MUX U1143 ( .IN0(n425), .IN1(n2951), .SEL(n2952), .F(n2823) );
  IV U1144 ( .A(n2953), .Z(n425) );
  MUX U1145 ( .IN0(n426), .IN1(n3116), .SEL(n3117), .F(n2981) );
  IV U1146 ( .A(n3118), .Z(n426) );
  XNOR U1147 ( .A(n3903), .B(n3208), .Z(n3212) );
  MUX U1148 ( .IN0(n427), .IN1(n868), .SEL(n869), .F(n831) );
  IV U1149 ( .A(n870), .Z(n427) );
  MUX U1150 ( .IN0(n946), .IN1(n428), .SEL(n945), .F(n906) );
  IV U1151 ( .A(n944), .Z(n428) );
  MUX U1152 ( .IN0(n1747), .IN1(n1749), .SEL(n1748), .F(n1656) );
  XOR U1153 ( .A(n1671), .B(n1762), .Z(n1672) );
  MUX U1154 ( .IN0(n2134), .IN1(n2136), .SEL(n2135), .F(n2029) );
  MUX U1155 ( .IN0(n2151), .IN1(n2153), .SEL(n2152), .F(n2046) );
  XOR U1156 ( .A(n2279), .B(n2393), .Z(n2280) );
  MUX U1157 ( .IN0(n2606), .IN1(n2608), .SEL(n2607), .F(n2484) );
  MUX U1158 ( .IN0(n2623), .IN1(n2625), .SEL(n2624), .F(n2501) );
  MUX U1159 ( .IN0(n2665), .IN1(n2667), .SEL(n2666), .F(n2541) );
  MUX U1160 ( .IN0(n3153), .IN1(n3155), .SEL(n3154), .F(n3018) );
  MUX U1161 ( .IN0(n3136), .IN1(n3138), .SEL(n3137), .F(n3001) );
  MUX U1162 ( .IN0(n3917), .IN1(n4355), .SEL(n3918), .F(n429) );
  MUX U1163 ( .IN0(n3099), .IN1(n430), .SEL(n3098), .F(n2961) );
  IV U1164 ( .A(n3097), .Z(n430) );
  XOR U1165 ( .A(n3180), .B(n3054), .Z(n3058) );
  AND U1166 ( .A(n824), .B(n823), .Z(n820) );
  MUX U1167 ( .IN0(n431), .IN1(n1103), .SEL(n1104), .F(n1041) );
  IV U1168 ( .A(n1105), .Z(n431) );
  MUX U1169 ( .IN0(n432), .IN1(n997), .SEL(n998), .F(n940) );
  IV U1170 ( .A(n999), .Z(n432) );
  XNOR U1171 ( .A(n1216), .B(n1156), .Z(n1162) );
  XOR U1172 ( .A(n1320), .B(n1253), .Z(n1257) );
  XNOR U1173 ( .A(n1403), .B(n1332), .Z(n1336) );
  MUX U1174 ( .IN0(n1786), .IN1(n433), .SEL(n1785), .F(n1685) );
  IV U1175 ( .A(n1784), .Z(n433) );
  NAND U1176 ( .A(n1459), .B(n1545), .Z(n1544) );
  MUX U1177 ( .IN0(n434), .IN1(n1555), .SEL(n1556), .F(n1470) );
  IV U1178 ( .A(n1557), .Z(n434) );
  XNOR U1179 ( .A(n1750), .B(n1662), .Z(n1666) );
  XNOR U1180 ( .A(n1700), .B(n1612), .Z(n1616) );
  MUX U1181 ( .IN0(n1915), .IN1(n435), .SEL(n1916), .F(n1818) );
  IV U1182 ( .A(n1917), .Z(n435) );
  MUX U1183 ( .IN0(n436), .IN1(n1932), .SEL(n1933), .F(n1835) );
  IV U1184 ( .A(n1934), .Z(n436) );
  MUX U1185 ( .IN0(n2084), .IN1(n2082), .SEL(n2083), .F(n437) );
  IV U1186 ( .A(n437), .Z(n1976) );
  XNOR U1187 ( .A(n2104), .B(n2002), .Z(n2006) );
  XNOR U1188 ( .A(n2154), .B(n2052), .Z(n2056) );
  MUX U1189 ( .IN0(n438), .IN1(n2371), .SEL(n2372), .F(n2255) );
  IV U1190 ( .A(n2373), .Z(n438) );
  XNOR U1191 ( .A(n2454), .B(n2336), .Z(n2340) );
  XNOR U1192 ( .A(n2544), .B(n2426), .Z(n2430) );
  MUX U1193 ( .IN0(n439), .IN1(n2532), .SEL(n2533), .F(n2411) );
  IV U1194 ( .A(n2534), .Z(n439) );
  XNOR U1195 ( .A(n2626), .B(n2507), .Z(n2511) );
  XOR U1196 ( .A(n2812), .B(n2691), .Z(n2692) );
  MUX U1197 ( .IN0(n2854), .IN1(n440), .SEL(n2855), .F(n2725) );
  IV U1198 ( .A(n2856), .Z(n440) );
  XNOR U1199 ( .A(n3021), .B(n2886), .Z(n2890) );
  XNOR U1200 ( .A(n2924), .B(n2798), .Z(n2802) );
  XNOR U1201 ( .A(n3106), .B(n2974), .Z(n2978) );
  MUX U1202 ( .IN0(n441), .IN1(n3100), .SEL(n3101), .F(n2967) );
  IV U1203 ( .A(n3102), .Z(n441) );
  XNOR U1204 ( .A(n3068), .B(n3067), .Z(n3050) );
  XNOR U1205 ( .A(n762), .B(n761), .Z(n757) );
  XNOR U1206 ( .A(n796), .B(n795), .Z(n787) );
  ANDN U1207 ( .A(n980), .B(n981), .Z(n979) );
  XNOR U1208 ( .A(n1235), .B(n1241), .Z(n1301) );
  MUX U1209 ( .IN0(n442), .IN1(n1713), .SEL(n1714), .F(n1622) );
  IV U1210 ( .A(n1715), .Z(n442) );
  XNOR U1211 ( .A(n1988), .B(n1987), .Z(n1979) );
  MUX U1212 ( .IN0(n443), .IN1(n2117), .SEL(n2118), .F(n2012) );
  IV U1213 ( .A(n2119), .Z(n443) );
  MUX U1214 ( .IN0(n444), .IN1(n2589), .SEL(n2590), .F(n2467) );
  IV U1215 ( .A(n2591), .Z(n444) );
  MUX U1216 ( .IN0(n445), .IN1(n2954), .SEL(n2955), .F(n2826) );
  IV U1217 ( .A(n2956), .Z(n445) );
  XNOR U1218 ( .A(n3029), .B(n3028), .Z(n3011) );
  MUX U1219 ( .IN0(n446), .IN1(n3119), .SEL(n3120), .F(n2984) );
  IV U1220 ( .A(n3121), .Z(n446) );
  AND U1221 ( .A(n802), .B(n803), .Z(n771) );
  XNOR U1222 ( .A(n862), .B(n861), .Z(n854) );
  XNOR U1223 ( .A(n900), .B(n899), .Z(n891) );
  AND U1224 ( .A(n1082), .B(n1083), .Z(n1024) );
  XNOR U1225 ( .A(n1058), .B(n1057), .Z(n1048) );
  XNOR U1226 ( .A(n1181), .B(n1180), .Z(n1170) );
  NOR U1227 ( .A(n1510), .B(n1511), .Z(n1509) );
  ANDN U1228 ( .A(n1674), .B(n1675), .Z(n1582) );
  ANDN U1229 ( .A(n2064), .B(n2065), .Z(n1959) );
  XNOR U1230 ( .A(n2450), .B(n2444), .Z(n2560) );
  ANDN U1231 ( .A(n2642), .B(n2641), .Z(n2519) );
  MUX U1232 ( .IN0(n2808), .IN1(n447), .SEL(n2809), .F(n2681) );
  IV U1233 ( .A(n2810), .Z(n447) );
  OR U1234 ( .A(n974), .B(n975), .Z(n930) );
  XOR U1235 ( .A(n1794), .B(n1791), .Z(n1870) );
  XOR U1236 ( .A(n2101), .B(n2098), .Z(n2178) );
  AND U1237 ( .A(n718), .B(n719), .Z(n714) );
  XNOR U1238 ( .A(n729), .B(n728), .Z(n747) );
  XNOR U1239 ( .A(n811), .B(n810), .Z(n848) );
  MUX U1240 ( .IN0(n448), .IN1(n1026), .SEL(n1027), .F(n968) );
  IV U1241 ( .A(o_reg[22]), .Z(n448) );
  XNOR U1242 ( .A(n1091), .B(n1090), .Z(n1148) );
  MUX U1243 ( .IN0(n1276), .IN1(n449), .SEL(n1277), .F(n1207) );
  IV U1244 ( .A(o_reg[18]), .Z(n449) );
  XOR U1245 ( .A(n1283), .B(n1282), .Z(n1349) );
  MUX U1246 ( .IN0(n1584), .IN1(n450), .SEL(n1585), .F(n1499) );
  IV U1247 ( .A(o_reg[14]), .Z(n450) );
  MUX U1248 ( .IN0(n1961), .IN1(n451), .SEL(n679), .F(n1864) );
  IV U1249 ( .A(o_reg[10]), .Z(n451) );
  MUX U1250 ( .IN0(n2400), .IN1(n452), .SEL(n683), .F(n2284) );
  IV U1251 ( .A(o_reg[6]), .Z(n452) );
  MUX U1252 ( .IN0(n453), .IN1(n2898), .SEL(n1146), .F(n2769) );
  IV U1253 ( .A(o_reg[2]), .Z(n453) );
  XOR U1254 ( .A(n691), .B(n726), .Z(n724) );
  XNOR U1255 ( .A(n3758), .B(n3723), .Z(n3727) );
  XOR U1256 ( .A(n3779), .B(n3744), .Z(n3748) );
  MUX U1257 ( .IN0(n454), .IN1(n4120), .SEL(n4121), .F(n4103) );
  IV U1258 ( .A(n4122), .Z(n454) );
  MUX U1259 ( .IN0(n455), .IN1(n3697), .SEL(n3698), .F(n3659) );
  IV U1260 ( .A(n3699), .Z(n455) );
  MUX U1261 ( .IN0(n456), .IN1(n4095), .SEL(n4096), .F(n4078) );
  IV U1262 ( .A(n4097), .Z(n456) );
  MUX U1263 ( .IN0(n457), .IN1(n4501), .SEL(n4502), .F(n4488) );
  IV U1264 ( .A(n4503), .Z(n457) );
  MUX U1265 ( .IN0(n458), .IN1(n3616), .SEL(n3617), .F(n3578) );
  IV U1266 ( .A(n3618), .Z(n458) );
  XNOR U1267 ( .A(n3644), .B(n3609), .Z(n3613) );
  MUX U1268 ( .IN0(n459), .IN1(n4508), .SEL(n4509), .F(n4495) );
  IV U1269 ( .A(n4510), .Z(n459) );
  MUX U1270 ( .IN0(n460), .IN1(n4106), .SEL(n3680), .F(n4089) );
  IV U1271 ( .A(n3678), .Z(n460) );
  MUX U1272 ( .IN0(n3633), .IN1(n3635), .SEL(n3634), .F(n3595) );
  MUX U1273 ( .IN0(n461), .IN1(n3591), .SEL(n3592), .F(n3553) );
  IV U1274 ( .A(n3593), .Z(n461) );
  MUX U1275 ( .IN0(n462), .IN1(n4052), .SEL(n4053), .F(n4035) );
  IV U1276 ( .A(n4054), .Z(n462) );
  MUX U1277 ( .IN0(n4067), .IN1(n4065), .SEL(n4066), .F(n4048) );
  MUX U1278 ( .IN0(n463), .IN1(n4027), .SEL(n4028), .F(n4010) );
  IV U1279 ( .A(n4029), .Z(n463) );
  MUX U1280 ( .IN0(n3586), .IN1(n464), .SEL(n3587), .F(n3548) );
  IV U1281 ( .A(n3588), .Z(n464) );
  XNOR U1282 ( .A(n3530), .B(n3495), .Z(n3499) );
  MUX U1283 ( .IN0(n4473), .IN1(n465), .SEL(n4058), .F(n4460) );
  IV U1284 ( .A(n4057), .Z(n465) );
  MUX U1285 ( .IN0(n466), .IN1(n3464), .SEL(n3465), .F(n3426) );
  IV U1286 ( .A(n3466), .Z(n466) );
  MUX U1287 ( .IN0(n467), .IN1(n4290), .SEL(n4291), .F(n4269) );
  IV U1288 ( .A(n4292), .Z(n467) );
  XOR U1289 ( .A(n4635), .B(n4627), .Z(n4308) );
  MUX U1290 ( .IN0(n468), .IN1(n4295), .SEL(n4296), .F(n4274) );
  IV U1291 ( .A(n4297), .Z(n468) );
  MUX U1292 ( .IN0(n469), .IN1(n4436), .SEL(n4437), .F(n4423) );
  IV U1293 ( .A(n4438), .Z(n469) );
  MUX U1294 ( .IN0(n470), .IN1(n4860), .SEL(n4861), .F(n4839) );
  IV U1295 ( .A(n4862), .Z(n470) );
  MUX U1296 ( .IN0(n471), .IN1(n4038), .SEL(n3528), .F(n4021) );
  IV U1297 ( .A(n3526), .Z(n471) );
  XOR U1298 ( .A(n3513), .B(n3478), .Z(n3482) );
  MUX U1299 ( .IN0(n472), .IN1(n3431), .SEL(n3432), .F(n3393) );
  IV U1300 ( .A(n3433), .Z(n472) );
  MUX U1301 ( .IN0(n473), .IN1(n4976), .SEL(n4977), .F(n4963) );
  IV U1302 ( .A(n4978), .Z(n473) );
  MUX U1303 ( .IN0(n474), .IN1(n4834), .SEL(n4835), .F(n4813) );
  IV U1304 ( .A(n4836), .Z(n474) );
  MUX U1305 ( .IN0(n475), .IN1(n4443), .SEL(n4444), .F(n4430) );
  IV U1306 ( .A(n4445), .Z(n475) );
  MUX U1307 ( .IN0(n3999), .IN1(n3997), .SEL(n3998), .F(n3980) );
  MUX U1308 ( .IN0(n3386), .IN1(n3384), .SEL(n3385), .F(n3346) );
  MUX U1309 ( .IN0(n476), .IN1(n3342), .SEL(n3343), .F(n3304) );
  IV U1310 ( .A(n3344), .Z(n476) );
  MUX U1311 ( .IN0(n477), .IN1(n3959), .SEL(n3960), .F(n3942) );
  IV U1312 ( .A(n3961), .Z(n477) );
  MUX U1313 ( .IN0(n3434), .IN1(n478), .SEL(n3435), .F(n3396) );
  IV U1314 ( .A(n3436), .Z(n478) );
  XOR U1315 ( .A(n4602), .B(n4594), .Z(n4245) );
  MUX U1316 ( .IN0(n4257), .IN1(n479), .SEL(n4258), .F(n4236) );
  IV U1317 ( .A(n4259), .Z(n479) );
  MUX U1318 ( .IN0(n4421), .IN1(n480), .SEL(n3990), .F(n4408) );
  IV U1319 ( .A(n3989), .Z(n480) );
  MUX U1320 ( .IN0(n4974), .IN1(n481), .SEL(n4831), .F(n4961) );
  IV U1321 ( .A(n4829), .Z(n481) );
  MUX U1322 ( .IN0(n482), .IN1(n3950), .SEL(n3951), .F(n3933) );
  IV U1323 ( .A(n3952), .Z(n482) );
  MUX U1324 ( .IN0(n3367), .IN1(n3369), .SEL(n3368), .F(n3329) );
  MUX U1325 ( .IN0(n483), .IN1(n3325), .SEL(n3326), .F(n3287) );
  IV U1326 ( .A(n3327), .Z(n483) );
  MUX U1327 ( .IN0(n3835), .IN1(n3849), .SEL(n3837), .F(n3819) );
  MUX U1328 ( .IN0(n484), .IN1(n4206), .SEL(n4207), .F(n4185) );
  IV U1329 ( .A(n4208), .Z(n484) );
  MUX U1330 ( .IN0(n4666), .IN1(n4681), .SEL(n4668), .F(n4643) );
  MUX U1331 ( .IN0(n4660), .IN1(n4675), .SEL(n4662), .F(n4649) );
  MUX U1332 ( .IN0(n485), .IN1(n4577), .SEL(n4578), .F(n4566) );
  IV U1333 ( .A(n4579), .Z(n485) );
  MUX U1334 ( .IN0(n486), .IN1(n4211), .SEL(n4212), .F(n4190) );
  IV U1335 ( .A(n4213), .Z(n486) );
  MUX U1336 ( .IN0(n5038), .IN1(n5053), .SEL(n5040), .F(n5015) );
  MUX U1337 ( .IN0(n5032), .IN1(n5047), .SEL(n5034), .F(n5021) );
  XOR U1338 ( .A(n4816), .B(n4798), .Z(n4802) );
  MUX U1339 ( .IN0(n487), .IN1(n4944), .SEL(n4945), .F(n4931) );
  IV U1340 ( .A(n4946), .Z(n487) );
  MUX U1341 ( .IN0(n488), .IN1(n3274), .SEL(n3275), .F(n3236) );
  IV U1342 ( .A(n3276), .Z(n488) );
  MUX U1343 ( .IN0(n489), .IN1(n3970), .SEL(n3376), .F(n3953) );
  IV U1344 ( .A(n3374), .Z(n489) );
  MUX U1345 ( .IN0(n3813), .IN1(n3828), .SEL(n3815), .F(n3802) );
  MUX U1346 ( .IN0(n490), .IN1(n3881), .SEL(n3882), .F(n3877) );
  IV U1347 ( .A(n3883), .Z(n490) );
  XNOR U1348 ( .A(n4713), .B(n4714), .Z(n4700) );
  MUX U1349 ( .IN0(n491), .IN1(n4571), .SEL(n4572), .F(n4560) );
  IV U1350 ( .A(n4573), .Z(n491) );
  NOR U1351 ( .A(\_MAC/_MULT/A__[0] ), .B(n5203), .Z(n5196) );
  XOR U1352 ( .A(n4372), .B(n4373), .Z(n3938) );
  MUX U1353 ( .IN0(n5124), .IN1(n5141), .SEL(n5126), .F(n5095) );
  XNOR U1354 ( .A(n5085), .B(n5086), .Z(n5072) );
  MUX U1355 ( .IN0(n492), .IN1(n4924), .SEL(n4925), .F(n4738) );
  IV U1356 ( .A(n4926), .Z(n492) );
  MUX U1357 ( .IN0(n493), .IN1(n4750), .SEL(n4751), .F(n4731) );
  IV U1358 ( .A(n4752), .Z(n493) );
  MUX U1359 ( .IN0(n494), .IN1(n3241), .SEL(n3242), .F(n3174) );
  IV U1360 ( .A(n3243), .Z(n494) );
  XNOR U1361 ( .A(n3264), .B(n3229), .Z(n3233) );
  XNOR U1362 ( .A(n3867), .B(n3868), .Z(n3853) );
  XNOR U1363 ( .A(n4334), .B(n4335), .Z(n4320) );
  XNOR U1364 ( .A(n5175), .B(n5176), .Z(n5162) );
  MUX U1365 ( .IN0(n5105), .IN1(n5115), .SEL(n5107), .F(n3149) );
  XNOR U1366 ( .A(n4899), .B(n4900), .Z(n4885) );
  MUX U1367 ( .IN0(n495), .IN1(n4378), .SEL(n4379), .F(n4362) );
  IV U1368 ( .A(n4380), .Z(n495) );
  XNOR U1369 ( .A(n3923), .B(n3906), .Z(n3910) );
  MUX U1370 ( .IN0(n3282), .IN1(n496), .SEL(n3283), .F(n3244) );
  IV U1371 ( .A(n3284), .Z(n496) );
  MUX U1372 ( .IN0(n4169), .IN1(n497), .SEL(n4170), .F(n4150) );
  IV U1373 ( .A(n4171), .Z(n497) );
  MUX U1374 ( .IN0(n4564), .IN1(n498), .SEL(n4182), .F(n4551) );
  IV U1375 ( .A(n4180), .Z(n498) );
  MUX U1376 ( .IN0(n499), .IN1(n937), .SEL(n938), .F(n895) );
  IV U1377 ( .A(n939), .Z(n499) );
  MUX U1378 ( .IN0(n500), .IN1(n1139), .SEL(n1140), .F(n1079) );
  IV U1379 ( .A(n1141), .Z(n500) );
  MUX U1380 ( .IN0(n501), .IN1(n1176), .SEL(n1177), .F(n1113) );
  IV U1381 ( .A(n1178), .Z(n501) );
  MUX U1382 ( .IN0(n502), .IN1(n1252), .SEL(n1253), .F(n1184) );
  IV U1383 ( .A(n1254), .Z(n502) );
  MUX U1384 ( .IN0(n503), .IN1(n1331), .SEL(n1332), .F(n1261) );
  IV U1385 ( .A(n1333), .Z(n503) );
  MUX U1386 ( .IN0(n504), .IN1(n1440), .SEL(n1441), .F(n1367) );
  IV U1387 ( .A(n1442), .Z(n504) );
  MUX U1388 ( .IN0(n505), .IN1(n1534), .SEL(n1535), .F(n1448) );
  IV U1389 ( .A(n1536), .Z(n505) );
  MUX U1390 ( .IN0(n506), .IN1(n1552), .SEL(n1553), .F(n1467) );
  IV U1391 ( .A(n1554), .Z(n506) );
  MUX U1392 ( .IN0(n507), .IN1(n1912), .SEL(n1913), .F(n1815) );
  IV U1393 ( .A(n1914), .Z(n507) );
  MUX U1394 ( .IN0(n508), .IN1(n1904), .SEL(n1905), .F(n1807) );
  IV U1395 ( .A(n1906), .Z(n508) );
  MUX U1396 ( .IN0(n509), .IN1(n1929), .SEL(n1930), .F(n1832) );
  IV U1397 ( .A(n1931), .Z(n509) );
  MUX U1398 ( .IN0(n510), .IN1(n2051), .SEL(n2052), .F(n1946) );
  IV U1399 ( .A(n2053), .Z(n510) );
  MUX U1400 ( .IN0(n511), .IN1(n2351), .SEL(n2352), .F(n2235) );
  IV U1401 ( .A(n2353), .Z(n511) );
  MUX U1402 ( .IN0(n512), .IN1(n2343), .SEL(n2344), .F(n2227) );
  IV U1403 ( .A(n2345), .Z(n512) );
  MUX U1404 ( .IN0(n513), .IN1(n2368), .SEL(n2369), .F(n2252) );
  IV U1405 ( .A(n2370), .Z(n513) );
  MUX U1406 ( .IN0(n514), .IN1(n2433), .SEL(n2434), .F(n2318) );
  IV U1407 ( .A(n2435), .Z(n514) );
  MUX U1408 ( .IN0(n515), .IN1(n2506), .SEL(n2507), .F(n2385) );
  IV U1409 ( .A(n2508), .Z(n515) );
  MUX U1410 ( .IN0(n516), .IN1(n2780), .SEL(n2781), .F(n2653) );
  IV U1411 ( .A(n2782), .Z(n516) );
  MUX U1412 ( .IN0(n517), .IN1(n2851), .SEL(n2852), .F(n2722) );
  IV U1413 ( .A(n2853), .Z(n517) );
  MUX U1414 ( .IN0(n518), .IN1(n2843), .SEL(n2844), .F(n2714) );
  IV U1415 ( .A(n2845), .Z(n518) );
  MUX U1416 ( .IN0(n519), .IN1(n2868), .SEL(n2869), .F(n2739) );
  IV U1417 ( .A(n2870), .Z(n519) );
  MUX U1418 ( .IN0(n520), .IN1(n3023), .SEL(n3024), .F(n2885) );
  IV U1419 ( .A(n3025), .Z(n520) );
  MUX U1420 ( .IN0(n521), .IN1(n2934), .SEL(n2935), .F(n2805) );
  IV U1421 ( .A(n2936), .Z(n521) );
  MUX U1422 ( .IN0(n522), .IN1(n3087), .SEL(n3088), .F(n2951) );
  IV U1423 ( .A(n3089), .Z(n522) );
  MUX U1424 ( .IN0(n523), .IN1(n3899), .SEL(n3900), .F(n3097) );
  IV U1425 ( .A(n3901), .Z(n523) );
  XNOR U1426 ( .A(n5192), .B(n5193), .Z(n3162) );
  XOR U1427 ( .A(n4753), .B(n4724), .Z(n4728) );
  XNOR U1428 ( .A(n3197), .B(n3196), .Z(n3179) );
  XOR U1429 ( .A(n3247), .B(n3183), .Z(n3187) );
  MUX U1430 ( .IN0(n1157), .IN1(n524), .SEL(n1156), .F(n1099) );
  IV U1431 ( .A(n1155), .Z(n524) );
  MUX U1432 ( .IN0(n1326), .IN1(n1328), .SEL(n1327), .F(n1256) );
  MUX U1433 ( .IN0(n1549), .IN1(n525), .SEL(n1548), .F(n1459) );
  IV U1434 ( .A(n1547), .Z(n525) );
  XOR U1435 ( .A(n1494), .B(n1577), .Z(n1495) );
  MUX U1436 ( .IN0(n526), .IN1(n2181), .SEL(n2182), .F(n2076) );
  IV U1437 ( .A(n2183), .Z(n526) );
  XOR U1438 ( .A(n4914), .B(n3133), .Z(n3137) );
  MUX U1439 ( .IN0(n3902), .IN1(n527), .SEL(n3224), .F(n3100) );
  IV U1440 ( .A(n3223), .Z(n527) );
  XNOR U1441 ( .A(n3766), .B(n3765), .Z(n3778) );
  XNOR U1442 ( .A(n866), .B(n832), .Z(n836) );
  XOR U1443 ( .A(n943), .B(n906), .Z(n904) );
  XNOR U1444 ( .A(n1010), .B(n955), .Z(n959) );
  XOR U1445 ( .A(n1119), .B(n1062), .Z(n1066) );
  XNOR U1446 ( .A(n1191), .B(n1131), .Z(n1135) );
  XNOR U1447 ( .A(n1355), .B(n1288), .Z(n1292) );
  MUX U1448 ( .IN0(n528), .IN1(n1788), .SEL(n1789), .F(n1691) );
  IV U1449 ( .A(n1790), .Z(n528) );
  XNOR U1450 ( .A(n1567), .B(n1485), .Z(n1489) );
  MUX U1451 ( .IN0(n1630), .IN1(n529), .SEL(n1631), .F(n1537) );
  IV U1452 ( .A(n1632), .Z(n529) );
  XNOR U1453 ( .A(n1609), .B(n1519), .Z(n1523) );
  XOR U1454 ( .A(n1650), .B(n1561), .Z(n1565) );
  XOR U1455 ( .A(n1821), .B(n1727), .Z(n1731) );
  XNOR U1456 ( .A(n1894), .B(n1800), .Z(n1804) );
  XOR U1457 ( .A(n1935), .B(n1841), .Z(n1845) );
  XNOR U1458 ( .A(n1980), .B(n1882), .Z(n1876) );
  XOR U1459 ( .A(n2128), .B(n2026), .Z(n2030) );
  XNOR U1460 ( .A(n2082), .B(n2187), .Z(n2083) );
  XOR U1461 ( .A(n2258), .B(n2148), .Z(n2152) );
  XNOR U1462 ( .A(n2217), .B(n2107), .Z(n2111) );
  MUX U1463 ( .IN0(n2238), .IN1(n530), .SEL(n2239), .F(n2125) );
  IV U1464 ( .A(n2240), .Z(n530) );
  XNOR U1465 ( .A(n2308), .B(n2199), .Z(n2203) );
  XOR U1466 ( .A(n2478), .B(n2360), .Z(n2364) );
  NAND U1467 ( .A(n2446), .B(n2565), .Z(n2564) );
  XOR U1468 ( .A(n2535), .B(n2417), .Z(n2421) );
  XNOR U1469 ( .A(n2576), .B(n2457), .Z(n2461) );
  XOR U1470 ( .A(n2617), .B(n2498), .Z(n2502) );
  MUX U1471 ( .IN0(n531), .IN1(n2656), .SEL(n2657), .F(n2532) );
  IV U1472 ( .A(n2658), .Z(n531) );
  XNOR U1473 ( .A(n2668), .B(n2547), .Z(n2551) );
  XOR U1474 ( .A(n2857), .B(n2731), .Z(n2735) );
  XNOR U1475 ( .A(n2971), .B(n2836), .Z(n2840) );
  XOR U1476 ( .A(n3012), .B(n2877), .Z(n2881) );
  XOR U1477 ( .A(n2915), .B(n2789), .Z(n2793) );
  XNOR U1478 ( .A(n2941), .B(n2820), .Z(n2814) );
  XNOR U1479 ( .A(n3060), .B(n2927), .Z(n2931) );
  XNOR U1480 ( .A(n3114), .B(n3113), .Z(n3129) );
  XNOR U1481 ( .A(n874), .B(n873), .Z(n862) );
  ANDN U1482 ( .A(n985), .B(n984), .Z(n983) );
  XOR U1483 ( .A(n1302), .B(n1309), .Z(n1373) );
  XNOR U1484 ( .A(n1575), .B(n1574), .Z(n1557) );
  XNOR U1485 ( .A(n1855), .B(n1854), .Z(n1837) );
  XNOR U1486 ( .A(n2164), .B(n2163), .Z(n2144) );
  XNOR U1487 ( .A(n2512), .B(n2511), .Z(n2494) );
  XNOR U1488 ( .A(n2891), .B(n2890), .Z(n2873) );
  MUX U1489 ( .IN0(n532), .IN1(n3090), .SEL(n3091), .F(n2954) );
  IV U1490 ( .A(n3092), .Z(n532) );
  XNOR U1491 ( .A(n3146), .B(n3145), .Z(n3121) );
  XNOR U1492 ( .A(n757), .B(n754), .Z(n753) );
  ANDN U1493 ( .A(n1274), .B(n1275), .Z(n1205) );
  XNOR U1494 ( .A(n1249), .B(n1248), .Z(n1232) );
  XNOR U1495 ( .A(n1393), .B(n1392), .Z(n1372) );
  XNOR U1496 ( .A(n1649), .B(n1648), .Z(n1624) );
  XNOR U1497 ( .A(n1740), .B(n1739), .Z(n1715) );
  XNOR U1498 ( .A(n1934), .B(n1933), .Z(n1909) );
  XNOR U1499 ( .A(n2039), .B(n2038), .Z(n2014) );
  XNOR U1500 ( .A(n2257), .B(n2256), .Z(n2232) );
  XNOR U1501 ( .A(n2297), .B(n2296), .Z(n2327) );
  XNOR U1502 ( .A(n2373), .B(n2372), .Z(n2348) );
  XNOR U1503 ( .A(n2572), .B(n2571), .Z(n2684) );
  XNOR U1504 ( .A(n2616), .B(n2615), .Z(n2591) );
  XNOR U1505 ( .A(n2744), .B(n2743), .Z(n2719) );
  MUX U1506 ( .IN0(n2937), .IN1(n533), .SEL(n2938), .F(n2808) );
  IV U1507 ( .A(n2939), .Z(n533) );
  ANDN U1508 ( .A(n717), .B(n716), .Z(n715) );
  XNOR U1509 ( .A(n782), .B(n781), .Z(n780) );
  XNOR U1510 ( .A(n891), .B(n890), .Z(n889) );
  XNOR U1511 ( .A(n991), .B(n990), .Z(n975) );
  XNOR U1512 ( .A(n1048), .B(n1047), .Z(n1033) );
  XNOR U1513 ( .A(n1170), .B(n1169), .Z(n1152) );
  XNOR U1514 ( .A(n1426), .B(n1510), .Z(n1505) );
  XOR U1515 ( .A(n1697), .B(n1694), .Z(n1775) );
  XOR U1516 ( .A(n1996), .B(n1993), .Z(n2071) );
  ANDN U1517 ( .A(n702), .B(n701), .Z(n695) );
  MUX U1518 ( .IN0(n3036), .IN1(n534), .SEL(n3037), .F(n2898) );
  IV U1519 ( .A(o_reg[1]), .Z(n534) );
  XOR U1520 ( .A(n744), .B(n748), .Z(n746) );
  XOR U1521 ( .A(n845), .B(n849), .Z(n847) );
  XOR U1522 ( .A(n968), .B(n972), .Z(n970) );
  XOR U1523 ( .A(n1144), .B(n1149), .Z(n1147) );
  XOR U1524 ( .A(n1346), .B(n1350), .Z(n1348) );
  XOR U1525 ( .A(n1584), .B(n1588), .Z(n1586) );
  XOR U1526 ( .A(n1864), .B(n1868), .Z(n1866) );
  XOR U1527 ( .A(n2173), .B(n2176), .Z(n2174) );
  XOR U1528 ( .A(n2521), .B(n2524), .Z(n2522) );
  XOR U1529 ( .A(n4528), .B(n4529), .Z(n4142) );
  MUX U1530 ( .IN0(n535), .IN1(n3692), .SEL(n3693), .F(n3654) );
  IV U1531 ( .A(n3694), .Z(n535) );
  MUX U1532 ( .IN0(n536), .IN1(n3684), .SEL(n3685), .F(n3646) );
  IV U1533 ( .A(n3686), .Z(n536) );
  MUX U1534 ( .IN0(n537), .IN1(n3705), .SEL(n3706), .F(n3667) );
  IV U1535 ( .A(n3707), .Z(n537) );
  MUX U1536 ( .IN0(n538), .IN1(n4103), .SEL(n4104), .F(n4086) );
  IV U1537 ( .A(n4105), .Z(n538) );
  MUX U1538 ( .IN0(n539), .IN1(n3659), .SEL(n3660), .F(n3621) );
  IV U1539 ( .A(n3661), .Z(n539) );
  MUX U1540 ( .IN0(n540), .IN1(n4123), .SEL(n3718), .F(n4106) );
  IV U1541 ( .A(n3716), .Z(n540) );
  MUX U1542 ( .IN0(n3700), .IN1(n541), .SEL(n3701), .F(n3662) );
  IV U1543 ( .A(n3702), .Z(n541) );
  MUX U1544 ( .IN0(n542), .IN1(n4488), .SEL(n4489), .F(n4475) );
  IV U1545 ( .A(n4490), .Z(n542) );
  XNOR U1546 ( .A(n3606), .B(n3571), .Z(n3575) );
  MUX U1547 ( .IN0(n543), .IN1(n3540), .SEL(n3541), .F(n3502) );
  IV U1548 ( .A(n3542), .Z(n543) );
  MUX U1549 ( .IN0(n544), .IN1(n4495), .SEL(n4496), .F(n4482) );
  IV U1550 ( .A(n4497), .Z(n544) );
  XNOR U1551 ( .A(n4076), .B(n4062), .Z(n4066) );
  MUX U1552 ( .IN0(n3595), .IN1(n3597), .SEL(n3596), .F(n3557) );
  MUX U1553 ( .IN0(n545), .IN1(n3553), .SEL(n3554), .F(n3515) );
  IV U1554 ( .A(n3555), .Z(n545) );
  MUX U1555 ( .IN0(n4486), .IN1(n546), .SEL(n4075), .F(n4473) );
  IV U1556 ( .A(n4074), .Z(n546) );
  MUX U1557 ( .IN0(n547), .IN1(n4035), .SEL(n4036), .F(n4018) );
  IV U1558 ( .A(n4037), .Z(n547) );
  MUX U1559 ( .IN0(n548), .IN1(n3507), .SEL(n3508), .F(n3469) );
  IV U1560 ( .A(n3509), .Z(n548) );
  MUX U1561 ( .IN0(n549), .IN1(n4876), .SEL(n4877), .F(n4855) );
  IV U1562 ( .A(n4878), .Z(n549) );
  MUX U1563 ( .IN0(n550), .IN1(n4055), .SEL(n3566), .F(n4038) );
  IV U1564 ( .A(n3564), .Z(n550) );
  MUX U1565 ( .IN0(n3548), .IN1(n551), .SEL(n3549), .F(n3510) );
  IV U1566 ( .A(n3550), .Z(n551) );
  XNOR U1567 ( .A(n3492), .B(n3457), .Z(n3461) );
  XOR U1568 ( .A(n4291), .B(n4292), .Z(n4301) );
  XOR U1569 ( .A(n4622), .B(n4623), .Z(n4306) );
  MUX U1570 ( .IN0(n552), .IN1(n4274), .SEL(n4275), .F(n4253) );
  IV U1571 ( .A(n4276), .Z(n552) );
  XOR U1572 ( .A(n4990), .B(n4991), .Z(n4871) );
  MUX U1573 ( .IN0(n553), .IN1(n3388), .SEL(n3389), .F(n3350) );
  IV U1574 ( .A(n3390), .Z(n553) );
  XNOR U1575 ( .A(n4008), .B(n3994), .Z(n3998) );
  MUX U1576 ( .IN0(n3443), .IN1(n3445), .SEL(n3444), .F(n3405) );
  MUX U1577 ( .IN0(n554), .IN1(n3401), .SEL(n3402), .F(n3363) );
  IV U1578 ( .A(n3403), .Z(n554) );
  MUX U1579 ( .IN0(n555), .IN1(n4248), .SEL(n4249), .F(n4227) );
  IV U1580 ( .A(n4250), .Z(n555) );
  MUX U1581 ( .IN0(n556), .IN1(n4599), .SEL(n4600), .F(n4588) );
  IV U1582 ( .A(n4601), .Z(n556) );
  MUX U1583 ( .IN0(n4434), .IN1(n557), .SEL(n4007), .F(n4421) );
  IV U1584 ( .A(n4006), .Z(n557) );
  MUX U1585 ( .IN0(n558), .IN1(n4410), .SEL(n4411), .F(n4397) );
  IV U1586 ( .A(n4412), .Z(n558) );
  XOR U1587 ( .A(n4977), .B(n4978), .Z(n4850) );
  MUX U1588 ( .IN0(n559), .IN1(n4970), .SEL(n4971), .F(n4957) );
  IV U1589 ( .A(n4972), .Z(n559) );
  MUX U1590 ( .IN0(n560), .IN1(n4430), .SEL(n4431), .F(n4417) );
  IV U1591 ( .A(n4432), .Z(n560) );
  MUX U1592 ( .IN0(n561), .IN1(n3967), .SEL(n3968), .F(n3950) );
  IV U1593 ( .A(n3969), .Z(n561) );
  MUX U1594 ( .IN0(n562), .IN1(n3355), .SEL(n3356), .F(n3317) );
  IV U1595 ( .A(n3357), .Z(n562) );
  XNOR U1596 ( .A(n3378), .B(n3343), .Z(n3347) );
  XOR U1597 ( .A(n4837), .B(n4819), .Z(n4823) );
  MUX U1598 ( .IN0(n563), .IN1(n4950), .SEL(n4951), .F(n4937) );
  IV U1599 ( .A(n4952), .Z(n563) );
  XOR U1600 ( .A(n4793), .B(n4794), .Z(n4803) );
  MUX U1601 ( .IN0(n564), .IN1(n3987), .SEL(n3414), .F(n3970) );
  IV U1602 ( .A(n3412), .Z(n564) );
  MUX U1603 ( .IN0(n3396), .IN1(n565), .SEL(n3397), .F(n3358) );
  IV U1604 ( .A(n3398), .Z(n565) );
  MUX U1605 ( .IN0(n4708), .IN1(n4711), .SEL(n4709), .F(n4692) );
  XOR U1606 ( .A(n4591), .B(n4583), .Z(n4224) );
  MUX U1607 ( .IN0(n5080), .IN1(n5083), .SEL(n5081), .F(n5064) );
  XOR U1608 ( .A(n4772), .B(n4773), .Z(n4782) );
  MUX U1609 ( .IN0(n566), .IN1(n4776), .SEL(n4777), .F(n4755) );
  IV U1610 ( .A(n4778), .Z(n566) );
  MUX U1611 ( .IN0(n567), .IN1(n3266), .SEL(n3267), .F(n3228) );
  IV U1612 ( .A(n3268), .Z(n567) );
  XNOR U1613 ( .A(n3310), .B(n3309), .Z(n3322) );
  MUX U1614 ( .IN0(n3819), .IN1(n3834), .SEL(n3821), .F(n3794) );
  MUX U1615 ( .IN0(n3862), .IN1(n3865), .SEL(n3863), .F(n3845) );
  MUX U1616 ( .IN0(n4649), .IN1(n4659), .SEL(n4651), .F(n4637) );
  XOR U1617 ( .A(n4230), .B(n4212), .Z(n4216) );
  MUX U1618 ( .IN0(n5170), .IN1(n5173), .SEL(n5171), .F(n5154) );
  MUX U1619 ( .IN0(n5021), .IN1(n5031), .SEL(n5023), .F(n5009) );
  MUX U1620 ( .IN0(n4948), .IN1(n568), .SEL(n4789), .F(n4935) );
  IV U1621 ( .A(n4787), .Z(n568) );
  XNOR U1622 ( .A(n3940), .B(n3926), .Z(n3930) );
  MUX U1623 ( .IN0(n3291), .IN1(n3293), .SEL(n3292), .F(n3253) );
  MUX U1624 ( .IN0(n569), .IN1(n3249), .SEL(n3250), .F(n3182) );
  IV U1625 ( .A(n3251), .Z(n569) );
  MUX U1626 ( .IN0(n570), .IN1(n4173), .SEL(n4174), .F(n4156) );
  IV U1627 ( .A(n4175), .Z(n570) );
  XOR U1628 ( .A(n4698), .B(n4699), .Z(n4347) );
  MUX U1629 ( .IN0(n571), .IN1(n4560), .SEL(n4561), .F(n4547) );
  IV U1630 ( .A(n4562), .Z(n571) );
  XOR U1631 ( .A(n4567), .B(n4568), .Z(n4201) );
  XOR U1632 ( .A(n5185), .B(g_input[3]), .Z(n5186) );
  MUX U1633 ( .IN0(n4382), .IN1(n572), .SEL(n3939), .F(n4369) );
  IV U1634 ( .A(n3938), .Z(n572) );
  MUX U1635 ( .IN0(n573), .IN1(n4366), .SEL(n4367), .F(n3899) );
  IV U1636 ( .A(n4368), .Z(n573) );
  XOR U1637 ( .A(n5070), .B(n5071), .Z(n4912) );
  MUX U1638 ( .IN0(n574), .IN1(n4918), .SEL(n4919), .F(n3132) );
  IV U1639 ( .A(n4920), .Z(n574) );
  MUX U1640 ( .IN0(n575), .IN1(n4731), .SEL(n4732), .F(n3116) );
  IV U1641 ( .A(n4733), .Z(n575) );
  MUX U1642 ( .IN0(n576), .IN1(n3199), .SEL(n3200), .F(n3070) );
  IV U1643 ( .A(n3201), .Z(n576) );
  MUX U1644 ( .IN0(n3234), .IN1(n3232), .SEL(n3233), .F(n3195) );
  MUX U1645 ( .IN0(n577), .IN1(n3215), .SEL(n3216), .F(n3087) );
  IV U1646 ( .A(n3217), .Z(n577) );
  XOR U1647 ( .A(n3851), .B(n3852), .Z(n3798) );
  XNOR U1648 ( .A(n4327), .B(n4317), .Z(n4321) );
  XOR U1649 ( .A(n4633), .B(n4634), .Z(n4325) );
  XOR U1650 ( .A(n4556), .B(n4557), .Z(n4180) );
  MUX U1651 ( .IN0(n578), .IN1(n1053), .SEL(n1054), .F(n994) );
  IV U1652 ( .A(n1055), .Z(n578) );
  MUX U1653 ( .IN0(n579), .IN1(n1227), .SEL(n1228), .F(n1165) );
  IV U1654 ( .A(n1229), .Z(n579) );
  MUX U1655 ( .IN0(n580), .IN1(n1314), .SEL(n1315), .F(n1244) );
  IV U1656 ( .A(n1316), .Z(n580) );
  MUX U1657 ( .IN0(n581), .IN1(n1526), .SEL(n1527), .F(n1440) );
  IV U1658 ( .A(n1528), .Z(n581) );
  MUX U1659 ( .IN0(n582), .IN1(n1560), .SEL(n1561), .F(n1475) );
  IV U1660 ( .A(n1562), .Z(n582) );
  MUX U1661 ( .IN0(n583), .IN1(n1569), .SEL(n1570), .F(n1484) );
  IV U1662 ( .A(n1571), .Z(n583) );
  MUX U1663 ( .IN0(n584), .IN1(n1627), .SEL(n1628), .F(n1534) );
  IV U1664 ( .A(n1629), .Z(n584) );
  MUX U1665 ( .IN0(n585), .IN1(n1644), .SEL(n1645), .F(n1552) );
  IV U1666 ( .A(n1646), .Z(n585) );
  MUX U1667 ( .IN0(n586), .IN1(n1896), .SEL(n1897), .F(n1799) );
  IV U1668 ( .A(n1898), .Z(n586) );
  MUX U1669 ( .IN0(n587), .IN1(n1946), .SEL(n1947), .F(n1849) );
  IV U1670 ( .A(n1948), .Z(n587) );
  MUX U1671 ( .IN0(n588), .IN1(n2034), .SEL(n2035), .F(n1929) );
  IV U1672 ( .A(n2036), .Z(n588) );
  MUX U1673 ( .IN0(n589), .IN1(n2017), .SEL(n2018), .F(n1912) );
  IV U1674 ( .A(n2019), .Z(n589) );
  MUX U1675 ( .IN0(n590), .IN1(n2318), .SEL(n2319), .F(n2206) );
  IV U1676 ( .A(n2320), .Z(n590) );
  MUX U1677 ( .IN0(n591), .IN1(n2335), .SEL(n2336), .F(n2219) );
  IV U1678 ( .A(n2337), .Z(n591) );
  MUX U1679 ( .IN0(n592), .IN1(n2385), .SEL(n2386), .F(n2269) );
  IV U1680 ( .A(n2387), .Z(n592) );
  MUX U1681 ( .IN0(n593), .IN1(n2408), .SEL(n2409), .F(n2292) );
  IV U1682 ( .A(n2410), .Z(n593) );
  MUX U1683 ( .IN0(n594), .IN1(n2489), .SEL(n2490), .F(n2368) );
  IV U1684 ( .A(n2491), .Z(n594) );
  MUX U1685 ( .IN0(n595), .IN1(n2472), .SEL(n2473), .F(n2351) );
  IV U1686 ( .A(n2474), .Z(n595) );
  MUX U1687 ( .IN0(n596), .IN1(n2835), .SEL(n2836), .F(n2706) );
  IV U1688 ( .A(n2837), .Z(n596) );
  MUX U1689 ( .IN0(n597), .IN1(n2885), .SEL(n2886), .F(n2756) );
  IV U1690 ( .A(n2887), .Z(n597) );
  MUX U1691 ( .IN0(n598), .IN1(n2989), .SEL(n2990), .F(n2851) );
  IV U1692 ( .A(n2991), .Z(n598) );
  MUX U1693 ( .IN0(n599), .IN1(n3006), .SEL(n3007), .F(n2868) );
  IV U1694 ( .A(n3008), .Z(n599) );
  MUX U1695 ( .IN0(n600), .IN1(n2926), .SEL(n2927), .F(n2797) );
  IV U1696 ( .A(n2928), .Z(n600) );
  MUX U1697 ( .IN0(n601), .IN1(n2909), .SEL(n2910), .F(n2780) );
  IV U1698 ( .A(n2911), .Z(n601) );
  XOR U1699 ( .A(n5160), .B(n5161), .Z(n5099) );
  XNOR U1700 ( .A(n4892), .B(n4882), .Z(n4886) );
  XOR U1701 ( .A(n5003), .B(n5004), .Z(n4890) );
  XOR U1702 ( .A(n4739), .B(n4740), .Z(n4745) );
  MUX U1703 ( .IN0(n4364), .IN1(n602), .SEL(n4363), .F(n4354) );
  IV U1704 ( .A(n4362), .Z(n602) );
  MUX U1705 ( .IN0(n603), .IN1(n3919), .SEL(n3262), .F(n3902) );
  IV U1706 ( .A(n3260), .Z(n603) );
  XOR U1707 ( .A(n3800), .B(n3782), .Z(n3786) );
  XNOR U1708 ( .A(n3875), .B(n3761), .Z(n3765) );
  XNOR U1709 ( .A(n4163), .B(n4147), .Z(n4153) );
  XOR U1710 ( .A(n4541), .B(n4542), .Z(n4161) );
  XOR U1711 ( .A(n2061), .B(n2166), .Z(n2062) );
  MUX U1712 ( .IN0(n604), .IN1(n2695), .SEL(n2696), .F(n2567) );
  IV U1713 ( .A(n2697), .Z(n604) );
  XOR U1714 ( .A(n2766), .B(n2893), .Z(n2767) );
  XNOR U1715 ( .A(n5183), .B(n3159), .Z(n3163) );
  XOR U1716 ( .A(n5101), .B(n3150), .Z(n3154) );
  XNOR U1717 ( .A(n4721), .B(n3109), .Z(n3113) );
  MUX U1718 ( .IN0(n3177), .IN1(n605), .SEL(n3178), .F(n3048) );
  IV U1719 ( .A(n3179), .Z(n605) );
  MUX U1720 ( .IN0(n606), .IN1(n831), .SEL(n832), .F(n789) );
  IV U1721 ( .A(n833), .Z(n606) );
  MUX U1722 ( .IN0(n607), .IN1(n857), .SEL(n858), .F(n823) );
  IV U1723 ( .A(n859), .Z(n607) );
  XNOR U1724 ( .A(n952), .B(n911), .Z(n915) );
  XOR U1725 ( .A(n1000), .B(n945), .Z(n950) );
  XNOR U1726 ( .A(n1128), .B(n1071), .Z(n1075) );
  XOR U1727 ( .A(n1182), .B(n1122), .Z(n1126) );
  XNOR U1728 ( .A(n1285), .B(n1220), .Z(n1224) );
  XNOR U1729 ( .A(n1329), .B(n1262), .Z(n1266) );
  NAND U1730 ( .A(n1308), .B(n1375), .Z(n1374) );
  XOR U1731 ( .A(n1394), .B(n1323), .Z(n1327) );
  XNOR U1732 ( .A(n1516), .B(n1433), .Z(n1437) );
  XOR U1733 ( .A(n1633), .B(n1548), .Z(n1542) );
  XOR U1734 ( .A(n1692), .B(n1693), .Z(n1687) );
  XOR U1735 ( .A(n1838), .B(n1744), .Z(n1748) );
  XOR U1736 ( .A(n1789), .B(n1790), .Z(n1786) );
  XOR U1737 ( .A(n1918), .B(n1824), .Z(n1828) );
  NAND U1738 ( .A(n1971), .B(n2074), .Z(n2073) );
  XNOR U1739 ( .A(n2085), .B(n1983), .Z(n1987) );
  XOR U1740 ( .A(n2145), .B(n2043), .Z(n2047) );
  XOR U1741 ( .A(n2241), .B(n2131), .Z(n2135) );
  NAND U1742 ( .A(n2192), .B(n2303), .Z(n2302) );
  XNOR U1743 ( .A(n2423), .B(n2311), .Z(n2315) );
  XOR U1744 ( .A(n2495), .B(n2377), .Z(n2381) );
  XOR U1745 ( .A(n2600), .B(n2481), .Z(n2485) );
  XOR U1746 ( .A(n2659), .B(n2538), .Z(n2542) );
  XOR U1747 ( .A(n2874), .B(n2748), .Z(n2752) );
  XOR U1748 ( .A(n2995), .B(n2860), .Z(n2864) );
  XOR U1749 ( .A(n3051), .B(n2918), .Z(n2922) );
  XNOR U1750 ( .A(n3077), .B(n2944), .Z(n2948) );
  MUX U1751 ( .IN0(n608), .IN1(n799), .SEL(n800), .F(n768) );
  IV U1752 ( .A(n801), .Z(n608) );
  XNOR U1753 ( .A(n837), .B(n836), .Z(n827) );
  AND U1754 ( .A(n986), .B(n987), .Z(n982) );
  XNOR U1755 ( .A(n960), .B(n959), .Z(n942) );
  XNOR U1756 ( .A(n1018), .B(n1017), .Z(n999) );
  XNOR U1757 ( .A(n1136), .B(n1135), .Z(n1118) );
  XNOR U1758 ( .A(n1199), .B(n1198), .Z(n1181) );
  XNOR U1759 ( .A(n1337), .B(n1336), .Z(n1319) );
  XNOR U1760 ( .A(n1365), .B(n1364), .Z(n1382) );
  XNOR U1761 ( .A(n1411), .B(n1410), .Z(n1393) );
  XNOR U1762 ( .A(n1667), .B(n1666), .Z(n1649) );
  XNOR U1763 ( .A(n1617), .B(n1616), .Z(n1632) );
  XNOR U1764 ( .A(n1805), .B(n1804), .Z(n1820) );
  XNOR U1765 ( .A(n1952), .B(n1951), .Z(n1934) );
  XNOR U1766 ( .A(n1902), .B(n1901), .Z(n1917) );
  XNOR U1767 ( .A(n2112), .B(n2111), .Z(n2127) );
  XNOR U1768 ( .A(n2225), .B(n2224), .Z(n2240) );
  XNOR U1769 ( .A(n2275), .B(n2274), .Z(n2257) );
  XNOR U1770 ( .A(n2431), .B(n2430), .Z(n2413) );
  XNOR U1771 ( .A(n2462), .B(n2461), .Z(n2477) );
  XNOR U1772 ( .A(n2552), .B(n2551), .Z(n2534) );
  XNOR U1773 ( .A(n2634), .B(n2633), .Z(n2616) );
  XNOR U1774 ( .A(n2584), .B(n2583), .Z(n2599) );
  XNOR U1775 ( .A(n2841), .B(n2840), .Z(n2856) );
  XNOR U1776 ( .A(n2803), .B(n2802), .Z(n2785) );
  XNOR U1777 ( .A(n2829), .B(n2957), .Z(n2830) );
  XNOR U1778 ( .A(n2979), .B(n2978), .Z(n2994) );
  XNOR U1779 ( .A(n2932), .B(n2931), .Z(n2914) );
  OR U1780 ( .A(n853), .B(n854), .Z(n812) );
  XOR U1781 ( .A(n1109), .B(n1106), .Z(n1153) );
  XNOR U1782 ( .A(n1472), .B(n1471), .Z(n1445) );
  ANDN U1783 ( .A(n1862), .B(n1863), .Z(n1767) );
  NANDN U1784 ( .B(n1891), .A(n1892), .Z(n1794) );
  XNOR U1785 ( .A(n1837), .B(n1836), .Z(n1812) );
  XNOR U1786 ( .A(n2144), .B(n2143), .Z(n2119) );
  XNOR U1787 ( .A(n2325), .B(n2439), .Z(n2326) );
  ANDN U1788 ( .A(n2519), .B(n2520), .Z(n2398) );
  XNOR U1789 ( .A(n2494), .B(n2493), .Z(n2469) );
  XNOR U1790 ( .A(n2658), .B(n2657), .Z(n2702) );
  XNOR U1791 ( .A(n2873), .B(n2872), .Z(n2848) );
  XNOR U1792 ( .A(n3011), .B(n3010), .Z(n2986) );
  MUX U1793 ( .IN0(n3073), .IN1(n609), .SEL(n3074), .F(n2937) );
  IV U1794 ( .A(n3075), .Z(n609) );
  MUX U1795 ( .IN0(n736), .IN1(n734), .SEL(n735), .F(n716) );
  XNOR U1796 ( .A(n731), .B(n730), .Z(n729) );
  XNOR U1797 ( .A(n1531), .B(n1530), .Z(n1514) );
  XNOR U1798 ( .A(n1715), .B(n1714), .Z(n1696) );
  XNOR U1799 ( .A(n2014), .B(n2013), .Z(n1995) );
  XNOR U1800 ( .A(n2348), .B(n2347), .Z(n2323) );
  XNOR U1801 ( .A(n2719), .B(n2718), .Z(n2683) );
  XNOR U1802 ( .A(n780), .B(n779), .Z(n807) );
  XNOR U1803 ( .A(n889), .B(n888), .Z(n927) );
  XNOR U1804 ( .A(n1033), .B(n1032), .Z(n1087) );
  XOR U1805 ( .A(n1214), .B(n1213), .Z(n1279) );
  XNOR U1806 ( .A(n688), .B(n689), .Z(n690) );
  XOR U1807 ( .A(n773), .B(n777), .Z(n775) );
  XOR U1808 ( .A(n882), .B(n886), .Z(n884) );
  XOR U1809 ( .A(n1026), .B(n1030), .Z(n1028) );
  XOR U1810 ( .A(n1207), .B(n1211), .Z(n1209) );
  XOR U1811 ( .A(n1420), .B(n1424), .Z(n1422) );
  XOR U1812 ( .A(n1676), .B(n1680), .Z(n1678) );
  XOR U1813 ( .A(n1961), .B(n1964), .Z(n1962) );
  XOR U1814 ( .A(n2284), .B(n2287), .Z(n2285) );
  XOR U1815 ( .A(n2643), .B(n2646), .Z(n2644) );
  MUX U1816 ( .IN0(n610), .IN1(n3722), .SEL(n3723), .F(n3684) );
  IV U1817 ( .A(n3724), .Z(n610) );
  MUX U1818 ( .IN0(n611), .IN1(n4112), .SEL(n4113), .F(n4095) );
  IV U1819 ( .A(n4114), .Z(n611) );
  XNOR U1820 ( .A(n3728), .B(n3727), .Z(n3740) );
  XNOR U1821 ( .A(n4135), .B(n4134), .Z(n3754) );
  XNOR U1822 ( .A(n3690), .B(n3689), .Z(n3702) );
  XNOR U1823 ( .A(n4118), .B(n4117), .Z(n3716) );
  XOR U1824 ( .A(n3703), .B(n3668), .Z(n3672) );
  MUX U1825 ( .IN0(n612), .IN1(n3621), .SEL(n3622), .F(n3583) );
  IV U1826 ( .A(n3623), .Z(n612) );
  XNOR U1827 ( .A(n3652), .B(n3651), .Z(n3664) );
  MUX U1828 ( .IN0(n613), .IN1(n3570), .SEL(n3571), .F(n3532) );
  IV U1829 ( .A(n3572), .Z(n613) );
  XNOR U1830 ( .A(n4101), .B(n4100), .Z(n3678) );
  XNOR U1831 ( .A(n3614), .B(n3613), .Z(n3626) );
  MUX U1832 ( .IN0(n4499), .IN1(n614), .SEL(n4092), .F(n4486) );
  IV U1833 ( .A(n4091), .Z(n614) );
  XNOR U1834 ( .A(n4084), .B(n4083), .Z(n3640) );
  MUX U1835 ( .IN0(n615), .IN1(n4044), .SEL(n4045), .F(n4027) );
  IV U1836 ( .A(n4046), .Z(n615) );
  XNOR U1837 ( .A(n3576), .B(n3575), .Z(n3588) );
  MUX U1838 ( .IN0(n616), .IN1(n4462), .SEL(n4463), .F(n4449) );
  IV U1839 ( .A(n4464), .Z(n616) );
  MUX U1840 ( .IN0(n617), .IN1(n4482), .SEL(n4483), .F(n4469) );
  IV U1841 ( .A(n4484), .Z(n617) );
  XNOR U1842 ( .A(n4067), .B(n4066), .Z(n3602) );
  XOR U1843 ( .A(n3589), .B(n3554), .Z(n3558) );
  XNOR U1844 ( .A(n3538), .B(n3537), .Z(n3550) );
  XNOR U1845 ( .A(n4050), .B(n4049), .Z(n3564) );
  MUX U1846 ( .IN0(n618), .IN1(n3469), .SEL(n3470), .F(n3431) );
  IV U1847 ( .A(n3471), .Z(n618) );
  XNOR U1848 ( .A(n3500), .B(n3499), .Z(n3512) );
  XOR U1849 ( .A(n4452), .B(n4444), .Z(n4024) );
  MUX U1850 ( .IN0(n619), .IN1(n4855), .SEL(n4856), .F(n4834) );
  IV U1851 ( .A(n4857), .Z(n619) );
  MUX U1852 ( .IN0(n620), .IN1(n3418), .SEL(n3419), .F(n3380) );
  IV U1853 ( .A(n3420), .Z(n620) );
  XNOR U1854 ( .A(n4033), .B(n4032), .Z(n3526) );
  XNOR U1855 ( .A(n3462), .B(n3461), .Z(n3474) );
  MUX U1856 ( .IN0(n621), .IN1(n4269), .SEL(n4270), .F(n4248) );
  IV U1857 ( .A(n4271), .Z(n621) );
  XOR U1858 ( .A(n4424), .B(n4425), .Z(n4006) );
  MUX U1859 ( .IN0(n622), .IN1(n4983), .SEL(n4984), .F(n4970) );
  IV U1860 ( .A(n4985), .Z(n622) );
  XNOR U1861 ( .A(n4016), .B(n4015), .Z(n3488) );
  XOR U1862 ( .A(n3475), .B(n3440), .Z(n3444) );
  MUX U1863 ( .IN0(n623), .IN1(n3976), .SEL(n3977), .F(n3959) );
  IV U1864 ( .A(n3978), .Z(n623) );
  XNOR U1865 ( .A(n3424), .B(n3423), .Z(n3436) );
  XOR U1866 ( .A(n4611), .B(n4612), .Z(n4285) );
  XOR U1867 ( .A(n4411), .B(n4412), .Z(n3989) );
  XOR U1868 ( .A(n4858), .B(n4840), .Z(n4844) );
  MUX U1869 ( .IN0(n624), .IN1(n4963), .SEL(n4964), .F(n4950) );
  IV U1870 ( .A(n4965), .Z(n624) );
  XNOR U1871 ( .A(n3999), .B(n3998), .Z(n3450) );
  XNOR U1872 ( .A(n3386), .B(n3385), .Z(n3398) );
  XOR U1873 ( .A(n4600), .B(n4601), .Z(n4264) );
  MUX U1874 ( .IN0(n625), .IN1(n5159), .SEL(n5160), .F(n5142) );
  IV U1875 ( .A(n5161), .Z(n625) );
  MUX U1876 ( .IN0(n626), .IN1(n3312), .SEL(n3313), .F(n3274) );
  IV U1877 ( .A(n3314), .Z(n626) );
  MUX U1878 ( .IN0(n627), .IN1(n4417), .SEL(n4418), .F(n4404) );
  IV U1879 ( .A(n4419), .Z(n627) );
  XNOR U1880 ( .A(n3982), .B(n3981), .Z(n3412) );
  MUX U1881 ( .IN0(n628), .IN1(n3317), .SEL(n3318), .F(n3279) );
  IV U1882 ( .A(n3319), .Z(n628) );
  XNOR U1883 ( .A(n3348), .B(n3347), .Z(n3360) );
  XNOR U1884 ( .A(n3340), .B(n3305), .Z(n3309) );
  MUX U1885 ( .IN0(n629), .IN1(n4582), .SEL(n4583), .F(n4571) );
  IV U1886 ( .A(n4584), .Z(n629) );
  XOR U1887 ( .A(n4251), .B(n4233), .Z(n4237) );
  MUX U1888 ( .IN0(n4961), .IN1(n630), .SEL(n4810), .F(n4948) );
  IV U1889 ( .A(n4808), .Z(n630) );
  MUX U1890 ( .IN0(n631), .IN1(n4771), .SEL(n4772), .F(n4750) );
  IV U1891 ( .A(n4773), .Z(n631) );
  XNOR U1892 ( .A(n3965), .B(n3964), .Z(n3374) );
  XOR U1893 ( .A(n3361), .B(n3326), .Z(n3330) );
  MUX U1894 ( .IN0(n632), .IN1(n4185), .SEL(n4186), .F(n4173) );
  IV U1895 ( .A(n4187), .Z(n632) );
  MUX U1896 ( .IN0(n4329), .IN1(n4332), .SEL(n4330), .F(n4316) );
  MUX U1897 ( .IN0(n4643), .IN1(n4665), .SEL(n4645), .F(n4632) );
  XOR U1898 ( .A(n4578), .B(n4579), .Z(n4222) );
  XOR U1899 ( .A(n4387), .B(n4379), .Z(n3939) );
  MUX U1900 ( .IN0(n633), .IN1(n4371), .SEL(n4372), .F(n4366) );
  IV U1901 ( .A(n4373), .Z(n633) );
  MUX U1902 ( .IN0(n5118), .IN1(n5133), .SEL(n5120), .F(n5105) );
  MUX U1903 ( .IN0(n4894), .IN1(n4897), .SEL(n4895), .F(n4881) );
  MUX U1904 ( .IN0(n5015), .IN1(n5037), .SEL(n5017), .F(n5002) );
  XOR U1905 ( .A(n4795), .B(n4777), .Z(n4781) );
  MUX U1906 ( .IN0(n634), .IN1(n4931), .SEL(n4932), .F(n4918) );
  IV U1907 ( .A(n4933), .Z(n634) );
  XNOR U1908 ( .A(n3948), .B(n3947), .Z(n3336) );
  MUX U1909 ( .IN0(n635), .IN1(n3905), .SEL(n3906), .F(n3207) );
  IV U1910 ( .A(n3907), .Z(n635) );
  MUX U1911 ( .IN0(n3794), .IN1(n3818), .SEL(n3796), .F(n3773) );
  MUX U1912 ( .IN0(n3802), .IN1(n3812), .SEL(n3804), .F(n3781) );
  XOR U1913 ( .A(n4706), .B(n4693), .Z(n4348) );
  MUX U1914 ( .IN0(n636), .IN1(n4555), .SEL(n4556), .F(n4540) );
  IV U1915 ( .A(n4557), .Z(n636) );
  MUX U1916 ( .IN0(g_input[1]), .IN1(n5203), .SEL(g_input[31]), .F(n3854) );
  XOR U1917 ( .A(n5078), .B(n5065), .Z(n4913) );
  XOR U1918 ( .A(n4925), .B(n4926), .Z(n4766) );
  MUX U1919 ( .IN0(e_input[1]), .IN1(n637), .SEL(e_input[31]), .F(n4352) );
  IV U1920 ( .A(n4719), .Z(n637) );
  XNOR U1921 ( .A(n3931), .B(n3930), .Z(n3298) );
  XOR U1922 ( .A(n3860), .B(n3846), .Z(n3799) );
  XNOR U1923 ( .A(n3882), .B(n3883), .Z(n3764) );
  XOR U1924 ( .A(n4647), .B(n4638), .Z(n4326) );
  XOR U1925 ( .A(n4188), .B(n4166), .Z(n4170) );
  MUX U1926 ( .IN0(n638), .IN1(n1113), .SEL(n1114), .F(n1053) );
  IV U1927 ( .A(n1115), .Z(n638) );
  MUX U1928 ( .IN0(n639), .IN1(n1202), .SEL(n1203), .F(n1139) );
  IV U1929 ( .A(n1204), .Z(n639) );
  MUX U1930 ( .IN0(n640), .IN1(n1219), .SEL(n1220), .F(n1155) );
  IV U1931 ( .A(n1221), .Z(n640) );
  MUX U1932 ( .IN0(n641), .IN1(n1388), .SEL(n1389), .F(n1314) );
  IV U1933 ( .A(n1390), .Z(n641) );
  MUX U1934 ( .IN0(n642), .IN1(n1735), .SEL(n1736), .F(n1644) );
  IV U1935 ( .A(n1737), .Z(n642) );
  MUX U1936 ( .IN0(n643), .IN1(n1752), .SEL(n1753), .F(n1661) );
  IV U1937 ( .A(n1754), .Z(n643) );
  MUX U1938 ( .IN0(n644), .IN1(n1702), .SEL(n1703), .F(n1611) );
  IV U1939 ( .A(n1704), .Z(n644) );
  MUX U1940 ( .IN0(n645), .IN1(n1718), .SEL(n1719), .F(n1627) );
  IV U1941 ( .A(n1720), .Z(n645) );
  MUX U1942 ( .IN0(n646), .IN1(n2087), .SEL(n2088), .F(n1982) );
  IV U1943 ( .A(n2089), .Z(n646) );
  MUX U1944 ( .IN0(n647), .IN1(n2122), .SEL(n2123), .F(n2017) );
  IV U1945 ( .A(n2124), .Z(n647) );
  MUX U1946 ( .IN0(n648), .IN1(n2106), .SEL(n2107), .F(n2001) );
  IV U1947 ( .A(n2108), .Z(n648) );
  MUX U1948 ( .IN0(n649), .IN1(n2156), .SEL(n2157), .F(n2051) );
  IV U1949 ( .A(n2158), .Z(n649) );
  MUX U1950 ( .IN0(n650), .IN1(n2139), .SEL(n2140), .F(n2034) );
  IV U1951 ( .A(n2141), .Z(n650) );
  MUX U1952 ( .IN0(n651), .IN1(n2227), .SEL(n2228), .F(n2114) );
  IV U1953 ( .A(n2229), .Z(n651) );
  MUX U1954 ( .IN0(n652), .IN1(n2546), .SEL(n2547), .F(n2425) );
  IV U1955 ( .A(n2548), .Z(n652) );
  MUX U1956 ( .IN0(n653), .IN1(n2554), .SEL(n2555), .F(n2433) );
  IV U1957 ( .A(n2556), .Z(n653) );
  MUX U1958 ( .IN0(n654), .IN1(n2529), .SEL(n2530), .F(n2408) );
  IV U1959 ( .A(n2531), .Z(n654) );
  MUX U1960 ( .IN0(n655), .IN1(n2594), .SEL(n2595), .F(n2472) );
  IV U1961 ( .A(n2596), .Z(n655) );
  MUX U1962 ( .IN0(n656), .IN1(n2578), .SEL(n2579), .F(n2456) );
  IV U1963 ( .A(n2580), .Z(n656) );
  MUX U1964 ( .IN0(n657), .IN1(n2628), .SEL(n2629), .F(n2506) );
  IV U1965 ( .A(n2630), .Z(n657) );
  MUX U1966 ( .IN0(n658), .IN1(n2611), .SEL(n2612), .F(n2489) );
  IV U1967 ( .A(n2613), .Z(n658) );
  MUX U1968 ( .IN0(n659), .IN1(n2981), .SEL(n2982), .F(n2843) );
  IV U1969 ( .A(n2983), .Z(n659) );
  MUX U1970 ( .IN0(g_input[9]), .IN1(n4995), .SEL(g_input[31]), .F(n2276) );
  MUX U1971 ( .IN0(e_input[24]), .IN1(n5181), .SEL(e_input[31]), .F(n1002) );
  MUX U1972 ( .IN0(e_input[25]), .IN1(n5182), .SEL(e_input[31]), .F(n948) );
  MUX U1973 ( .IN0(g_input[8]), .IN1(n5007), .SEL(g_input[31]), .F(n2392) );
  MUX U1974 ( .IN0(e_input[27]), .IN1(n5166), .SEL(e_input[31]), .F(n660) );
  IV U1975 ( .A(n660), .Z(n856) );
  MUX U1976 ( .IN0(g_input[6]), .IN1(n5116), .SEL(g_input[31]), .F(n2635) );
  MUX U1977 ( .IN0(e_input[26]), .IN1(n5167), .SEL(e_input[31]), .F(n894) );
  MUX U1978 ( .IN0(g_input[7]), .IN1(n5104), .SEL(g_input[31]), .F(n2513) );
  MUX U1979 ( .IN0(n661), .IN1(n3141), .SEL(n3142), .F(n3006) );
  IV U1980 ( .A(n3143), .Z(n661) );
  MUX U1981 ( .IN0(g_input[2]), .IN1(n5195), .SEL(g_input[31]), .F(n3165) );
  MUX U1982 ( .IN0(g_input[3]), .IN1(n5186), .SEL(g_input[31]), .F(n662) );
  IV U1983 ( .A(n662), .Z(n3030) );
  MUX U1984 ( .IN0(g_input[5]), .IN1(n5135), .SEL(g_input[31]), .F(n2763) );
  MUX U1985 ( .IN0(n663), .IN1(n3158), .SEL(n3159), .F(n3023) );
  IV U1986 ( .A(n3160), .Z(n663) );
  MUX U1987 ( .IN0(g_input[4]), .IN1(n5152), .SEL(g_input[31]), .F(n664) );
  IV U1988 ( .A(n664), .Z(n2892) );
  MUX U1989 ( .IN0(g_input[10]), .IN1(n4981), .SEL(g_input[31]), .F(n2165) );
  MUX U1990 ( .IN0(g_input[11]), .IN1(n4969), .SEL(g_input[31]), .F(n2058) );
  MUX U1991 ( .IN0(e_input[20]), .IN1(n4905), .SEL(e_input[31]), .F(n1218) );
  MUX U1992 ( .IN0(g_input[13]), .IN1(n4943), .SEL(g_input[31]), .F(n1856) );
  MUX U1993 ( .IN0(n665), .IN1(n3108), .SEL(n3109), .F(n2973) );
  IV U1994 ( .A(n3110), .Z(n665) );
  MUX U1995 ( .IN0(e_input[21]), .IN1(n4906), .SEL(e_input[31]), .F(n1158) );
  MUX U1996 ( .IN0(g_input[12]), .IN1(n4955), .SEL(g_input[31]), .F(n1953) );
  MUX U1997 ( .IN0(g_input[14]), .IN1(n4929), .SEL(g_input[31]), .F(n1761) );
  MUX U1998 ( .IN0(g_input[15]), .IN1(n4917), .SEL(g_input[31]), .F(n1668) );
  MUX U1999 ( .IN0(n666), .IN1(n3124), .SEL(n3125), .F(n2989) );
  IV U2000 ( .A(n3126), .Z(n666) );
  MUX U2001 ( .IN0(g_input[17]), .IN1(n4533), .SEL(g_input[31]), .F(n1491) );
  MUX U2002 ( .IN0(e_input[16]), .IN1(n5091), .SEL(e_input[31]), .F(n1546) );
  MUX U2003 ( .IN0(e_input[17]), .IN1(n5092), .SEL(e_input[31]), .F(n1457) );
  MUX U2004 ( .IN0(g_input[16]), .IN1(n4545), .SEL(g_input[31]), .F(n1576) );
  MUX U2005 ( .IN0(g_input[19]), .IN1(n4507), .SEL(g_input[31]), .F(n1338) );
  MUX U2006 ( .IN0(n667), .IN1(n3070), .SEL(n3071), .F(n2934) );
  IV U2007 ( .A(n3072), .Z(n667) );
  MUX U2008 ( .IN0(g_input[18]), .IN1(n4519), .SEL(g_input[31]), .F(n1412) );
  MUX U2009 ( .IN0(e_input[12]), .IN1(n3888), .SEL(e_input[31]), .F(n1880) );
  MUX U2010 ( .IN0(g_input[21]), .IN1(n4481), .SEL(g_input[31]), .F(n1200) );
  MUX U2011 ( .IN0(n668), .IN1(n3062), .SEL(n3063), .F(n2926) );
  IV U2012 ( .A(n3064), .Z(n668) );
  MUX U2013 ( .IN0(g_input[20]), .IN1(n4493), .SEL(g_input[31]), .F(n1268) );
  MUX U2014 ( .IN0(g_input[23]), .IN1(n4455), .SEL(g_input[31]), .F(n1077) );
  MUX U2015 ( .IN0(n669), .IN1(n3045), .SEL(n3046), .F(n2909) );
  IV U2016 ( .A(n3047), .Z(n669) );
  MUX U2017 ( .IN0(g_input[22]), .IN1(n4467), .SEL(g_input[31]), .F(n1137) );
  MUX U2018 ( .IN0(e_input[8]), .IN1(n3873), .SEL(e_input[31]), .F(n2304) );
  MUX U2019 ( .IN0(g_input[25]), .IN1(n4429), .SEL(g_input[31]), .F(n961) );
  MUX U2020 ( .IN0(n670), .IN1(n3053), .SEL(n3054), .F(n2917) );
  IV U2021 ( .A(n3055), .Z(n670) );
  MUX U2022 ( .IN0(e_input[9]), .IN1(n3874), .SEL(e_input[31]), .F(n2190) );
  MUX U2023 ( .IN0(g_input[24]), .IN1(n4441), .SEL(g_input[31]), .F(n1019) );
  MUX U2024 ( .IN0(e_input[4]), .IN1(n4340), .SEL(e_input[31]), .F(n2818) );
  MUX U2025 ( .IN0(g_input[26]), .IN1(n4415), .SEL(g_input[31]), .F(n917) );
  MUX U2026 ( .IN0(g_input[27]), .IN1(n4403), .SEL(g_input[31]), .F(n875) );
  XOR U2027 ( .A(n5168), .B(n5155), .Z(n5100) );
  XOR U2028 ( .A(n5019), .B(n5010), .Z(n4891) );
  MUX U2029 ( .IN0(n3197), .IN1(n3195), .SEL(n3196), .F(n3066) );
  MUX U2030 ( .IN0(n3186), .IN1(n3188), .SEL(n3187), .F(n3057) );
  XNOR U2031 ( .A(n3911), .B(n3910), .Z(n3260) );
  MUX U2032 ( .IN0(n3244), .IN1(n671), .SEL(n3245), .F(n3177) );
  IV U2033 ( .A(n3246), .Z(n671) );
  XNOR U2034 ( .A(n4322), .B(n4321), .Z(n3895) );
  XOR U2035 ( .A(n4558), .B(n4548), .Z(n4162) );
  MUX U2036 ( .IN0(e_input[28]), .IN1(n5200), .SEL(e_input[31]), .F(n830) );
  MUX U2037 ( .IN0(e_input[29]), .IN1(n5201), .SEL(e_input[31]), .F(n793) );
  MUX U2038 ( .IN0(n672), .IN1(n877), .SEL(n878), .F(n840) );
  IV U2039 ( .A(n879), .Z(n672) );
  MUX U2040 ( .IN0(g_input[28]), .IN1(n4389), .SEL(g_input[31]), .F(n838) );
  MUX U2041 ( .IN0(n673), .IN1(n895), .SEL(n896), .F(n857) );
  IV U2042 ( .A(n897), .Z(n673) );
  MUX U2043 ( .IN0(e_input[22]), .IN1(n4911), .SEL(e_input[31]), .F(n1102) );
  MUX U2044 ( .IN0(e_input[23]), .IN1(n4910), .SEL(e_input[31]), .F(n674) );
  IV U2045 ( .A(n674), .Z(n1040) );
  MUX U2046 ( .IN0(e_input[19]), .IN1(n5077), .SEL(e_input[31]), .F(n1306) );
  MUX U2047 ( .IN0(e_input[18]), .IN1(n5076), .SEL(e_input[31]), .F(n1376) );
  MUX U2048 ( .IN0(e_input[13]), .IN1(n3889), .SEL(e_input[31]), .F(n1781) );
  MUX U2049 ( .IN0(n1902), .IN1(n1900), .SEL(n1901), .F(n1803) );
  XOR U2050 ( .A(n1859), .B(n1954), .Z(n1860) );
  MUX U2051 ( .IN0(n1952), .IN1(n1950), .SEL(n1951), .F(n1853) );
  MUX U2052 ( .IN0(e_input[11]), .IN1(n3859), .SEL(e_input[31]), .F(n1974) );
  MUX U2053 ( .IN0(e_input[10]), .IN1(n3858), .SEL(e_input[31]), .F(n2075) );
  MUX U2054 ( .IN0(e_input[6]), .IN1(n4345), .SEL(e_input[31]), .F(n2566) );
  MUX U2055 ( .IN0(n2584), .IN1(n2582), .SEL(n2583), .F(n2460) );
  XOR U2056 ( .A(n2516), .B(n2636), .Z(n2517) );
  MUX U2057 ( .IN0(n2634), .IN1(n2632), .SEL(n2633), .F(n2510) );
  MUX U2058 ( .IN0(e_input[5]), .IN1(n4341), .SEL(e_input[31]), .F(n2688) );
  MUX U2059 ( .IN0(n2821), .IN1(n675), .SEL(n2820), .F(n2690) );
  IV U2060 ( .A(n2819), .Z(n675) );
  MUX U2061 ( .IN0(e_input[3]), .IN1(n4705), .SEL(e_input[31]), .F(n2964) );
  XOR U2062 ( .A(n3033), .B(n3166), .Z(n3034) );
  MUX U2063 ( .IN0(n3164), .IN1(n3162), .SEL(n3163), .F(n3027) );
  MUX U2064 ( .IN0(n3114), .IN1(n3112), .SEL(n3113), .F(n2977) );
  MUX U2065 ( .IN0(e_input[2]), .IN1(n4704), .SEL(e_input[31]), .F(n3096) );
  XNOR U2066 ( .A(n4887), .B(n4886), .Z(n4734) );
  XNOR U2067 ( .A(n3213), .B(n3212), .Z(n3223) );
  XNOR U2068 ( .A(n4154), .B(n4153), .Z(n3790) );
  MUX U2069 ( .IN0(g_input[29]), .IN1(n4377), .SEL(g_input[31]), .F(n797) );
  OR U2070 ( .A(n906), .B(n907), .Z(n901) );
  XNOR U2071 ( .A(n908), .B(n869), .Z(n873) );
  XNOR U2072 ( .A(n1068), .B(n1013), .Z(n1017) );
  XOR U2073 ( .A(n1059), .B(n1004), .Z(n1008) );
  XOR U2074 ( .A(n1250), .B(n1185), .Z(n1189) );
  XNOR U2075 ( .A(n1259), .B(n1194), .Z(n1198) );
  XOR U2076 ( .A(n1378), .B(n1379), .Z(n1385) );
  XNOR U2077 ( .A(n1430), .B(n1358), .Z(n1364) );
  XNOR U2078 ( .A(n1482), .B(n1406), .Z(n1410) );
  XOR U2079 ( .A(n1473), .B(n1397), .Z(n1401) );
  MUX U2080 ( .IN0(e_input[14]), .IN1(n3893), .SEL(e_input[31]), .F(n1690) );
  XOR U2081 ( .A(n1449), .B(n1450), .Z(n1464) );
  XOR U2082 ( .A(n1741), .B(n1653), .Z(n1657) );
  XOR U2083 ( .A(n1724), .B(n1636), .Z(n1640) );
  XOR U2084 ( .A(n1874), .B(n1784), .Z(n1785) );
  MUX U2085 ( .IN0(n2078), .IN1(n676), .SEL(n2077), .F(n1971) );
  IV U2086 ( .A(n2076), .Z(n676) );
  XOR U2087 ( .A(n2040), .B(n1938), .Z(n1942) );
  XOR U2088 ( .A(n2023), .B(n1921), .Z(n1925) );
  XOR U2089 ( .A(n2357), .B(n2244), .Z(n2248) );
  XOR U2090 ( .A(n2374), .B(n2261), .Z(n2265) );
  XOR U2091 ( .A(n2414), .B(n2306), .Z(n2300) );
  MUX U2092 ( .IN0(e_input[7]), .IN1(n4346), .SEL(e_input[31]), .F(n2443) );
  XOR U2093 ( .A(n2568), .B(n2569), .Z(n2563) );
  XOR U2094 ( .A(n2745), .B(n2620), .Z(n2624) );
  XOR U2095 ( .A(n2728), .B(n2603), .Z(n2607) );
  XOR U2096 ( .A(n2786), .B(n2662), .Z(n2666) );
  XOR U2097 ( .A(n2696), .B(n2697), .Z(n2693) );
  XOR U2098 ( .A(n3147), .B(n3015), .Z(n3019) );
  XOR U2099 ( .A(n3130), .B(n2998), .Z(n3002) );
  NAND U2100 ( .A(n2961), .B(n3095), .Z(n3094) );
  XNOR U2101 ( .A(n3085), .B(n3084), .Z(n3102) );
  XNOR U2102 ( .A(n3778), .B(n3777), .Z(n3202) );
  MUX U2103 ( .IN0(g_input[30]), .IN1(n4359), .SEL(g_input[31]), .F(n765) );
  MUX U2104 ( .IN0(e_input[30]), .IN1(n5206), .SEL(e_input[31]), .F(n767) );
  XNOR U2105 ( .A(n916), .B(n915), .Z(n900) );
  XNOR U2106 ( .A(n985), .B(n984), .Z(n981) );
  XNOR U2107 ( .A(n1076), .B(n1075), .Z(n1058) );
  XNOR U2108 ( .A(n1039), .B(n1038), .Z(n1050) );
  XNOR U2109 ( .A(n1097), .B(n1096), .Z(n1110) );
  XNOR U2110 ( .A(n1163), .B(n1162), .Z(n1173) );
  XNOR U2111 ( .A(n1225), .B(n1224), .Z(n1239) );
  XNOR U2112 ( .A(n1267), .B(n1266), .Z(n1249) );
  XNOR U2113 ( .A(n1293), .B(n1292), .Z(n1311) );
  MUX U2114 ( .IN0(n677), .IN1(n1691), .SEL(n1692), .F(n1604) );
  IV U2115 ( .A(n1693), .Z(n677) );
  XNOR U2116 ( .A(n1438), .B(n1437), .Z(n1453) );
  XNOR U2117 ( .A(n1490), .B(n1489), .Z(n1472) );
  XNOR U2118 ( .A(n1524), .B(n1523), .Z(n1539) );
  MUX U2119 ( .IN0(e_input[15]), .IN1(n3894), .SEL(e_input[31]), .F(n1596) );
  XNOR U2120 ( .A(n1760), .B(n1759), .Z(n1740) );
  XNOR U2121 ( .A(n1708), .B(n1707), .Z(n1723) );
  XNOR U2122 ( .A(n1877), .B(n1876), .Z(n1873) );
  XNOR U2123 ( .A(n2007), .B(n2006), .Z(n2022) );
  XNOR U2124 ( .A(n2057), .B(n2056), .Z(n2039) );
  XNOR U2125 ( .A(n2093), .B(n2092), .Z(n2081) );
  XNOR U2126 ( .A(n2204), .B(n2203), .Z(n2186) );
  XNOR U2127 ( .A(n2316), .B(n2315), .Z(n2297) );
  XNOR U2128 ( .A(n2391), .B(n2390), .Z(n2373) );
  XNOR U2129 ( .A(n2341), .B(n2340), .Z(n2356) );
  XNOR U2130 ( .A(n2676), .B(n2675), .Z(n2658) );
  XNOR U2131 ( .A(n2712), .B(n2711), .Z(n2727) );
  XNOR U2132 ( .A(n2762), .B(n2761), .Z(n2744) );
  XNOR U2133 ( .A(n2815), .B(n2814), .Z(n2831) );
  XNOR U2134 ( .A(n2949), .B(n2948), .Z(n2969) );
  XNOR U2135 ( .A(n3050), .B(n3049), .Z(n3092) );
  MUX U2136 ( .IN0(n762), .IN1(n760), .SEL(n761), .F(n734) );
  XNOR U2137 ( .A(n733), .B(n732), .Z(n731) );
  XNOR U2138 ( .A(n827), .B(n826), .Z(n815) );
  XNOR U2139 ( .A(n942), .B(n941), .Z(n934) );
  XNOR U2140 ( .A(n1118), .B(n1117), .Z(n1108) );
  XNOR U2141 ( .A(n1319), .B(n1318), .Z(n1300) );
  XNOR U2142 ( .A(n1557), .B(n1556), .Z(n1531) );
  NANDN U2143 ( .B(n1591), .A(n1592), .Z(n1510) );
  NANDN U2144 ( .B(n1996), .A(n1997), .Z(n1891) );
  XNOR U2145 ( .A(n2413), .B(n2412), .Z(n2452) );
  XNOR U2146 ( .A(n2534), .B(n2533), .Z(n2574) );
  XNOR U2147 ( .A(n2785), .B(n2784), .Z(n2828) );
  XNOR U2148 ( .A(n2914), .B(n2913), .Z(n2956) );
  XNOR U2149 ( .A(n3121), .B(n3120), .Z(n3075) );
  MUX U2150 ( .IN0(n678), .IN1(n739), .SEL(n740), .F(n718) );
  IV U2151 ( .A(n741), .Z(n678) );
  XNOR U2152 ( .A(n1624), .B(n1623), .Z(n1607) );
  XNOR U2153 ( .A(n1812), .B(n1811), .Z(n1793) );
  XNOR U2154 ( .A(n1909), .B(n1908), .Z(n1890) );
  XNOR U2155 ( .A(n2119), .B(n2118), .Z(n2100) );
  XNOR U2156 ( .A(n2232), .B(n2231), .Z(n2211) );
  XNOR U2157 ( .A(n2469), .B(n2468), .Z(n2438) );
  XNOR U2158 ( .A(n2591), .B(n2590), .Z(n2559) );
  XNOR U2159 ( .A(n2848), .B(n2847), .Z(n2810) );
  XNOR U2160 ( .A(n2986), .B(n2985), .Z(n2939) );
  XNOR U2161 ( .A(n702), .B(n701), .Z(n725) );
  XNOR U2162 ( .A(n751), .B(n750), .Z(n776) );
  XNOR U2163 ( .A(n852), .B(n851), .Z(n885) );
  XNOR U2164 ( .A(n975), .B(n974), .Z(n1029) );
  XNOR U2165 ( .A(n1152), .B(n1151), .Z(n1210) );
  XOR U2166 ( .A(n1353), .B(n1352), .Z(n1423) );
  XOR U2167 ( .A(n804), .B(n808), .Z(n806) );
  XOR U2168 ( .A(n924), .B(n928), .Z(n926) );
  XOR U2169 ( .A(n1084), .B(n1088), .Z(n1086) );
  XOR U2170 ( .A(n1276), .B(n1280), .Z(n1278) );
  XOR U2171 ( .A(n1499), .B(n1503), .Z(n1501) );
  XOR U2172 ( .A(n1769), .B(n1773), .Z(n1771) );
  XOR U2173 ( .A(n2066), .B(n2069), .Z(n2067) );
  XOR U2174 ( .A(n2400), .B(n2403), .Z(n2401) );
  XOR U2175 ( .A(n2769), .B(n2772), .Z(n2770) );
  MUX U2176 ( .IN0(n686), .IN1(o[30]), .SEL(n687), .F(o[31]) );
  XOR U2177 ( .A(n679), .B(o_reg[10]), .Z(o[9]) );
  XOR U2178 ( .A(n680), .B(o_reg[9]), .Z(o[8]) );
  XOR U2179 ( .A(n681), .B(o_reg[8]), .Z(o[7]) );
  XOR U2180 ( .A(n682), .B(o_reg[7]), .Z(o[6]) );
  XOR U2181 ( .A(n683), .B(o_reg[6]), .Z(o[5]) );
  XOR U2182 ( .A(n684), .B(o_reg[5]), .Z(o[4]) );
  XNOR U2183 ( .A(n685), .B(o_reg[4]), .Z(o[3]) );
  XNOR U2184 ( .A(o_reg[31]), .B(n688), .Z(n687) );
  XNOR U2185 ( .A(n690), .B(o_reg[31]), .Z(o[30]) );
  XOR U2186 ( .A(n693), .B(n694), .Z(n688) );
  XOR U2187 ( .A(n695), .B(n696), .Z(n694) );
  AND U2188 ( .A(n697), .B(n698), .Z(n696) );
  XNOR U2189 ( .A(n703), .B(n701), .Z(n693) );
  XOR U2190 ( .A(n704), .B(n705), .Z(n703) );
  XOR U2191 ( .A(n706), .B(n707), .Z(n705) );
  XOR U2192 ( .A(n708), .B(n709), .Z(n707) );
  XOR U2193 ( .A(n714), .B(n715), .Z(n706) );
  XOR U2194 ( .A(n720), .B(n721), .Z(n704) );
  XNOR U2195 ( .A(n710), .B(n722), .Z(n721) );
  XOR U2196 ( .A(n718), .B(n716), .Z(n720) );
  XNOR U2197 ( .A(n723), .B(o_reg[3]), .Z(o[2]) );
  XNOR U2198 ( .A(o_reg[30]), .B(n692), .Z(o[29]) );
  XNOR U2199 ( .A(n724), .B(n725), .Z(n692) );
  AND U2200 ( .A(n697), .B(n727), .Z(n726) );
  XOR U2201 ( .A(n700), .B(n725), .Z(n727) );
  XNOR U2202 ( .A(n699), .B(n725), .Z(n700) );
  XOR U2203 ( .A(n713), .B(n722), .Z(n711) );
  IV U2204 ( .A(n712), .Z(n722) );
  XOR U2205 ( .A(n718), .B(n719), .Z(n717) );
  OR U2206 ( .A(n737), .B(n738), .Z(n719) );
  XNOR U2207 ( .A(o_reg[29]), .B(n745), .Z(o[28]) );
  XNOR U2208 ( .A(n746), .B(n747), .Z(n745) );
  AND U2209 ( .A(n697), .B(n749), .Z(n748) );
  XOR U2210 ( .A(n743), .B(n747), .Z(n749) );
  XNOR U2211 ( .A(n742), .B(n747), .Z(n743) );
  XOR U2212 ( .A(n754), .B(n755), .Z(n732) );
  ANDN U2213 ( .A(n756), .B(n754), .Z(n755) );
  XOR U2214 ( .A(n754), .B(n757), .Z(n756) );
  XOR U2215 ( .A(n758), .B(n759), .Z(n735) );
  IV U2216 ( .A(n734), .Z(n759) );
  XNOR U2217 ( .A(n740), .B(n741), .Z(n736) );
  NANDN U2218 ( .B(n737), .A(n765), .Z(n741) );
  XNOR U2219 ( .A(n739), .B(n766), .Z(n740) );
  ANDN U2220 ( .A(n767), .B(n738), .Z(n766) );
  XNOR U2221 ( .A(o_reg[28]), .B(n774), .Z(o[27]) );
  XNOR U2222 ( .A(n775), .B(n776), .Z(n774) );
  AND U2223 ( .A(n697), .B(n778), .Z(n777) );
  XOR U2224 ( .A(n772), .B(n776), .Z(n778) );
  XNOR U2225 ( .A(n771), .B(n776), .Z(n772) );
  XOR U2226 ( .A(n783), .B(n784), .Z(n754) );
  ANDN U2227 ( .A(n785), .B(n786), .Z(n784) );
  XOR U2228 ( .A(n783), .B(n787), .Z(n785) );
  XOR U2229 ( .A(n792), .B(n764), .Z(n788) );
  NANDN U2230 ( .B(n738), .A(n793), .Z(n764) );
  IV U2231 ( .A(n760), .Z(n792) );
  XNOR U2232 ( .A(n769), .B(n770), .Z(n762) );
  NANDN U2233 ( .B(n737), .A(n797), .Z(n770) );
  XNOR U2234 ( .A(n768), .B(n798), .Z(n769) );
  AND U2235 ( .A(n765), .B(n767), .Z(n798) );
  XNOR U2236 ( .A(o_reg[27]), .B(n805), .Z(o[26]) );
  XNOR U2237 ( .A(n806), .B(n807), .Z(n805) );
  AND U2238 ( .A(n697), .B(n809), .Z(n808) );
  XOR U2239 ( .A(n803), .B(n807), .Z(n809) );
  XNOR U2240 ( .A(n802), .B(n807), .Z(n803) );
  XOR U2241 ( .A(n812), .B(n813), .Z(n781) );
  ANDN U2242 ( .A(n814), .B(n812), .Z(n813) );
  XOR U2243 ( .A(n812), .B(n815), .Z(n814) );
  XNOR U2244 ( .A(n787), .B(n786), .Z(n782) );
  XOR U2245 ( .A(n816), .B(n817), .Z(n786) );
  XOR U2246 ( .A(n818), .B(n819), .Z(n817) );
  XOR U2247 ( .A(n820), .B(n821), .Z(n819) );
  XNOR U2248 ( .A(n789), .B(n829), .Z(n790) );
  ANDN U2249 ( .A(n830), .B(n738), .Z(n829) );
  XOR U2250 ( .A(n834), .B(n791), .Z(n828) );
  NAND U2251 ( .A(n793), .B(n765), .Z(n791) );
  IV U2252 ( .A(n794), .Z(n834) );
  XNOR U2253 ( .A(n800), .B(n801), .Z(n796) );
  NANDN U2254 ( .B(n737), .A(n838), .Z(n801) );
  XNOR U2255 ( .A(n799), .B(n839), .Z(n800) );
  AND U2256 ( .A(n797), .B(n767), .Z(n839) );
  XNOR U2257 ( .A(o_reg[26]), .B(n846), .Z(o[25]) );
  XNOR U2258 ( .A(n847), .B(n848), .Z(n846) );
  AND U2259 ( .A(n697), .B(n850), .Z(n849) );
  XOR U2260 ( .A(n844), .B(n848), .Z(n850) );
  XNOR U2261 ( .A(n843), .B(n848), .Z(n844) );
  XNOR U2262 ( .A(n855), .B(n822), .Z(n826) );
  XOR U2263 ( .A(n823), .B(n824), .Z(n822) );
  OR U2264 ( .A(n738), .B(n856), .Z(n824) );
  XNOR U2265 ( .A(n818), .B(n825), .Z(n855) );
  XNOR U2266 ( .A(n831), .B(n867), .Z(n832) );
  AND U2267 ( .A(n765), .B(n830), .Z(n867) );
  XOR U2268 ( .A(n871), .B(n833), .Z(n866) );
  NAND U2269 ( .A(n793), .B(n797), .Z(n833) );
  IV U2270 ( .A(n835), .Z(n871) );
  XNOR U2271 ( .A(n841), .B(n842), .Z(n837) );
  NANDN U2272 ( .B(n737), .A(n875), .Z(n842) );
  XNOR U2273 ( .A(n840), .B(n876), .Z(n841) );
  AND U2274 ( .A(n838), .B(n767), .Z(n876) );
  XNOR U2275 ( .A(o_reg[25]), .B(n883), .Z(o[24]) );
  XNOR U2276 ( .A(n884), .B(n885), .Z(n883) );
  AND U2277 ( .A(n697), .B(n887), .Z(n886) );
  XOR U2278 ( .A(n881), .B(n885), .Z(n887) );
  XNOR U2279 ( .A(n880), .B(n885), .Z(n881) );
  XNOR U2280 ( .A(n892), .B(n865), .Z(n861) );
  XNOR U2281 ( .A(n858), .B(n859), .Z(n865) );
  NANDN U2282 ( .B(n856), .A(n765), .Z(n859) );
  XNOR U2283 ( .A(n857), .B(n893), .Z(n858) );
  ANDN U2284 ( .A(n894), .B(n738), .Z(n893) );
  XNOR U2285 ( .A(n864), .B(n860), .Z(n892) );
  XNOR U2286 ( .A(n901), .B(n902), .Z(n864) );
  IV U2287 ( .A(n863), .Z(n902) );
  XNOR U2288 ( .A(n868), .B(n909), .Z(n869) );
  AND U2289 ( .A(n797), .B(n830), .Z(n909) );
  XOR U2290 ( .A(n913), .B(n870), .Z(n908) );
  NAND U2291 ( .A(n793), .B(n838), .Z(n870) );
  IV U2292 ( .A(n872), .Z(n913) );
  XNOR U2293 ( .A(n878), .B(n879), .Z(n874) );
  NANDN U2294 ( .B(n737), .A(n917), .Z(n879) );
  XNOR U2295 ( .A(n877), .B(n918), .Z(n878) );
  AND U2296 ( .A(n875), .B(n767), .Z(n918) );
  XNOR U2297 ( .A(o_reg[24]), .B(n925), .Z(o[23]) );
  XNOR U2298 ( .A(n926), .B(n927), .Z(n925) );
  AND U2299 ( .A(n697), .B(n929), .Z(n928) );
  XOR U2300 ( .A(n923), .B(n927), .Z(n929) );
  XNOR U2301 ( .A(n922), .B(n927), .Z(n923) );
  XNOR U2302 ( .A(n935), .B(n905), .Z(n899) );
  XNOR U2303 ( .A(n896), .B(n897), .Z(n905) );
  NANDN U2304 ( .B(n856), .A(n797), .Z(n897) );
  XNOR U2305 ( .A(n895), .B(n936), .Z(n896) );
  AND U2306 ( .A(n765), .B(n894), .Z(n936) );
  XNOR U2307 ( .A(n904), .B(n898), .Z(n935) );
  XOR U2308 ( .A(n947), .B(n907), .Z(n943) );
  NANDN U2309 ( .B(n738), .A(n948), .Z(n907) );
  IV U2310 ( .A(n903), .Z(n947) );
  XNOR U2311 ( .A(n910), .B(n953), .Z(n911) );
  AND U2312 ( .A(n838), .B(n830), .Z(n953) );
  XOR U2313 ( .A(n957), .B(n912), .Z(n952) );
  NAND U2314 ( .A(n793), .B(n875), .Z(n912) );
  IV U2315 ( .A(n914), .Z(n957) );
  XNOR U2316 ( .A(n920), .B(n921), .Z(n916) );
  NANDN U2317 ( .B(n737), .A(n961), .Z(n921) );
  XNOR U2318 ( .A(n919), .B(n962), .Z(n920) );
  AND U2319 ( .A(n917), .B(n767), .Z(n962) );
  XNOR U2320 ( .A(o_reg[23]), .B(n969), .Z(o[22]) );
  XNOR U2321 ( .A(n970), .B(n971), .Z(n969) );
  AND U2322 ( .A(n697), .B(n973), .Z(n972) );
  XOR U2323 ( .A(n967), .B(n971), .Z(n973) );
  XNOR U2324 ( .A(n966), .B(n971), .Z(n967) );
  XNOR U2325 ( .A(n934), .B(n933), .Z(n931) );
  XOR U2326 ( .A(n976), .B(n977), .Z(n933) );
  XOR U2327 ( .A(n978), .B(n979), .Z(n977) );
  XOR U2328 ( .A(n982), .B(n983), .Z(n978) );
  XOR U2329 ( .A(n988), .B(n932), .Z(n976) );
  XOR U2330 ( .A(n986), .B(n984), .Z(n988) );
  XNOR U2331 ( .A(n992), .B(n951), .Z(n941) );
  XNOR U2332 ( .A(n938), .B(n939), .Z(n951) );
  NANDN U2333 ( .B(n856), .A(n838), .Z(n939) );
  XNOR U2334 ( .A(n937), .B(n993), .Z(n938) );
  AND U2335 ( .A(n797), .B(n894), .Z(n993) );
  XNOR U2336 ( .A(n950), .B(n940), .Z(n992) );
  XNOR U2337 ( .A(n944), .B(n1001), .Z(n945) );
  ANDN U2338 ( .A(n1002), .B(n738), .Z(n1001) );
  XOR U2339 ( .A(n1006), .B(n946), .Z(n1000) );
  NAND U2340 ( .A(n948), .B(n765), .Z(n946) );
  IV U2341 ( .A(n949), .Z(n1006) );
  XNOR U2342 ( .A(n954), .B(n1011), .Z(n955) );
  AND U2343 ( .A(n875), .B(n830), .Z(n1011) );
  XOR U2344 ( .A(n1015), .B(n956), .Z(n1010) );
  NAND U2345 ( .A(n793), .B(n917), .Z(n956) );
  IV U2346 ( .A(n958), .Z(n1015) );
  XNOR U2347 ( .A(n964), .B(n965), .Z(n960) );
  NANDN U2348 ( .B(n737), .A(n1019), .Z(n965) );
  XNOR U2349 ( .A(n963), .B(n1020), .Z(n964) );
  AND U2350 ( .A(n961), .B(n767), .Z(n1020) );
  XNOR U2351 ( .A(o_reg[22]), .B(n1027), .Z(o[21]) );
  XNOR U2352 ( .A(n1028), .B(n1029), .Z(n1027) );
  AND U2353 ( .A(n697), .B(n1031), .Z(n1030) );
  XOR U2354 ( .A(n1025), .B(n1029), .Z(n1031) );
  XNOR U2355 ( .A(n1024), .B(n1029), .Z(n1025) );
  XNOR U2356 ( .A(n1034), .B(n981), .Z(n990) );
  XOR U2357 ( .A(n1035), .B(n1036), .Z(n984) );
  ANDN U2358 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR U2359 ( .A(n1035), .B(n1039), .Z(n1037) );
  XOR U2360 ( .A(n986), .B(n987), .Z(n985) );
  OR U2361 ( .A(n738), .B(n1040), .Z(n987) );
  XNOR U2362 ( .A(n980), .B(n989), .Z(n1034) );
  XOR U2363 ( .A(n1044), .B(n1045), .Z(n989) );
  ANDN U2364 ( .A(n1046), .B(n1047), .Z(n1045) );
  XNOR U2365 ( .A(n1044), .B(n1048), .Z(n1046) );
  XNOR U2366 ( .A(n1051), .B(n1009), .Z(n998) );
  XNOR U2367 ( .A(n995), .B(n996), .Z(n1009) );
  NANDN U2368 ( .B(n856), .A(n875), .Z(n996) );
  XNOR U2369 ( .A(n994), .B(n1052), .Z(n995) );
  AND U2370 ( .A(n838), .B(n894), .Z(n1052) );
  XNOR U2371 ( .A(n1008), .B(n997), .Z(n1051) );
  XNOR U2372 ( .A(n1003), .B(n1060), .Z(n1004) );
  AND U2373 ( .A(n765), .B(n1002), .Z(n1060) );
  XOR U2374 ( .A(n1064), .B(n1005), .Z(n1059) );
  NAND U2375 ( .A(n948), .B(n797), .Z(n1005) );
  IV U2376 ( .A(n1007), .Z(n1064) );
  XNOR U2377 ( .A(n1012), .B(n1069), .Z(n1013) );
  AND U2378 ( .A(n917), .B(n830), .Z(n1069) );
  XOR U2379 ( .A(n1073), .B(n1014), .Z(n1068) );
  NAND U2380 ( .A(n793), .B(n961), .Z(n1014) );
  IV U2381 ( .A(n1016), .Z(n1073) );
  XNOR U2382 ( .A(n1022), .B(n1023), .Z(n1018) );
  NANDN U2383 ( .B(n737), .A(n1077), .Z(n1023) );
  XNOR U2384 ( .A(n1021), .B(n1078), .Z(n1022) );
  AND U2385 ( .A(n1019), .B(n767), .Z(n1078) );
  XNOR U2386 ( .A(o_reg[21]), .B(n1085), .Z(o[20]) );
  XNOR U2387 ( .A(n1086), .B(n1087), .Z(n1085) );
  AND U2388 ( .A(n697), .B(n1089), .Z(n1088) );
  XOR U2389 ( .A(n1083), .B(n1087), .Z(n1089) );
  XNOR U2390 ( .A(n1082), .B(n1087), .Z(n1083) );
  XNOR U2391 ( .A(n1092), .B(n1050), .Z(n1047) );
  XOR U2392 ( .A(n1093), .B(n1094), .Z(n1038) );
  IV U2393 ( .A(n1035), .Z(n1094) );
  XNOR U2394 ( .A(n1042), .B(n1043), .Z(n1039) );
  NANDN U2395 ( .B(n1040), .A(n765), .Z(n1043) );
  XNOR U2396 ( .A(n1041), .B(n1101), .Z(n1042) );
  ANDN U2397 ( .A(n1102), .B(n738), .Z(n1101) );
  XNOR U2398 ( .A(n1111), .B(n1067), .Z(n1057) );
  XNOR U2399 ( .A(n1054), .B(n1055), .Z(n1067) );
  NANDN U2400 ( .B(n856), .A(n917), .Z(n1055) );
  XNOR U2401 ( .A(n1053), .B(n1112), .Z(n1054) );
  AND U2402 ( .A(n875), .B(n894), .Z(n1112) );
  XNOR U2403 ( .A(n1066), .B(n1056), .Z(n1111) );
  XNOR U2404 ( .A(n1061), .B(n1120), .Z(n1062) );
  AND U2405 ( .A(n797), .B(n1002), .Z(n1120) );
  XOR U2406 ( .A(n1124), .B(n1063), .Z(n1119) );
  NAND U2407 ( .A(n948), .B(n838), .Z(n1063) );
  IV U2408 ( .A(n1065), .Z(n1124) );
  XNOR U2409 ( .A(n1070), .B(n1129), .Z(n1071) );
  AND U2410 ( .A(n961), .B(n830), .Z(n1129) );
  XOR U2411 ( .A(n1133), .B(n1072), .Z(n1128) );
  NAND U2412 ( .A(n793), .B(n1019), .Z(n1072) );
  IV U2413 ( .A(n1074), .Z(n1133) );
  XNOR U2414 ( .A(n1080), .B(n1081), .Z(n1076) );
  NANDN U2415 ( .B(n737), .A(n1137), .Z(n1081) );
  XNOR U2416 ( .A(n1079), .B(n1138), .Z(n1080) );
  AND U2417 ( .A(n1077), .B(n767), .Z(n1138) );
  XNOR U2418 ( .A(n1146), .B(o_reg[2]), .Z(o[1]) );
  XNOR U2419 ( .A(o_reg[20]), .B(n1145), .Z(o[19]) );
  XNOR U2420 ( .A(n1147), .B(n1148), .Z(n1145) );
  AND U2421 ( .A(n697), .B(n1150), .Z(n1149) );
  XOR U2422 ( .A(n1143), .B(n1148), .Z(n1150) );
  XNOR U2423 ( .A(n1142), .B(n1148), .Z(n1143) );
  XNOR U2424 ( .A(n1153), .B(n1110), .Z(n1107) );
  XOR U2425 ( .A(n1154), .B(n1098), .Z(n1096) );
  IV U2426 ( .A(n1099), .Z(n1098) );
  NANDN U2427 ( .B(n738), .A(n1158), .Z(n1100) );
  XOR U2428 ( .A(n1159), .B(n1160), .Z(n1095) );
  ANDN U2429 ( .A(n1161), .B(n1162), .Z(n1160) );
  XOR U2430 ( .A(n1159), .B(n1163), .Z(n1161) );
  XNOR U2431 ( .A(n1104), .B(n1105), .Z(n1097) );
  NANDN U2432 ( .B(n1040), .A(n797), .Z(n1105) );
  XNOR U2433 ( .A(n1103), .B(n1164), .Z(n1104) );
  AND U2434 ( .A(n765), .B(n1102), .Z(n1164) );
  XNOR U2435 ( .A(n1174), .B(n1127), .Z(n1117) );
  XNOR U2436 ( .A(n1114), .B(n1115), .Z(n1127) );
  NANDN U2437 ( .B(n856), .A(n961), .Z(n1115) );
  XNOR U2438 ( .A(n1113), .B(n1175), .Z(n1114) );
  AND U2439 ( .A(n917), .B(n894), .Z(n1175) );
  XNOR U2440 ( .A(n1126), .B(n1116), .Z(n1174) );
  XNOR U2441 ( .A(n1121), .B(n1183), .Z(n1122) );
  AND U2442 ( .A(n838), .B(n1002), .Z(n1183) );
  XOR U2443 ( .A(n1187), .B(n1123), .Z(n1182) );
  NAND U2444 ( .A(n948), .B(n875), .Z(n1123) );
  IV U2445 ( .A(n1125), .Z(n1187) );
  XNOR U2446 ( .A(n1130), .B(n1192), .Z(n1131) );
  AND U2447 ( .A(n1019), .B(n830), .Z(n1192) );
  XOR U2448 ( .A(n1196), .B(n1132), .Z(n1191) );
  NAND U2449 ( .A(n793), .B(n1077), .Z(n1132) );
  IV U2450 ( .A(n1134), .Z(n1196) );
  XNOR U2451 ( .A(n1140), .B(n1141), .Z(n1136) );
  NANDN U2452 ( .B(n737), .A(n1200), .Z(n1141) );
  XNOR U2453 ( .A(n1139), .B(n1201), .Z(n1140) );
  AND U2454 ( .A(n1137), .B(n767), .Z(n1201) );
  XNOR U2455 ( .A(o_reg[19]), .B(n1208), .Z(o[18]) );
  XNOR U2456 ( .A(n1209), .B(n1210), .Z(n1208) );
  AND U2457 ( .A(n697), .B(n1212), .Z(n1211) );
  XOR U2458 ( .A(n1206), .B(n1210), .Z(n1212) );
  XNOR U2459 ( .A(n1205), .B(n1210), .Z(n1206) );
  XNOR U2460 ( .A(n1215), .B(n1173), .Z(n1169) );
  XNOR U2461 ( .A(n1155), .B(n1217), .Z(n1156) );
  ANDN U2462 ( .A(n1218), .B(n738), .Z(n1217) );
  XOR U2463 ( .A(n1222), .B(n1157), .Z(n1216) );
  NAND U2464 ( .A(n1158), .B(n765), .Z(n1157) );
  IV U2465 ( .A(n1159), .Z(n1222) );
  XNOR U2466 ( .A(n1166), .B(n1167), .Z(n1163) );
  NANDN U2467 ( .B(n1040), .A(n838), .Z(n1167) );
  XNOR U2468 ( .A(n1165), .B(n1226), .Z(n1166) );
  AND U2469 ( .A(n797), .B(n1102), .Z(n1226) );
  XNOR U2470 ( .A(n1172), .B(n1168), .Z(n1215) );
  XNOR U2471 ( .A(n1233), .B(n1234), .Z(n1172) );
  IV U2472 ( .A(n1171), .Z(n1234) );
  XOR U2473 ( .A(n1235), .B(n1236), .Z(n1171) );
  ANDN U2474 ( .A(n1237), .B(n1238), .Z(n1236) );
  XOR U2475 ( .A(n1235), .B(n1239), .Z(n1237) );
  XNOR U2476 ( .A(n1242), .B(n1190), .Z(n1180) );
  XNOR U2477 ( .A(n1177), .B(n1178), .Z(n1190) );
  NANDN U2478 ( .B(n856), .A(n1019), .Z(n1178) );
  XNOR U2479 ( .A(n1176), .B(n1243), .Z(n1177) );
  AND U2480 ( .A(n961), .B(n894), .Z(n1243) );
  XNOR U2481 ( .A(n1189), .B(n1179), .Z(n1242) );
  XNOR U2482 ( .A(n1184), .B(n1251), .Z(n1185) );
  AND U2483 ( .A(n875), .B(n1002), .Z(n1251) );
  XOR U2484 ( .A(n1255), .B(n1186), .Z(n1250) );
  NAND U2485 ( .A(n948), .B(n917), .Z(n1186) );
  IV U2486 ( .A(n1188), .Z(n1255) );
  XNOR U2487 ( .A(n1193), .B(n1260), .Z(n1194) );
  AND U2488 ( .A(n1077), .B(n830), .Z(n1260) );
  XOR U2489 ( .A(n1264), .B(n1195), .Z(n1259) );
  NAND U2490 ( .A(n793), .B(n1137), .Z(n1195) );
  IV U2491 ( .A(n1197), .Z(n1264) );
  XNOR U2492 ( .A(n1203), .B(n1204), .Z(n1199) );
  NANDN U2493 ( .B(n737), .A(n1268), .Z(n1204) );
  XNOR U2494 ( .A(n1202), .B(n1269), .Z(n1203) );
  AND U2495 ( .A(n1200), .B(n767), .Z(n1269) );
  ANDN U2496 ( .A(n1270), .B(n1271), .Z(n1202) );
  NANDN U2497 ( .B(n1272), .A(n1273), .Z(n1270) );
  XOR U2498 ( .A(n1277), .B(o_reg[18]), .Z(o[17]) );
  XNOR U2499 ( .A(n1278), .B(n1279), .Z(n1277) );
  AND U2500 ( .A(n697), .B(n1281), .Z(n1280) );
  XOR U2501 ( .A(n1275), .B(n1279), .Z(n1281) );
  XNOR U2502 ( .A(n1274), .B(n1279), .Z(n1275) );
  XNOR U2503 ( .A(n1232), .B(n1231), .Z(n1214) );
  XOR U2504 ( .A(n1284), .B(n1239), .Z(n1231) );
  XNOR U2505 ( .A(n1219), .B(n1286), .Z(n1220) );
  AND U2506 ( .A(n765), .B(n1218), .Z(n1286) );
  XOR U2507 ( .A(n1290), .B(n1221), .Z(n1285) );
  NAND U2508 ( .A(n1158), .B(n797), .Z(n1221) );
  IV U2509 ( .A(n1223), .Z(n1290) );
  XNOR U2510 ( .A(n1228), .B(n1229), .Z(n1225) );
  NANDN U2511 ( .B(n1040), .A(n875), .Z(n1229) );
  XNOR U2512 ( .A(n1227), .B(n1294), .Z(n1228) );
  AND U2513 ( .A(n838), .B(n1102), .Z(n1294) );
  XNOR U2514 ( .A(n1238), .B(n1230), .Z(n1284) );
  XOR U2515 ( .A(n1301), .B(n1240), .Z(n1238) );
  NAND U2516 ( .A(n1304), .B(n1305), .Z(n1241) );
  NANDN U2517 ( .B(n738), .A(n1306), .Z(n1305) );
  OR U2518 ( .A(n1307), .B(n1308), .Z(n1304) );
  XNOR U2519 ( .A(n1312), .B(n1258), .Z(n1248) );
  XNOR U2520 ( .A(n1245), .B(n1246), .Z(n1258) );
  NANDN U2521 ( .B(n856), .A(n1077), .Z(n1246) );
  XNOR U2522 ( .A(n1244), .B(n1313), .Z(n1245) );
  AND U2523 ( .A(n1019), .B(n894), .Z(n1313) );
  XNOR U2524 ( .A(n1257), .B(n1247), .Z(n1312) );
  XNOR U2525 ( .A(n1252), .B(n1321), .Z(n1253) );
  AND U2526 ( .A(n917), .B(n1002), .Z(n1321) );
  XOR U2527 ( .A(n1325), .B(n1254), .Z(n1320) );
  NAND U2528 ( .A(n948), .B(n961), .Z(n1254) );
  IV U2529 ( .A(n1256), .Z(n1325) );
  XNOR U2530 ( .A(n1261), .B(n1330), .Z(n1262) );
  AND U2531 ( .A(n1137), .B(n830), .Z(n1330) );
  XOR U2532 ( .A(n1334), .B(n1263), .Z(n1329) );
  NAND U2533 ( .A(n793), .B(n1200), .Z(n1263) );
  IV U2534 ( .A(n1265), .Z(n1334) );
  XNOR U2535 ( .A(n1272), .B(n1273), .Z(n1267) );
  NANDN U2536 ( .B(n737), .A(n1338), .Z(n1273) );
  XOR U2537 ( .A(n1271), .B(n1339), .Z(n1272) );
  AND U2538 ( .A(n1268), .B(n767), .Z(n1339) );
  NAND U2539 ( .A(n1340), .B(n1341), .Z(n1271) );
  NANDN U2540 ( .B(n1342), .A(n1343), .Z(n1340) );
  XOR U2541 ( .A(n1347), .B(o_reg[17]), .Z(o[16]) );
  XNOR U2542 ( .A(n1348), .B(n1349), .Z(n1347) );
  AND U2543 ( .A(n697), .B(n1351), .Z(n1350) );
  XOR U2544 ( .A(n1345), .B(n1349), .Z(n1351) );
  XNOR U2545 ( .A(n1344), .B(n1349), .Z(n1345) );
  XNOR U2546 ( .A(n1300), .B(n1299), .Z(n1283) );
  XOR U2547 ( .A(n1354), .B(n1311), .Z(n1299) );
  XNOR U2548 ( .A(n1287), .B(n1356), .Z(n1288) );
  AND U2549 ( .A(n797), .B(n1218), .Z(n1356) );
  XOR U2550 ( .A(n1360), .B(n1289), .Z(n1355) );
  NAND U2551 ( .A(n1158), .B(n838), .Z(n1289) );
  IV U2552 ( .A(n1291), .Z(n1360) );
  XOR U2553 ( .A(n1361), .B(n1362), .Z(n1291) );
  ANDN U2554 ( .A(n1363), .B(n1364), .Z(n1362) );
  XOR U2555 ( .A(n1361), .B(n1365), .Z(n1363) );
  XNOR U2556 ( .A(n1296), .B(n1297), .Z(n1293) );
  NANDN U2557 ( .B(n1040), .A(n917), .Z(n1297) );
  XNOR U2558 ( .A(n1295), .B(n1366), .Z(n1296) );
  AND U2559 ( .A(n875), .B(n1102), .Z(n1366) );
  XNOR U2560 ( .A(n1310), .B(n1298), .Z(n1354) );
  XNOR U2561 ( .A(n1373), .B(n1303), .Z(n1310) );
  XOR U2562 ( .A(n1374), .B(n1307), .Z(n1303) );
  NAND U2563 ( .A(n1306), .B(n765), .Z(n1307) );
  NANDN U2564 ( .B(n738), .A(n1376), .Z(n1375) );
  XNOR U2565 ( .A(n1386), .B(n1328), .Z(n1318) );
  XNOR U2566 ( .A(n1315), .B(n1316), .Z(n1328) );
  NANDN U2567 ( .B(n856), .A(n1137), .Z(n1316) );
  XNOR U2568 ( .A(n1314), .B(n1387), .Z(n1315) );
  AND U2569 ( .A(n1077), .B(n894), .Z(n1387) );
  XNOR U2570 ( .A(n1327), .B(n1317), .Z(n1386) );
  XNOR U2571 ( .A(n1322), .B(n1395), .Z(n1323) );
  AND U2572 ( .A(n961), .B(n1002), .Z(n1395) );
  XOR U2573 ( .A(n1399), .B(n1324), .Z(n1394) );
  NAND U2574 ( .A(n948), .B(n1019), .Z(n1324) );
  IV U2575 ( .A(n1326), .Z(n1399) );
  XNOR U2576 ( .A(n1331), .B(n1404), .Z(n1332) );
  AND U2577 ( .A(n1200), .B(n830), .Z(n1404) );
  XOR U2578 ( .A(n1408), .B(n1333), .Z(n1403) );
  NAND U2579 ( .A(n793), .B(n1268), .Z(n1333) );
  IV U2580 ( .A(n1335), .Z(n1408) );
  XNOR U2581 ( .A(n1342), .B(n1343), .Z(n1337) );
  NANDN U2582 ( .B(n737), .A(n1412), .Z(n1343) );
  XNOR U2583 ( .A(n1341), .B(n1413), .Z(n1342) );
  AND U2584 ( .A(n1338), .B(n767), .Z(n1413) );
  AND U2585 ( .A(n1414), .B(n1415), .Z(n1341) );
  NANDN U2586 ( .B(n1416), .A(n1417), .Z(n1414) );
  XOR U2587 ( .A(n1421), .B(o_reg[16]), .Z(o[15]) );
  XNOR U2588 ( .A(n1422), .B(n1423), .Z(n1421) );
  AND U2589 ( .A(n697), .B(n1425), .Z(n1424) );
  XOR U2590 ( .A(n1419), .B(n1423), .Z(n1425) );
  XNOR U2591 ( .A(n1418), .B(n1423), .Z(n1419) );
  XNOR U2592 ( .A(n1372), .B(n1371), .Z(n1353) );
  XOR U2593 ( .A(n1429), .B(n1382), .Z(n1371) );
  XNOR U2594 ( .A(n1357), .B(n1431), .Z(n1358) );
  AND U2595 ( .A(n838), .B(n1218), .Z(n1431) );
  XOR U2596 ( .A(n1435), .B(n1359), .Z(n1430) );
  NAND U2597 ( .A(n1158), .B(n875), .Z(n1359) );
  IV U2598 ( .A(n1361), .Z(n1435) );
  XNOR U2599 ( .A(n1368), .B(n1369), .Z(n1365) );
  NANDN U2600 ( .B(n1040), .A(n961), .Z(n1369) );
  XNOR U2601 ( .A(n1367), .B(n1439), .Z(n1368) );
  AND U2602 ( .A(n917), .B(n1102), .Z(n1439) );
  XNOR U2603 ( .A(n1381), .B(n1370), .Z(n1429) );
  XNOR U2604 ( .A(n1446), .B(n1385), .Z(n1381) );
  NAND U2605 ( .A(n1306), .B(n797), .Z(n1379) );
  XNOR U2606 ( .A(n1377), .B(n1447), .Z(n1378) );
  AND U2607 ( .A(n765), .B(n1376), .Z(n1447) );
  XNOR U2608 ( .A(n1384), .B(n1380), .Z(n1446) );
  AND U2609 ( .A(n1455), .B(n1456), .Z(n1454) );
  NANDN U2610 ( .B(n738), .A(n1457), .Z(n1456) );
  OR U2611 ( .A(n1458), .B(n1459), .Z(n1455) );
  XNOR U2612 ( .A(n1460), .B(n1461), .Z(n1383) );
  ANDN U2613 ( .A(n1462), .B(n1463), .Z(n1461) );
  XOR U2614 ( .A(n1460), .B(n1464), .Z(n1462) );
  XNOR U2615 ( .A(n1465), .B(n1402), .Z(n1392) );
  XNOR U2616 ( .A(n1389), .B(n1390), .Z(n1402) );
  NANDN U2617 ( .B(n856), .A(n1200), .Z(n1390) );
  XNOR U2618 ( .A(n1388), .B(n1466), .Z(n1389) );
  AND U2619 ( .A(n1137), .B(n894), .Z(n1466) );
  XNOR U2620 ( .A(n1401), .B(n1391), .Z(n1465) );
  XNOR U2621 ( .A(n1396), .B(n1474), .Z(n1397) );
  AND U2622 ( .A(n1019), .B(n1002), .Z(n1474) );
  XOR U2623 ( .A(n1478), .B(n1398), .Z(n1473) );
  NAND U2624 ( .A(n948), .B(n1077), .Z(n1398) );
  IV U2625 ( .A(n1400), .Z(n1478) );
  XNOR U2626 ( .A(n1405), .B(n1483), .Z(n1406) );
  AND U2627 ( .A(n1268), .B(n830), .Z(n1483) );
  XOR U2628 ( .A(n1487), .B(n1407), .Z(n1482) );
  NAND U2629 ( .A(n793), .B(n1338), .Z(n1407) );
  IV U2630 ( .A(n1409), .Z(n1487) );
  XNOR U2631 ( .A(n1416), .B(n1417), .Z(n1411) );
  NANDN U2632 ( .B(n737), .A(n1491), .Z(n1417) );
  XNOR U2633 ( .A(n1415), .B(n1492), .Z(n1416) );
  AND U2634 ( .A(n1412), .B(n767), .Z(n1492) );
  ANDN U2635 ( .A(n1493), .B(n1494), .Z(n1415) );
  NANDN U2636 ( .B(n1495), .A(n1496), .Z(n1493) );
  XOR U2637 ( .A(n1500), .B(o_reg[15]), .Z(o[14]) );
  XNOR U2638 ( .A(n1501), .B(n1502), .Z(n1500) );
  AND U2639 ( .A(n697), .B(n1504), .Z(n1503) );
  XOR U2640 ( .A(n1498), .B(n1502), .Z(n1504) );
  XNOR U2641 ( .A(n1497), .B(n1502), .Z(n1498) );
  XOR U2642 ( .A(n1428), .B(n1427), .Z(n1502) );
  XOR U2643 ( .A(n1505), .B(n1506), .Z(n1427) );
  XOR U2644 ( .A(n1507), .B(n1508), .Z(n1506) );
  XOR U2645 ( .A(n1509), .B(n1507), .Z(n1508) );
  XNOR U2646 ( .A(n1445), .B(n1444), .Z(n1428) );
  XOR U2647 ( .A(n1515), .B(n1453), .Z(n1444) );
  XNOR U2648 ( .A(n1432), .B(n1517), .Z(n1433) );
  AND U2649 ( .A(n875), .B(n1218), .Z(n1517) );
  XOR U2650 ( .A(n1521), .B(n1434), .Z(n1516) );
  NAND U2651 ( .A(n1158), .B(n917), .Z(n1434) );
  IV U2652 ( .A(n1436), .Z(n1521) );
  XNOR U2653 ( .A(n1441), .B(n1442), .Z(n1438) );
  NANDN U2654 ( .B(n1040), .A(n1019), .Z(n1442) );
  XNOR U2655 ( .A(n1440), .B(n1525), .Z(n1441) );
  AND U2656 ( .A(n961), .B(n1102), .Z(n1525) );
  XNOR U2657 ( .A(n1452), .B(n1443), .Z(n1515) );
  XNOR U2658 ( .A(n1532), .B(n1464), .Z(n1452) );
  NAND U2659 ( .A(n1306), .B(n838), .Z(n1450) );
  XNOR U2660 ( .A(n1448), .B(n1533), .Z(n1449) );
  AND U2661 ( .A(n797), .B(n1376), .Z(n1533) );
  XNOR U2662 ( .A(n1463), .B(n1451), .Z(n1532) );
  XNOR U2663 ( .A(n1540), .B(n1460), .Z(n1463) );
  XNOR U2664 ( .A(n1544), .B(n1458), .Z(n1540) );
  NAND U2665 ( .A(n1457), .B(n765), .Z(n1458) );
  NANDN U2666 ( .B(n738), .A(n1546), .Z(n1545) );
  XNOR U2667 ( .A(n1550), .B(n1481), .Z(n1471) );
  XNOR U2668 ( .A(n1468), .B(n1469), .Z(n1481) );
  NANDN U2669 ( .B(n856), .A(n1268), .Z(n1469) );
  XNOR U2670 ( .A(n1467), .B(n1551), .Z(n1468) );
  AND U2671 ( .A(n1200), .B(n894), .Z(n1551) );
  XNOR U2672 ( .A(n1480), .B(n1470), .Z(n1550) );
  XNOR U2673 ( .A(n1475), .B(n1559), .Z(n1476) );
  AND U2674 ( .A(n1077), .B(n1002), .Z(n1559) );
  XOR U2675 ( .A(n1563), .B(n1477), .Z(n1558) );
  NAND U2676 ( .A(n948), .B(n1137), .Z(n1477) );
  IV U2677 ( .A(n1479), .Z(n1563) );
  XNOR U2678 ( .A(n1484), .B(n1568), .Z(n1485) );
  AND U2679 ( .A(n1338), .B(n830), .Z(n1568) );
  XOR U2680 ( .A(n1572), .B(n1486), .Z(n1567) );
  NAND U2681 ( .A(n793), .B(n1412), .Z(n1486) );
  IV U2682 ( .A(n1488), .Z(n1572) );
  XNOR U2683 ( .A(n1495), .B(n1496), .Z(n1490) );
  NANDN U2684 ( .B(n737), .A(n1576), .Z(n1496) );
  AND U2685 ( .A(n1491), .B(n767), .Z(n1577) );
  NAND U2686 ( .A(n1578), .B(n1579), .Z(n1494) );
  NANDN U2687 ( .B(n1580), .A(n1581), .Z(n1578) );
  XOR U2688 ( .A(n1585), .B(o_reg[14]), .Z(o[13]) );
  XNOR U2689 ( .A(n1586), .B(n1587), .Z(n1585) );
  AND U2690 ( .A(n697), .B(n1589), .Z(n1588) );
  XOR U2691 ( .A(n1583), .B(n1587), .Z(n1589) );
  XNOR U2692 ( .A(n1582), .B(n1587), .Z(n1583) );
  XNOR U2693 ( .A(n1514), .B(n1513), .Z(n1587) );
  XNOR U2694 ( .A(n1590), .B(n1510), .Z(n1513) );
  NAND U2695 ( .A(n1507), .B(n1593), .Z(n1511) );
  AND U2696 ( .A(n1594), .B(n1595), .Z(n1593) );
  NANDN U2697 ( .B(n738), .A(n1596), .Z(n1595) );
  NANDN U2698 ( .B(n1597), .A(n1598), .Z(n1594) );
  AND U2699 ( .A(n1599), .B(n1600), .Z(n1507) );
  NANDN U2700 ( .B(n1601), .A(n1602), .Z(n1600) );
  NANDN U2701 ( .B(n1603), .A(n1604), .Z(n1599) );
  XNOR U2702 ( .A(n1608), .B(n1539), .Z(n1530) );
  XNOR U2703 ( .A(n1518), .B(n1610), .Z(n1519) );
  AND U2704 ( .A(n917), .B(n1218), .Z(n1610) );
  XOR U2705 ( .A(n1614), .B(n1520), .Z(n1609) );
  NAND U2706 ( .A(n1158), .B(n961), .Z(n1520) );
  IV U2707 ( .A(n1522), .Z(n1614) );
  XNOR U2708 ( .A(n1527), .B(n1528), .Z(n1524) );
  NANDN U2709 ( .B(n1040), .A(n1077), .Z(n1528) );
  XNOR U2710 ( .A(n1526), .B(n1618), .Z(n1527) );
  AND U2711 ( .A(n1019), .B(n1102), .Z(n1618) );
  XNOR U2712 ( .A(n1538), .B(n1529), .Z(n1608) );
  XOR U2713 ( .A(n1625), .B(n1543), .Z(n1538) );
  XNOR U2714 ( .A(n1535), .B(n1536), .Z(n1543) );
  NAND U2715 ( .A(n1306), .B(n875), .Z(n1536) );
  XNOR U2716 ( .A(n1534), .B(n1626), .Z(n1535) );
  AND U2717 ( .A(n838), .B(n1376), .Z(n1626) );
  XNOR U2718 ( .A(n1542), .B(n1537), .Z(n1625) );
  XNOR U2719 ( .A(n1547), .B(n1634), .Z(n1548) );
  AND U2720 ( .A(n765), .B(n1546), .Z(n1634) );
  XOR U2721 ( .A(n1638), .B(n1549), .Z(n1633) );
  NAND U2722 ( .A(n1457), .B(n797), .Z(n1549) );
  IV U2723 ( .A(n1541), .Z(n1638) );
  XNOR U2724 ( .A(n1642), .B(n1566), .Z(n1556) );
  XNOR U2725 ( .A(n1553), .B(n1554), .Z(n1566) );
  NANDN U2726 ( .B(n856), .A(n1338), .Z(n1554) );
  XNOR U2727 ( .A(n1552), .B(n1643), .Z(n1553) );
  AND U2728 ( .A(n1268), .B(n894), .Z(n1643) );
  XNOR U2729 ( .A(n1565), .B(n1555), .Z(n1642) );
  XNOR U2730 ( .A(n1560), .B(n1651), .Z(n1561) );
  AND U2731 ( .A(n1137), .B(n1002), .Z(n1651) );
  XOR U2732 ( .A(n1655), .B(n1562), .Z(n1650) );
  NAND U2733 ( .A(n948), .B(n1200), .Z(n1562) );
  IV U2734 ( .A(n1564), .Z(n1655) );
  XNOR U2735 ( .A(n1569), .B(n1660), .Z(n1570) );
  AND U2736 ( .A(n1412), .B(n830), .Z(n1660) );
  XOR U2737 ( .A(n1664), .B(n1571), .Z(n1659) );
  NAND U2738 ( .A(n793), .B(n1491), .Z(n1571) );
  IV U2739 ( .A(n1573), .Z(n1664) );
  XNOR U2740 ( .A(n1580), .B(n1581), .Z(n1575) );
  NANDN U2741 ( .B(n737), .A(n1668), .Z(n1581) );
  XNOR U2742 ( .A(n1579), .B(n1669), .Z(n1580) );
  AND U2743 ( .A(n1576), .B(n767), .Z(n1669) );
  ANDN U2744 ( .A(n1670), .B(n1671), .Z(n1579) );
  NANDN U2745 ( .B(n1672), .A(n1673), .Z(n1670) );
  XOR U2746 ( .A(n1677), .B(o_reg[13]), .Z(o[12]) );
  XNOR U2747 ( .A(n1678), .B(n1679), .Z(n1677) );
  AND U2748 ( .A(n697), .B(n1681), .Z(n1680) );
  XOR U2749 ( .A(n1675), .B(n1679), .Z(n1681) );
  XNOR U2750 ( .A(n1674), .B(n1679), .Z(n1675) );
  XNOR U2751 ( .A(n1607), .B(n1606), .Z(n1679) );
  XNOR U2752 ( .A(n1682), .B(n1592), .Z(n1606) );
  XNOR U2753 ( .A(n1598), .B(n1597), .Z(n1592) );
  OR U2754 ( .A(n1683), .B(n1684), .Z(n1597) );
  XNOR U2755 ( .A(n1601), .B(n1602), .Z(n1598) );
  XOR U2756 ( .A(n1688), .B(n1603), .Z(n1601) );
  NAND U2757 ( .A(n765), .B(n1596), .Z(n1603) );
  NANDN U2758 ( .B(n1604), .A(n1689), .Z(n1688) );
  NANDN U2759 ( .B(n738), .A(n1690), .Z(n1689) );
  XNOR U2760 ( .A(n1699), .B(n1632), .Z(n1623) );
  XNOR U2761 ( .A(n1611), .B(n1701), .Z(n1612) );
  AND U2762 ( .A(n961), .B(n1218), .Z(n1701) );
  XOR U2763 ( .A(n1705), .B(n1613), .Z(n1700) );
  NAND U2764 ( .A(n1158), .B(n1019), .Z(n1613) );
  IV U2765 ( .A(n1615), .Z(n1705) );
  XNOR U2766 ( .A(n1620), .B(n1621), .Z(n1617) );
  NANDN U2767 ( .B(n1040), .A(n1137), .Z(n1621) );
  XNOR U2768 ( .A(n1619), .B(n1709), .Z(n1620) );
  AND U2769 ( .A(n1077), .B(n1102), .Z(n1709) );
  XNOR U2770 ( .A(n1631), .B(n1622), .Z(n1699) );
  XOR U2771 ( .A(n1716), .B(n1641), .Z(n1631) );
  XNOR U2772 ( .A(n1628), .B(n1629), .Z(n1641) );
  NAND U2773 ( .A(n1306), .B(n917), .Z(n1629) );
  XNOR U2774 ( .A(n1627), .B(n1717), .Z(n1628) );
  AND U2775 ( .A(n875), .B(n1376), .Z(n1717) );
  XNOR U2776 ( .A(n1640), .B(n1630), .Z(n1716) );
  XNOR U2777 ( .A(n1635), .B(n1725), .Z(n1636) );
  AND U2778 ( .A(n797), .B(n1546), .Z(n1725) );
  XOR U2779 ( .A(n1729), .B(n1637), .Z(n1724) );
  NAND U2780 ( .A(n1457), .B(n838), .Z(n1637) );
  IV U2781 ( .A(n1639), .Z(n1729) );
  XNOR U2782 ( .A(n1733), .B(n1658), .Z(n1648) );
  XNOR U2783 ( .A(n1645), .B(n1646), .Z(n1658) );
  NANDN U2784 ( .B(n856), .A(n1412), .Z(n1646) );
  XNOR U2785 ( .A(n1644), .B(n1734), .Z(n1645) );
  AND U2786 ( .A(n1338), .B(n894), .Z(n1734) );
  XNOR U2787 ( .A(n1657), .B(n1647), .Z(n1733) );
  XNOR U2788 ( .A(n1652), .B(n1742), .Z(n1653) );
  AND U2789 ( .A(n1200), .B(n1002), .Z(n1742) );
  XOR U2790 ( .A(n1746), .B(n1654), .Z(n1741) );
  NAND U2791 ( .A(n948), .B(n1268), .Z(n1654) );
  IV U2792 ( .A(n1656), .Z(n1746) );
  XNOR U2793 ( .A(n1661), .B(n1751), .Z(n1662) );
  AND U2794 ( .A(n1491), .B(n830), .Z(n1751) );
  XOR U2795 ( .A(n1755), .B(n1663), .Z(n1750) );
  NAND U2796 ( .A(n793), .B(n1576), .Z(n1663) );
  IV U2797 ( .A(n1665), .Z(n1755) );
  XOR U2798 ( .A(n1756), .B(n1757), .Z(n1665) );
  ANDN U2799 ( .A(n1758), .B(n1759), .Z(n1757) );
  XOR U2800 ( .A(n1756), .B(n1760), .Z(n1758) );
  XNOR U2801 ( .A(n1672), .B(n1673), .Z(n1667) );
  NANDN U2802 ( .B(n737), .A(n1761), .Z(n1673) );
  AND U2803 ( .A(n1668), .B(n767), .Z(n1762) );
  NAND U2804 ( .A(n1763), .B(n1764), .Z(n1671) );
  NANDN U2805 ( .B(n1765), .A(n1766), .Z(n1763) );
  XOR U2806 ( .A(n1770), .B(o_reg[12]), .Z(o[11]) );
  XNOR U2807 ( .A(n1771), .B(n1772), .Z(n1770) );
  AND U2808 ( .A(n697), .B(n1774), .Z(n1773) );
  XOR U2809 ( .A(n1768), .B(n1772), .Z(n1774) );
  XNOR U2810 ( .A(n1767), .B(n1772), .Z(n1768) );
  XNOR U2811 ( .A(n1696), .B(n1695), .Z(n1772) );
  XNOR U2812 ( .A(n1775), .B(n1698), .Z(n1695) );
  XOR U2813 ( .A(n1684), .B(n1683), .Z(n1698) );
  NANDN U2814 ( .B(n1776), .A(n1777), .Z(n1683) );
  XOR U2815 ( .A(n1687), .B(n1686), .Z(n1684) );
  XOR U2816 ( .A(n1685), .B(n1778), .Z(n1686) );
  AND U2817 ( .A(n1779), .B(n1780), .Z(n1778) );
  NANDN U2818 ( .B(n738), .A(n1781), .Z(n1780) );
  OR U2819 ( .A(n1782), .B(n1783), .Z(n1779) );
  NAND U2820 ( .A(n797), .B(n1596), .Z(n1693) );
  XNOR U2821 ( .A(n1691), .B(n1787), .Z(n1692) );
  AND U2822 ( .A(n1690), .B(n765), .Z(n1787) );
  XNOR U2823 ( .A(n1796), .B(n1723), .Z(n1714) );
  XNOR U2824 ( .A(n1702), .B(n1798), .Z(n1703) );
  AND U2825 ( .A(n1019), .B(n1218), .Z(n1798) );
  XOR U2826 ( .A(n1802), .B(n1704), .Z(n1797) );
  NAND U2827 ( .A(n1158), .B(n1077), .Z(n1704) );
  IV U2828 ( .A(n1706), .Z(n1802) );
  XNOR U2829 ( .A(n1711), .B(n1712), .Z(n1708) );
  NANDN U2830 ( .B(n1040), .A(n1200), .Z(n1712) );
  XNOR U2831 ( .A(n1710), .B(n1806), .Z(n1711) );
  AND U2832 ( .A(n1137), .B(n1102), .Z(n1806) );
  XNOR U2833 ( .A(n1722), .B(n1713), .Z(n1796) );
  XOR U2834 ( .A(n1813), .B(n1732), .Z(n1722) );
  XNOR U2835 ( .A(n1719), .B(n1720), .Z(n1732) );
  NAND U2836 ( .A(n1306), .B(n961), .Z(n1720) );
  XNOR U2837 ( .A(n1718), .B(n1814), .Z(n1719) );
  AND U2838 ( .A(n917), .B(n1376), .Z(n1814) );
  XNOR U2839 ( .A(n1731), .B(n1721), .Z(n1813) );
  XNOR U2840 ( .A(n1726), .B(n1822), .Z(n1727) );
  AND U2841 ( .A(n838), .B(n1546), .Z(n1822) );
  XOR U2842 ( .A(n1826), .B(n1728), .Z(n1821) );
  NAND U2843 ( .A(n1457), .B(n875), .Z(n1728) );
  IV U2844 ( .A(n1730), .Z(n1826) );
  XNOR U2845 ( .A(n1830), .B(n1749), .Z(n1739) );
  XNOR U2846 ( .A(n1736), .B(n1737), .Z(n1749) );
  NANDN U2847 ( .B(n856), .A(n1491), .Z(n1737) );
  XNOR U2848 ( .A(n1735), .B(n1831), .Z(n1736) );
  AND U2849 ( .A(n1412), .B(n894), .Z(n1831) );
  XNOR U2850 ( .A(n1748), .B(n1738), .Z(n1830) );
  XNOR U2851 ( .A(n1743), .B(n1839), .Z(n1744) );
  AND U2852 ( .A(n1268), .B(n1002), .Z(n1839) );
  XOR U2853 ( .A(n1843), .B(n1745), .Z(n1838) );
  NAND U2854 ( .A(n948), .B(n1338), .Z(n1745) );
  IV U2855 ( .A(n1747), .Z(n1843) );
  XNOR U2856 ( .A(n1752), .B(n1848), .Z(n1753) );
  AND U2857 ( .A(n1576), .B(n830), .Z(n1848) );
  XOR U2858 ( .A(n1852), .B(n1754), .Z(n1847) );
  NAND U2859 ( .A(n793), .B(n1668), .Z(n1754) );
  IV U2860 ( .A(n1756), .Z(n1852) );
  XNOR U2861 ( .A(n1765), .B(n1766), .Z(n1760) );
  NANDN U2862 ( .B(n737), .A(n1856), .Z(n1766) );
  XNOR U2863 ( .A(n1764), .B(n1857), .Z(n1765) );
  AND U2864 ( .A(n1761), .B(n767), .Z(n1857) );
  ANDN U2865 ( .A(n1858), .B(n1859), .Z(n1764) );
  NANDN U2866 ( .B(n1860), .A(n1861), .Z(n1858) );
  XOR U2867 ( .A(n1865), .B(o_reg[11]), .Z(o[10]) );
  XNOR U2868 ( .A(n1866), .B(n1867), .Z(n1865) );
  AND U2869 ( .A(n697), .B(n1869), .Z(n1868) );
  XOR U2870 ( .A(n1863), .B(n1867), .Z(n1869) );
  XNOR U2871 ( .A(n1862), .B(n1867), .Z(n1863) );
  XNOR U2872 ( .A(n1793), .B(n1792), .Z(n1867) );
  XNOR U2873 ( .A(n1870), .B(n1795), .Z(n1792) );
  XNOR U2874 ( .A(n1776), .B(n1777), .Z(n1795) );
  XOR U2875 ( .A(n1786), .B(n1785), .Z(n1776) );
  XNOR U2876 ( .A(n1878), .B(n1782), .Z(n1874) );
  NAND U2877 ( .A(n765), .B(n1781), .Z(n1782) );
  NANDN U2878 ( .B(n738), .A(n1880), .Z(n1879) );
  NAND U2879 ( .A(n838), .B(n1596), .Z(n1790) );
  XNOR U2880 ( .A(n1788), .B(n1884), .Z(n1789) );
  AND U2881 ( .A(n1690), .B(n797), .Z(n1884) );
  XNOR U2882 ( .A(n1893), .B(n1820), .Z(n1811) );
  XNOR U2883 ( .A(n1799), .B(n1895), .Z(n1800) );
  AND U2884 ( .A(n1077), .B(n1218), .Z(n1895) );
  XOR U2885 ( .A(n1899), .B(n1801), .Z(n1894) );
  NAND U2886 ( .A(n1158), .B(n1137), .Z(n1801) );
  IV U2887 ( .A(n1803), .Z(n1899) );
  XNOR U2888 ( .A(n1808), .B(n1809), .Z(n1805) );
  NANDN U2889 ( .B(n1040), .A(n1268), .Z(n1809) );
  XNOR U2890 ( .A(n1807), .B(n1903), .Z(n1808) );
  AND U2891 ( .A(n1200), .B(n1102), .Z(n1903) );
  XNOR U2892 ( .A(n1819), .B(n1810), .Z(n1893) );
  XOR U2893 ( .A(n1910), .B(n1829), .Z(n1819) );
  XNOR U2894 ( .A(n1816), .B(n1817), .Z(n1829) );
  NAND U2895 ( .A(n1306), .B(n1019), .Z(n1817) );
  XNOR U2896 ( .A(n1815), .B(n1911), .Z(n1816) );
  AND U2897 ( .A(n961), .B(n1376), .Z(n1911) );
  XNOR U2898 ( .A(n1828), .B(n1818), .Z(n1910) );
  XNOR U2899 ( .A(n1823), .B(n1919), .Z(n1824) );
  AND U2900 ( .A(n875), .B(n1546), .Z(n1919) );
  XOR U2901 ( .A(n1923), .B(n1825), .Z(n1918) );
  NAND U2902 ( .A(n1457), .B(n917), .Z(n1825) );
  IV U2903 ( .A(n1827), .Z(n1923) );
  XNOR U2904 ( .A(n1927), .B(n1846), .Z(n1836) );
  XNOR U2905 ( .A(n1833), .B(n1834), .Z(n1846) );
  NANDN U2906 ( .B(n856), .A(n1576), .Z(n1834) );
  XNOR U2907 ( .A(n1832), .B(n1928), .Z(n1833) );
  AND U2908 ( .A(n1491), .B(n894), .Z(n1928) );
  XNOR U2909 ( .A(n1845), .B(n1835), .Z(n1927) );
  XNOR U2910 ( .A(n1840), .B(n1936), .Z(n1841) );
  AND U2911 ( .A(n1338), .B(n1002), .Z(n1936) );
  XOR U2912 ( .A(n1940), .B(n1842), .Z(n1935) );
  NAND U2913 ( .A(n948), .B(n1412), .Z(n1842) );
  IV U2914 ( .A(n1844), .Z(n1940) );
  XNOR U2915 ( .A(n1849), .B(n1945), .Z(n1850) );
  AND U2916 ( .A(n1668), .B(n830), .Z(n1945) );
  XOR U2917 ( .A(n1949), .B(n1851), .Z(n1944) );
  NAND U2918 ( .A(n793), .B(n1761), .Z(n1851) );
  IV U2919 ( .A(n1853), .Z(n1949) );
  XNOR U2920 ( .A(n1860), .B(n1861), .Z(n1855) );
  NANDN U2921 ( .B(n737), .A(n1953), .Z(n1861) );
  AND U2922 ( .A(n1856), .B(n767), .Z(n1954) );
  NAND U2923 ( .A(n1955), .B(n1956), .Z(n1859) );
  NANDN U2924 ( .B(n1957), .A(n1958), .Z(n1955) );
  XNOR U2925 ( .A(n1962), .B(n1963), .Z(n679) );
  AND U2926 ( .A(n697), .B(n1965), .Z(n1964) );
  XOR U2927 ( .A(n1960), .B(n1963), .Z(n1965) );
  XNOR U2928 ( .A(n1959), .B(n1963), .Z(n1960) );
  XNOR U2929 ( .A(n1890), .B(n1889), .Z(n1963) );
  XNOR U2930 ( .A(n1966), .B(n1892), .Z(n1889) );
  XNOR U2931 ( .A(n1873), .B(n1872), .Z(n1892) );
  XNOR U2932 ( .A(n1871), .B(n1967), .Z(n1872) );
  AND U2933 ( .A(n1968), .B(n1969), .Z(n1967) );
  OR U2934 ( .A(n1970), .B(n1971), .Z(n1969) );
  AND U2935 ( .A(n1972), .B(n1973), .Z(n1968) );
  NANDN U2936 ( .B(n738), .A(n1974), .Z(n1973) );
  NAND U2937 ( .A(n1975), .B(n1976), .Z(n1972) );
  XNOR U2938 ( .A(n1881), .B(n1981), .Z(n1882) );
  AND U2939 ( .A(n1880), .B(n765), .Z(n1981) );
  XOR U2940 ( .A(n1985), .B(n1883), .Z(n1980) );
  NAND U2941 ( .A(n797), .B(n1781), .Z(n1883) );
  IV U2942 ( .A(n1875), .Z(n1985) );
  XNOR U2943 ( .A(n1886), .B(n1887), .Z(n1877) );
  NAND U2944 ( .A(n875), .B(n1596), .Z(n1887) );
  XNOR U2945 ( .A(n1885), .B(n1989), .Z(n1886) );
  AND U2946 ( .A(n1690), .B(n838), .Z(n1989) );
  XNOR U2947 ( .A(n1998), .B(n1917), .Z(n1908) );
  XNOR U2948 ( .A(n1896), .B(n2000), .Z(n1897) );
  AND U2949 ( .A(n1137), .B(n1218), .Z(n2000) );
  XOR U2950 ( .A(n2004), .B(n1898), .Z(n1999) );
  NAND U2951 ( .A(n1158), .B(n1200), .Z(n1898) );
  IV U2952 ( .A(n1900), .Z(n2004) );
  XNOR U2953 ( .A(n1905), .B(n1906), .Z(n1902) );
  NANDN U2954 ( .B(n1040), .A(n1338), .Z(n1906) );
  XNOR U2955 ( .A(n1904), .B(n2008), .Z(n1905) );
  AND U2956 ( .A(n1268), .B(n1102), .Z(n2008) );
  XNOR U2957 ( .A(n1916), .B(n1907), .Z(n1998) );
  XOR U2958 ( .A(n2015), .B(n1926), .Z(n1916) );
  XNOR U2959 ( .A(n1913), .B(n1914), .Z(n1926) );
  NAND U2960 ( .A(n1306), .B(n1077), .Z(n1914) );
  XNOR U2961 ( .A(n1912), .B(n2016), .Z(n1913) );
  AND U2962 ( .A(n1019), .B(n1376), .Z(n2016) );
  XNOR U2963 ( .A(n1925), .B(n1915), .Z(n2015) );
  XNOR U2964 ( .A(n1920), .B(n2024), .Z(n1921) );
  AND U2965 ( .A(n917), .B(n1546), .Z(n2024) );
  XOR U2966 ( .A(n2028), .B(n1922), .Z(n2023) );
  NAND U2967 ( .A(n1457), .B(n961), .Z(n1922) );
  IV U2968 ( .A(n1924), .Z(n2028) );
  XNOR U2969 ( .A(n2032), .B(n1943), .Z(n1933) );
  XNOR U2970 ( .A(n1930), .B(n1931), .Z(n1943) );
  NANDN U2971 ( .B(n856), .A(n1668), .Z(n1931) );
  XNOR U2972 ( .A(n1929), .B(n2033), .Z(n1930) );
  AND U2973 ( .A(n1576), .B(n894), .Z(n2033) );
  XNOR U2974 ( .A(n1942), .B(n1932), .Z(n2032) );
  XNOR U2975 ( .A(n1937), .B(n2041), .Z(n1938) );
  AND U2976 ( .A(n1412), .B(n1002), .Z(n2041) );
  XOR U2977 ( .A(n2045), .B(n1939), .Z(n2040) );
  NAND U2978 ( .A(n948), .B(n1491), .Z(n1939) );
  IV U2979 ( .A(n1941), .Z(n2045) );
  XNOR U2980 ( .A(n1946), .B(n2050), .Z(n1947) );
  AND U2981 ( .A(n1761), .B(n830), .Z(n2050) );
  XOR U2982 ( .A(n2054), .B(n1948), .Z(n2049) );
  NAND U2983 ( .A(n793), .B(n1856), .Z(n1948) );
  IV U2984 ( .A(n1950), .Z(n2054) );
  XNOR U2985 ( .A(n1957), .B(n1958), .Z(n1952) );
  NANDN U2986 ( .B(n737), .A(n2058), .Z(n1958) );
  XNOR U2987 ( .A(n1956), .B(n2059), .Z(n1957) );
  AND U2988 ( .A(n1953), .B(n767), .Z(n2059) );
  ANDN U2989 ( .A(n2060), .B(n2061), .Z(n1956) );
  NANDN U2990 ( .B(n2062), .A(n2063), .Z(n2060) );
  XNOR U2991 ( .A(n2067), .B(n2068), .Z(n680) );
  AND U2992 ( .A(n697), .B(n2070), .Z(n2069) );
  XOR U2993 ( .A(n2065), .B(n2068), .Z(n2070) );
  XNOR U2994 ( .A(n2064), .B(n2068), .Z(n2065) );
  XNOR U2995 ( .A(n1995), .B(n1994), .Z(n2068) );
  XNOR U2996 ( .A(n2071), .B(n1997), .Z(n1994) );
  XNOR U2997 ( .A(n1979), .B(n1978), .Z(n1997) );
  XNOR U2998 ( .A(n2072), .B(n1975), .Z(n1978) );
  XNOR U2999 ( .A(n2073), .B(n1970), .Z(n1975) );
  NAND U3000 ( .A(n765), .B(n1974), .Z(n1970) );
  NANDN U3001 ( .B(n738), .A(n2075), .Z(n2074) );
  XNOR U3002 ( .A(n1976), .B(n1977), .Z(n2072) );
  XNOR U3003 ( .A(n1982), .B(n2086), .Z(n1983) );
  AND U3004 ( .A(n1880), .B(n797), .Z(n2086) );
  XOR U3005 ( .A(n2090), .B(n1984), .Z(n2085) );
  NAND U3006 ( .A(n838), .B(n1781), .Z(n1984) );
  IV U3007 ( .A(n1986), .Z(n2090) );
  XNOR U3008 ( .A(n1991), .B(n1992), .Z(n1988) );
  NAND U3009 ( .A(n917), .B(n1596), .Z(n1992) );
  XNOR U3010 ( .A(n1990), .B(n2094), .Z(n1991) );
  AND U3011 ( .A(n1690), .B(n875), .Z(n2094) );
  XNOR U3012 ( .A(n2103), .B(n2022), .Z(n2013) );
  XNOR U3013 ( .A(n2001), .B(n2105), .Z(n2002) );
  AND U3014 ( .A(n1200), .B(n1218), .Z(n2105) );
  XOR U3015 ( .A(n2109), .B(n2003), .Z(n2104) );
  NAND U3016 ( .A(n1158), .B(n1268), .Z(n2003) );
  IV U3017 ( .A(n2005), .Z(n2109) );
  XNOR U3018 ( .A(n2010), .B(n2011), .Z(n2007) );
  NANDN U3019 ( .B(n1040), .A(n1412), .Z(n2011) );
  XNOR U3020 ( .A(n2009), .B(n2113), .Z(n2010) );
  AND U3021 ( .A(n1338), .B(n1102), .Z(n2113) );
  XNOR U3022 ( .A(n2021), .B(n2012), .Z(n2103) );
  XOR U3023 ( .A(n2120), .B(n2031), .Z(n2021) );
  XNOR U3024 ( .A(n2018), .B(n2019), .Z(n2031) );
  NAND U3025 ( .A(n1306), .B(n1137), .Z(n2019) );
  XNOR U3026 ( .A(n2017), .B(n2121), .Z(n2018) );
  AND U3027 ( .A(n1077), .B(n1376), .Z(n2121) );
  XNOR U3028 ( .A(n2030), .B(n2020), .Z(n2120) );
  XNOR U3029 ( .A(n2025), .B(n2129), .Z(n2026) );
  AND U3030 ( .A(n961), .B(n1546), .Z(n2129) );
  XOR U3031 ( .A(n2133), .B(n2027), .Z(n2128) );
  NAND U3032 ( .A(n1457), .B(n1019), .Z(n2027) );
  IV U3033 ( .A(n2029), .Z(n2133) );
  XNOR U3034 ( .A(n2137), .B(n2048), .Z(n2038) );
  XNOR U3035 ( .A(n2035), .B(n2036), .Z(n2048) );
  NANDN U3036 ( .B(n856), .A(n1761), .Z(n2036) );
  XNOR U3037 ( .A(n2034), .B(n2138), .Z(n2035) );
  AND U3038 ( .A(n1668), .B(n894), .Z(n2138) );
  XNOR U3039 ( .A(n2047), .B(n2037), .Z(n2137) );
  XNOR U3040 ( .A(n2042), .B(n2146), .Z(n2043) );
  AND U3041 ( .A(n1491), .B(n1002), .Z(n2146) );
  XOR U3042 ( .A(n2150), .B(n2044), .Z(n2145) );
  NAND U3043 ( .A(n948), .B(n1576), .Z(n2044) );
  IV U3044 ( .A(n2046), .Z(n2150) );
  XNOR U3045 ( .A(n2051), .B(n2155), .Z(n2052) );
  AND U3046 ( .A(n1856), .B(n830), .Z(n2155) );
  XOR U3047 ( .A(n2159), .B(n2053), .Z(n2154) );
  NAND U3048 ( .A(n793), .B(n1953), .Z(n2053) );
  IV U3049 ( .A(n2055), .Z(n2159) );
  XOR U3050 ( .A(n2160), .B(n2161), .Z(n2055) );
  ANDN U3051 ( .A(n2162), .B(n2163), .Z(n2161) );
  XOR U3052 ( .A(n2160), .B(n2164), .Z(n2162) );
  XNOR U3053 ( .A(n2062), .B(n2063), .Z(n2057) );
  NANDN U3054 ( .B(n737), .A(n2165), .Z(n2063) );
  AND U3055 ( .A(n2058), .B(n767), .Z(n2166) );
  NAND U3056 ( .A(n2167), .B(n2168), .Z(n2061) );
  NANDN U3057 ( .B(n2169), .A(n2170), .Z(n2167) );
  XNOR U3058 ( .A(n2174), .B(n2175), .Z(n681) );
  AND U3059 ( .A(n697), .B(n2177), .Z(n2176) );
  XOR U3060 ( .A(n2172), .B(n2175), .Z(n2177) );
  XNOR U3061 ( .A(n2171), .B(n2175), .Z(n2172) );
  XNOR U3062 ( .A(n2100), .B(n2099), .Z(n2175) );
  XNOR U3063 ( .A(n2178), .B(n2102), .Z(n2099) );
  XNOR U3064 ( .A(n2081), .B(n2080), .Z(n2102) );
  XNOR U3065 ( .A(n2179), .B(n2084), .Z(n2080) );
  XNOR U3066 ( .A(n2077), .B(n2078), .Z(n2084) );
  NAND U3067 ( .A(n797), .B(n1974), .Z(n2078) );
  XNOR U3068 ( .A(n2076), .B(n2180), .Z(n2077) );
  AND U3069 ( .A(n2075), .B(n765), .Z(n2180) );
  XNOR U3070 ( .A(n2083), .B(n2079), .Z(n2179) );
  AND U3071 ( .A(n2188), .B(n2189), .Z(n2187) );
  NANDN U3072 ( .B(n738), .A(n2190), .Z(n2189) );
  OR U3073 ( .A(n2191), .B(n2192), .Z(n2188) );
  XNOR U3074 ( .A(n2087), .B(n2197), .Z(n2088) );
  AND U3075 ( .A(n1880), .B(n838), .Z(n2197) );
  XOR U3076 ( .A(n2201), .B(n2089), .Z(n2196) );
  NAND U3077 ( .A(n875), .B(n1781), .Z(n2089) );
  IV U3078 ( .A(n2091), .Z(n2201) );
  XNOR U3079 ( .A(n2096), .B(n2097), .Z(n2093) );
  NAND U3080 ( .A(n961), .B(n1596), .Z(n2097) );
  XNOR U3081 ( .A(n2095), .B(n2205), .Z(n2096) );
  AND U3082 ( .A(n1690), .B(n917), .Z(n2205) );
  XNOR U3083 ( .A(n2215), .B(n2212), .Z(n2214) );
  XNOR U3084 ( .A(n2216), .B(n2127), .Z(n2118) );
  XNOR U3085 ( .A(n2106), .B(n2218), .Z(n2107) );
  AND U3086 ( .A(n1268), .B(n1218), .Z(n2218) );
  XOR U3087 ( .A(n2222), .B(n2108), .Z(n2217) );
  NAND U3088 ( .A(n1158), .B(n1338), .Z(n2108) );
  IV U3089 ( .A(n2110), .Z(n2222) );
  XNOR U3090 ( .A(n2115), .B(n2116), .Z(n2112) );
  NANDN U3091 ( .B(n1040), .A(n1491), .Z(n2116) );
  XNOR U3092 ( .A(n2114), .B(n2226), .Z(n2115) );
  AND U3093 ( .A(n1412), .B(n1102), .Z(n2226) );
  XNOR U3094 ( .A(n2126), .B(n2117), .Z(n2216) );
  XOR U3095 ( .A(n2233), .B(n2136), .Z(n2126) );
  XNOR U3096 ( .A(n2123), .B(n2124), .Z(n2136) );
  NAND U3097 ( .A(n1306), .B(n1200), .Z(n2124) );
  XNOR U3098 ( .A(n2122), .B(n2234), .Z(n2123) );
  AND U3099 ( .A(n1137), .B(n1376), .Z(n2234) );
  XNOR U3100 ( .A(n2135), .B(n2125), .Z(n2233) );
  XNOR U3101 ( .A(n2130), .B(n2242), .Z(n2131) );
  AND U3102 ( .A(n1019), .B(n1546), .Z(n2242) );
  XOR U3103 ( .A(n2246), .B(n2132), .Z(n2241) );
  NAND U3104 ( .A(n1457), .B(n1077), .Z(n2132) );
  IV U3105 ( .A(n2134), .Z(n2246) );
  XNOR U3106 ( .A(n2250), .B(n2153), .Z(n2143) );
  XNOR U3107 ( .A(n2140), .B(n2141), .Z(n2153) );
  NANDN U3108 ( .B(n856), .A(n1856), .Z(n2141) );
  XNOR U3109 ( .A(n2139), .B(n2251), .Z(n2140) );
  AND U3110 ( .A(n1761), .B(n894), .Z(n2251) );
  XNOR U3111 ( .A(n2152), .B(n2142), .Z(n2250) );
  XNOR U3112 ( .A(n2147), .B(n2259), .Z(n2148) );
  AND U3113 ( .A(n1576), .B(n1002), .Z(n2259) );
  XOR U3114 ( .A(n2263), .B(n2149), .Z(n2258) );
  NAND U3115 ( .A(n948), .B(n1668), .Z(n2149) );
  IV U3116 ( .A(n2151), .Z(n2263) );
  XNOR U3117 ( .A(n2156), .B(n2268), .Z(n2157) );
  AND U3118 ( .A(n1953), .B(n830), .Z(n2268) );
  XOR U3119 ( .A(n2272), .B(n2158), .Z(n2267) );
  NAND U3120 ( .A(n793), .B(n2058), .Z(n2158) );
  IV U3121 ( .A(n2160), .Z(n2272) );
  XNOR U3122 ( .A(n2169), .B(n2170), .Z(n2164) );
  NANDN U3123 ( .B(n737), .A(n2276), .Z(n2170) );
  XNOR U3124 ( .A(n2168), .B(n2277), .Z(n2169) );
  AND U3125 ( .A(n2165), .B(n767), .Z(n2277) );
  ANDN U3126 ( .A(n2278), .B(n2279), .Z(n2168) );
  NANDN U3127 ( .B(n2280), .A(n2281), .Z(n2278) );
  XNOR U3128 ( .A(n2285), .B(n2286), .Z(n682) );
  AND U3129 ( .A(n697), .B(n2288), .Z(n2287) );
  XOR U3130 ( .A(n2283), .B(n2286), .Z(n2288) );
  XNOR U3131 ( .A(n2282), .B(n2286), .Z(n2283) );
  XNOR U3132 ( .A(n2211), .B(n2210), .Z(n2286) );
  XNOR U3133 ( .A(n2289), .B(n2215), .Z(n2210) );
  XNOR U3134 ( .A(n2186), .B(n2185), .Z(n2215) );
  XNOR U3135 ( .A(n2290), .B(n2195), .Z(n2185) );
  XNOR U3136 ( .A(n2182), .B(n2183), .Z(n2195) );
  NAND U3137 ( .A(n838), .B(n1974), .Z(n2183) );
  XNOR U3138 ( .A(n2181), .B(n2291), .Z(n2182) );
  AND U3139 ( .A(n2075), .B(n797), .Z(n2291) );
  XNOR U3140 ( .A(n2194), .B(n2184), .Z(n2290) );
  XNOR U3141 ( .A(n2298), .B(n2193), .Z(n2194) );
  XNOR U3142 ( .A(n2302), .B(n2191), .Z(n2298) );
  NAND U3143 ( .A(n765), .B(n2190), .Z(n2191) );
  NANDN U3144 ( .B(n738), .A(n2304), .Z(n2303) );
  XNOR U3145 ( .A(n2198), .B(n2309), .Z(n2199) );
  AND U3146 ( .A(n1880), .B(n875), .Z(n2309) );
  XOR U3147 ( .A(n2313), .B(n2200), .Z(n2308) );
  NAND U3148 ( .A(n917), .B(n1781), .Z(n2200) );
  IV U3149 ( .A(n2202), .Z(n2313) );
  XNOR U3150 ( .A(n2207), .B(n2208), .Z(n2204) );
  NAND U3151 ( .A(n1019), .B(n1596), .Z(n2208) );
  XNOR U3152 ( .A(n2206), .B(n2317), .Z(n2207) );
  AND U3153 ( .A(n1690), .B(n961), .Z(n2317) );
  XNOR U3154 ( .A(n2213), .B(n2209), .Z(n2289) );
  XOR U3155 ( .A(n2328), .B(n2329), .Z(n2324) );
  NANDN U3156 ( .B(n2330), .A(n2331), .Z(n2328) );
  XNOR U3157 ( .A(n2332), .B(n2240), .Z(n2231) );
  XNOR U3158 ( .A(n2219), .B(n2334), .Z(n2220) );
  AND U3159 ( .A(n1338), .B(n1218), .Z(n2334) );
  XOR U3160 ( .A(n2338), .B(n2221), .Z(n2333) );
  NAND U3161 ( .A(n1158), .B(n1412), .Z(n2221) );
  IV U3162 ( .A(n2223), .Z(n2338) );
  XNOR U3163 ( .A(n2228), .B(n2229), .Z(n2225) );
  NANDN U3164 ( .B(n1040), .A(n1576), .Z(n2229) );
  XNOR U3165 ( .A(n2227), .B(n2342), .Z(n2228) );
  AND U3166 ( .A(n1491), .B(n1102), .Z(n2342) );
  XNOR U3167 ( .A(n2239), .B(n2230), .Z(n2332) );
  XOR U3168 ( .A(n2349), .B(n2249), .Z(n2239) );
  XNOR U3169 ( .A(n2236), .B(n2237), .Z(n2249) );
  NAND U3170 ( .A(n1306), .B(n1268), .Z(n2237) );
  XNOR U3171 ( .A(n2235), .B(n2350), .Z(n2236) );
  AND U3172 ( .A(n1200), .B(n1376), .Z(n2350) );
  XNOR U3173 ( .A(n2248), .B(n2238), .Z(n2349) );
  XNOR U3174 ( .A(n2243), .B(n2358), .Z(n2244) );
  AND U3175 ( .A(n1077), .B(n1546), .Z(n2358) );
  XOR U3176 ( .A(n2362), .B(n2245), .Z(n2357) );
  NAND U3177 ( .A(n1457), .B(n1137), .Z(n2245) );
  IV U3178 ( .A(n2247), .Z(n2362) );
  XNOR U3179 ( .A(n2366), .B(n2266), .Z(n2256) );
  XNOR U3180 ( .A(n2253), .B(n2254), .Z(n2266) );
  NANDN U3181 ( .B(n856), .A(n1953), .Z(n2254) );
  XNOR U3182 ( .A(n2252), .B(n2367), .Z(n2253) );
  AND U3183 ( .A(n1856), .B(n894), .Z(n2367) );
  XNOR U3184 ( .A(n2265), .B(n2255), .Z(n2366) );
  XNOR U3185 ( .A(n2260), .B(n2375), .Z(n2261) );
  AND U3186 ( .A(n1668), .B(n1002), .Z(n2375) );
  XOR U3187 ( .A(n2379), .B(n2262), .Z(n2374) );
  NAND U3188 ( .A(n948), .B(n1761), .Z(n2262) );
  IV U3189 ( .A(n2264), .Z(n2379) );
  XNOR U3190 ( .A(n2269), .B(n2384), .Z(n2270) );
  AND U3191 ( .A(n2058), .B(n830), .Z(n2384) );
  XOR U3192 ( .A(n2388), .B(n2271), .Z(n2383) );
  NAND U3193 ( .A(n793), .B(n2165), .Z(n2271) );
  IV U3194 ( .A(n2273), .Z(n2388) );
  XNOR U3195 ( .A(n2280), .B(n2281), .Z(n2275) );
  NANDN U3196 ( .B(n737), .A(n2392), .Z(n2281) );
  AND U3197 ( .A(n2276), .B(n767), .Z(n2393) );
  NAND U3198 ( .A(n2394), .B(n2395), .Z(n2279) );
  NANDN U3199 ( .B(n2396), .A(n2397), .Z(n2394) );
  XNOR U3200 ( .A(n2401), .B(n2402), .Z(n683) );
  AND U3201 ( .A(n697), .B(n2404), .Z(n2403) );
  XOR U3202 ( .A(n2399), .B(n2402), .Z(n2404) );
  XNOR U3203 ( .A(n2398), .B(n2402), .Z(n2399) );
  XNOR U3204 ( .A(n2323), .B(n2322), .Z(n2402) );
  XNOR U3205 ( .A(n2405), .B(n2327), .Z(n2322) );
  XNOR U3206 ( .A(n2406), .B(n2301), .Z(n2296) );
  XNOR U3207 ( .A(n2293), .B(n2294), .Z(n2301) );
  NAND U3208 ( .A(n875), .B(n1974), .Z(n2294) );
  XNOR U3209 ( .A(n2292), .B(n2407), .Z(n2293) );
  AND U3210 ( .A(n2075), .B(n838), .Z(n2407) );
  XNOR U3211 ( .A(n2300), .B(n2295), .Z(n2406) );
  XNOR U3212 ( .A(n2305), .B(n2415), .Z(n2306) );
  AND U3213 ( .A(n2304), .B(n765), .Z(n2415) );
  XOR U3214 ( .A(n2419), .B(n2307), .Z(n2414) );
  NAND U3215 ( .A(n797), .B(n2190), .Z(n2307) );
  IV U3216 ( .A(n2299), .Z(n2419) );
  XNOR U3217 ( .A(n2310), .B(n2424), .Z(n2311) );
  AND U3218 ( .A(n1880), .B(n917), .Z(n2424) );
  XOR U3219 ( .A(n2428), .B(n2312), .Z(n2423) );
  NAND U3220 ( .A(n961), .B(n1781), .Z(n2312) );
  IV U3221 ( .A(n2314), .Z(n2428) );
  XNOR U3222 ( .A(n2319), .B(n2320), .Z(n2316) );
  NAND U3223 ( .A(n1077), .B(n1596), .Z(n2320) );
  XNOR U3224 ( .A(n2318), .B(n2432), .Z(n2319) );
  AND U3225 ( .A(n1690), .B(n1019), .Z(n2432) );
  XNOR U3226 ( .A(n2326), .B(n2321), .Z(n2405) );
  AND U3227 ( .A(n2329), .B(n2440), .Z(n2439) );
  AND U3228 ( .A(n2441), .B(n2442), .Z(n2440) );
  NANDN U3229 ( .B(n738), .A(n2443), .Z(n2442) );
  NANDN U3230 ( .B(n2444), .A(n2445), .Z(n2441) );
  ANDN U3231 ( .A(n2331), .B(n2330), .Z(n2329) );
  NOR U3232 ( .A(n2446), .B(n2447), .Z(n2330) );
  NANDN U3233 ( .B(n2448), .A(n2449), .Z(n2331) );
  XNOR U3234 ( .A(n2453), .B(n2356), .Z(n2347) );
  XNOR U3235 ( .A(n2335), .B(n2455), .Z(n2336) );
  AND U3236 ( .A(n1412), .B(n1218), .Z(n2455) );
  XOR U3237 ( .A(n2459), .B(n2337), .Z(n2454) );
  NAND U3238 ( .A(n1158), .B(n1491), .Z(n2337) );
  IV U3239 ( .A(n2339), .Z(n2459) );
  XNOR U3240 ( .A(n2344), .B(n2345), .Z(n2341) );
  NANDN U3241 ( .B(n1040), .A(n1668), .Z(n2345) );
  XNOR U3242 ( .A(n2343), .B(n2463), .Z(n2344) );
  AND U3243 ( .A(n1576), .B(n1102), .Z(n2463) );
  XNOR U3244 ( .A(n2355), .B(n2346), .Z(n2453) );
  XOR U3245 ( .A(n2470), .B(n2365), .Z(n2355) );
  XNOR U3246 ( .A(n2352), .B(n2353), .Z(n2365) );
  NAND U3247 ( .A(n1306), .B(n1338), .Z(n2353) );
  XNOR U3248 ( .A(n2351), .B(n2471), .Z(n2352) );
  AND U3249 ( .A(n1268), .B(n1376), .Z(n2471) );
  XNOR U3250 ( .A(n2364), .B(n2354), .Z(n2470) );
  XNOR U3251 ( .A(n2359), .B(n2479), .Z(n2360) );
  AND U3252 ( .A(n1137), .B(n1546), .Z(n2479) );
  XOR U3253 ( .A(n2483), .B(n2361), .Z(n2478) );
  NAND U3254 ( .A(n1457), .B(n1200), .Z(n2361) );
  IV U3255 ( .A(n2363), .Z(n2483) );
  XNOR U3256 ( .A(n2487), .B(n2382), .Z(n2372) );
  XNOR U3257 ( .A(n2369), .B(n2370), .Z(n2382) );
  NANDN U3258 ( .B(n856), .A(n2058), .Z(n2370) );
  XNOR U3259 ( .A(n2368), .B(n2488), .Z(n2369) );
  AND U3260 ( .A(n1953), .B(n894), .Z(n2488) );
  XNOR U3261 ( .A(n2381), .B(n2371), .Z(n2487) );
  XNOR U3262 ( .A(n2376), .B(n2496), .Z(n2377) );
  AND U3263 ( .A(n1761), .B(n1002), .Z(n2496) );
  XOR U3264 ( .A(n2500), .B(n2378), .Z(n2495) );
  NAND U3265 ( .A(n948), .B(n1856), .Z(n2378) );
  IV U3266 ( .A(n2380), .Z(n2500) );
  XNOR U3267 ( .A(n2385), .B(n2505), .Z(n2386) );
  AND U3268 ( .A(n2165), .B(n830), .Z(n2505) );
  XOR U3269 ( .A(n2509), .B(n2387), .Z(n2504) );
  NAND U3270 ( .A(n793), .B(n2276), .Z(n2387) );
  IV U3271 ( .A(n2389), .Z(n2509) );
  XNOR U3272 ( .A(n2396), .B(n2397), .Z(n2391) );
  NANDN U3273 ( .B(n737), .A(n2513), .Z(n2397) );
  XNOR U3274 ( .A(n2395), .B(n2514), .Z(n2396) );
  AND U3275 ( .A(n2392), .B(n767), .Z(n2514) );
  ANDN U3276 ( .A(n2515), .B(n2516), .Z(n2395) );
  NANDN U3277 ( .B(n2517), .A(n2518), .Z(n2515) );
  XNOR U3278 ( .A(n2522), .B(n2523), .Z(n684) );
  AND U3279 ( .A(n697), .B(n2525), .Z(n2524) );
  XOR U3280 ( .A(n2520), .B(n2523), .Z(n2525) );
  XNOR U3281 ( .A(n2519), .B(n2523), .Z(n2520) );
  XNOR U3282 ( .A(n2438), .B(n2437), .Z(n2523) );
  XNOR U3283 ( .A(n2526), .B(n2452), .Z(n2437) );
  XNOR U3284 ( .A(n2527), .B(n2422), .Z(n2412) );
  XNOR U3285 ( .A(n2409), .B(n2410), .Z(n2422) );
  NAND U3286 ( .A(n917), .B(n1974), .Z(n2410) );
  XNOR U3287 ( .A(n2408), .B(n2528), .Z(n2409) );
  AND U3288 ( .A(n2075), .B(n875), .Z(n2528) );
  XNOR U3289 ( .A(n2421), .B(n2411), .Z(n2527) );
  XNOR U3290 ( .A(n2416), .B(n2536), .Z(n2417) );
  AND U3291 ( .A(n2304), .B(n797), .Z(n2536) );
  XOR U3292 ( .A(n2540), .B(n2418), .Z(n2535) );
  NAND U3293 ( .A(n838), .B(n2190), .Z(n2418) );
  IV U3294 ( .A(n2420), .Z(n2540) );
  XNOR U3295 ( .A(n2425), .B(n2545), .Z(n2426) );
  AND U3296 ( .A(n1880), .B(n961), .Z(n2545) );
  XOR U3297 ( .A(n2549), .B(n2427), .Z(n2544) );
  NAND U3298 ( .A(n1019), .B(n1781), .Z(n2427) );
  IV U3299 ( .A(n2429), .Z(n2549) );
  XNOR U3300 ( .A(n2434), .B(n2435), .Z(n2431) );
  NAND U3301 ( .A(n1137), .B(n1596), .Z(n2435) );
  XNOR U3302 ( .A(n2433), .B(n2553), .Z(n2434) );
  AND U3303 ( .A(n1690), .B(n1077), .Z(n2553) );
  XNOR U3304 ( .A(n2451), .B(n2436), .Z(n2526) );
  XOR U3305 ( .A(n2560), .B(n2445), .Z(n2451) );
  XNOR U3306 ( .A(n2448), .B(n2449), .Z(n2445) );
  XOR U3307 ( .A(n2564), .B(n2447), .Z(n2448) );
  NAND U3308 ( .A(n765), .B(n2443), .Z(n2447) );
  NANDN U3309 ( .B(n738), .A(n2566), .Z(n2565) );
  OR U3310 ( .A(n2570), .B(n2571), .Z(n2444) );
  XNOR U3311 ( .A(n2575), .B(n2477), .Z(n2468) );
  XNOR U3312 ( .A(n2456), .B(n2577), .Z(n2457) );
  AND U3313 ( .A(n1491), .B(n1218), .Z(n2577) );
  XOR U3314 ( .A(n2581), .B(n2458), .Z(n2576) );
  NAND U3315 ( .A(n1158), .B(n1576), .Z(n2458) );
  IV U3316 ( .A(n2460), .Z(n2581) );
  XNOR U3317 ( .A(n2465), .B(n2466), .Z(n2462) );
  NANDN U3318 ( .B(n1040), .A(n1761), .Z(n2466) );
  XNOR U3319 ( .A(n2464), .B(n2585), .Z(n2465) );
  AND U3320 ( .A(n1668), .B(n1102), .Z(n2585) );
  XNOR U3321 ( .A(n2476), .B(n2467), .Z(n2575) );
  XOR U3322 ( .A(n2592), .B(n2486), .Z(n2476) );
  XNOR U3323 ( .A(n2473), .B(n2474), .Z(n2486) );
  NAND U3324 ( .A(n1306), .B(n1412), .Z(n2474) );
  XNOR U3325 ( .A(n2472), .B(n2593), .Z(n2473) );
  AND U3326 ( .A(n1338), .B(n1376), .Z(n2593) );
  XNOR U3327 ( .A(n2485), .B(n2475), .Z(n2592) );
  XNOR U3328 ( .A(n2480), .B(n2601), .Z(n2481) );
  AND U3329 ( .A(n1200), .B(n1546), .Z(n2601) );
  XOR U3330 ( .A(n2605), .B(n2482), .Z(n2600) );
  NAND U3331 ( .A(n1457), .B(n1268), .Z(n2482) );
  IV U3332 ( .A(n2484), .Z(n2605) );
  XNOR U3333 ( .A(n2609), .B(n2503), .Z(n2493) );
  XNOR U3334 ( .A(n2490), .B(n2491), .Z(n2503) );
  NANDN U3335 ( .B(n856), .A(n2165), .Z(n2491) );
  XNOR U3336 ( .A(n2489), .B(n2610), .Z(n2490) );
  AND U3337 ( .A(n2058), .B(n894), .Z(n2610) );
  XNOR U3338 ( .A(n2502), .B(n2492), .Z(n2609) );
  XNOR U3339 ( .A(n2497), .B(n2618), .Z(n2498) );
  AND U3340 ( .A(n1856), .B(n1002), .Z(n2618) );
  XOR U3341 ( .A(n2622), .B(n2499), .Z(n2617) );
  NAND U3342 ( .A(n948), .B(n1953), .Z(n2499) );
  IV U3343 ( .A(n2501), .Z(n2622) );
  XNOR U3344 ( .A(n2506), .B(n2627), .Z(n2507) );
  AND U3345 ( .A(n2276), .B(n830), .Z(n2627) );
  XOR U3346 ( .A(n2631), .B(n2508), .Z(n2626) );
  NAND U3347 ( .A(n793), .B(n2392), .Z(n2508) );
  IV U3348 ( .A(n2510), .Z(n2631) );
  XNOR U3349 ( .A(n2517), .B(n2518), .Z(n2512) );
  NANDN U3350 ( .B(n737), .A(n2635), .Z(n2518) );
  AND U3351 ( .A(n2513), .B(n767), .Z(n2636) );
  NAND U3352 ( .A(n2637), .B(n2638), .Z(n2516) );
  NANDN U3353 ( .B(n2639), .A(n2640), .Z(n2637) );
  XOR U3354 ( .A(n2644), .B(n2645), .Z(n685) );
  AND U3355 ( .A(n697), .B(n2647), .Z(n2646) );
  XNOR U3356 ( .A(n2642), .B(n2645), .Z(n2647) );
  XNOR U3357 ( .A(n2645), .B(n2641), .Z(n2642) );
  OR U3358 ( .A(n2648), .B(n2649), .Z(n2641) );
  XNOR U3359 ( .A(n2559), .B(n2558), .Z(n2645) );
  XNOR U3360 ( .A(n2650), .B(n2574), .Z(n2558) );
  XNOR U3361 ( .A(n2651), .B(n2543), .Z(n2533) );
  XNOR U3362 ( .A(n2530), .B(n2531), .Z(n2543) );
  NAND U3363 ( .A(n961), .B(n1974), .Z(n2531) );
  XNOR U3364 ( .A(n2529), .B(n2652), .Z(n2530) );
  AND U3365 ( .A(n2075), .B(n917), .Z(n2652) );
  XNOR U3366 ( .A(n2542), .B(n2532), .Z(n2651) );
  XNOR U3367 ( .A(n2537), .B(n2660), .Z(n2538) );
  AND U3368 ( .A(n2304), .B(n838), .Z(n2660) );
  XOR U3369 ( .A(n2664), .B(n2539), .Z(n2659) );
  NAND U3370 ( .A(n875), .B(n2190), .Z(n2539) );
  IV U3371 ( .A(n2541), .Z(n2664) );
  XNOR U3372 ( .A(n2546), .B(n2669), .Z(n2547) );
  AND U3373 ( .A(n1880), .B(n1019), .Z(n2669) );
  XOR U3374 ( .A(n2673), .B(n2548), .Z(n2668) );
  NAND U3375 ( .A(n1077), .B(n1781), .Z(n2548) );
  IV U3376 ( .A(n2550), .Z(n2673) );
  XNOR U3377 ( .A(n2555), .B(n2556), .Z(n2552) );
  NAND U3378 ( .A(n1200), .B(n1596), .Z(n2556) );
  XNOR U3379 ( .A(n2554), .B(n2677), .Z(n2555) );
  AND U3380 ( .A(n1690), .B(n1137), .Z(n2677) );
  XNOR U3381 ( .A(n2573), .B(n2557), .Z(n2650) );
  XNOR U3382 ( .A(n2684), .B(n2570), .Z(n2573) );
  XOR U3383 ( .A(n2563), .B(n2562), .Z(n2570) );
  XOR U3384 ( .A(n2561), .B(n2685), .Z(n2562) );
  AND U3385 ( .A(n2686), .B(n2687), .Z(n2685) );
  NANDN U3386 ( .B(n738), .A(n2688), .Z(n2687) );
  OR U3387 ( .A(n2689), .B(n2690), .Z(n2686) );
  NAND U3388 ( .A(n797), .B(n2443), .Z(n2569) );
  XNOR U3389 ( .A(n2567), .B(n2694), .Z(n2568) );
  AND U3390 ( .A(n2566), .B(n765), .Z(n2694) );
  NANDN U3391 ( .B(n2698), .A(n2699), .Z(n2571) );
  XNOR U3392 ( .A(n2703), .B(n2599), .Z(n2590) );
  XNOR U3393 ( .A(n2578), .B(n2705), .Z(n2579) );
  AND U3394 ( .A(n1576), .B(n1218), .Z(n2705) );
  XOR U3395 ( .A(n2709), .B(n2580), .Z(n2704) );
  NAND U3396 ( .A(n1158), .B(n1668), .Z(n2580) );
  IV U3397 ( .A(n2582), .Z(n2709) );
  XNOR U3398 ( .A(n2587), .B(n2588), .Z(n2584) );
  NANDN U3399 ( .B(n1040), .A(n1856), .Z(n2588) );
  XNOR U3400 ( .A(n2586), .B(n2713), .Z(n2587) );
  AND U3401 ( .A(n1761), .B(n1102), .Z(n2713) );
  XNOR U3402 ( .A(n2598), .B(n2589), .Z(n2703) );
  XOR U3403 ( .A(n2720), .B(n2608), .Z(n2598) );
  XNOR U3404 ( .A(n2595), .B(n2596), .Z(n2608) );
  NAND U3405 ( .A(n1306), .B(n1491), .Z(n2596) );
  XNOR U3406 ( .A(n2594), .B(n2721), .Z(n2595) );
  AND U3407 ( .A(n1412), .B(n1376), .Z(n2721) );
  XNOR U3408 ( .A(n2607), .B(n2597), .Z(n2720) );
  XNOR U3409 ( .A(n2602), .B(n2729), .Z(n2603) );
  AND U3410 ( .A(n1268), .B(n1546), .Z(n2729) );
  XOR U3411 ( .A(n2733), .B(n2604), .Z(n2728) );
  NAND U3412 ( .A(n1457), .B(n1338), .Z(n2604) );
  IV U3413 ( .A(n2606), .Z(n2733) );
  XNOR U3414 ( .A(n2737), .B(n2625), .Z(n2615) );
  XNOR U3415 ( .A(n2612), .B(n2613), .Z(n2625) );
  NANDN U3416 ( .B(n856), .A(n2276), .Z(n2613) );
  XNOR U3417 ( .A(n2611), .B(n2738), .Z(n2612) );
  AND U3418 ( .A(n2165), .B(n894), .Z(n2738) );
  XNOR U3419 ( .A(n2624), .B(n2614), .Z(n2737) );
  XNOR U3420 ( .A(n2619), .B(n2746), .Z(n2620) );
  AND U3421 ( .A(n1953), .B(n1002), .Z(n2746) );
  XOR U3422 ( .A(n2750), .B(n2621), .Z(n2745) );
  NAND U3423 ( .A(n948), .B(n2058), .Z(n2621) );
  IV U3424 ( .A(n2623), .Z(n2750) );
  XNOR U3425 ( .A(n2628), .B(n2755), .Z(n2629) );
  AND U3426 ( .A(n2392), .B(n830), .Z(n2755) );
  XOR U3427 ( .A(n2759), .B(n2630), .Z(n2754) );
  NAND U3428 ( .A(n793), .B(n2513), .Z(n2630) );
  IV U3429 ( .A(n2632), .Z(n2759) );
  XNOR U3430 ( .A(n2639), .B(n2640), .Z(n2634) );
  NANDN U3431 ( .B(n737), .A(n2763), .Z(n2640) );
  XNOR U3432 ( .A(n2638), .B(n2764), .Z(n2639) );
  AND U3433 ( .A(n2635), .B(n767), .Z(n2764) );
  ANDN U3434 ( .A(n2765), .B(n2766), .Z(n2638) );
  NANDN U3435 ( .B(n2767), .A(n2768), .Z(n2765) );
  XNOR U3436 ( .A(n2770), .B(n2771), .Z(n723) );
  AND U3437 ( .A(n697), .B(n2773), .Z(n2772) );
  XOR U3438 ( .A(n2648), .B(n2774), .Z(n2773) );
  XOR U3439 ( .A(n2774), .B(n2649), .Z(n2648) );
  OR U3440 ( .A(n2775), .B(n2776), .Z(n2649) );
  IV U3441 ( .A(n2771), .Z(n2774) );
  XOR U3442 ( .A(n2683), .B(n2682), .Z(n2771) );
  XNOR U3443 ( .A(n2777), .B(n2702), .Z(n2682) );
  XNOR U3444 ( .A(n2778), .B(n2667), .Z(n2657) );
  XNOR U3445 ( .A(n2654), .B(n2655), .Z(n2667) );
  NAND U3446 ( .A(n1019), .B(n1974), .Z(n2655) );
  XNOR U3447 ( .A(n2653), .B(n2779), .Z(n2654) );
  AND U3448 ( .A(n2075), .B(n961), .Z(n2779) );
  XNOR U3449 ( .A(n2666), .B(n2656), .Z(n2778) );
  XNOR U3450 ( .A(n2661), .B(n2787), .Z(n2662) );
  AND U3451 ( .A(n2304), .B(n875), .Z(n2787) );
  XOR U3452 ( .A(n2791), .B(n2663), .Z(n2786) );
  NAND U3453 ( .A(n917), .B(n2190), .Z(n2663) );
  IV U3454 ( .A(n2665), .Z(n2791) );
  XNOR U3455 ( .A(n2670), .B(n2796), .Z(n2671) );
  AND U3456 ( .A(n1880), .B(n1077), .Z(n2796) );
  XOR U3457 ( .A(n2800), .B(n2672), .Z(n2795) );
  NAND U3458 ( .A(n1137), .B(n1781), .Z(n2672) );
  IV U3459 ( .A(n2674), .Z(n2800) );
  XNOR U3460 ( .A(n2679), .B(n2680), .Z(n2676) );
  NAND U3461 ( .A(n1268), .B(n1596), .Z(n2680) );
  XNOR U3462 ( .A(n2678), .B(n2804), .Z(n2679) );
  AND U3463 ( .A(n1690), .B(n1200), .Z(n2804) );
  XNOR U3464 ( .A(n2701), .B(n2681), .Z(n2777) );
  XNOR U3465 ( .A(n2811), .B(n2698), .Z(n2701) );
  XOR U3466 ( .A(n2693), .B(n2692), .Z(n2698) );
  XNOR U3467 ( .A(n2816), .B(n2689), .Z(n2812) );
  NAND U3468 ( .A(n765), .B(n2688), .Z(n2689) );
  NANDN U3469 ( .B(n738), .A(n2818), .Z(n2817) );
  NAND U3470 ( .A(n838), .B(n2443), .Z(n2697) );
  XNOR U3471 ( .A(n2695), .B(n2822), .Z(n2696) );
  AND U3472 ( .A(n2566), .B(n797), .Z(n2822) );
  XNOR U3473 ( .A(n2699), .B(n2700), .Z(n2811) );
  XNOR U3474 ( .A(n2832), .B(n2727), .Z(n2718) );
  XNOR U3475 ( .A(n2706), .B(n2834), .Z(n2707) );
  AND U3476 ( .A(n1668), .B(n1218), .Z(n2834) );
  XOR U3477 ( .A(n2838), .B(n2708), .Z(n2833) );
  NAND U3478 ( .A(n1158), .B(n1761), .Z(n2708) );
  IV U3479 ( .A(n2710), .Z(n2838) );
  XNOR U3480 ( .A(n2715), .B(n2716), .Z(n2712) );
  NANDN U3481 ( .B(n1040), .A(n1953), .Z(n2716) );
  XNOR U3482 ( .A(n2714), .B(n2842), .Z(n2715) );
  AND U3483 ( .A(n1856), .B(n1102), .Z(n2842) );
  XNOR U3484 ( .A(n2726), .B(n2717), .Z(n2832) );
  XOR U3485 ( .A(n2849), .B(n2736), .Z(n2726) );
  XNOR U3486 ( .A(n2723), .B(n2724), .Z(n2736) );
  NAND U3487 ( .A(n1306), .B(n1576), .Z(n2724) );
  XNOR U3488 ( .A(n2722), .B(n2850), .Z(n2723) );
  AND U3489 ( .A(n1491), .B(n1376), .Z(n2850) );
  XNOR U3490 ( .A(n2735), .B(n2725), .Z(n2849) );
  XNOR U3491 ( .A(n2730), .B(n2858), .Z(n2731) );
  AND U3492 ( .A(n1338), .B(n1546), .Z(n2858) );
  XOR U3493 ( .A(n2862), .B(n2732), .Z(n2857) );
  NAND U3494 ( .A(n1457), .B(n1412), .Z(n2732) );
  IV U3495 ( .A(n2734), .Z(n2862) );
  XNOR U3496 ( .A(n2866), .B(n2753), .Z(n2743) );
  XNOR U3497 ( .A(n2740), .B(n2741), .Z(n2753) );
  NANDN U3498 ( .B(n856), .A(n2392), .Z(n2741) );
  XNOR U3499 ( .A(n2739), .B(n2867), .Z(n2740) );
  AND U3500 ( .A(n2276), .B(n894), .Z(n2867) );
  XNOR U3501 ( .A(n2752), .B(n2742), .Z(n2866) );
  XNOR U3502 ( .A(n2747), .B(n2875), .Z(n2748) );
  AND U3503 ( .A(n2058), .B(n1002), .Z(n2875) );
  XOR U3504 ( .A(n2879), .B(n2749), .Z(n2874) );
  NAND U3505 ( .A(n948), .B(n2165), .Z(n2749) );
  IV U3506 ( .A(n2751), .Z(n2879) );
  XNOR U3507 ( .A(n2756), .B(n2884), .Z(n2757) );
  AND U3508 ( .A(n2513), .B(n830), .Z(n2884) );
  XOR U3509 ( .A(n2888), .B(n2758), .Z(n2883) );
  NAND U3510 ( .A(n793), .B(n2635), .Z(n2758) );
  IV U3511 ( .A(n2760), .Z(n2888) );
  XNOR U3512 ( .A(n2767), .B(n2768), .Z(n2762) );
  OR U3513 ( .A(n2892), .B(n737), .Z(n2768) );
  AND U3514 ( .A(n2763), .B(n767), .Z(n2893) );
  NAND U3515 ( .A(n2894), .B(n2895), .Z(n2766) );
  NANDN U3516 ( .B(n2896), .A(n2897), .Z(n2894) );
  XNOR U3517 ( .A(n2899), .B(n2900), .Z(n1146) );
  XOR U3518 ( .A(n2898), .B(n2901), .Z(n2899) );
  AND U3519 ( .A(n697), .B(n2902), .Z(n2901) );
  XOR U3520 ( .A(n2775), .B(n2903), .Z(n2902) );
  XOR U3521 ( .A(n2903), .B(n2776), .Z(n2775) );
  NANDN U3522 ( .B(n2904), .A(n2905), .Z(n2776) );
  IV U3523 ( .A(n2900), .Z(n2903) );
  XOR U3524 ( .A(n2810), .B(n2809), .Z(n2900) );
  XNOR U3525 ( .A(n2906), .B(n2828), .Z(n2809) );
  XNOR U3526 ( .A(n2907), .B(n2794), .Z(n2784) );
  XNOR U3527 ( .A(n2781), .B(n2782), .Z(n2794) );
  NAND U3528 ( .A(n1077), .B(n1974), .Z(n2782) );
  XNOR U3529 ( .A(n2780), .B(n2908), .Z(n2781) );
  AND U3530 ( .A(n2075), .B(n1019), .Z(n2908) );
  XNOR U3531 ( .A(n2793), .B(n2783), .Z(n2907) );
  XNOR U3532 ( .A(n2788), .B(n2916), .Z(n2789) );
  AND U3533 ( .A(n2304), .B(n917), .Z(n2916) );
  XOR U3534 ( .A(n2920), .B(n2790), .Z(n2915) );
  NAND U3535 ( .A(n961), .B(n2190), .Z(n2790) );
  IV U3536 ( .A(n2792), .Z(n2920) );
  XNOR U3537 ( .A(n2797), .B(n2925), .Z(n2798) );
  AND U3538 ( .A(n1880), .B(n1137), .Z(n2925) );
  XOR U3539 ( .A(n2929), .B(n2799), .Z(n2924) );
  NAND U3540 ( .A(n1200), .B(n1781), .Z(n2799) );
  IV U3541 ( .A(n2801), .Z(n2929) );
  XNOR U3542 ( .A(n2806), .B(n2807), .Z(n2803) );
  NAND U3543 ( .A(n1338), .B(n1596), .Z(n2807) );
  XNOR U3544 ( .A(n2805), .B(n2933), .Z(n2806) );
  AND U3545 ( .A(n1690), .B(n1268), .Z(n2933) );
  XNOR U3546 ( .A(n2827), .B(n2808), .Z(n2906) );
  XOR U3547 ( .A(n2940), .B(n2831), .Z(n2827) );
  XNOR U3548 ( .A(n2819), .B(n2942), .Z(n2820) );
  AND U3549 ( .A(n2818), .B(n765), .Z(n2942) );
  XOR U3550 ( .A(n2946), .B(n2821), .Z(n2941) );
  NAND U3551 ( .A(n797), .B(n2688), .Z(n2821) );
  IV U3552 ( .A(n2813), .Z(n2946) );
  XNOR U3553 ( .A(n2824), .B(n2825), .Z(n2815) );
  NAND U3554 ( .A(n875), .B(n2443), .Z(n2825) );
  XNOR U3555 ( .A(n2823), .B(n2950), .Z(n2824) );
  AND U3556 ( .A(n2566), .B(n838), .Z(n2950) );
  XNOR U3557 ( .A(n2830), .B(n2826), .Z(n2940) );
  AND U3558 ( .A(n2958), .B(n2959), .Z(n2957) );
  OR U3559 ( .A(n2960), .B(n2961), .Z(n2959) );
  AND U3560 ( .A(n2962), .B(n2963), .Z(n2958) );
  NANDN U3561 ( .B(n738), .A(n2964), .Z(n2963) );
  NANDN U3562 ( .B(n2965), .A(n2966), .Z(n2962) );
  XNOR U3563 ( .A(n2970), .B(n2856), .Z(n2847) );
  XNOR U3564 ( .A(n2835), .B(n2972), .Z(n2836) );
  AND U3565 ( .A(n1761), .B(n1218), .Z(n2972) );
  XOR U3566 ( .A(n2976), .B(n2837), .Z(n2971) );
  NAND U3567 ( .A(n1158), .B(n1856), .Z(n2837) );
  IV U3568 ( .A(n2839), .Z(n2976) );
  XNOR U3569 ( .A(n2844), .B(n2845), .Z(n2841) );
  NANDN U3570 ( .B(n1040), .A(n2058), .Z(n2845) );
  XNOR U3571 ( .A(n2843), .B(n2980), .Z(n2844) );
  AND U3572 ( .A(n1953), .B(n1102), .Z(n2980) );
  XNOR U3573 ( .A(n2855), .B(n2846), .Z(n2970) );
  XOR U3574 ( .A(n2987), .B(n2865), .Z(n2855) );
  XNOR U3575 ( .A(n2852), .B(n2853), .Z(n2865) );
  NAND U3576 ( .A(n1306), .B(n1668), .Z(n2853) );
  XNOR U3577 ( .A(n2851), .B(n2988), .Z(n2852) );
  AND U3578 ( .A(n1576), .B(n1376), .Z(n2988) );
  XNOR U3579 ( .A(n2864), .B(n2854), .Z(n2987) );
  XNOR U3580 ( .A(n2859), .B(n2996), .Z(n2860) );
  AND U3581 ( .A(n1412), .B(n1546), .Z(n2996) );
  XOR U3582 ( .A(n3000), .B(n2861), .Z(n2995) );
  NAND U3583 ( .A(n1457), .B(n1491), .Z(n2861) );
  IV U3584 ( .A(n2863), .Z(n3000) );
  XNOR U3585 ( .A(n3004), .B(n2882), .Z(n2872) );
  XNOR U3586 ( .A(n2869), .B(n2870), .Z(n2882) );
  NANDN U3587 ( .B(n856), .A(n2513), .Z(n2870) );
  XNOR U3588 ( .A(n2868), .B(n3005), .Z(n2869) );
  AND U3589 ( .A(n2392), .B(n894), .Z(n3005) );
  XNOR U3590 ( .A(n2881), .B(n2871), .Z(n3004) );
  XNOR U3591 ( .A(n2876), .B(n3013), .Z(n2877) );
  AND U3592 ( .A(n2165), .B(n1002), .Z(n3013) );
  XOR U3593 ( .A(n3017), .B(n2878), .Z(n3012) );
  NAND U3594 ( .A(n948), .B(n2276), .Z(n2878) );
  IV U3595 ( .A(n2880), .Z(n3017) );
  XNOR U3596 ( .A(n2885), .B(n3022), .Z(n2886) );
  AND U3597 ( .A(n2635), .B(n830), .Z(n3022) );
  XOR U3598 ( .A(n3026), .B(n2887), .Z(n3021) );
  NAND U3599 ( .A(n793), .B(n2763), .Z(n2887) );
  IV U3600 ( .A(n2889), .Z(n3026) );
  XNOR U3601 ( .A(n2896), .B(n2897), .Z(n2891) );
  OR U3602 ( .A(n3030), .B(n737), .Z(n2897) );
  XNOR U3603 ( .A(n2895), .B(n3031), .Z(n2896) );
  ANDN U3604 ( .A(n767), .B(n2892), .Z(n3031) );
  ANDN U3605 ( .A(n3032), .B(n3033), .Z(n2895) );
  NANDN U3606 ( .B(n3034), .A(n3035), .Z(n3032) );
  XOR U3607 ( .A(n3037), .B(o_reg[1]), .Z(o[0]) );
  XOR U3608 ( .A(n3038), .B(n3039), .Z(n3037) );
  XNOR U3609 ( .A(n3040), .B(n3036), .Z(n3038) );
  NANDN U3610 ( .B(n2905), .A(o_reg[0]), .Z(n3036) );
  NAND U3611 ( .A(n3041), .B(n697), .Z(n3040) );
  XOR U3612 ( .A(e_input[31]), .B(g_input[31]), .Z(n697) );
  XNOR U3613 ( .A(n2904), .B(n3039), .Z(n3041) );
  XOR U3614 ( .A(n2905), .B(n3039), .Z(n2904) );
  XOR U3615 ( .A(n2939), .B(n2938), .Z(n3039) );
  XNOR U3616 ( .A(n3042), .B(n2956), .Z(n2938) );
  XNOR U3617 ( .A(n3043), .B(n2923), .Z(n2913) );
  XNOR U3618 ( .A(n2910), .B(n2911), .Z(n2923) );
  NAND U3619 ( .A(n1137), .B(n1974), .Z(n2911) );
  XNOR U3620 ( .A(n2909), .B(n3044), .Z(n2910) );
  AND U3621 ( .A(n2075), .B(n1077), .Z(n3044) );
  XNOR U3622 ( .A(n2922), .B(n2912), .Z(n3043) );
  XNOR U3623 ( .A(n2917), .B(n3052), .Z(n2918) );
  AND U3624 ( .A(n2304), .B(n961), .Z(n3052) );
  XOR U3625 ( .A(n3056), .B(n2919), .Z(n3051) );
  NAND U3626 ( .A(n1019), .B(n2190), .Z(n2919) );
  IV U3627 ( .A(n2921), .Z(n3056) );
  XNOR U3628 ( .A(n2926), .B(n3061), .Z(n2927) );
  AND U3629 ( .A(n1880), .B(n1200), .Z(n3061) );
  XOR U3630 ( .A(n3065), .B(n2928), .Z(n3060) );
  NAND U3631 ( .A(n1268), .B(n1781), .Z(n2928) );
  IV U3632 ( .A(n2930), .Z(n3065) );
  XNOR U3633 ( .A(n2935), .B(n2936), .Z(n2932) );
  NAND U3634 ( .A(n1412), .B(n1596), .Z(n2936) );
  XNOR U3635 ( .A(n2934), .B(n3069), .Z(n2935) );
  AND U3636 ( .A(n1690), .B(n1338), .Z(n3069) );
  XNOR U3637 ( .A(n2955), .B(n2937), .Z(n3042) );
  XOR U3638 ( .A(n3076), .B(n2969), .Z(n2955) );
  XNOR U3639 ( .A(n2943), .B(n3078), .Z(n2944) );
  AND U3640 ( .A(n2818), .B(n797), .Z(n3078) );
  XOR U3641 ( .A(n3082), .B(n2945), .Z(n3077) );
  NAND U3642 ( .A(n838), .B(n2688), .Z(n2945) );
  IV U3643 ( .A(n2947), .Z(n3082) );
  XNOR U3644 ( .A(n2952), .B(n2953), .Z(n2949) );
  NAND U3645 ( .A(n917), .B(n2443), .Z(n2953) );
  XNOR U3646 ( .A(n2951), .B(n3086), .Z(n2952) );
  AND U3647 ( .A(n2566), .B(n875), .Z(n3086) );
  XNOR U3648 ( .A(n2968), .B(n2954), .Z(n3076) );
  XNOR U3649 ( .A(n3093), .B(n2965), .Z(n2968) );
  XOR U3650 ( .A(n3094), .B(n2960), .Z(n2965) );
  NAND U3651 ( .A(n765), .B(n2964), .Z(n2960) );
  NANDN U3652 ( .B(n738), .A(n3096), .Z(n3095) );
  XNOR U3653 ( .A(n2966), .B(n2967), .Z(n3093) );
  XNOR U3654 ( .A(n3105), .B(n2994), .Z(n2985) );
  XNOR U3655 ( .A(n2973), .B(n3107), .Z(n2974) );
  AND U3656 ( .A(n1856), .B(n1218), .Z(n3107) );
  XOR U3657 ( .A(n3111), .B(n2975), .Z(n3106) );
  NAND U3658 ( .A(n1158), .B(n1953), .Z(n2975) );
  IV U3659 ( .A(n2977), .Z(n3111) );
  XNOR U3660 ( .A(n2982), .B(n2983), .Z(n2979) );
  NANDN U3661 ( .B(n1040), .A(n2165), .Z(n2983) );
  XNOR U3662 ( .A(n2981), .B(n3115), .Z(n2982) );
  AND U3663 ( .A(n2058), .B(n1102), .Z(n3115) );
  XNOR U3664 ( .A(n2993), .B(n2984), .Z(n3105) );
  XOR U3665 ( .A(n3122), .B(n3003), .Z(n2993) );
  XNOR U3666 ( .A(n2990), .B(n2991), .Z(n3003) );
  NAND U3667 ( .A(n1306), .B(n1761), .Z(n2991) );
  XNOR U3668 ( .A(n2989), .B(n3123), .Z(n2990) );
  AND U3669 ( .A(n1668), .B(n1376), .Z(n3123) );
  XNOR U3670 ( .A(n3002), .B(n2992), .Z(n3122) );
  XNOR U3671 ( .A(n2997), .B(n3131), .Z(n2998) );
  AND U3672 ( .A(n1491), .B(n1546), .Z(n3131) );
  XOR U3673 ( .A(n3135), .B(n2999), .Z(n3130) );
  NAND U3674 ( .A(n1457), .B(n1576), .Z(n2999) );
  IV U3675 ( .A(n3001), .Z(n3135) );
  XNOR U3676 ( .A(n3139), .B(n3020), .Z(n3010) );
  XNOR U3677 ( .A(n3007), .B(n3008), .Z(n3020) );
  NANDN U3678 ( .B(n856), .A(n2635), .Z(n3008) );
  XNOR U3679 ( .A(n3006), .B(n3140), .Z(n3007) );
  AND U3680 ( .A(n2513), .B(n894), .Z(n3140) );
  XNOR U3681 ( .A(n3019), .B(n3009), .Z(n3139) );
  XNOR U3682 ( .A(n3014), .B(n3148), .Z(n3015) );
  AND U3683 ( .A(n2276), .B(n1002), .Z(n3148) );
  XOR U3684 ( .A(n3152), .B(n3016), .Z(n3147) );
  NAND U3685 ( .A(n948), .B(n2392), .Z(n3016) );
  IV U3686 ( .A(n3018), .Z(n3152) );
  XNOR U3687 ( .A(n3023), .B(n3157), .Z(n3024) );
  AND U3688 ( .A(n2763), .B(n830), .Z(n3157) );
  XOR U3689 ( .A(n3161), .B(n3025), .Z(n3156) );
  NANDN U3690 ( .B(n2892), .A(n793), .Z(n3025) );
  IV U3691 ( .A(n3027), .Z(n3161) );
  XNOR U3692 ( .A(n3034), .B(n3035), .Z(n3029) );
  NANDN U3693 ( .B(n737), .A(n3165), .Z(n3035) );
  ANDN U3694 ( .A(n767), .B(n3030), .Z(n3166) );
  NAND U3695 ( .A(n3167), .B(n3168), .Z(n3033) );
  NANDN U3696 ( .B(n3169), .A(n3170), .Z(n3167) );
  XOR U3697 ( .A(n3075), .B(n3074), .Z(n2905) );
  XNOR U3698 ( .A(n3171), .B(n3092), .Z(n3074) );
  XNOR U3699 ( .A(n3172), .B(n3059), .Z(n3049) );
  XNOR U3700 ( .A(n3046), .B(n3047), .Z(n3059) );
  NAND U3701 ( .A(n1200), .B(n1974), .Z(n3047) );
  XNOR U3702 ( .A(n3045), .B(n3173), .Z(n3046) );
  AND U3703 ( .A(n2075), .B(n1137), .Z(n3173) );
  XNOR U3704 ( .A(n3058), .B(n3048), .Z(n3172) );
  XNOR U3705 ( .A(n3053), .B(n3181), .Z(n3054) );
  AND U3706 ( .A(n2304), .B(n1019), .Z(n3181) );
  XOR U3707 ( .A(n3185), .B(n3055), .Z(n3180) );
  NAND U3708 ( .A(n1077), .B(n2190), .Z(n3055) );
  IV U3709 ( .A(n3057), .Z(n3185) );
  XNOR U3710 ( .A(n3062), .B(n3190), .Z(n3063) );
  AND U3711 ( .A(n1880), .B(n1268), .Z(n3190) );
  XOR U3712 ( .A(n3194), .B(n3064), .Z(n3189) );
  NAND U3713 ( .A(n1338), .B(n1781), .Z(n3064) );
  IV U3714 ( .A(n3066), .Z(n3194) );
  XNOR U3715 ( .A(n3071), .B(n3072), .Z(n3068) );
  NAND U3716 ( .A(n1491), .B(n1596), .Z(n3072) );
  XNOR U3717 ( .A(n3070), .B(n3198), .Z(n3071) );
  AND U3718 ( .A(n1690), .B(n1412), .Z(n3198) );
  XNOR U3719 ( .A(n3091), .B(n3073), .Z(n3171) );
  XOR U3720 ( .A(n3202), .B(n3203), .Z(n3073) );
  XOR U3721 ( .A(n3204), .B(n3102), .Z(n3091) );
  XNOR U3722 ( .A(n3079), .B(n3206), .Z(n3080) );
  AND U3723 ( .A(n2818), .B(n838), .Z(n3206) );
  XOR U3724 ( .A(n3210), .B(n3081), .Z(n3205) );
  NAND U3725 ( .A(n875), .B(n2688), .Z(n3081) );
  IV U3726 ( .A(n3083), .Z(n3210) );
  XNOR U3727 ( .A(n3088), .B(n3089), .Z(n3085) );
  NAND U3728 ( .A(n961), .B(n2443), .Z(n3089) );
  XNOR U3729 ( .A(n3087), .B(n3214), .Z(n3088) );
  AND U3730 ( .A(n2566), .B(n917), .Z(n3214) );
  XNOR U3731 ( .A(n3101), .B(n3090), .Z(n3204) );
  XOR U3732 ( .A(n3218), .B(n3219), .Z(n3090) );
  AND U3733 ( .A(n3220), .B(n3221), .Z(n3219) );
  XNOR U3734 ( .A(n3222), .B(n3223), .Z(n3221) );
  XOR U3735 ( .A(n3224), .B(n3218), .Z(n3222) );
  XOR U3736 ( .A(n3178), .B(n3225), .Z(n3220) );
  XNOR U3737 ( .A(n3218), .B(n3179), .Z(n3225) );
  XNOR U3738 ( .A(n3191), .B(n3227), .Z(n3192) );
  AND U3739 ( .A(n1880), .B(n1338), .Z(n3227) );
  XOR U3740 ( .A(n3231), .B(n3193), .Z(n3226) );
  NAND U3741 ( .A(n1412), .B(n1781), .Z(n3193) );
  IV U3742 ( .A(n3195), .Z(n3231) );
  XNOR U3743 ( .A(n3200), .B(n3201), .Z(n3197) );
  NAND U3744 ( .A(n1596), .B(n1576), .Z(n3201) );
  XNOR U3745 ( .A(n3199), .B(n3235), .Z(n3200) );
  AND U3746 ( .A(n1690), .B(n1491), .Z(n3235) );
  XOR U3747 ( .A(n3239), .B(n3188), .Z(n3178) );
  XNOR U3748 ( .A(n3175), .B(n3176), .Z(n3188) );
  NAND U3749 ( .A(n1268), .B(n1974), .Z(n3176) );
  XNOR U3750 ( .A(n3174), .B(n3240), .Z(n3175) );
  AND U3751 ( .A(n2075), .B(n1200), .Z(n3240) );
  XNOR U3752 ( .A(n3187), .B(n3177), .Z(n3239) );
  XNOR U3753 ( .A(n3182), .B(n3248), .Z(n3183) );
  AND U3754 ( .A(n2304), .B(n1077), .Z(n3248) );
  XOR U3755 ( .A(n3252), .B(n3184), .Z(n3247) );
  NAND U3756 ( .A(n1137), .B(n2190), .Z(n3184) );
  IV U3757 ( .A(n3186), .Z(n3252) );
  XOR U3758 ( .A(n3256), .B(n3257), .Z(n3218) );
  AND U3759 ( .A(n3258), .B(n3259), .Z(n3257) );
  XNOR U3760 ( .A(n3260), .B(n3261), .Z(n3259) );
  XNOR U3761 ( .A(n3256), .B(n3262), .Z(n3261) );
  XOR U3762 ( .A(n3245), .B(n3263), .Z(n3258) );
  XNOR U3763 ( .A(n3256), .B(n3246), .Z(n3263) );
  XNOR U3764 ( .A(n3228), .B(n3265), .Z(n3229) );
  AND U3765 ( .A(n1880), .B(n1412), .Z(n3265) );
  XOR U3766 ( .A(n3269), .B(n3230), .Z(n3264) );
  NAND U3767 ( .A(n1491), .B(n1781), .Z(n3230) );
  IV U3768 ( .A(n3232), .Z(n3269) );
  XNOR U3769 ( .A(n3237), .B(n3238), .Z(n3234) );
  NAND U3770 ( .A(n1596), .B(n1668), .Z(n3238) );
  XNOR U3771 ( .A(n3236), .B(n3273), .Z(n3237) );
  AND U3772 ( .A(n1576), .B(n1690), .Z(n3273) );
  XOR U3773 ( .A(n3277), .B(n3255), .Z(n3245) );
  XNOR U3774 ( .A(n3242), .B(n3243), .Z(n3255) );
  NAND U3775 ( .A(n1338), .B(n1974), .Z(n3243) );
  XNOR U3776 ( .A(n3241), .B(n3278), .Z(n3242) );
  AND U3777 ( .A(n2075), .B(n1268), .Z(n3278) );
  XNOR U3778 ( .A(n3254), .B(n3244), .Z(n3277) );
  XNOR U3779 ( .A(n3249), .B(n3286), .Z(n3250) );
  AND U3780 ( .A(n2304), .B(n1137), .Z(n3286) );
  XOR U3781 ( .A(n3290), .B(n3251), .Z(n3285) );
  NAND U3782 ( .A(n1200), .B(n2190), .Z(n3251) );
  IV U3783 ( .A(n3253), .Z(n3290) );
  XOR U3784 ( .A(n3294), .B(n3295), .Z(n3256) );
  AND U3785 ( .A(n3296), .B(n3297), .Z(n3295) );
  XNOR U3786 ( .A(n3298), .B(n3299), .Z(n3297) );
  XNOR U3787 ( .A(n3294), .B(n3300), .Z(n3299) );
  XOR U3788 ( .A(n3283), .B(n3301), .Z(n3296) );
  XNOR U3789 ( .A(n3294), .B(n3284), .Z(n3301) );
  XNOR U3790 ( .A(n3266), .B(n3303), .Z(n3267) );
  AND U3791 ( .A(n1880), .B(n1491), .Z(n3303) );
  XOR U3792 ( .A(n3307), .B(n3268), .Z(n3302) );
  NAND U3793 ( .A(n1781), .B(n1576), .Z(n3268) );
  IV U3794 ( .A(n3270), .Z(n3307) );
  XNOR U3795 ( .A(n3275), .B(n3276), .Z(n3272) );
  NAND U3796 ( .A(n1596), .B(n1761), .Z(n3276) );
  XNOR U3797 ( .A(n3274), .B(n3311), .Z(n3275) );
  AND U3798 ( .A(n1668), .B(n1690), .Z(n3311) );
  XOR U3799 ( .A(n3315), .B(n3293), .Z(n3283) );
  XNOR U3800 ( .A(n3280), .B(n3281), .Z(n3293) );
  NAND U3801 ( .A(n1412), .B(n1974), .Z(n3281) );
  XNOR U3802 ( .A(n3279), .B(n3316), .Z(n3280) );
  AND U3803 ( .A(n2075), .B(n1338), .Z(n3316) );
  XNOR U3804 ( .A(n3292), .B(n3282), .Z(n3315) );
  XNOR U3805 ( .A(n3287), .B(n3324), .Z(n3288) );
  AND U3806 ( .A(n2304), .B(n1200), .Z(n3324) );
  XOR U3807 ( .A(n3328), .B(n3289), .Z(n3323) );
  NAND U3808 ( .A(n1268), .B(n2190), .Z(n3289) );
  IV U3809 ( .A(n3291), .Z(n3328) );
  XOR U3810 ( .A(n3332), .B(n3333), .Z(n3294) );
  AND U3811 ( .A(n3334), .B(n3335), .Z(n3333) );
  XNOR U3812 ( .A(n3336), .B(n3337), .Z(n3335) );
  XNOR U3813 ( .A(n3332), .B(n3338), .Z(n3337) );
  XOR U3814 ( .A(n3321), .B(n3339), .Z(n3334) );
  XNOR U3815 ( .A(n3332), .B(n3322), .Z(n3339) );
  XNOR U3816 ( .A(n3304), .B(n3341), .Z(n3305) );
  AND U3817 ( .A(n1576), .B(n1880), .Z(n3341) );
  XOR U3818 ( .A(n3345), .B(n3306), .Z(n3340) );
  NAND U3819 ( .A(n1781), .B(n1668), .Z(n3306) );
  IV U3820 ( .A(n3308), .Z(n3345) );
  XNOR U3821 ( .A(n3313), .B(n3314), .Z(n3310) );
  NAND U3822 ( .A(n1596), .B(n1856), .Z(n3314) );
  XNOR U3823 ( .A(n3312), .B(n3349), .Z(n3313) );
  AND U3824 ( .A(n1761), .B(n1690), .Z(n3349) );
  XOR U3825 ( .A(n3353), .B(n3331), .Z(n3321) );
  XNOR U3826 ( .A(n3318), .B(n3319), .Z(n3331) );
  NAND U3827 ( .A(n1491), .B(n1974), .Z(n3319) );
  XNOR U3828 ( .A(n3317), .B(n3354), .Z(n3318) );
  AND U3829 ( .A(n2075), .B(n1412), .Z(n3354) );
  XNOR U3830 ( .A(n3330), .B(n3320), .Z(n3353) );
  XNOR U3831 ( .A(n3325), .B(n3362), .Z(n3326) );
  AND U3832 ( .A(n2304), .B(n1268), .Z(n3362) );
  XOR U3833 ( .A(n3366), .B(n3327), .Z(n3361) );
  NAND U3834 ( .A(n1338), .B(n2190), .Z(n3327) );
  IV U3835 ( .A(n3329), .Z(n3366) );
  XOR U3836 ( .A(n3370), .B(n3371), .Z(n3332) );
  AND U3837 ( .A(n3372), .B(n3373), .Z(n3371) );
  XNOR U3838 ( .A(n3374), .B(n3375), .Z(n3373) );
  XNOR U3839 ( .A(n3370), .B(n3376), .Z(n3375) );
  XOR U3840 ( .A(n3359), .B(n3377), .Z(n3372) );
  XNOR U3841 ( .A(n3370), .B(n3360), .Z(n3377) );
  XNOR U3842 ( .A(n3342), .B(n3379), .Z(n3343) );
  AND U3843 ( .A(n1668), .B(n1880), .Z(n3379) );
  XOR U3844 ( .A(n3383), .B(n3344), .Z(n3378) );
  NAND U3845 ( .A(n1781), .B(n1761), .Z(n3344) );
  IV U3846 ( .A(n3346), .Z(n3383) );
  XNOR U3847 ( .A(n3351), .B(n3352), .Z(n3348) );
  NAND U3848 ( .A(n1596), .B(n1953), .Z(n3352) );
  XNOR U3849 ( .A(n3350), .B(n3387), .Z(n3351) );
  AND U3850 ( .A(n1856), .B(n1690), .Z(n3387) );
  XOR U3851 ( .A(n3391), .B(n3369), .Z(n3359) );
  XNOR U3852 ( .A(n3356), .B(n3357), .Z(n3369) );
  NAND U3853 ( .A(n1974), .B(n1576), .Z(n3357) );
  XNOR U3854 ( .A(n3355), .B(n3392), .Z(n3356) );
  AND U3855 ( .A(n2075), .B(n1491), .Z(n3392) );
  XNOR U3856 ( .A(n3368), .B(n3358), .Z(n3391) );
  XNOR U3857 ( .A(n3363), .B(n3400), .Z(n3364) );
  AND U3858 ( .A(n2304), .B(n1338), .Z(n3400) );
  XOR U3859 ( .A(n3404), .B(n3365), .Z(n3399) );
  NAND U3860 ( .A(n1412), .B(n2190), .Z(n3365) );
  IV U3861 ( .A(n3367), .Z(n3404) );
  XOR U3862 ( .A(n3408), .B(n3409), .Z(n3370) );
  AND U3863 ( .A(n3410), .B(n3411), .Z(n3409) );
  XNOR U3864 ( .A(n3412), .B(n3413), .Z(n3411) );
  XNOR U3865 ( .A(n3408), .B(n3414), .Z(n3413) );
  XOR U3866 ( .A(n3397), .B(n3415), .Z(n3410) );
  XNOR U3867 ( .A(n3408), .B(n3398), .Z(n3415) );
  XNOR U3868 ( .A(n3380), .B(n3417), .Z(n3381) );
  AND U3869 ( .A(n1761), .B(n1880), .Z(n3417) );
  XOR U3870 ( .A(n3421), .B(n3382), .Z(n3416) );
  NAND U3871 ( .A(n1781), .B(n1856), .Z(n3382) );
  IV U3872 ( .A(n3384), .Z(n3421) );
  XNOR U3873 ( .A(n3389), .B(n3390), .Z(n3386) );
  NAND U3874 ( .A(n1596), .B(n2058), .Z(n3390) );
  XNOR U3875 ( .A(n3388), .B(n3425), .Z(n3389) );
  AND U3876 ( .A(n1953), .B(n1690), .Z(n3425) );
  XOR U3877 ( .A(n3429), .B(n3407), .Z(n3397) );
  XNOR U3878 ( .A(n3394), .B(n3395), .Z(n3407) );
  NAND U3879 ( .A(n1974), .B(n1668), .Z(n3395) );
  XNOR U3880 ( .A(n3393), .B(n3430), .Z(n3394) );
  AND U3881 ( .A(n1576), .B(n2075), .Z(n3430) );
  XNOR U3882 ( .A(n3406), .B(n3396), .Z(n3429) );
  XNOR U3883 ( .A(n3401), .B(n3438), .Z(n3402) );
  AND U3884 ( .A(n2304), .B(n1412), .Z(n3438) );
  XOR U3885 ( .A(n3442), .B(n3403), .Z(n3437) );
  NAND U3886 ( .A(n1491), .B(n2190), .Z(n3403) );
  IV U3887 ( .A(n3405), .Z(n3442) );
  XOR U3888 ( .A(n3446), .B(n3447), .Z(n3408) );
  AND U3889 ( .A(n3448), .B(n3449), .Z(n3447) );
  XNOR U3890 ( .A(n3450), .B(n3451), .Z(n3449) );
  XNOR U3891 ( .A(n3446), .B(n3452), .Z(n3451) );
  XOR U3892 ( .A(n3435), .B(n3453), .Z(n3448) );
  XNOR U3893 ( .A(n3446), .B(n3436), .Z(n3453) );
  XNOR U3894 ( .A(n3418), .B(n3455), .Z(n3419) );
  AND U3895 ( .A(n1856), .B(n1880), .Z(n3455) );
  XOR U3896 ( .A(n3459), .B(n3420), .Z(n3454) );
  NAND U3897 ( .A(n1781), .B(n1953), .Z(n3420) );
  IV U3898 ( .A(n3422), .Z(n3459) );
  XNOR U3899 ( .A(n3427), .B(n3428), .Z(n3424) );
  NAND U3900 ( .A(n1596), .B(n2165), .Z(n3428) );
  XNOR U3901 ( .A(n3426), .B(n3463), .Z(n3427) );
  AND U3902 ( .A(n2058), .B(n1690), .Z(n3463) );
  XOR U3903 ( .A(n3467), .B(n3445), .Z(n3435) );
  XNOR U3904 ( .A(n3432), .B(n3433), .Z(n3445) );
  NAND U3905 ( .A(n1974), .B(n1761), .Z(n3433) );
  XNOR U3906 ( .A(n3431), .B(n3468), .Z(n3432) );
  AND U3907 ( .A(n1668), .B(n2075), .Z(n3468) );
  XNOR U3908 ( .A(n3444), .B(n3434), .Z(n3467) );
  XNOR U3909 ( .A(n3439), .B(n3476), .Z(n3440) );
  AND U3910 ( .A(n2304), .B(n1491), .Z(n3476) );
  XOR U3911 ( .A(n3480), .B(n3441), .Z(n3475) );
  NAND U3912 ( .A(n2190), .B(n1576), .Z(n3441) );
  IV U3913 ( .A(n3443), .Z(n3480) );
  XOR U3914 ( .A(n3484), .B(n3485), .Z(n3446) );
  AND U3915 ( .A(n3486), .B(n3487), .Z(n3485) );
  XNOR U3916 ( .A(n3488), .B(n3489), .Z(n3487) );
  XNOR U3917 ( .A(n3484), .B(n3490), .Z(n3489) );
  XOR U3918 ( .A(n3473), .B(n3491), .Z(n3486) );
  XNOR U3919 ( .A(n3484), .B(n3474), .Z(n3491) );
  XNOR U3920 ( .A(n3456), .B(n3493), .Z(n3457) );
  AND U3921 ( .A(n1953), .B(n1880), .Z(n3493) );
  XOR U3922 ( .A(n3497), .B(n3458), .Z(n3492) );
  NAND U3923 ( .A(n1781), .B(n2058), .Z(n3458) );
  IV U3924 ( .A(n3460), .Z(n3497) );
  XNOR U3925 ( .A(n3465), .B(n3466), .Z(n3462) );
  NAND U3926 ( .A(n1596), .B(n2276), .Z(n3466) );
  XNOR U3927 ( .A(n3464), .B(n3501), .Z(n3465) );
  AND U3928 ( .A(n2165), .B(n1690), .Z(n3501) );
  XOR U3929 ( .A(n3505), .B(n3483), .Z(n3473) );
  XNOR U3930 ( .A(n3470), .B(n3471), .Z(n3483) );
  NAND U3931 ( .A(n1974), .B(n1856), .Z(n3471) );
  XNOR U3932 ( .A(n3469), .B(n3506), .Z(n3470) );
  AND U3933 ( .A(n1761), .B(n2075), .Z(n3506) );
  XNOR U3934 ( .A(n3482), .B(n3472), .Z(n3505) );
  XNOR U3935 ( .A(n3477), .B(n3514), .Z(n3478) );
  AND U3936 ( .A(n1576), .B(n2304), .Z(n3514) );
  XOR U3937 ( .A(n3518), .B(n3479), .Z(n3513) );
  NAND U3938 ( .A(n2190), .B(n1668), .Z(n3479) );
  IV U3939 ( .A(n3481), .Z(n3518) );
  XOR U3940 ( .A(n3522), .B(n3523), .Z(n3484) );
  AND U3941 ( .A(n3524), .B(n3525), .Z(n3523) );
  XNOR U3942 ( .A(n3526), .B(n3527), .Z(n3525) );
  XNOR U3943 ( .A(n3522), .B(n3528), .Z(n3527) );
  XOR U3944 ( .A(n3511), .B(n3529), .Z(n3524) );
  XNOR U3945 ( .A(n3522), .B(n3512), .Z(n3529) );
  XNOR U3946 ( .A(n3494), .B(n3531), .Z(n3495) );
  AND U3947 ( .A(n2058), .B(n1880), .Z(n3531) );
  XOR U3948 ( .A(n3535), .B(n3496), .Z(n3530) );
  NAND U3949 ( .A(n1781), .B(n2165), .Z(n3496) );
  IV U3950 ( .A(n3498), .Z(n3535) );
  XNOR U3951 ( .A(n3503), .B(n3504), .Z(n3500) );
  NAND U3952 ( .A(n1596), .B(n2392), .Z(n3504) );
  XNOR U3953 ( .A(n3502), .B(n3539), .Z(n3503) );
  AND U3954 ( .A(n2276), .B(n1690), .Z(n3539) );
  XOR U3955 ( .A(n3543), .B(n3521), .Z(n3511) );
  XNOR U3956 ( .A(n3508), .B(n3509), .Z(n3521) );
  NAND U3957 ( .A(n1974), .B(n1953), .Z(n3509) );
  XNOR U3958 ( .A(n3507), .B(n3544), .Z(n3508) );
  AND U3959 ( .A(n1856), .B(n2075), .Z(n3544) );
  XNOR U3960 ( .A(n3520), .B(n3510), .Z(n3543) );
  XNOR U3961 ( .A(n3515), .B(n3552), .Z(n3516) );
  AND U3962 ( .A(n1668), .B(n2304), .Z(n3552) );
  XOR U3963 ( .A(n3556), .B(n3517), .Z(n3551) );
  NAND U3964 ( .A(n2190), .B(n1761), .Z(n3517) );
  IV U3965 ( .A(n3519), .Z(n3556) );
  XOR U3966 ( .A(n3560), .B(n3561), .Z(n3522) );
  AND U3967 ( .A(n3562), .B(n3563), .Z(n3561) );
  XNOR U3968 ( .A(n3564), .B(n3565), .Z(n3563) );
  XNOR U3969 ( .A(n3560), .B(n3566), .Z(n3565) );
  XOR U3970 ( .A(n3549), .B(n3567), .Z(n3562) );
  XNOR U3971 ( .A(n3560), .B(n3550), .Z(n3567) );
  XNOR U3972 ( .A(n3532), .B(n3569), .Z(n3533) );
  AND U3973 ( .A(n2165), .B(n1880), .Z(n3569) );
  XOR U3974 ( .A(n3573), .B(n3534), .Z(n3568) );
  NAND U3975 ( .A(n1781), .B(n2276), .Z(n3534) );
  IV U3976 ( .A(n3536), .Z(n3573) );
  XNOR U3977 ( .A(n3541), .B(n3542), .Z(n3538) );
  NAND U3978 ( .A(n1596), .B(n2513), .Z(n3542) );
  XNOR U3979 ( .A(n3540), .B(n3577), .Z(n3541) );
  AND U3980 ( .A(n2392), .B(n1690), .Z(n3577) );
  XOR U3981 ( .A(n3581), .B(n3559), .Z(n3549) );
  XNOR U3982 ( .A(n3546), .B(n3547), .Z(n3559) );
  NAND U3983 ( .A(n1974), .B(n2058), .Z(n3547) );
  XNOR U3984 ( .A(n3545), .B(n3582), .Z(n3546) );
  AND U3985 ( .A(n1953), .B(n2075), .Z(n3582) );
  XNOR U3986 ( .A(n3558), .B(n3548), .Z(n3581) );
  XNOR U3987 ( .A(n3553), .B(n3590), .Z(n3554) );
  AND U3988 ( .A(n1761), .B(n2304), .Z(n3590) );
  XOR U3989 ( .A(n3594), .B(n3555), .Z(n3589) );
  NAND U3990 ( .A(n2190), .B(n1856), .Z(n3555) );
  IV U3991 ( .A(n3557), .Z(n3594) );
  XOR U3992 ( .A(n3598), .B(n3599), .Z(n3560) );
  AND U3993 ( .A(n3600), .B(n3601), .Z(n3599) );
  XNOR U3994 ( .A(n3602), .B(n3603), .Z(n3601) );
  XNOR U3995 ( .A(n3598), .B(n3604), .Z(n3603) );
  XOR U3996 ( .A(n3587), .B(n3605), .Z(n3600) );
  XNOR U3997 ( .A(n3598), .B(n3588), .Z(n3605) );
  XNOR U3998 ( .A(n3570), .B(n3607), .Z(n3571) );
  AND U3999 ( .A(n2276), .B(n1880), .Z(n3607) );
  XOR U4000 ( .A(n3611), .B(n3572), .Z(n3606) );
  NAND U4001 ( .A(n1781), .B(n2392), .Z(n3572) );
  IV U4002 ( .A(n3574), .Z(n3611) );
  XNOR U4003 ( .A(n3579), .B(n3580), .Z(n3576) );
  NAND U4004 ( .A(n1596), .B(n2635), .Z(n3580) );
  XNOR U4005 ( .A(n3578), .B(n3615), .Z(n3579) );
  AND U4006 ( .A(n2513), .B(n1690), .Z(n3615) );
  XOR U4007 ( .A(n3619), .B(n3597), .Z(n3587) );
  XNOR U4008 ( .A(n3584), .B(n3585), .Z(n3597) );
  NAND U4009 ( .A(n1974), .B(n2165), .Z(n3585) );
  XNOR U4010 ( .A(n3583), .B(n3620), .Z(n3584) );
  AND U4011 ( .A(n2058), .B(n2075), .Z(n3620) );
  XNOR U4012 ( .A(n3596), .B(n3586), .Z(n3619) );
  XNOR U4013 ( .A(n3591), .B(n3628), .Z(n3592) );
  AND U4014 ( .A(n1856), .B(n2304), .Z(n3628) );
  XOR U4015 ( .A(n3632), .B(n3593), .Z(n3627) );
  NAND U4016 ( .A(n2190), .B(n1953), .Z(n3593) );
  IV U4017 ( .A(n3595), .Z(n3632) );
  XOR U4018 ( .A(n3636), .B(n3637), .Z(n3598) );
  AND U4019 ( .A(n3638), .B(n3639), .Z(n3637) );
  XNOR U4020 ( .A(n3640), .B(n3641), .Z(n3639) );
  XNOR U4021 ( .A(n3636), .B(n3642), .Z(n3641) );
  XOR U4022 ( .A(n3625), .B(n3643), .Z(n3638) );
  XNOR U4023 ( .A(n3636), .B(n3626), .Z(n3643) );
  XNOR U4024 ( .A(n3608), .B(n3645), .Z(n3609) );
  AND U4025 ( .A(n2392), .B(n1880), .Z(n3645) );
  XOR U4026 ( .A(n3649), .B(n3610), .Z(n3644) );
  NAND U4027 ( .A(n1781), .B(n2513), .Z(n3610) );
  IV U4028 ( .A(n3612), .Z(n3649) );
  XNOR U4029 ( .A(n3617), .B(n3618), .Z(n3614) );
  NAND U4030 ( .A(n1596), .B(n2763), .Z(n3618) );
  XNOR U4031 ( .A(n3616), .B(n3653), .Z(n3617) );
  AND U4032 ( .A(n2635), .B(n1690), .Z(n3653) );
  XOR U4033 ( .A(n3657), .B(n3635), .Z(n3625) );
  XNOR U4034 ( .A(n3622), .B(n3623), .Z(n3635) );
  NAND U4035 ( .A(n1974), .B(n2276), .Z(n3623) );
  XNOR U4036 ( .A(n3621), .B(n3658), .Z(n3622) );
  AND U4037 ( .A(n2165), .B(n2075), .Z(n3658) );
  XNOR U4038 ( .A(n3634), .B(n3624), .Z(n3657) );
  XNOR U4039 ( .A(n3629), .B(n3666), .Z(n3630) );
  AND U4040 ( .A(n1953), .B(n2304), .Z(n3666) );
  XOR U4041 ( .A(n3670), .B(n3631), .Z(n3665) );
  NAND U4042 ( .A(n2190), .B(n2058), .Z(n3631) );
  IV U4043 ( .A(n3633), .Z(n3670) );
  XOR U4044 ( .A(n3674), .B(n3675), .Z(n3636) );
  AND U4045 ( .A(n3676), .B(n3677), .Z(n3675) );
  XNOR U4046 ( .A(n3678), .B(n3679), .Z(n3677) );
  XNOR U4047 ( .A(n3674), .B(n3680), .Z(n3679) );
  XOR U4048 ( .A(n3663), .B(n3681), .Z(n3676) );
  XNOR U4049 ( .A(n3674), .B(n3664), .Z(n3681) );
  XNOR U4050 ( .A(n3646), .B(n3683), .Z(n3647) );
  AND U4051 ( .A(n2513), .B(n1880), .Z(n3683) );
  XOR U4052 ( .A(n3687), .B(n3648), .Z(n3682) );
  NAND U4053 ( .A(n1781), .B(n2635), .Z(n3648) );
  IV U4054 ( .A(n3650), .Z(n3687) );
  XNOR U4055 ( .A(n3655), .B(n3656), .Z(n3652) );
  NANDN U4056 ( .B(n2892), .A(n1596), .Z(n3656) );
  XNOR U4057 ( .A(n3654), .B(n3691), .Z(n3655) );
  AND U4058 ( .A(n2763), .B(n1690), .Z(n3691) );
  XOR U4059 ( .A(n3695), .B(n3673), .Z(n3663) );
  XNOR U4060 ( .A(n3660), .B(n3661), .Z(n3673) );
  NAND U4061 ( .A(n1974), .B(n2392), .Z(n3661) );
  XNOR U4062 ( .A(n3659), .B(n3696), .Z(n3660) );
  AND U4063 ( .A(n2276), .B(n2075), .Z(n3696) );
  XNOR U4064 ( .A(n3672), .B(n3662), .Z(n3695) );
  XNOR U4065 ( .A(n3667), .B(n3704), .Z(n3668) );
  AND U4066 ( .A(n2058), .B(n2304), .Z(n3704) );
  XOR U4067 ( .A(n3708), .B(n3669), .Z(n3703) );
  NAND U4068 ( .A(n2190), .B(n2165), .Z(n3669) );
  IV U4069 ( .A(n3671), .Z(n3708) );
  XOR U4070 ( .A(n3712), .B(n3713), .Z(n3674) );
  AND U4071 ( .A(n3714), .B(n3715), .Z(n3713) );
  XNOR U4072 ( .A(n3716), .B(n3717), .Z(n3715) );
  XNOR U4073 ( .A(n3712), .B(n3718), .Z(n3717) );
  XOR U4074 ( .A(n3701), .B(n3719), .Z(n3714) );
  XNOR U4075 ( .A(n3712), .B(n3702), .Z(n3719) );
  XNOR U4076 ( .A(n3684), .B(n3721), .Z(n3685) );
  AND U4077 ( .A(n2635), .B(n1880), .Z(n3721) );
  XOR U4078 ( .A(n3725), .B(n3686), .Z(n3720) );
  NAND U4079 ( .A(n1781), .B(n2763), .Z(n3686) );
  IV U4080 ( .A(n3688), .Z(n3725) );
  XNOR U4081 ( .A(n3693), .B(n3694), .Z(n3690) );
  NANDN U4082 ( .B(n3030), .A(n1596), .Z(n3694) );
  XNOR U4083 ( .A(n3692), .B(n3729), .Z(n3693) );
  ANDN U4084 ( .A(n1690), .B(n2892), .Z(n3729) );
  XOR U4085 ( .A(n3733), .B(n3711), .Z(n3701) );
  XNOR U4086 ( .A(n3698), .B(n3699), .Z(n3711) );
  NAND U4087 ( .A(n1974), .B(n2513), .Z(n3699) );
  XNOR U4088 ( .A(n3697), .B(n3734), .Z(n3698) );
  AND U4089 ( .A(n2392), .B(n2075), .Z(n3734) );
  XNOR U4090 ( .A(n3710), .B(n3700), .Z(n3733) );
  XNOR U4091 ( .A(n3705), .B(n3742), .Z(n3706) );
  AND U4092 ( .A(n2165), .B(n2304), .Z(n3742) );
  XOR U4093 ( .A(n3746), .B(n3707), .Z(n3741) );
  NAND U4094 ( .A(n2190), .B(n2276), .Z(n3707) );
  IV U4095 ( .A(n3709), .Z(n3746) );
  XOR U4096 ( .A(n3750), .B(n3751), .Z(n3712) );
  AND U4097 ( .A(n3752), .B(n3753), .Z(n3751) );
  XNOR U4098 ( .A(n3754), .B(n3755), .Z(n3753) );
  XNOR U4099 ( .A(n3750), .B(n3756), .Z(n3755) );
  XOR U4100 ( .A(n3739), .B(n3757), .Z(n3752) );
  XNOR U4101 ( .A(n3750), .B(n3740), .Z(n3757) );
  XNOR U4102 ( .A(n3722), .B(n3759), .Z(n3723) );
  AND U4103 ( .A(n2763), .B(n1880), .Z(n3759) );
  XOR U4104 ( .A(n3763), .B(n3724), .Z(n3758) );
  NANDN U4105 ( .B(n2892), .A(n1781), .Z(n3724) );
  IV U4106 ( .A(n3726), .Z(n3763) );
  XNOR U4107 ( .A(n3731), .B(n3732), .Z(n3728) );
  NAND U4108 ( .A(n1596), .B(n3165), .Z(n3732) );
  XNOR U4109 ( .A(n3730), .B(n3767), .Z(n3731) );
  ANDN U4110 ( .A(n1690), .B(n3030), .Z(n3767) );
  XOR U4111 ( .A(n3771), .B(n3749), .Z(n3739) );
  XNOR U4112 ( .A(n3736), .B(n3737), .Z(n3749) );
  NAND U4113 ( .A(n1974), .B(n2635), .Z(n3737) );
  XNOR U4114 ( .A(n3735), .B(n3772), .Z(n3736) );
  AND U4115 ( .A(n2513), .B(n2075), .Z(n3772) );
  XNOR U4116 ( .A(n3748), .B(n3738), .Z(n3771) );
  XNOR U4117 ( .A(n3743), .B(n3780), .Z(n3744) );
  AND U4118 ( .A(n2276), .B(n2304), .Z(n3780) );
  XOR U4119 ( .A(n3784), .B(n3745), .Z(n3779) );
  NAND U4120 ( .A(n2190), .B(n2392), .Z(n3745) );
  IV U4121 ( .A(n3747), .Z(n3784) );
  XNOR U4122 ( .A(n3789), .B(n3790), .Z(n3203) );
  XOR U4123 ( .A(n3791), .B(n3788), .Z(n3789) );
  XNOR U4124 ( .A(n3792), .B(n3787), .Z(n3777) );
  XNOR U4125 ( .A(n3774), .B(n3775), .Z(n3787) );
  NAND U4126 ( .A(n1974), .B(n2763), .Z(n3775) );
  XNOR U4127 ( .A(n3773), .B(n3793), .Z(n3774) );
  AND U4128 ( .A(n2635), .B(n2075), .Z(n3793) );
  XNOR U4129 ( .A(n3797), .B(n3794), .Z(n3796) );
  XNOR U4130 ( .A(n3786), .B(n3776), .Z(n3792) );
  XOR U4131 ( .A(n3798), .B(n3799), .Z(n3776) );
  XNOR U4132 ( .A(n3781), .B(n3801), .Z(n3782) );
  AND U4133 ( .A(n2392), .B(n2304), .Z(n3801) );
  XNOR U4134 ( .A(n3805), .B(n3802), .Z(n3804) );
  XOR U4135 ( .A(n3806), .B(n3783), .Z(n3800) );
  NAND U4136 ( .A(n2190), .B(n2513), .Z(n3783) );
  IV U4137 ( .A(n3785), .Z(n3806) );
  XNOR U4138 ( .A(n3807), .B(n3808), .Z(n3785) );
  AND U4139 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U4140 ( .A(n3803), .B(n3811), .Z(n3810) );
  XNOR U4141 ( .A(n3805), .B(n3807), .Z(n3811) );
  NAND U4142 ( .A(n2190), .B(n2635), .Z(n3805) );
  XOR U4143 ( .A(n3802), .B(n3812), .Z(n3803) );
  AND U4144 ( .A(n2513), .B(n2304), .Z(n3812) );
  XNOR U4145 ( .A(n3816), .B(n3813), .Z(n3815) );
  XOR U4146 ( .A(n3795), .B(n3817), .Z(n3809) );
  XNOR U4147 ( .A(n3797), .B(n3807), .Z(n3817) );
  NANDN U4148 ( .B(n2892), .A(n1974), .Z(n3797) );
  XOR U4149 ( .A(n3794), .B(n3818), .Z(n3795) );
  AND U4150 ( .A(n2763), .B(n2075), .Z(n3818) );
  XNOR U4151 ( .A(n3822), .B(n3819), .Z(n3821) );
  XOR U4152 ( .A(n3823), .B(n3824), .Z(n3807) );
  AND U4153 ( .A(n3825), .B(n3826), .Z(n3824) );
  XOR U4154 ( .A(n3814), .B(n3827), .Z(n3826) );
  XNOR U4155 ( .A(n3816), .B(n3823), .Z(n3827) );
  NAND U4156 ( .A(n2190), .B(n2763), .Z(n3816) );
  XOR U4157 ( .A(n3813), .B(n3828), .Z(n3814) );
  AND U4158 ( .A(n2635), .B(n2304), .Z(n3828) );
  XNOR U4159 ( .A(n3832), .B(n3829), .Z(n3831) );
  XOR U4160 ( .A(n3820), .B(n3833), .Z(n3825) );
  XNOR U4161 ( .A(n3822), .B(n3823), .Z(n3833) );
  NANDN U4162 ( .B(n3030), .A(n1974), .Z(n3822) );
  XOR U4163 ( .A(n3819), .B(n3834), .Z(n3820) );
  ANDN U4164 ( .A(n2075), .B(n2892), .Z(n3834) );
  XNOR U4165 ( .A(n3838), .B(n3835), .Z(n3837) );
  XOR U4166 ( .A(n3839), .B(n3840), .Z(n3823) );
  AND U4167 ( .A(n3841), .B(n3842), .Z(n3840) );
  XOR U4168 ( .A(n3830), .B(n3843), .Z(n3842) );
  XNOR U4169 ( .A(n3832), .B(n3839), .Z(n3843) );
  NANDN U4170 ( .B(n2892), .A(n2190), .Z(n3832) );
  XOR U4171 ( .A(n3829), .B(n3844), .Z(n3830) );
  AND U4172 ( .A(n2763), .B(n2304), .Z(n3844) );
  XOR U4173 ( .A(n3836), .B(n3848), .Z(n3841) );
  XNOR U4174 ( .A(n3838), .B(n3839), .Z(n3848) );
  NAND U4175 ( .A(n1974), .B(n3165), .Z(n3838) );
  XOR U4176 ( .A(n3835), .B(n3849), .Z(n3836) );
  ANDN U4177 ( .A(n2075), .B(n3030), .Z(n3849) );
  NAND U4178 ( .A(n1974), .B(n3854), .Z(n3852) );
  XNOR U4179 ( .A(n3850), .B(n3855), .Z(n3851) );
  AND U4180 ( .A(n3165), .B(n2075), .Z(n3855) );
  AND U4181 ( .A(n3856), .B(\_MAC/_MULT/A__[0] ), .Z(n3850) );
  NANDN U4182 ( .B(n1974), .A(n3857), .Z(n3856) );
  NAND U4183 ( .A(n3854), .B(n2075), .Z(n3857) );
  XNOR U4184 ( .A(n3845), .B(n3861), .Z(n3846) );
  ANDN U4185 ( .A(n2304), .B(n2892), .Z(n3861) );
  XOR U4186 ( .A(n3864), .B(n3862), .Z(n3863) );
  ANDN U4187 ( .A(n2304), .B(n3030), .Z(n3864) );
  AND U4188 ( .A(n3165), .B(n2190), .Z(n3865) );
  XOR U4189 ( .A(n3869), .B(n3847), .Z(n3860) );
  NANDN U4190 ( .B(n3030), .A(n2190), .Z(n3847) );
  IV U4191 ( .A(n3853), .Z(n3869) );
  NAND U4192 ( .A(n2190), .B(n3854), .Z(n3868) );
  XNOR U4193 ( .A(n3866), .B(n3870), .Z(n3867) );
  AND U4194 ( .A(n3165), .B(n2304), .Z(n3870) );
  AND U4195 ( .A(n3871), .B(\_MAC/_MULT/A__[0] ), .Z(n3866) );
  NANDN U4196 ( .B(n2190), .A(n3872), .Z(n3871) );
  NAND U4197 ( .A(n3854), .B(n2304), .Z(n3872) );
  XNOR U4198 ( .A(n3760), .B(n3876), .Z(n3761) );
  ANDN U4199 ( .A(n1880), .B(n2892), .Z(n3876) );
  XOR U4200 ( .A(n3879), .B(n3877), .Z(n3878) );
  ANDN U4201 ( .A(n1880), .B(n3030), .Z(n3879) );
  AND U4202 ( .A(n3165), .B(n1781), .Z(n3880) );
  XOR U4203 ( .A(n3884), .B(n3762), .Z(n3875) );
  NANDN U4204 ( .B(n3030), .A(n1781), .Z(n3762) );
  IV U4205 ( .A(n3764), .Z(n3884) );
  NAND U4206 ( .A(n1781), .B(n3854), .Z(n3883) );
  XNOR U4207 ( .A(n3881), .B(n3885), .Z(n3882) );
  AND U4208 ( .A(n3165), .B(n1880), .Z(n3885) );
  AND U4209 ( .A(n3886), .B(\_MAC/_MULT/A__[0] ), .Z(n3881) );
  NANDN U4210 ( .B(n1781), .A(n3887), .Z(n3886) );
  NAND U4211 ( .A(n3854), .B(n1880), .Z(n3887) );
  XNOR U4212 ( .A(n3769), .B(n3770), .Z(n3766) );
  NAND U4213 ( .A(n1596), .B(n3854), .Z(n3770) );
  XNOR U4214 ( .A(n3768), .B(n3890), .Z(n3769) );
  AND U4215 ( .A(n3165), .B(n1690), .Z(n3890) );
  AND U4216 ( .A(n3891), .B(\_MAC/_MULT/A__[0] ), .Z(n3768) );
  NANDN U4217 ( .B(n1596), .A(n3892), .Z(n3891) );
  NAND U4218 ( .A(n3854), .B(n1690), .Z(n3892) );
  XOR U4219 ( .A(n3895), .B(n3896), .Z(n3788) );
  XNOR U4220 ( .A(n3897), .B(n3104), .Z(n3101) );
  NAND U4221 ( .A(n797), .B(n2964), .Z(n3099) );
  XNOR U4222 ( .A(n3097), .B(n3898), .Z(n3098) );
  AND U4223 ( .A(n3096), .B(n765), .Z(n3898) );
  XNOR U4224 ( .A(n3103), .B(n3100), .Z(n3897) );
  XNOR U4225 ( .A(n3207), .B(n3904), .Z(n3208) );
  AND U4226 ( .A(n2818), .B(n875), .Z(n3904) );
  XOR U4227 ( .A(n3908), .B(n3209), .Z(n3903) );
  NAND U4228 ( .A(n917), .B(n2688), .Z(n3209) );
  IV U4229 ( .A(n3211), .Z(n3908) );
  XNOR U4230 ( .A(n3216), .B(n3217), .Z(n3213) );
  NAND U4231 ( .A(n1019), .B(n2443), .Z(n3217) );
  XNOR U4232 ( .A(n3215), .B(n3912), .Z(n3216) );
  AND U4233 ( .A(n2566), .B(n961), .Z(n3912) );
  XOR U4234 ( .A(n3916), .B(n3917), .Z(n3224) );
  XNOR U4235 ( .A(n3918), .B(n3902), .Z(n3916) );
  XOR U4236 ( .A(n3920), .B(n3921), .Z(n3262) );
  XNOR U4237 ( .A(n3922), .B(n3919), .Z(n3920) );
  XNOR U4238 ( .A(n3905), .B(n3924), .Z(n3906) );
  AND U4239 ( .A(n2818), .B(n917), .Z(n3924) );
  XOR U4240 ( .A(n3928), .B(n3907), .Z(n3923) );
  NAND U4241 ( .A(n961), .B(n2688), .Z(n3907) );
  IV U4242 ( .A(n3909), .Z(n3928) );
  XNOR U4243 ( .A(n3914), .B(n3915), .Z(n3911) );
  NAND U4244 ( .A(n1077), .B(n2443), .Z(n3915) );
  XNOR U4245 ( .A(n3913), .B(n3932), .Z(n3914) );
  AND U4246 ( .A(n2566), .B(n1019), .Z(n3932) );
  XOR U4247 ( .A(n3937), .B(n3938), .Z(n3300) );
  XNOR U4248 ( .A(n3939), .B(n3936), .Z(n3937) );
  XNOR U4249 ( .A(n3925), .B(n3941), .Z(n3926) );
  AND U4250 ( .A(n2818), .B(n961), .Z(n3941) );
  XOR U4251 ( .A(n3945), .B(n3927), .Z(n3940) );
  NAND U4252 ( .A(n1019), .B(n2688), .Z(n3927) );
  IV U4253 ( .A(n3929), .Z(n3945) );
  XNOR U4254 ( .A(n3934), .B(n3935), .Z(n3931) );
  NAND U4255 ( .A(n1137), .B(n2443), .Z(n3935) );
  XNOR U4256 ( .A(n3933), .B(n3949), .Z(n3934) );
  AND U4257 ( .A(n2566), .B(n1077), .Z(n3949) );
  XOR U4258 ( .A(n3954), .B(n3955), .Z(n3338) );
  XNOR U4259 ( .A(n3956), .B(n3953), .Z(n3954) );
  XNOR U4260 ( .A(n3942), .B(n3958), .Z(n3943) );
  AND U4261 ( .A(n2818), .B(n1019), .Z(n3958) );
  XOR U4262 ( .A(n3962), .B(n3944), .Z(n3957) );
  NAND U4263 ( .A(n1077), .B(n2688), .Z(n3944) );
  IV U4264 ( .A(n3946), .Z(n3962) );
  XNOR U4265 ( .A(n3951), .B(n3952), .Z(n3948) );
  NAND U4266 ( .A(n1200), .B(n2443), .Z(n3952) );
  XNOR U4267 ( .A(n3950), .B(n3966), .Z(n3951) );
  AND U4268 ( .A(n2566), .B(n1137), .Z(n3966) );
  XOR U4269 ( .A(n3971), .B(n3972), .Z(n3376) );
  XNOR U4270 ( .A(n3973), .B(n3970), .Z(n3971) );
  XNOR U4271 ( .A(n3959), .B(n3975), .Z(n3960) );
  AND U4272 ( .A(n2818), .B(n1077), .Z(n3975) );
  XOR U4273 ( .A(n3979), .B(n3961), .Z(n3974) );
  NAND U4274 ( .A(n1137), .B(n2688), .Z(n3961) );
  IV U4275 ( .A(n3963), .Z(n3979) );
  XNOR U4276 ( .A(n3968), .B(n3969), .Z(n3965) );
  NAND U4277 ( .A(n1268), .B(n2443), .Z(n3969) );
  XNOR U4278 ( .A(n3967), .B(n3983), .Z(n3968) );
  AND U4279 ( .A(n2566), .B(n1200), .Z(n3983) );
  XOR U4280 ( .A(n3988), .B(n3989), .Z(n3414) );
  XNOR U4281 ( .A(n3990), .B(n3987), .Z(n3988) );
  XNOR U4282 ( .A(n3976), .B(n3992), .Z(n3977) );
  AND U4283 ( .A(n2818), .B(n1137), .Z(n3992) );
  XOR U4284 ( .A(n3996), .B(n3978), .Z(n3991) );
  NAND U4285 ( .A(n1200), .B(n2688), .Z(n3978) );
  IV U4286 ( .A(n3980), .Z(n3996) );
  XNOR U4287 ( .A(n3985), .B(n3986), .Z(n3982) );
  NAND U4288 ( .A(n1338), .B(n2443), .Z(n3986) );
  XNOR U4289 ( .A(n3984), .B(n4000), .Z(n3985) );
  AND U4290 ( .A(n2566), .B(n1268), .Z(n4000) );
  XOR U4291 ( .A(n4005), .B(n4006), .Z(n3452) );
  XNOR U4292 ( .A(n4007), .B(n4004), .Z(n4005) );
  XNOR U4293 ( .A(n3993), .B(n4009), .Z(n3994) );
  AND U4294 ( .A(n2818), .B(n1200), .Z(n4009) );
  XOR U4295 ( .A(n4013), .B(n3995), .Z(n4008) );
  NAND U4296 ( .A(n1268), .B(n2688), .Z(n3995) );
  IV U4297 ( .A(n3997), .Z(n4013) );
  XNOR U4298 ( .A(n4002), .B(n4003), .Z(n3999) );
  NAND U4299 ( .A(n1412), .B(n2443), .Z(n4003) );
  XNOR U4300 ( .A(n4001), .B(n4017), .Z(n4002) );
  AND U4301 ( .A(n2566), .B(n1338), .Z(n4017) );
  XOR U4302 ( .A(n4022), .B(n4023), .Z(n3490) );
  XNOR U4303 ( .A(n4024), .B(n4021), .Z(n4022) );
  XNOR U4304 ( .A(n4010), .B(n4026), .Z(n4011) );
  AND U4305 ( .A(n2818), .B(n1268), .Z(n4026) );
  XOR U4306 ( .A(n4030), .B(n4012), .Z(n4025) );
  NAND U4307 ( .A(n1338), .B(n2688), .Z(n4012) );
  IV U4308 ( .A(n4014), .Z(n4030) );
  XNOR U4309 ( .A(n4019), .B(n4020), .Z(n4016) );
  NAND U4310 ( .A(n1491), .B(n2443), .Z(n4020) );
  XNOR U4311 ( .A(n4018), .B(n4034), .Z(n4019) );
  AND U4312 ( .A(n2566), .B(n1412), .Z(n4034) );
  XOR U4313 ( .A(n4039), .B(n4040), .Z(n3528) );
  XNOR U4314 ( .A(n4041), .B(n4038), .Z(n4039) );
  XNOR U4315 ( .A(n4027), .B(n4043), .Z(n4028) );
  AND U4316 ( .A(n2818), .B(n1338), .Z(n4043) );
  XOR U4317 ( .A(n4047), .B(n4029), .Z(n4042) );
  NAND U4318 ( .A(n1412), .B(n2688), .Z(n4029) );
  IV U4319 ( .A(n4031), .Z(n4047) );
  XNOR U4320 ( .A(n4036), .B(n4037), .Z(n4033) );
  NAND U4321 ( .A(n1576), .B(n2443), .Z(n4037) );
  XNOR U4322 ( .A(n4035), .B(n4051), .Z(n4036) );
  AND U4323 ( .A(n2566), .B(n1491), .Z(n4051) );
  XOR U4324 ( .A(n4056), .B(n4057), .Z(n3566) );
  XNOR U4325 ( .A(n4058), .B(n4055), .Z(n4056) );
  XNOR U4326 ( .A(n4044), .B(n4060), .Z(n4045) );
  AND U4327 ( .A(n2818), .B(n1412), .Z(n4060) );
  XOR U4328 ( .A(n4064), .B(n4046), .Z(n4059) );
  NAND U4329 ( .A(n1491), .B(n2688), .Z(n4046) );
  IV U4330 ( .A(n4048), .Z(n4064) );
  XNOR U4331 ( .A(n4053), .B(n4054), .Z(n4050) );
  NAND U4332 ( .A(n1668), .B(n2443), .Z(n4054) );
  XNOR U4333 ( .A(n4052), .B(n4068), .Z(n4053) );
  AND U4334 ( .A(n2566), .B(n1576), .Z(n4068) );
  XOR U4335 ( .A(n4073), .B(n4074), .Z(n3604) );
  XNOR U4336 ( .A(n4075), .B(n4072), .Z(n4073) );
  XNOR U4337 ( .A(n4061), .B(n4077), .Z(n4062) );
  AND U4338 ( .A(n2818), .B(n1491), .Z(n4077) );
  XOR U4339 ( .A(n4081), .B(n4063), .Z(n4076) );
  NAND U4340 ( .A(n1576), .B(n2688), .Z(n4063) );
  IV U4341 ( .A(n4065), .Z(n4081) );
  XNOR U4342 ( .A(n4070), .B(n4071), .Z(n4067) );
  NAND U4343 ( .A(n1761), .B(n2443), .Z(n4071) );
  XNOR U4344 ( .A(n4069), .B(n4085), .Z(n4070) );
  AND U4345 ( .A(n2566), .B(n1668), .Z(n4085) );
  XOR U4346 ( .A(n4090), .B(n4091), .Z(n3642) );
  XNOR U4347 ( .A(n4092), .B(n4089), .Z(n4090) );
  XNOR U4348 ( .A(n4078), .B(n4094), .Z(n4079) );
  AND U4349 ( .A(n2818), .B(n1576), .Z(n4094) );
  XOR U4350 ( .A(n4098), .B(n4080), .Z(n4093) );
  NAND U4351 ( .A(n1668), .B(n2688), .Z(n4080) );
  IV U4352 ( .A(n4082), .Z(n4098) );
  XNOR U4353 ( .A(n4087), .B(n4088), .Z(n4084) );
  NAND U4354 ( .A(n1856), .B(n2443), .Z(n4088) );
  XNOR U4355 ( .A(n4086), .B(n4102), .Z(n4087) );
  AND U4356 ( .A(n2566), .B(n1761), .Z(n4102) );
  XOR U4357 ( .A(n4107), .B(n4108), .Z(n3680) );
  XNOR U4358 ( .A(n4109), .B(n4106), .Z(n4107) );
  XNOR U4359 ( .A(n4095), .B(n4111), .Z(n4096) );
  AND U4360 ( .A(n2818), .B(n1668), .Z(n4111) );
  XOR U4361 ( .A(n4115), .B(n4097), .Z(n4110) );
  NAND U4362 ( .A(n1761), .B(n2688), .Z(n4097) );
  IV U4363 ( .A(n4099), .Z(n4115) );
  XNOR U4364 ( .A(n4104), .B(n4105), .Z(n4101) );
  NAND U4365 ( .A(n1953), .B(n2443), .Z(n4105) );
  XNOR U4366 ( .A(n4103), .B(n4119), .Z(n4104) );
  AND U4367 ( .A(n2566), .B(n1856), .Z(n4119) );
  XOR U4368 ( .A(n4124), .B(n4125), .Z(n3718) );
  XNOR U4369 ( .A(n4126), .B(n4123), .Z(n4124) );
  XNOR U4370 ( .A(n4112), .B(n4128), .Z(n4113) );
  AND U4371 ( .A(n2818), .B(n1761), .Z(n4128) );
  XOR U4372 ( .A(n4132), .B(n4114), .Z(n4127) );
  NAND U4373 ( .A(n1856), .B(n2688), .Z(n4114) );
  IV U4374 ( .A(n4116), .Z(n4132) );
  XNOR U4375 ( .A(n4121), .B(n4122), .Z(n4118) );
  NAND U4376 ( .A(n2058), .B(n2443), .Z(n4122) );
  XNOR U4377 ( .A(n4120), .B(n4136), .Z(n4121) );
  AND U4378 ( .A(n2566), .B(n1953), .Z(n4136) );
  XOR U4379 ( .A(n4141), .B(n4142), .Z(n3756) );
  XNOR U4380 ( .A(n4143), .B(n4140), .Z(n4141) );
  XNOR U4381 ( .A(n4129), .B(n4145), .Z(n4130) );
  AND U4382 ( .A(n2818), .B(n1856), .Z(n4145) );
  XOR U4383 ( .A(n4149), .B(n4131), .Z(n4144) );
  NAND U4384 ( .A(n1953), .B(n2688), .Z(n4131) );
  IV U4385 ( .A(n4133), .Z(n4149) );
  XOR U4386 ( .A(n4150), .B(n4151), .Z(n4133) );
  ANDN U4387 ( .A(n4152), .B(n4153), .Z(n4151) );
  XOR U4388 ( .A(n4150), .B(n4154), .Z(n4152) );
  XNOR U4389 ( .A(n4138), .B(n4139), .Z(n4135) );
  NAND U4390 ( .A(n2165), .B(n2443), .Z(n4139) );
  XNOR U4391 ( .A(n4137), .B(n4155), .Z(n4138) );
  AND U4392 ( .A(n2566), .B(n2058), .Z(n4155) );
  XOR U4393 ( .A(n4160), .B(n4161), .Z(n3791) );
  XNOR U4394 ( .A(n4162), .B(n4159), .Z(n4160) );
  XNOR U4395 ( .A(n4146), .B(n4164), .Z(n4147) );
  AND U4396 ( .A(n2818), .B(n1953), .Z(n4164) );
  XOR U4397 ( .A(n4168), .B(n4148), .Z(n4163) );
  NAND U4398 ( .A(n2058), .B(n2688), .Z(n4148) );
  IV U4399 ( .A(n4150), .Z(n4168) );
  XNOR U4400 ( .A(n4157), .B(n4158), .Z(n4154) );
  NAND U4401 ( .A(n2276), .B(n2443), .Z(n4158) );
  XNOR U4402 ( .A(n4156), .B(n4172), .Z(n4157) );
  AND U4403 ( .A(n2566), .B(n2165), .Z(n4172) );
  XOR U4404 ( .A(n4176), .B(n4177), .Z(n4159) );
  AND U4405 ( .A(n4178), .B(n4179), .Z(n4177) );
  XOR U4406 ( .A(n4180), .B(n4181), .Z(n4179) );
  XOR U4407 ( .A(n4176), .B(n4182), .Z(n4181) );
  XOR U4408 ( .A(n4170), .B(n4183), .Z(n4178) );
  XOR U4409 ( .A(n4176), .B(n4171), .Z(n4183) );
  NAND U4410 ( .A(n2443), .B(n2392), .Z(n4175) );
  XNOR U4411 ( .A(n4173), .B(n4184), .Z(n4174) );
  AND U4412 ( .A(n2566), .B(n2276), .Z(n4184) );
  XNOR U4413 ( .A(n4165), .B(n4189), .Z(n4166) );
  AND U4414 ( .A(n2818), .B(n2058), .Z(n4189) );
  XOR U4415 ( .A(n4193), .B(n4167), .Z(n4188) );
  NAND U4416 ( .A(n2165), .B(n2688), .Z(n4167) );
  IV U4417 ( .A(n4169), .Z(n4193) );
  XOR U4418 ( .A(n4197), .B(n4198), .Z(n4176) );
  AND U4419 ( .A(n4199), .B(n4200), .Z(n4198) );
  XOR U4420 ( .A(n4201), .B(n4202), .Z(n4200) );
  XOR U4421 ( .A(n4197), .B(n4203), .Z(n4202) );
  XOR U4422 ( .A(n4195), .B(n4204), .Z(n4199) );
  XOR U4423 ( .A(n4197), .B(n4196), .Z(n4204) );
  NAND U4424 ( .A(n2443), .B(n2513), .Z(n4187) );
  XNOR U4425 ( .A(n4185), .B(n4205), .Z(n4186) );
  AND U4426 ( .A(n2392), .B(n2566), .Z(n4205) );
  XNOR U4427 ( .A(n4190), .B(n4210), .Z(n4191) );
  AND U4428 ( .A(n2818), .B(n2165), .Z(n4210) );
  XOR U4429 ( .A(n4214), .B(n4192), .Z(n4209) );
  NAND U4430 ( .A(n2276), .B(n2688), .Z(n4192) );
  IV U4431 ( .A(n4194), .Z(n4214) );
  XOR U4432 ( .A(n4218), .B(n4219), .Z(n4197) );
  AND U4433 ( .A(n4220), .B(n4221), .Z(n4219) );
  XOR U4434 ( .A(n4222), .B(n4223), .Z(n4221) );
  XOR U4435 ( .A(n4218), .B(n4224), .Z(n4223) );
  XOR U4436 ( .A(n4216), .B(n4225), .Z(n4220) );
  XOR U4437 ( .A(n4218), .B(n4217), .Z(n4225) );
  NAND U4438 ( .A(n2443), .B(n2635), .Z(n4208) );
  XNOR U4439 ( .A(n4206), .B(n4226), .Z(n4207) );
  AND U4440 ( .A(n2513), .B(n2566), .Z(n4226) );
  XNOR U4441 ( .A(n4211), .B(n4231), .Z(n4212) );
  AND U4442 ( .A(n2818), .B(n2276), .Z(n4231) );
  XOR U4443 ( .A(n4235), .B(n4213), .Z(n4230) );
  NAND U4444 ( .A(n2688), .B(n2392), .Z(n4213) );
  IV U4445 ( .A(n4215), .Z(n4235) );
  XOR U4446 ( .A(n4239), .B(n4240), .Z(n4218) );
  AND U4447 ( .A(n4241), .B(n4242), .Z(n4240) );
  XOR U4448 ( .A(n4243), .B(n4244), .Z(n4242) );
  XOR U4449 ( .A(n4239), .B(n4245), .Z(n4244) );
  XOR U4450 ( .A(n4237), .B(n4246), .Z(n4241) );
  XOR U4451 ( .A(n4239), .B(n4238), .Z(n4246) );
  NAND U4452 ( .A(n2443), .B(n2763), .Z(n4229) );
  XNOR U4453 ( .A(n4227), .B(n4247), .Z(n4228) );
  AND U4454 ( .A(n2635), .B(n2566), .Z(n4247) );
  XNOR U4455 ( .A(n4232), .B(n4252), .Z(n4233) );
  AND U4456 ( .A(n2392), .B(n2818), .Z(n4252) );
  XOR U4457 ( .A(n4256), .B(n4234), .Z(n4251) );
  NAND U4458 ( .A(n2688), .B(n2513), .Z(n4234) );
  IV U4459 ( .A(n4236), .Z(n4256) );
  XOR U4460 ( .A(n4260), .B(n4261), .Z(n4239) );
  AND U4461 ( .A(n4262), .B(n4263), .Z(n4261) );
  XOR U4462 ( .A(n4264), .B(n4265), .Z(n4263) );
  XOR U4463 ( .A(n4260), .B(n4266), .Z(n4265) );
  XOR U4464 ( .A(n4258), .B(n4267), .Z(n4262) );
  XOR U4465 ( .A(n4260), .B(n4259), .Z(n4267) );
  NANDN U4466 ( .B(n2892), .A(n2443), .Z(n4250) );
  XNOR U4467 ( .A(n4248), .B(n4268), .Z(n4249) );
  AND U4468 ( .A(n2763), .B(n2566), .Z(n4268) );
  XNOR U4469 ( .A(n4253), .B(n4273), .Z(n4254) );
  AND U4470 ( .A(n2513), .B(n2818), .Z(n4273) );
  XOR U4471 ( .A(n4277), .B(n4255), .Z(n4272) );
  NAND U4472 ( .A(n2688), .B(n2635), .Z(n4255) );
  IV U4473 ( .A(n4257), .Z(n4277) );
  XOR U4474 ( .A(n4281), .B(n4282), .Z(n4260) );
  AND U4475 ( .A(n4283), .B(n4284), .Z(n4282) );
  XOR U4476 ( .A(n4285), .B(n4286), .Z(n4284) );
  XOR U4477 ( .A(n4281), .B(n4287), .Z(n4286) );
  XOR U4478 ( .A(n4279), .B(n4288), .Z(n4283) );
  XOR U4479 ( .A(n4281), .B(n4280), .Z(n4288) );
  NANDN U4480 ( .B(n3030), .A(n2443), .Z(n4271) );
  XNOR U4481 ( .A(n4269), .B(n4289), .Z(n4270) );
  ANDN U4482 ( .A(n2566), .B(n2892), .Z(n4289) );
  XNOR U4483 ( .A(n4274), .B(n4294), .Z(n4275) );
  AND U4484 ( .A(n2635), .B(n2818), .Z(n4294) );
  XOR U4485 ( .A(n4298), .B(n4276), .Z(n4293) );
  NAND U4486 ( .A(n2688), .B(n2763), .Z(n4276) );
  IV U4487 ( .A(n4278), .Z(n4298) );
  XOR U4488 ( .A(n4302), .B(n4303), .Z(n4281) );
  AND U4489 ( .A(n4304), .B(n4305), .Z(n4303) );
  XOR U4490 ( .A(n4306), .B(n4307), .Z(n4305) );
  XOR U4491 ( .A(n4302), .B(n4308), .Z(n4307) );
  XOR U4492 ( .A(n4300), .B(n4309), .Z(n4304) );
  XOR U4493 ( .A(n4302), .B(n4301), .Z(n4309) );
  NAND U4494 ( .A(n2443), .B(n3165), .Z(n4292) );
  XNOR U4495 ( .A(n4290), .B(n4310), .Z(n4291) );
  ANDN U4496 ( .A(n2566), .B(n3030), .Z(n4310) );
  XNOR U4497 ( .A(n4295), .B(n4315), .Z(n4296) );
  AND U4498 ( .A(n2763), .B(n2818), .Z(n4315) );
  XOR U4499 ( .A(n4319), .B(n4297), .Z(n4314) );
  NANDN U4500 ( .B(n2892), .A(n2688), .Z(n4297) );
  IV U4501 ( .A(n4299), .Z(n4319) );
  XOR U4502 ( .A(n4324), .B(n4325), .Z(n3896) );
  XNOR U4503 ( .A(n4326), .B(n4323), .Z(n4324) );
  XNOR U4504 ( .A(n4316), .B(n4328), .Z(n4317) );
  ANDN U4505 ( .A(n2818), .B(n2892), .Z(n4328) );
  XOR U4506 ( .A(n4331), .B(n4329), .Z(n4330) );
  ANDN U4507 ( .A(n2818), .B(n3030), .Z(n4331) );
  AND U4508 ( .A(n3165), .B(n2688), .Z(n4332) );
  XOR U4509 ( .A(n4336), .B(n4318), .Z(n4327) );
  NANDN U4510 ( .B(n3030), .A(n2688), .Z(n4318) );
  IV U4511 ( .A(n4320), .Z(n4336) );
  NAND U4512 ( .A(n2688), .B(n3854), .Z(n4335) );
  XNOR U4513 ( .A(n4333), .B(n4337), .Z(n4334) );
  AND U4514 ( .A(n3165), .B(n2818), .Z(n4337) );
  AND U4515 ( .A(n4338), .B(\_MAC/_MULT/A__[0] ), .Z(n4333) );
  NANDN U4516 ( .B(n2688), .A(n4339), .Z(n4338) );
  NAND U4517 ( .A(n3854), .B(n2818), .Z(n4339) );
  XNOR U4518 ( .A(n4312), .B(n4313), .Z(n4322) );
  NAND U4519 ( .A(n2443), .B(n3854), .Z(n4313) );
  XNOR U4520 ( .A(n4311), .B(n4342), .Z(n4312) );
  AND U4521 ( .A(n3165), .B(n2566), .Z(n4342) );
  AND U4522 ( .A(n4343), .B(\_MAC/_MULT/A__[0] ), .Z(n4311) );
  NANDN U4523 ( .B(n2443), .A(n4344), .Z(n4343) );
  NAND U4524 ( .A(n3854), .B(n2566), .Z(n4344) );
  XOR U4525 ( .A(n4347), .B(n4348), .Z(n4323) );
  AND U4526 ( .A(n4350), .B(n4351), .Z(n4349) );
  NANDN U4527 ( .B(n738), .A(n4352), .Z(n4351) );
  OR U4528 ( .A(n4353), .B(n4354), .Z(n4350) );
  XNOR U4529 ( .A(n4356), .B(n4355), .Z(n3918) );
  XNOR U4530 ( .A(n4357), .B(n4353), .Z(n4356) );
  NAND U4531 ( .A(n765), .B(n4352), .Z(n4353) );
  NANDN U4532 ( .B(n738), .A(\_MAC/_MULT/X__[0] ), .Z(n4358) );
  NANDN U4533 ( .B(n4359), .A(n4360), .Z(n738) );
  AND U4534 ( .A(n4361), .B(g_input[31]), .Z(n4360) );
  NAND U4535 ( .A(n838), .B(n2964), .Z(n3901) );
  XNOR U4536 ( .A(n3899), .B(n4365), .Z(n3900) );
  AND U4537 ( .A(n3096), .B(n797), .Z(n4365) );
  NAND U4538 ( .A(n875), .B(n2964), .Z(n4368) );
  XNOR U4539 ( .A(n4366), .B(n4370), .Z(n4367) );
  AND U4540 ( .A(n3096), .B(n838), .Z(n4370) );
  XNOR U4541 ( .A(n4362), .B(n4375), .Z(n4363) );
  AND U4542 ( .A(n765), .B(\_MAC/_MULT/X__[0] ), .Z(n4375) );
  XNOR U4543 ( .A(n4361), .B(g_input[30]), .Z(n4359) );
  NOR U4544 ( .A(n4376), .B(n4377), .Z(n4361) );
  XOR U4545 ( .A(n4381), .B(n4364), .Z(n4374) );
  NAND U4546 ( .A(n797), .B(n4352), .Z(n4364) );
  IV U4547 ( .A(n4369), .Z(n4381) );
  NAND U4548 ( .A(n917), .B(n2964), .Z(n4373) );
  XNOR U4549 ( .A(n4371), .B(n4383), .Z(n4372) );
  AND U4550 ( .A(n3096), .B(n875), .Z(n4383) );
  XNOR U4551 ( .A(n4378), .B(n4388), .Z(n4379) );
  AND U4552 ( .A(n797), .B(\_MAC/_MULT/X__[0] ), .Z(n4388) );
  XOR U4553 ( .A(n4376), .B(g_input[29]), .Z(n4377) );
  NANDN U4554 ( .B(n4389), .A(n4390), .Z(n4376) );
  XOR U4555 ( .A(n4394), .B(n4380), .Z(n4387) );
  NAND U4556 ( .A(n838), .B(n4352), .Z(n4380) );
  IV U4557 ( .A(n4382), .Z(n4394) );
  NAND U4558 ( .A(n961), .B(n2964), .Z(n4386) );
  XNOR U4559 ( .A(n4384), .B(n4396), .Z(n4385) );
  AND U4560 ( .A(n3096), .B(n917), .Z(n4396) );
  XNOR U4561 ( .A(n4391), .B(n4401), .Z(n4392) );
  AND U4562 ( .A(n838), .B(\_MAC/_MULT/X__[0] ), .Z(n4401) );
  XNOR U4563 ( .A(n4390), .B(g_input[28]), .Z(n4389) );
  NOR U4564 ( .A(n4402), .B(n4403), .Z(n4390) );
  XOR U4565 ( .A(n4407), .B(n4393), .Z(n4400) );
  NAND U4566 ( .A(n875), .B(n4352), .Z(n4393) );
  IV U4567 ( .A(n4395), .Z(n4407) );
  NAND U4568 ( .A(n1019), .B(n2964), .Z(n4399) );
  XNOR U4569 ( .A(n4397), .B(n4409), .Z(n4398) );
  AND U4570 ( .A(n3096), .B(n961), .Z(n4409) );
  XNOR U4571 ( .A(n4404), .B(n4414), .Z(n4405) );
  AND U4572 ( .A(n875), .B(\_MAC/_MULT/X__[0] ), .Z(n4414) );
  XOR U4573 ( .A(n4402), .B(g_input[27]), .Z(n4403) );
  NANDN U4574 ( .B(n4415), .A(n4416), .Z(n4402) );
  XOR U4575 ( .A(n4420), .B(n4406), .Z(n4413) );
  NAND U4576 ( .A(n917), .B(n4352), .Z(n4406) );
  IV U4577 ( .A(n4408), .Z(n4420) );
  NAND U4578 ( .A(n1077), .B(n2964), .Z(n4412) );
  XNOR U4579 ( .A(n4410), .B(n4422), .Z(n4411) );
  AND U4580 ( .A(n3096), .B(n1019), .Z(n4422) );
  XNOR U4581 ( .A(n4417), .B(n4427), .Z(n4418) );
  AND U4582 ( .A(n917), .B(\_MAC/_MULT/X__[0] ), .Z(n4427) );
  XNOR U4583 ( .A(n4416), .B(g_input[26]), .Z(n4415) );
  NOR U4584 ( .A(n4428), .B(n4429), .Z(n4416) );
  XOR U4585 ( .A(n4433), .B(n4419), .Z(n4426) );
  NAND U4586 ( .A(n961), .B(n4352), .Z(n4419) );
  IV U4587 ( .A(n4421), .Z(n4433) );
  NAND U4588 ( .A(n1137), .B(n2964), .Z(n4425) );
  XNOR U4589 ( .A(n4423), .B(n4435), .Z(n4424) );
  AND U4590 ( .A(n3096), .B(n1077), .Z(n4435) );
  XNOR U4591 ( .A(n4430), .B(n4440), .Z(n4431) );
  AND U4592 ( .A(n961), .B(\_MAC/_MULT/X__[0] ), .Z(n4440) );
  XOR U4593 ( .A(n4428), .B(g_input[25]), .Z(n4429) );
  NANDN U4594 ( .B(n4441), .A(n4442), .Z(n4428) );
  XOR U4595 ( .A(n4446), .B(n4432), .Z(n4439) );
  NAND U4596 ( .A(n1019), .B(n4352), .Z(n4432) );
  IV U4597 ( .A(n4434), .Z(n4446) );
  NAND U4598 ( .A(n1200), .B(n2964), .Z(n4438) );
  XNOR U4599 ( .A(n4436), .B(n4448), .Z(n4437) );
  AND U4600 ( .A(n3096), .B(n1137), .Z(n4448) );
  XNOR U4601 ( .A(n4443), .B(n4453), .Z(n4444) );
  AND U4602 ( .A(n1019), .B(\_MAC/_MULT/X__[0] ), .Z(n4453) );
  XNOR U4603 ( .A(n4442), .B(g_input[24]), .Z(n4441) );
  NOR U4604 ( .A(n4454), .B(n4455), .Z(n4442) );
  XOR U4605 ( .A(n4459), .B(n4445), .Z(n4452) );
  NAND U4606 ( .A(n1077), .B(n4352), .Z(n4445) );
  IV U4607 ( .A(n4447), .Z(n4459) );
  NAND U4608 ( .A(n1268), .B(n2964), .Z(n4451) );
  XNOR U4609 ( .A(n4449), .B(n4461), .Z(n4450) );
  AND U4610 ( .A(n3096), .B(n1200), .Z(n4461) );
  XNOR U4611 ( .A(n4456), .B(n4466), .Z(n4457) );
  AND U4612 ( .A(n1077), .B(\_MAC/_MULT/X__[0] ), .Z(n4466) );
  XOR U4613 ( .A(n4454), .B(g_input[23]), .Z(n4455) );
  NANDN U4614 ( .B(n4467), .A(n4468), .Z(n4454) );
  XOR U4615 ( .A(n4472), .B(n4458), .Z(n4465) );
  NAND U4616 ( .A(n1137), .B(n4352), .Z(n4458) );
  IV U4617 ( .A(n4460), .Z(n4472) );
  NAND U4618 ( .A(n1338), .B(n2964), .Z(n4464) );
  XNOR U4619 ( .A(n4462), .B(n4474), .Z(n4463) );
  AND U4620 ( .A(n3096), .B(n1268), .Z(n4474) );
  XNOR U4621 ( .A(n4469), .B(n4479), .Z(n4470) );
  AND U4622 ( .A(n1137), .B(\_MAC/_MULT/X__[0] ), .Z(n4479) );
  XNOR U4623 ( .A(n4468), .B(g_input[22]), .Z(n4467) );
  NOR U4624 ( .A(n4480), .B(n4481), .Z(n4468) );
  XOR U4625 ( .A(n4485), .B(n4471), .Z(n4478) );
  NAND U4626 ( .A(n1200), .B(n4352), .Z(n4471) );
  IV U4627 ( .A(n4473), .Z(n4485) );
  NAND U4628 ( .A(n1412), .B(n2964), .Z(n4477) );
  XNOR U4629 ( .A(n4475), .B(n4487), .Z(n4476) );
  AND U4630 ( .A(n3096), .B(n1338), .Z(n4487) );
  XNOR U4631 ( .A(n4482), .B(n4492), .Z(n4483) );
  AND U4632 ( .A(n1200), .B(\_MAC/_MULT/X__[0] ), .Z(n4492) );
  XOR U4633 ( .A(n4480), .B(g_input[21]), .Z(n4481) );
  NANDN U4634 ( .B(n4493), .A(n4494), .Z(n4480) );
  XOR U4635 ( .A(n4498), .B(n4484), .Z(n4491) );
  NAND U4636 ( .A(n1268), .B(n4352), .Z(n4484) );
  IV U4637 ( .A(n4486), .Z(n4498) );
  NAND U4638 ( .A(n1491), .B(n2964), .Z(n4490) );
  XNOR U4639 ( .A(n4488), .B(n4500), .Z(n4489) );
  AND U4640 ( .A(n3096), .B(n1412), .Z(n4500) );
  XNOR U4641 ( .A(n4495), .B(n4505), .Z(n4496) );
  AND U4642 ( .A(n1268), .B(\_MAC/_MULT/X__[0] ), .Z(n4505) );
  XNOR U4643 ( .A(n4494), .B(g_input[20]), .Z(n4493) );
  NOR U4644 ( .A(n4506), .B(n4507), .Z(n4494) );
  XOR U4645 ( .A(n4511), .B(n4497), .Z(n4504) );
  NAND U4646 ( .A(n1338), .B(n4352), .Z(n4497) );
  IV U4647 ( .A(n4499), .Z(n4511) );
  NAND U4648 ( .A(n1576), .B(n2964), .Z(n4503) );
  XNOR U4649 ( .A(n4501), .B(n4513), .Z(n4502) );
  AND U4650 ( .A(n3096), .B(n1491), .Z(n4513) );
  XNOR U4651 ( .A(n4508), .B(n4518), .Z(n4509) );
  AND U4652 ( .A(n1338), .B(\_MAC/_MULT/X__[0] ), .Z(n4518) );
  XOR U4653 ( .A(n4506), .B(g_input[19]), .Z(n4507) );
  NANDN U4654 ( .B(n4519), .A(n4520), .Z(n4506) );
  XOR U4655 ( .A(n4524), .B(n4510), .Z(n4517) );
  NAND U4656 ( .A(n1412), .B(n4352), .Z(n4510) );
  IV U4657 ( .A(n4512), .Z(n4524) );
  NAND U4658 ( .A(n1668), .B(n2964), .Z(n4516) );
  XNOR U4659 ( .A(n4514), .B(n4526), .Z(n4515) );
  AND U4660 ( .A(n3096), .B(n1576), .Z(n4526) );
  XNOR U4661 ( .A(n4521), .B(n4531), .Z(n4522) );
  AND U4662 ( .A(n1412), .B(\_MAC/_MULT/X__[0] ), .Z(n4531) );
  XNOR U4663 ( .A(n4520), .B(g_input[18]), .Z(n4519) );
  NOR U4664 ( .A(n4532), .B(n4533), .Z(n4520) );
  XOR U4665 ( .A(n4537), .B(n4523), .Z(n4530) );
  NAND U4666 ( .A(n1491), .B(n4352), .Z(n4523) );
  IV U4667 ( .A(n4525), .Z(n4537) );
  NAND U4668 ( .A(n1761), .B(n2964), .Z(n4529) );
  XNOR U4669 ( .A(n4527), .B(n4539), .Z(n4528) );
  AND U4670 ( .A(n3096), .B(n1668), .Z(n4539) );
  XNOR U4671 ( .A(n4534), .B(n4544), .Z(n4535) );
  AND U4672 ( .A(n1491), .B(\_MAC/_MULT/X__[0] ), .Z(n4544) );
  XOR U4673 ( .A(n4532), .B(g_input[17]), .Z(n4533) );
  NANDN U4674 ( .B(n4545), .A(n4546), .Z(n4532) );
  XOR U4675 ( .A(n4550), .B(n4536), .Z(n4543) );
  NAND U4676 ( .A(n1576), .B(n4352), .Z(n4536) );
  IV U4677 ( .A(n4538), .Z(n4550) );
  XOR U4678 ( .A(n4551), .B(n4552), .Z(n4538) );
  AND U4679 ( .A(n4162), .B(n4553), .Z(n4552) );
  XNOR U4680 ( .A(n4551), .B(n4161), .Z(n4553) );
  NAND U4681 ( .A(n1856), .B(n2964), .Z(n4542) );
  XNOR U4682 ( .A(n4540), .B(n4554), .Z(n4541) );
  AND U4683 ( .A(n3096), .B(n1761), .Z(n4554) );
  XNOR U4684 ( .A(n4547), .B(n4559), .Z(n4548) );
  AND U4685 ( .A(n1576), .B(\_MAC/_MULT/X__[0] ), .Z(n4559) );
  XOR U4686 ( .A(n4563), .B(n4549), .Z(n4558) );
  NAND U4687 ( .A(n1668), .B(n4352), .Z(n4549) );
  IV U4688 ( .A(n4551), .Z(n4563) );
  NAND U4689 ( .A(n1953), .B(n2964), .Z(n4557) );
  XNOR U4690 ( .A(n4555), .B(n4565), .Z(n4556) );
  AND U4691 ( .A(n3096), .B(n1856), .Z(n4565) );
  XNOR U4692 ( .A(n4560), .B(n4570), .Z(n4561) );
  AND U4693 ( .A(n1668), .B(\_MAC/_MULT/X__[0] ), .Z(n4570) );
  XOR U4694 ( .A(n4574), .B(n4562), .Z(n4569) );
  NAND U4695 ( .A(n1761), .B(n4352), .Z(n4562) );
  IV U4696 ( .A(n4564), .Z(n4574) );
  NAND U4697 ( .A(n2058), .B(n2964), .Z(n4568) );
  XNOR U4698 ( .A(n4566), .B(n4576), .Z(n4567) );
  AND U4699 ( .A(n3096), .B(n1953), .Z(n4576) );
  XNOR U4700 ( .A(n4571), .B(n4581), .Z(n4572) );
  AND U4701 ( .A(n1761), .B(\_MAC/_MULT/X__[0] ), .Z(n4581) );
  XOR U4702 ( .A(n4585), .B(n4573), .Z(n4580) );
  NAND U4703 ( .A(n1856), .B(n4352), .Z(n4573) );
  IV U4704 ( .A(n4575), .Z(n4585) );
  NAND U4705 ( .A(n2165), .B(n2964), .Z(n4579) );
  XNOR U4706 ( .A(n4577), .B(n4587), .Z(n4578) );
  AND U4707 ( .A(n3096), .B(n2058), .Z(n4587) );
  XNOR U4708 ( .A(n4582), .B(n4592), .Z(n4583) );
  AND U4709 ( .A(n1856), .B(\_MAC/_MULT/X__[0] ), .Z(n4592) );
  XOR U4710 ( .A(n4596), .B(n4584), .Z(n4591) );
  NAND U4711 ( .A(n1953), .B(n4352), .Z(n4584) );
  IV U4712 ( .A(n4586), .Z(n4596) );
  NAND U4713 ( .A(n2276), .B(n2964), .Z(n4590) );
  XNOR U4714 ( .A(n4588), .B(n4598), .Z(n4589) );
  AND U4715 ( .A(n3096), .B(n2165), .Z(n4598) );
  XNOR U4716 ( .A(n4593), .B(n4603), .Z(n4594) );
  AND U4717 ( .A(n1953), .B(\_MAC/_MULT/X__[0] ), .Z(n4603) );
  XOR U4718 ( .A(n4607), .B(n4595), .Z(n4602) );
  NAND U4719 ( .A(n2058), .B(n4352), .Z(n4595) );
  IV U4720 ( .A(n4597), .Z(n4607) );
  NAND U4721 ( .A(n2392), .B(n2964), .Z(n4601) );
  XNOR U4722 ( .A(n4599), .B(n4609), .Z(n4600) );
  AND U4723 ( .A(n3096), .B(n2276), .Z(n4609) );
  XNOR U4724 ( .A(n4604), .B(n4614), .Z(n4605) );
  AND U4725 ( .A(n2058), .B(\_MAC/_MULT/X__[0] ), .Z(n4614) );
  XOR U4726 ( .A(n4618), .B(n4606), .Z(n4613) );
  NAND U4727 ( .A(n2165), .B(n4352), .Z(n4606) );
  IV U4728 ( .A(n4608), .Z(n4618) );
  NAND U4729 ( .A(n2513), .B(n2964), .Z(n4612) );
  XNOR U4730 ( .A(n4610), .B(n4620), .Z(n4611) );
  AND U4731 ( .A(n3096), .B(n2392), .Z(n4620) );
  XNOR U4732 ( .A(n4615), .B(n4625), .Z(n4616) );
  AND U4733 ( .A(n2165), .B(\_MAC/_MULT/X__[0] ), .Z(n4625) );
  XOR U4734 ( .A(n4629), .B(n4617), .Z(n4624) );
  NAND U4735 ( .A(n2276), .B(n4352), .Z(n4617) );
  IV U4736 ( .A(n4619), .Z(n4629) );
  NAND U4737 ( .A(n2635), .B(n2964), .Z(n4623) );
  XNOR U4738 ( .A(n4621), .B(n4631), .Z(n4622) );
  AND U4739 ( .A(n3096), .B(n2513), .Z(n4631) );
  XNOR U4740 ( .A(n4626), .B(n4636), .Z(n4627) );
  AND U4741 ( .A(n2276), .B(\_MAC/_MULT/X__[0] ), .Z(n4636) );
  XOR U4742 ( .A(n4640), .B(n4628), .Z(n4635) );
  NAND U4743 ( .A(n2392), .B(n4352), .Z(n4628) );
  IV U4744 ( .A(n4630), .Z(n4640) );
  NAND U4745 ( .A(n2763), .B(n2964), .Z(n4634) );
  XNOR U4746 ( .A(n4632), .B(n4642), .Z(n4633) );
  AND U4747 ( .A(n3096), .B(n2635), .Z(n4642) );
  XNOR U4748 ( .A(n4646), .B(n4643), .Z(n4645) );
  XNOR U4749 ( .A(n4637), .B(n4648), .Z(n4638) );
  AND U4750 ( .A(n2392), .B(\_MAC/_MULT/X__[0] ), .Z(n4648) );
  XNOR U4751 ( .A(n4652), .B(n4649), .Z(n4651) );
  XOR U4752 ( .A(n4653), .B(n4639), .Z(n4647) );
  NAND U4753 ( .A(n2513), .B(n4352), .Z(n4639) );
  IV U4754 ( .A(n4641), .Z(n4653) );
  XNOR U4755 ( .A(n4654), .B(n4655), .Z(n4641) );
  AND U4756 ( .A(n4656), .B(n4657), .Z(n4655) );
  XOR U4757 ( .A(n4650), .B(n4658), .Z(n4657) );
  XNOR U4758 ( .A(n4652), .B(n4654), .Z(n4658) );
  NAND U4759 ( .A(n2635), .B(n4352), .Z(n4652) );
  XOR U4760 ( .A(n4649), .B(n4659), .Z(n4650) );
  AND U4761 ( .A(n2513), .B(\_MAC/_MULT/X__[0] ), .Z(n4659) );
  XNOR U4762 ( .A(n4663), .B(n4660), .Z(n4662) );
  XOR U4763 ( .A(n4644), .B(n4664), .Z(n4656) );
  XNOR U4764 ( .A(n4646), .B(n4654), .Z(n4664) );
  NANDN U4765 ( .B(n2892), .A(n2964), .Z(n4646) );
  XOR U4766 ( .A(n4643), .B(n4665), .Z(n4644) );
  AND U4767 ( .A(n3096), .B(n2763), .Z(n4665) );
  XNOR U4768 ( .A(n4669), .B(n4666), .Z(n4668) );
  XOR U4769 ( .A(n4670), .B(n4671), .Z(n4654) );
  AND U4770 ( .A(n4672), .B(n4673), .Z(n4671) );
  XOR U4771 ( .A(n4661), .B(n4674), .Z(n4673) );
  XNOR U4772 ( .A(n4663), .B(n4670), .Z(n4674) );
  NAND U4773 ( .A(n2763), .B(n4352), .Z(n4663) );
  XOR U4774 ( .A(n4660), .B(n4675), .Z(n4661) );
  AND U4775 ( .A(n2635), .B(\_MAC/_MULT/X__[0] ), .Z(n4675) );
  XNOR U4776 ( .A(n4679), .B(n4676), .Z(n4678) );
  XOR U4777 ( .A(n4667), .B(n4680), .Z(n4672) );
  XNOR U4778 ( .A(n4669), .B(n4670), .Z(n4680) );
  NANDN U4779 ( .B(n3030), .A(n2964), .Z(n4669) );
  XOR U4780 ( .A(n4666), .B(n4681), .Z(n4667) );
  ANDN U4781 ( .A(n3096), .B(n2892), .Z(n4681) );
  XNOR U4782 ( .A(n4685), .B(n4682), .Z(n4684) );
  XOR U4783 ( .A(n4686), .B(n4687), .Z(n4670) );
  AND U4784 ( .A(n4688), .B(n4689), .Z(n4687) );
  XOR U4785 ( .A(n4677), .B(n4690), .Z(n4689) );
  XNOR U4786 ( .A(n4679), .B(n4686), .Z(n4690) );
  NANDN U4787 ( .B(n2892), .A(n4352), .Z(n4679) );
  XOR U4788 ( .A(n4676), .B(n4691), .Z(n4677) );
  AND U4789 ( .A(n2763), .B(\_MAC/_MULT/X__[0] ), .Z(n4691) );
  XOR U4790 ( .A(n4683), .B(n4695), .Z(n4688) );
  XNOR U4791 ( .A(n4685), .B(n4686), .Z(n4695) );
  NAND U4792 ( .A(n2964), .B(n3165), .Z(n4685) );
  XOR U4793 ( .A(n4682), .B(n4696), .Z(n4683) );
  ANDN U4794 ( .A(n3096), .B(n3030), .Z(n4696) );
  NAND U4795 ( .A(n2964), .B(n3854), .Z(n4699) );
  XNOR U4796 ( .A(n4697), .B(n4701), .Z(n4698) );
  AND U4797 ( .A(n3165), .B(n3096), .Z(n4701) );
  AND U4798 ( .A(n4702), .B(\_MAC/_MULT/A__[0] ), .Z(n4697) );
  NANDN U4799 ( .B(n2964), .A(n4703), .Z(n4702) );
  NAND U4800 ( .A(n3854), .B(n3096), .Z(n4703) );
  XNOR U4801 ( .A(n4692), .B(n4707), .Z(n4693) );
  ANDN U4802 ( .A(\_MAC/_MULT/X__[0] ), .B(n2892), .Z(n4707) );
  XOR U4803 ( .A(n4710), .B(n4708), .Z(n4709) );
  ANDN U4804 ( .A(\_MAC/_MULT/X__[0] ), .B(n3030), .Z(n4710) );
  AND U4805 ( .A(n4352), .B(n3165), .Z(n4711) );
  XOR U4806 ( .A(n4715), .B(n4694), .Z(n4706) );
  NANDN U4807 ( .B(n3030), .A(n4352), .Z(n4694) );
  IV U4808 ( .A(n4700), .Z(n4715) );
  NAND U4809 ( .A(n4352), .B(n3854), .Z(n4714) );
  XNOR U4810 ( .A(n4712), .B(n4716), .Z(n4713) );
  AND U4811 ( .A(n3165), .B(\_MAC/_MULT/X__[0] ), .Z(n4716) );
  AND U4812 ( .A(n4717), .B(\_MAC/_MULT/A__[0] ), .Z(n4712) );
  NANDN U4813 ( .B(n4352), .A(n4718), .Z(n4717) );
  NAND U4814 ( .A(n3854), .B(\_MAC/_MULT/X__[0] ), .Z(n4718) );
  XNOR U4815 ( .A(n4720), .B(n3129), .Z(n3120) );
  XNOR U4816 ( .A(n3108), .B(n4722), .Z(n3109) );
  AND U4817 ( .A(n1953), .B(n1218), .Z(n4722) );
  XOR U4818 ( .A(n4726), .B(n3110), .Z(n4721) );
  NAND U4819 ( .A(n1158), .B(n2058), .Z(n3110) );
  IV U4820 ( .A(n3112), .Z(n4726) );
  XNOR U4821 ( .A(n3117), .B(n3118), .Z(n3114) );
  NANDN U4822 ( .B(n1040), .A(n2276), .Z(n3118) );
  XNOR U4823 ( .A(n3116), .B(n4730), .Z(n3117) );
  AND U4824 ( .A(n2165), .B(n1102), .Z(n4730) );
  XNOR U4825 ( .A(n3128), .B(n3119), .Z(n4720) );
  XOR U4826 ( .A(n4734), .B(n4735), .Z(n3119) );
  XOR U4827 ( .A(n4736), .B(n3138), .Z(n3128) );
  XNOR U4828 ( .A(n3125), .B(n3126), .Z(n3138) );
  NAND U4829 ( .A(n1306), .B(n1856), .Z(n3126) );
  XNOR U4830 ( .A(n3124), .B(n4737), .Z(n3125) );
  AND U4831 ( .A(n1761), .B(n1376), .Z(n4737) );
  XNOR U4832 ( .A(n3137), .B(n3127), .Z(n4736) );
  XOR U4833 ( .A(n4741), .B(n4742), .Z(n3127) );
  AND U4834 ( .A(n4743), .B(n4744), .Z(n4742) );
  XOR U4835 ( .A(n4745), .B(n4746), .Z(n4744) );
  XOR U4836 ( .A(n4741), .B(n4747), .Z(n4746) );
  XOR U4837 ( .A(n4728), .B(n4748), .Z(n4743) );
  XOR U4838 ( .A(n4741), .B(n4729), .Z(n4748) );
  NANDN U4839 ( .B(n1040), .A(n2392), .Z(n4733) );
  XNOR U4840 ( .A(n4731), .B(n4749), .Z(n4732) );
  AND U4841 ( .A(n2276), .B(n1102), .Z(n4749) );
  XNOR U4842 ( .A(n4723), .B(n4754), .Z(n4724) );
  AND U4843 ( .A(n2058), .B(n1218), .Z(n4754) );
  XOR U4844 ( .A(n4758), .B(n4725), .Z(n4753) );
  NAND U4845 ( .A(n1158), .B(n2165), .Z(n4725) );
  IV U4846 ( .A(n4727), .Z(n4758) );
  XOR U4847 ( .A(n4762), .B(n4763), .Z(n4741) );
  AND U4848 ( .A(n4764), .B(n4765), .Z(n4763) );
  XOR U4849 ( .A(n4766), .B(n4767), .Z(n4765) );
  XOR U4850 ( .A(n4762), .B(n4768), .Z(n4767) );
  XOR U4851 ( .A(n4760), .B(n4769), .Z(n4764) );
  XOR U4852 ( .A(n4762), .B(n4761), .Z(n4769) );
  NANDN U4853 ( .B(n1040), .A(n2513), .Z(n4752) );
  XNOR U4854 ( .A(n4750), .B(n4770), .Z(n4751) );
  AND U4855 ( .A(n2392), .B(n1102), .Z(n4770) );
  XNOR U4856 ( .A(n4755), .B(n4775), .Z(n4756) );
  AND U4857 ( .A(n2165), .B(n1218), .Z(n4775) );
  XOR U4858 ( .A(n4779), .B(n4757), .Z(n4774) );
  NAND U4859 ( .A(n1158), .B(n2276), .Z(n4757) );
  IV U4860 ( .A(n4759), .Z(n4779) );
  XOR U4861 ( .A(n4783), .B(n4784), .Z(n4762) );
  AND U4862 ( .A(n4785), .B(n4786), .Z(n4784) );
  XOR U4863 ( .A(n4787), .B(n4788), .Z(n4786) );
  XOR U4864 ( .A(n4783), .B(n4789), .Z(n4788) );
  XOR U4865 ( .A(n4781), .B(n4790), .Z(n4785) );
  XOR U4866 ( .A(n4783), .B(n4782), .Z(n4790) );
  NANDN U4867 ( .B(n1040), .A(n2635), .Z(n4773) );
  XNOR U4868 ( .A(n4771), .B(n4791), .Z(n4772) );
  AND U4869 ( .A(n2513), .B(n1102), .Z(n4791) );
  XNOR U4870 ( .A(n4776), .B(n4796), .Z(n4777) );
  AND U4871 ( .A(n2276), .B(n1218), .Z(n4796) );
  XOR U4872 ( .A(n4800), .B(n4778), .Z(n4795) );
  NAND U4873 ( .A(n1158), .B(n2392), .Z(n4778) );
  IV U4874 ( .A(n4780), .Z(n4800) );
  XOR U4875 ( .A(n4804), .B(n4805), .Z(n4783) );
  AND U4876 ( .A(n4806), .B(n4807), .Z(n4805) );
  XOR U4877 ( .A(n4808), .B(n4809), .Z(n4807) );
  XOR U4878 ( .A(n4804), .B(n4810), .Z(n4809) );
  XOR U4879 ( .A(n4802), .B(n4811), .Z(n4806) );
  XOR U4880 ( .A(n4804), .B(n4803), .Z(n4811) );
  NANDN U4881 ( .B(n1040), .A(n2763), .Z(n4794) );
  XNOR U4882 ( .A(n4792), .B(n4812), .Z(n4793) );
  AND U4883 ( .A(n2635), .B(n1102), .Z(n4812) );
  XNOR U4884 ( .A(n4797), .B(n4817), .Z(n4798) );
  AND U4885 ( .A(n2392), .B(n1218), .Z(n4817) );
  XOR U4886 ( .A(n4821), .B(n4799), .Z(n4816) );
  NAND U4887 ( .A(n1158), .B(n2513), .Z(n4799) );
  IV U4888 ( .A(n4801), .Z(n4821) );
  XOR U4889 ( .A(n4825), .B(n4826), .Z(n4804) );
  AND U4890 ( .A(n4827), .B(n4828), .Z(n4826) );
  XOR U4891 ( .A(n4829), .B(n4830), .Z(n4828) );
  XOR U4892 ( .A(n4825), .B(n4831), .Z(n4830) );
  XOR U4893 ( .A(n4823), .B(n4832), .Z(n4827) );
  XOR U4894 ( .A(n4825), .B(n4824), .Z(n4832) );
  OR U4895 ( .A(n1040), .B(n2892), .Z(n4815) );
  XNOR U4896 ( .A(n4813), .B(n4833), .Z(n4814) );
  AND U4897 ( .A(n2763), .B(n1102), .Z(n4833) );
  XNOR U4898 ( .A(n4818), .B(n4838), .Z(n4819) );
  AND U4899 ( .A(n2513), .B(n1218), .Z(n4838) );
  XOR U4900 ( .A(n4842), .B(n4820), .Z(n4837) );
  NAND U4901 ( .A(n1158), .B(n2635), .Z(n4820) );
  IV U4902 ( .A(n4822), .Z(n4842) );
  XOR U4903 ( .A(n4846), .B(n4847), .Z(n4825) );
  AND U4904 ( .A(n4848), .B(n4849), .Z(n4847) );
  XOR U4905 ( .A(n4850), .B(n4851), .Z(n4849) );
  XOR U4906 ( .A(n4846), .B(n4852), .Z(n4851) );
  XOR U4907 ( .A(n4844), .B(n4853), .Z(n4848) );
  XOR U4908 ( .A(n4846), .B(n4845), .Z(n4853) );
  OR U4909 ( .A(n1040), .B(n3030), .Z(n4836) );
  XNOR U4910 ( .A(n4834), .B(n4854), .Z(n4835) );
  ANDN U4911 ( .A(n1102), .B(n2892), .Z(n4854) );
  XNOR U4912 ( .A(n4839), .B(n4859), .Z(n4840) );
  AND U4913 ( .A(n2635), .B(n1218), .Z(n4859) );
  XOR U4914 ( .A(n4863), .B(n4841), .Z(n4858) );
  NAND U4915 ( .A(n1158), .B(n2763), .Z(n4841) );
  IV U4916 ( .A(n4843), .Z(n4863) );
  XOR U4917 ( .A(n4867), .B(n4868), .Z(n4846) );
  AND U4918 ( .A(n4869), .B(n4870), .Z(n4868) );
  XOR U4919 ( .A(n4871), .B(n4872), .Z(n4870) );
  XOR U4920 ( .A(n4867), .B(n4873), .Z(n4872) );
  XOR U4921 ( .A(n4865), .B(n4874), .Z(n4869) );
  XOR U4922 ( .A(n4867), .B(n4866), .Z(n4874) );
  NANDN U4923 ( .B(n1040), .A(n3165), .Z(n4857) );
  XNOR U4924 ( .A(n4855), .B(n4875), .Z(n4856) );
  ANDN U4925 ( .A(n1102), .B(n3030), .Z(n4875) );
  XNOR U4926 ( .A(n4860), .B(n4880), .Z(n4861) );
  AND U4927 ( .A(n2763), .B(n1218), .Z(n4880) );
  XOR U4928 ( .A(n4884), .B(n4862), .Z(n4879) );
  NANDN U4929 ( .B(n2892), .A(n1158), .Z(n4862) );
  IV U4930 ( .A(n4864), .Z(n4884) );
  XOR U4931 ( .A(n4889), .B(n4890), .Z(n4735) );
  XNOR U4932 ( .A(n4891), .B(n4888), .Z(n4889) );
  XNOR U4933 ( .A(n4881), .B(n4893), .Z(n4882) );
  ANDN U4934 ( .A(n1218), .B(n2892), .Z(n4893) );
  XOR U4935 ( .A(n4896), .B(n4894), .Z(n4895) );
  ANDN U4936 ( .A(n1218), .B(n3030), .Z(n4896) );
  AND U4937 ( .A(n3165), .B(n1158), .Z(n4897) );
  XOR U4938 ( .A(n4901), .B(n4883), .Z(n4892) );
  NANDN U4939 ( .B(n3030), .A(n1158), .Z(n4883) );
  IV U4940 ( .A(n4885), .Z(n4901) );
  NAND U4941 ( .A(n1158), .B(n3854), .Z(n4900) );
  XNOR U4942 ( .A(n4898), .B(n4902), .Z(n4899) );
  AND U4943 ( .A(n3165), .B(n1218), .Z(n4902) );
  AND U4944 ( .A(n4903), .B(\_MAC/_MULT/A__[0] ), .Z(n4898) );
  NANDN U4945 ( .B(n1158), .A(n4904), .Z(n4903) );
  NAND U4946 ( .A(n3854), .B(n1218), .Z(n4904) );
  XNOR U4947 ( .A(n4877), .B(n4878), .Z(n4887) );
  NANDN U4948 ( .B(n1040), .A(n3854), .Z(n4878) );
  XNOR U4949 ( .A(n4876), .B(n4907), .Z(n4877) );
  AND U4950 ( .A(n3165), .B(n1102), .Z(n4907) );
  AND U4951 ( .A(n4908), .B(\_MAC/_MULT/A__[0] ), .Z(n4876) );
  NAND U4952 ( .A(n4909), .B(n1040), .Z(n4908) );
  NAND U4953 ( .A(n3854), .B(n1102), .Z(n4909) );
  XOR U4954 ( .A(n4912), .B(n4913), .Z(n4888) );
  XNOR U4955 ( .A(n3132), .B(n4915), .Z(n3133) );
  AND U4956 ( .A(n1576), .B(n1546), .Z(n4915) );
  XNOR U4957 ( .A(n4546), .B(g_input[16]), .Z(n4545) );
  NOR U4958 ( .A(n4916), .B(n4917), .Z(n4546) );
  XOR U4959 ( .A(n4921), .B(n3134), .Z(n4914) );
  NAND U4960 ( .A(n1457), .B(n1668), .Z(n3134) );
  IV U4961 ( .A(n3136), .Z(n4921) );
  NAND U4962 ( .A(n1306), .B(n1953), .Z(n4740) );
  XNOR U4963 ( .A(n4738), .B(n4923), .Z(n4739) );
  AND U4964 ( .A(n1856), .B(n1376), .Z(n4923) );
  XNOR U4965 ( .A(n4918), .B(n4928), .Z(n4919) );
  AND U4966 ( .A(n1668), .B(n1546), .Z(n4928) );
  XOR U4967 ( .A(n4916), .B(g_input[15]), .Z(n4917) );
  NANDN U4968 ( .B(n4929), .A(n4930), .Z(n4916) );
  XOR U4969 ( .A(n4934), .B(n4920), .Z(n4927) );
  NAND U4970 ( .A(n1457), .B(n1761), .Z(n4920) );
  IV U4971 ( .A(n4922), .Z(n4934) );
  NAND U4972 ( .A(n1306), .B(n2058), .Z(n4926) );
  XNOR U4973 ( .A(n4924), .B(n4936), .Z(n4925) );
  AND U4974 ( .A(n1953), .B(n1376), .Z(n4936) );
  XNOR U4975 ( .A(n4931), .B(n4941), .Z(n4932) );
  AND U4976 ( .A(n1761), .B(n1546), .Z(n4941) );
  XNOR U4977 ( .A(n4930), .B(g_input[14]), .Z(n4929) );
  NOR U4978 ( .A(n4942), .B(n4943), .Z(n4930) );
  XOR U4979 ( .A(n4947), .B(n4933), .Z(n4940) );
  NAND U4980 ( .A(n1457), .B(n1856), .Z(n4933) );
  IV U4981 ( .A(n4935), .Z(n4947) );
  NAND U4982 ( .A(n1306), .B(n2165), .Z(n4939) );
  XNOR U4983 ( .A(n4937), .B(n4949), .Z(n4938) );
  AND U4984 ( .A(n2058), .B(n1376), .Z(n4949) );
  XNOR U4985 ( .A(n4944), .B(n4954), .Z(n4945) );
  AND U4986 ( .A(n1856), .B(n1546), .Z(n4954) );
  XOR U4987 ( .A(n4942), .B(g_input[13]), .Z(n4943) );
  NANDN U4988 ( .B(n4955), .A(n4956), .Z(n4942) );
  XOR U4989 ( .A(n4960), .B(n4946), .Z(n4953) );
  NAND U4990 ( .A(n1457), .B(n1953), .Z(n4946) );
  IV U4991 ( .A(n4948), .Z(n4960) );
  NAND U4992 ( .A(n1306), .B(n2276), .Z(n4952) );
  XNOR U4993 ( .A(n4950), .B(n4962), .Z(n4951) );
  AND U4994 ( .A(n2165), .B(n1376), .Z(n4962) );
  XNOR U4995 ( .A(n4957), .B(n4967), .Z(n4958) );
  AND U4996 ( .A(n1953), .B(n1546), .Z(n4967) );
  XNOR U4997 ( .A(n4956), .B(g_input[12]), .Z(n4955) );
  NOR U4998 ( .A(n4968), .B(n4969), .Z(n4956) );
  XOR U4999 ( .A(n4973), .B(n4959), .Z(n4966) );
  NAND U5000 ( .A(n1457), .B(n2058), .Z(n4959) );
  IV U5001 ( .A(n4961), .Z(n4973) );
  NAND U5002 ( .A(n1306), .B(n2392), .Z(n4965) );
  XNOR U5003 ( .A(n4963), .B(n4975), .Z(n4964) );
  AND U5004 ( .A(n2276), .B(n1376), .Z(n4975) );
  XNOR U5005 ( .A(n4970), .B(n4980), .Z(n4971) );
  AND U5006 ( .A(n2058), .B(n1546), .Z(n4980) );
  XOR U5007 ( .A(n4968), .B(g_input[11]), .Z(n4969) );
  NANDN U5008 ( .B(n4981), .A(n4982), .Z(n4968) );
  XOR U5009 ( .A(n4986), .B(n4972), .Z(n4979) );
  NAND U5010 ( .A(n1457), .B(n2165), .Z(n4972) );
  IV U5011 ( .A(n4974), .Z(n4986) );
  NAND U5012 ( .A(n1306), .B(n2513), .Z(n4978) );
  XNOR U5013 ( .A(n4976), .B(n4988), .Z(n4977) );
  AND U5014 ( .A(n2392), .B(n1376), .Z(n4988) );
  XNOR U5015 ( .A(n4983), .B(n4993), .Z(n4984) );
  AND U5016 ( .A(n2165), .B(n1546), .Z(n4993) );
  XNOR U5017 ( .A(n4982), .B(g_input[10]), .Z(n4981) );
  NOR U5018 ( .A(n4994), .B(n4995), .Z(n4982) );
  XOR U5019 ( .A(n4999), .B(n4985), .Z(n4992) );
  NAND U5020 ( .A(n1457), .B(n2276), .Z(n4985) );
  IV U5021 ( .A(n4987), .Z(n4999) );
  NAND U5022 ( .A(n1306), .B(n2635), .Z(n4991) );
  XNOR U5023 ( .A(n4989), .B(n5001), .Z(n4990) );
  AND U5024 ( .A(n2513), .B(n1376), .Z(n5001) );
  XNOR U5025 ( .A(n4996), .B(n5006), .Z(n4997) );
  AND U5026 ( .A(n2276), .B(n1546), .Z(n5006) );
  XOR U5027 ( .A(n4994), .B(g_input[9]), .Z(n4995) );
  NANDN U5028 ( .B(n5007), .A(n5008), .Z(n4994) );
  XOR U5029 ( .A(n5012), .B(n4998), .Z(n5005) );
  NAND U5030 ( .A(n1457), .B(n2392), .Z(n4998) );
  IV U5031 ( .A(n5000), .Z(n5012) );
  NAND U5032 ( .A(n1306), .B(n2763), .Z(n5004) );
  XNOR U5033 ( .A(n5002), .B(n5014), .Z(n5003) );
  AND U5034 ( .A(n2635), .B(n1376), .Z(n5014) );
  XNOR U5035 ( .A(n5018), .B(n5015), .Z(n5017) );
  XNOR U5036 ( .A(n5009), .B(n5020), .Z(n5010) );
  AND U5037 ( .A(n2392), .B(n1546), .Z(n5020) );
  XNOR U5038 ( .A(n5024), .B(n5021), .Z(n5023) );
  XOR U5039 ( .A(n5025), .B(n5011), .Z(n5019) );
  NAND U5040 ( .A(n1457), .B(n2513), .Z(n5011) );
  IV U5041 ( .A(n5013), .Z(n5025) );
  XNOR U5042 ( .A(n5026), .B(n5027), .Z(n5013) );
  AND U5043 ( .A(n5028), .B(n5029), .Z(n5027) );
  XOR U5044 ( .A(n5022), .B(n5030), .Z(n5029) );
  XNOR U5045 ( .A(n5024), .B(n5026), .Z(n5030) );
  NAND U5046 ( .A(n1457), .B(n2635), .Z(n5024) );
  XOR U5047 ( .A(n5021), .B(n5031), .Z(n5022) );
  AND U5048 ( .A(n2513), .B(n1546), .Z(n5031) );
  XNOR U5049 ( .A(n5035), .B(n5032), .Z(n5034) );
  XOR U5050 ( .A(n5016), .B(n5036), .Z(n5028) );
  XNOR U5051 ( .A(n5018), .B(n5026), .Z(n5036) );
  NANDN U5052 ( .B(n2892), .A(n1306), .Z(n5018) );
  XOR U5053 ( .A(n5015), .B(n5037), .Z(n5016) );
  AND U5054 ( .A(n2763), .B(n1376), .Z(n5037) );
  XNOR U5055 ( .A(n5041), .B(n5038), .Z(n5040) );
  XOR U5056 ( .A(n5042), .B(n5043), .Z(n5026) );
  AND U5057 ( .A(n5044), .B(n5045), .Z(n5043) );
  XOR U5058 ( .A(n5033), .B(n5046), .Z(n5045) );
  XNOR U5059 ( .A(n5035), .B(n5042), .Z(n5046) );
  NAND U5060 ( .A(n1457), .B(n2763), .Z(n5035) );
  XOR U5061 ( .A(n5032), .B(n5047), .Z(n5033) );
  AND U5062 ( .A(n2635), .B(n1546), .Z(n5047) );
  XNOR U5063 ( .A(n5051), .B(n5048), .Z(n5050) );
  XOR U5064 ( .A(n5039), .B(n5052), .Z(n5044) );
  XNOR U5065 ( .A(n5041), .B(n5042), .Z(n5052) );
  NANDN U5066 ( .B(n3030), .A(n1306), .Z(n5041) );
  XOR U5067 ( .A(n5038), .B(n5053), .Z(n5039) );
  ANDN U5068 ( .A(n1376), .B(n2892), .Z(n5053) );
  XNOR U5069 ( .A(n5057), .B(n5054), .Z(n5056) );
  XOR U5070 ( .A(n5058), .B(n5059), .Z(n5042) );
  AND U5071 ( .A(n5060), .B(n5061), .Z(n5059) );
  XOR U5072 ( .A(n5049), .B(n5062), .Z(n5061) );
  XNOR U5073 ( .A(n5051), .B(n5058), .Z(n5062) );
  NANDN U5074 ( .B(n2892), .A(n1457), .Z(n5051) );
  XOR U5075 ( .A(n5048), .B(n5063), .Z(n5049) );
  AND U5076 ( .A(n2763), .B(n1546), .Z(n5063) );
  XOR U5077 ( .A(n5055), .B(n5067), .Z(n5060) );
  XNOR U5078 ( .A(n5057), .B(n5058), .Z(n5067) );
  NAND U5079 ( .A(n1306), .B(n3165), .Z(n5057) );
  XOR U5080 ( .A(n5054), .B(n5068), .Z(n5055) );
  ANDN U5081 ( .A(n1376), .B(n3030), .Z(n5068) );
  NAND U5082 ( .A(n1306), .B(n3854), .Z(n5071) );
  XNOR U5083 ( .A(n5069), .B(n5073), .Z(n5070) );
  AND U5084 ( .A(n3165), .B(n1376), .Z(n5073) );
  AND U5085 ( .A(n5074), .B(\_MAC/_MULT/A__[0] ), .Z(n5069) );
  NANDN U5086 ( .B(n1306), .A(n5075), .Z(n5074) );
  NAND U5087 ( .A(n3854), .B(n1376), .Z(n5075) );
  XNOR U5088 ( .A(n5064), .B(n5079), .Z(n5065) );
  ANDN U5089 ( .A(n1546), .B(n2892), .Z(n5079) );
  XOR U5090 ( .A(n5082), .B(n5080), .Z(n5081) );
  ANDN U5091 ( .A(n1546), .B(n3030), .Z(n5082) );
  AND U5092 ( .A(n3165), .B(n1457), .Z(n5083) );
  XOR U5093 ( .A(n5087), .B(n5066), .Z(n5078) );
  NANDN U5094 ( .B(n3030), .A(n1457), .Z(n5066) );
  IV U5095 ( .A(n5072), .Z(n5087) );
  NAND U5096 ( .A(n1457), .B(n3854), .Z(n5086) );
  XNOR U5097 ( .A(n5084), .B(n5088), .Z(n5085) );
  AND U5098 ( .A(n3165), .B(n1546), .Z(n5088) );
  AND U5099 ( .A(n5089), .B(\_MAC/_MULT/A__[0] ), .Z(n5084) );
  NANDN U5100 ( .B(n1457), .A(n5090), .Z(n5089) );
  NAND U5101 ( .A(n3854), .B(n1546), .Z(n5090) );
  XNOR U5102 ( .A(n5093), .B(n3155), .Z(n3145) );
  XNOR U5103 ( .A(n3142), .B(n3143), .Z(n3155) );
  NANDN U5104 ( .B(n856), .A(n2763), .Z(n3143) );
  XNOR U5105 ( .A(n3141), .B(n5094), .Z(n3142) );
  AND U5106 ( .A(n2635), .B(n894), .Z(n5094) );
  XNOR U5107 ( .A(n5098), .B(n5095), .Z(n5097) );
  XNOR U5108 ( .A(n3154), .B(n3144), .Z(n5093) );
  XOR U5109 ( .A(n5099), .B(n5100), .Z(n3144) );
  XNOR U5110 ( .A(n3149), .B(n5102), .Z(n3150) );
  AND U5111 ( .A(n2392), .B(n1002), .Z(n5102) );
  XNOR U5112 ( .A(n5008), .B(g_input[8]), .Z(n5007) );
  NOR U5113 ( .A(n5103), .B(n5104), .Z(n5008) );
  XNOR U5114 ( .A(n5108), .B(n5105), .Z(n5107) );
  XOR U5115 ( .A(n5109), .B(n3151), .Z(n5101) );
  NAND U5116 ( .A(n948), .B(n2513), .Z(n3151) );
  IV U5117 ( .A(n3153), .Z(n5109) );
  XNOR U5118 ( .A(n5110), .B(n5111), .Z(n3153) );
  AND U5119 ( .A(n5112), .B(n5113), .Z(n5111) );
  XOR U5120 ( .A(n5106), .B(n5114), .Z(n5113) );
  XNOR U5121 ( .A(n5108), .B(n5110), .Z(n5114) );
  NAND U5122 ( .A(n948), .B(n2635), .Z(n5108) );
  XOR U5123 ( .A(n5105), .B(n5115), .Z(n5106) );
  AND U5124 ( .A(n2513), .B(n1002), .Z(n5115) );
  XOR U5125 ( .A(n5103), .B(g_input[7]), .Z(n5104) );
  NANDN U5126 ( .B(n5116), .A(n5117), .Z(n5103) );
  XNOR U5127 ( .A(n5121), .B(n5118), .Z(n5120) );
  XOR U5128 ( .A(n5096), .B(n5122), .Z(n5112) );
  XNOR U5129 ( .A(n5098), .B(n5110), .Z(n5122) );
  OR U5130 ( .A(n856), .B(n2892), .Z(n5098) );
  XOR U5131 ( .A(n5095), .B(n5123), .Z(n5096) );
  AND U5132 ( .A(n2763), .B(n894), .Z(n5123) );
  XNOR U5133 ( .A(n5127), .B(n5124), .Z(n5126) );
  XOR U5134 ( .A(n5128), .B(n5129), .Z(n5110) );
  AND U5135 ( .A(n5130), .B(n5131), .Z(n5129) );
  XOR U5136 ( .A(n5119), .B(n5132), .Z(n5131) );
  XNOR U5137 ( .A(n5121), .B(n5128), .Z(n5132) );
  NAND U5138 ( .A(n948), .B(n2763), .Z(n5121) );
  XOR U5139 ( .A(n5118), .B(n5133), .Z(n5119) );
  AND U5140 ( .A(n2635), .B(n1002), .Z(n5133) );
  XNOR U5141 ( .A(n5117), .B(g_input[6]), .Z(n5116) );
  NOR U5142 ( .A(n5134), .B(n5135), .Z(n5117) );
  XNOR U5143 ( .A(n5139), .B(n5136), .Z(n5138) );
  XOR U5144 ( .A(n5125), .B(n5140), .Z(n5130) );
  XNOR U5145 ( .A(n5127), .B(n5128), .Z(n5140) );
  OR U5146 ( .A(n856), .B(n3030), .Z(n5127) );
  XOR U5147 ( .A(n5124), .B(n5141), .Z(n5125) );
  ANDN U5148 ( .A(n894), .B(n2892), .Z(n5141) );
  XNOR U5149 ( .A(n5145), .B(n5142), .Z(n5144) );
  XOR U5150 ( .A(n5146), .B(n5147), .Z(n5128) );
  AND U5151 ( .A(n5148), .B(n5149), .Z(n5147) );
  XOR U5152 ( .A(n5137), .B(n5150), .Z(n5149) );
  XNOR U5153 ( .A(n5139), .B(n5146), .Z(n5150) );
  NANDN U5154 ( .B(n2892), .A(n948), .Z(n5139) );
  XOR U5155 ( .A(n5136), .B(n5151), .Z(n5137) );
  AND U5156 ( .A(n2763), .B(n1002), .Z(n5151) );
  XOR U5157 ( .A(n5134), .B(g_input[5]), .Z(n5135) );
  NANDN U5158 ( .B(n5152), .A(n5153), .Z(n5134) );
  XOR U5159 ( .A(n5143), .B(n5157), .Z(n5148) );
  XNOR U5160 ( .A(n5145), .B(n5146), .Z(n5157) );
  NANDN U5161 ( .B(n856), .A(n3165), .Z(n5145) );
  XOR U5162 ( .A(n5142), .B(n5158), .Z(n5143) );
  ANDN U5163 ( .A(n894), .B(n3030), .Z(n5158) );
  NANDN U5164 ( .B(n856), .A(n3854), .Z(n5161) );
  XNOR U5165 ( .A(n5159), .B(n5163), .Z(n5160) );
  AND U5166 ( .A(n3165), .B(n894), .Z(n5163) );
  AND U5167 ( .A(n5164), .B(\_MAC/_MULT/A__[0] ), .Z(n5159) );
  NAND U5168 ( .A(n5165), .B(n856), .Z(n5164) );
  NAND U5169 ( .A(n3854), .B(n894), .Z(n5165) );
  XNOR U5170 ( .A(n5154), .B(n5169), .Z(n5155) );
  ANDN U5171 ( .A(n1002), .B(n2892), .Z(n5169) );
  XOR U5172 ( .A(n5172), .B(n5170), .Z(n5171) );
  ANDN U5173 ( .A(n1002), .B(n3030), .Z(n5172) );
  AND U5174 ( .A(n3165), .B(n948), .Z(n5173) );
  XOR U5175 ( .A(n5177), .B(n5156), .Z(n5168) );
  NANDN U5176 ( .B(n3030), .A(n948), .Z(n5156) );
  IV U5177 ( .A(n5162), .Z(n5177) );
  NAND U5178 ( .A(n948), .B(n3854), .Z(n5176) );
  XNOR U5179 ( .A(n5174), .B(n5178), .Z(n5175) );
  AND U5180 ( .A(n3165), .B(n1002), .Z(n5178) );
  AND U5181 ( .A(n5179), .B(\_MAC/_MULT/A__[0] ), .Z(n5174) );
  NANDN U5182 ( .B(n948), .A(n5180), .Z(n5179) );
  NAND U5183 ( .A(n3854), .B(n1002), .Z(n5180) );
  XNOR U5184 ( .A(n3158), .B(n5184), .Z(n3159) );
  ANDN U5185 ( .A(n830), .B(n2892), .Z(n5184) );
  XNOR U5186 ( .A(n5153), .B(g_input[4]), .Z(n5152) );
  NOR U5187 ( .A(n5185), .B(n5186), .Z(n5153) );
  XOR U5188 ( .A(n5189), .B(n5187), .Z(n5188) );
  ANDN U5189 ( .A(n830), .B(n3030), .Z(n5189) );
  AND U5190 ( .A(n3165), .B(n793), .Z(n5190) );
  XOR U5191 ( .A(n5194), .B(n3160), .Z(n5183) );
  NANDN U5192 ( .B(n3030), .A(n793), .Z(n3160) );
  NANDN U5193 ( .B(n5195), .A(n5196), .Z(n5185) );
  IV U5194 ( .A(n3162), .Z(n5194) );
  NAND U5195 ( .A(n793), .B(n3854), .Z(n5193) );
  XNOR U5196 ( .A(n5191), .B(n5197), .Z(n5192) );
  AND U5197 ( .A(n3165), .B(n830), .Z(n5197) );
  AND U5198 ( .A(n5198), .B(\_MAC/_MULT/A__[0] ), .Z(n5191) );
  NANDN U5199 ( .B(n793), .A(n5199), .Z(n5198) );
  NAND U5200 ( .A(n3854), .B(n830), .Z(n5199) );
  XNOR U5201 ( .A(n3169), .B(n3170), .Z(n3164) );
  NANDN U5202 ( .B(n737), .A(n3854), .Z(n3170) );
  XNOR U5203 ( .A(n3168), .B(n5202), .Z(n3169) );
  AND U5204 ( .A(n3165), .B(n767), .Z(n5202) );
  XNOR U5205 ( .A(n5196), .B(g_input[2]), .Z(n5195) );
  AND U5206 ( .A(n5204), .B(\_MAC/_MULT/A__[0] ), .Z(n3168) );
  NAND U5207 ( .A(n5205), .B(n737), .Z(n5204) );
  NANDN U5208 ( .B(n5206), .A(n5207), .Z(n737) );
  ANDN U5209 ( .A(e_input[31]), .B(n5208), .Z(n5207) );
  NAND U5210 ( .A(n3854), .B(n767), .Z(n5205) );
  XOR U5211 ( .A(n5208), .B(e_input[30]), .Z(n5206) );
  OR U5212 ( .A(n5201), .B(n5209), .Z(n5208) );
  XOR U5213 ( .A(n5209), .B(e_input[29]), .Z(n5201) );
  OR U5214 ( .A(n5200), .B(n5210), .Z(n5209) );
  XOR U5215 ( .A(n5210), .B(e_input[28]), .Z(n5200) );
  OR U5216 ( .A(n5166), .B(n5211), .Z(n5210) );
  XOR U5217 ( .A(n5211), .B(e_input[27]), .Z(n5166) );
  OR U5218 ( .A(n5167), .B(n5212), .Z(n5211) );
  XOR U5219 ( .A(n5212), .B(e_input[26]), .Z(n5167) );
  OR U5220 ( .A(n5182), .B(n5213), .Z(n5212) );
  XOR U5221 ( .A(n5213), .B(e_input[25]), .Z(n5182) );
  OR U5222 ( .A(n5181), .B(n5214), .Z(n5213) );
  XOR U5223 ( .A(n5214), .B(e_input[24]), .Z(n5181) );
  OR U5224 ( .A(n4910), .B(n5215), .Z(n5214) );
  XOR U5225 ( .A(n5215), .B(e_input[23]), .Z(n4910) );
  OR U5226 ( .A(n4911), .B(n5216), .Z(n5215) );
  XOR U5227 ( .A(n5216), .B(e_input[22]), .Z(n4911) );
  OR U5228 ( .A(n4906), .B(n5217), .Z(n5216) );
  XOR U5229 ( .A(n5217), .B(e_input[21]), .Z(n4906) );
  OR U5230 ( .A(n4905), .B(n5218), .Z(n5217) );
  XOR U5231 ( .A(n5218), .B(e_input[20]), .Z(n4905) );
  OR U5232 ( .A(n5077), .B(n5219), .Z(n5218) );
  XOR U5233 ( .A(n5219), .B(e_input[19]), .Z(n5077) );
  OR U5234 ( .A(n5076), .B(n5220), .Z(n5219) );
  XOR U5235 ( .A(n5220), .B(e_input[18]), .Z(n5076) );
  OR U5236 ( .A(n5092), .B(n5221), .Z(n5220) );
  XOR U5237 ( .A(n5221), .B(e_input[17]), .Z(n5092) );
  OR U5238 ( .A(n5091), .B(n5222), .Z(n5221) );
  XOR U5239 ( .A(n5222), .B(e_input[16]), .Z(n5091) );
  OR U5240 ( .A(n3894), .B(n5223), .Z(n5222) );
  XOR U5241 ( .A(n5223), .B(e_input[15]), .Z(n3894) );
  OR U5242 ( .A(n3893), .B(n5224), .Z(n5223) );
  XOR U5243 ( .A(n5224), .B(e_input[14]), .Z(n3893) );
  OR U5244 ( .A(n3889), .B(n5225), .Z(n5224) );
  XOR U5245 ( .A(n5225), .B(e_input[13]), .Z(n3889) );
  OR U5246 ( .A(n3888), .B(n5226), .Z(n5225) );
  XOR U5247 ( .A(n5226), .B(e_input[12]), .Z(n3888) );
  OR U5248 ( .A(n3859), .B(n5227), .Z(n5226) );
  XOR U5249 ( .A(n5227), .B(e_input[11]), .Z(n3859) );
  OR U5250 ( .A(n3858), .B(n5228), .Z(n5227) );
  XOR U5251 ( .A(n5228), .B(e_input[10]), .Z(n3858) );
  OR U5252 ( .A(n3874), .B(n5229), .Z(n5228) );
  XOR U5253 ( .A(n5229), .B(e_input[9]), .Z(n3874) );
  OR U5254 ( .A(n3873), .B(n5230), .Z(n5229) );
  XOR U5255 ( .A(n5230), .B(e_input[8]), .Z(n3873) );
  OR U5256 ( .A(n4346), .B(n5231), .Z(n5230) );
  XOR U5257 ( .A(n5231), .B(e_input[7]), .Z(n4346) );
  OR U5258 ( .A(n4345), .B(n5232), .Z(n5231) );
  XOR U5259 ( .A(n5232), .B(e_input[6]), .Z(n4345) );
  OR U5260 ( .A(n4341), .B(n5233), .Z(n5232) );
  XOR U5261 ( .A(n5233), .B(e_input[5]), .Z(n4341) );
  OR U5262 ( .A(n4340), .B(n5234), .Z(n5233) );
  XOR U5263 ( .A(n5234), .B(e_input[4]), .Z(n4340) );
  OR U5264 ( .A(n4705), .B(n5235), .Z(n5234) );
  XOR U5265 ( .A(n5235), .B(e_input[3]), .Z(n4705) );
  OR U5266 ( .A(n4704), .B(n5236), .Z(n5235) );
  XOR U5267 ( .A(n5236), .B(e_input[2]), .Z(n4704) );
  NANDN U5268 ( .B(\_MAC/_MULT/X__[0] ), .A(n4719), .Z(n5236) );
  XNOR U5269 ( .A(\_MAC/_MULT/X__[0] ), .B(e_input[1]), .Z(n4719) );
  XOR U5270 ( .A(\_MAC/_MULT/A__[0] ), .B(g_input[1]), .Z(n5203) );
endmodule

