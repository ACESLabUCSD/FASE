
module MxM_TG_W8_N10000 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n64 , \_MxM/n61 , \_MxM/n58 , \_MxM/n55 , \_MxM/n52 ,
         \_MxM/n49 , \_MxM/n46 , \_MxM/n43 , \_MxM/N31 , \_MxM/N30 ,
         \_MxM/N29 , \_MxM/N28 , \_MxM/N27 , \_MxM/N26 , \_MxM/N25 ,
         \_MxM/N24 , \_MxM/N23 , \_MxM/N22 , \_MxM/N21 , \_MxM/N20 ,
         \_MxM/N19 , \_MxM/N18 , \_MxM/N16 , \_MxM/N15 , \_MxM/N14 ,
         \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 ,
         \_MxM/N7 , \_MxM/N6 , \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/n[10] , \_MxM/n[11] ,
         \_MxM/n[12] , \_MxM/n[13] , \_MxM/Y1[0] , \_MxM/Y1[1] , \_MxM/Y1[2] ,
         \_MxM/Y1[3] , \_MxM/Y1[4] , \_MxM/Y1[5] , \_MxM/Y1[6] , \_MxM/Y1[7] ,
         \_MxM/Y0[7] , \_MxM/Y0[6] , \_MxM/Y0[5] , \_MxM/Y0[4] , \_MxM/Y0[3] ,
         \_MxM/Y0[2] , \_MxM/Y0[1] , \_MxM/Y0[0] , \_MxM/add_43/carry[13] ,
         \_MxM/add_43/carry[12] , \_MxM/add_43/carry[11] ,
         \_MxM/add_43/carry[10] , \_MxM/add_43/carry[9] ,
         \_MxM/add_43/carry[8] , \_MxM/add_43/carry[7] ,
         \_MxM/add_43/carry[6] , \_MxM/add_43/carry[5] ,
         \_MxM/add_43/carry[4] , \_MxM/add_43/carry[3] ,
         \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374;

  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n43 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n46 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n49 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n52 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n55 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n58 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n61 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n64 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[13]  ( .D(\_MxM/N31 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[13] ) );
  DFF \_MxM/n_reg[12]  ( .D(\_MxM/N30 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[12] ) );
  DFF \_MxM/n_reg[11]  ( .D(\_MxM/N29 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[11] ) );
  DFF \_MxM/n_reg[10]  ( .D(\_MxM/N28 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[10] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N27 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N26 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N25 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N24 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_43/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_43/carry[6] ), .COUT(\_MxM/add_43/carry[7] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_43/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_43/carry[7] ), .COUT(\_MxM/add_43/carry[8] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_43/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_43/carry[8] ), .COUT(\_MxM/add_43/carry[9] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_43/U1_1_9  ( .IN0(\_MxM/n[9] ), .IN1(\_MxM/add_43/carry[9] ), .COUT(\_MxM/add_43/carry[10] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_43/U1_1_10  ( .IN0(\_MxM/n[10] ), .IN1(
        \_MxM/add_43/carry[10] ), .COUT(\_MxM/add_43/carry[11] ), .SUM(
        \_MxM/N14 ) );
  HADDER \_MxM/add_43/U1_1_11  ( .IN0(\_MxM/n[11] ), .IN1(
        \_MxM/add_43/carry[11] ), .COUT(\_MxM/add_43/carry[12] ), .SUM(
        \_MxM/N15 ) );
  HADDER \_MxM/add_43/U1_1_12  ( .IN0(\_MxM/n[12] ), .IN1(
        \_MxM/add_43/carry[12] ), .COUT(\_MxM/add_43/carry[13] ), .SUM(
        \_MxM/N16 ) );
  MUX U1 ( .IN0(n1), .IN1(n227), .SEL(n228), .F(n273) );
  IV U2 ( .A(n295), .Z(n1) );
  MUX U3 ( .IN0(n243), .IN1(n258), .SEL(n245), .F(n237) );
  XOR U4 ( .A(n177), .B(n215), .Z(n178) );
  MUX U5 ( .IN0(e_input[5]), .IN1(n352), .SEL(e_input[7]), .F(n94) );
  XNOR U6 ( .A(n120), .B(n121), .Z(n119) );
  NAND U7 ( .A(n152), .B(n188), .Z(n187) );
  MUX U8 ( .IN0(n2), .IN1(n105), .SEL(n106), .F(n79) );
  IV U9 ( .A(\_MxM/Y0[3] ), .Z(n2) );
  XOR U10 ( .A(n329), .B(g_input[3]), .Z(n330) );
  XNOR U11 ( .A(n198), .B(n229), .Z(n199) );
  MUX U12 ( .IN0(e_input[3]), .IN1(n303), .SEL(e_input[7]), .F(n155) );
  MUX U13 ( .IN0(e_input[6]), .IN1(n357), .SEL(e_input[7]), .F(n77) );
  XNOR U14 ( .A(n161), .B(n131), .Z(n123) );
  MUX U15 ( .IN0(n158), .IN1(n3), .SEL(n159), .F(n115) );
  IV U16 ( .A(n160), .Z(n3) );
  MUX U17 ( .IN0(n4), .IN1(n79), .SEL(n80), .F(n50) );
  IV U18 ( .A(\_MxM/Y0[4] ), .Z(n4) );
  XNOR U19 ( .A(n316), .B(n317), .Z(n295) );
  MUX U20 ( .IN0(n249), .IN1(n267), .SEL(n251), .F(n222) );
  XOR U21 ( .A(n102), .B(n134), .Z(n103) );
  MUX U22 ( .IN0(n200), .IN1(n198), .SEL(n199), .F(n5) );
  IV U23 ( .A(n5), .Z(n157) );
  XNOR U24 ( .A(n213), .B(n212), .Z(n197) );
  NAND U25 ( .A(n96), .B(n126), .Z(n125) );
  XNOR U26 ( .A(n173), .B(n172), .Z(n160) );
  XNOR U27 ( .A(n124), .B(n123), .Z(n117) );
  XNOR U28 ( .A(n50), .B(n51), .Z(n32) );
  NOR U29 ( .A(g_input[0]), .B(n354), .Z(n344) );
  XOR U30 ( .A(n293), .B(n294), .Z(n227) );
  XNOR U31 ( .A(n325), .B(n206), .Z(n212) );
  MUX U32 ( .IN0(n98), .IN1(n119), .SEL(n97), .F(n66) );
  MUX U33 ( .IN0(g_input[6]), .IN1(n233), .SEL(g_input[7]), .F(n78) );
  MUX U34 ( .IN0(n6), .IN1(n117), .SEL(n116), .F(n90) );
  IV U35 ( .A(n115), .Z(n6) );
  MUX U36 ( .IN0(n7), .IN1(n139), .SEL(n140), .F(n105) );
  IV U37 ( .A(\_MxM/Y0[2] ), .Z(n7) );
  MUX U38 ( .IN0(\_MxM/Y0[6] ), .IN1(n32), .SEL(n31), .F(n29) );
  MUX U39 ( .IN0(g_input[1]), .IN1(n354), .SEL(g_input[7]), .F(n296) );
  MUX U40 ( .IN0(g_input[2]), .IN1(n343), .SEL(g_input[7]), .F(n214) );
  MUX U41 ( .IN0(g_input[3]), .IN1(n330), .SEL(g_input[7]), .F(n8) );
  IV U42 ( .A(n8), .Z(n174) );
  XNOR U43 ( .A(n201), .B(n166), .Z(n172) );
  MUX U44 ( .IN0(n192), .IN1(n9), .SEL(n191), .F(n152) );
  IV U45 ( .A(n190), .Z(n9) );
  AND U46 ( .A(n72), .B(n41), .Z(n71) );
  MUX U47 ( .IN0(n10), .IN1(n180), .SEL(n181), .F(n139) );
  IV U48 ( .A(\_MxM/Y0[1] ), .Z(n10) );
  XNOR U49 ( .A(n89), .B(n90), .Z(n109) );
  MUX U50 ( .IN0(\_MxM/Y0[7] ), .IN1(n29), .SEL(n30), .F(n11) );
  IV U51 ( .A(n11), .Z(n26) );
  MUX U52 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n12), .F(\_MxM/n64 ) );
  MUX U53 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n12), .F(\_MxM/n61 ) );
  MUX U54 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n12), .F(\_MxM/n58 ) );
  MUX U55 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n12), .F(\_MxM/n55 ) );
  MUX U56 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n12), .F(\_MxM/n52 ) );
  MUX U57 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n12), .F(\_MxM/n49 ) );
  IV U58 ( .A(n13), .Z(n12) );
  MUX U59 ( .IN0(o[6]), .IN1(\_MxM/Y1[6] ), .SEL(n13), .F(\_MxM/n46 ) );
  MUX U60 ( .IN0(o[7]), .IN1(\_MxM/Y1[7] ), .SEL(n13), .F(\_MxM/n43 ) );
  AND U61 ( .A(n14), .B(n15), .Z(n13) );
  AND U62 ( .A(n16), .B(n17), .Z(n15) );
  ANDN U63 ( .A(n18), .B(\_MxM/n[3] ), .Z(n17) );
  NOR U64 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n18) );
  ANDN U65 ( .A(n19), .B(\_MxM/n[13] ), .Z(n16) );
  NOR U66 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n19) );
  AND U67 ( .A(n20), .B(n21), .Z(n14) );
  ANDN U68 ( .A(n22), .B(\_MxM/n[10] ), .Z(n21) );
  ANDN U69 ( .A(n23), .B(n24), .Z(n20) );
  NOR U70 ( .A(\_MxM/n[0] ), .B(n25), .Z(n23) );
  XNOR U71 ( .A(n26), .B(n27), .Z(\_MxM/Y1[7] ) );
  XNOR U72 ( .A(\_MxM/Y0[7] ), .B(n28), .Z(n27) );
  XNOR U73 ( .A(n30), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XOR U74 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U75 ( .A(n31), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XOR U76 ( .A(n32), .B(n33), .Z(n31) );
  ANDN U77 ( .A(n28), .B(n34), .Z(n33) );
  NANDN U78 ( .B(n35), .A(n36), .Z(n28) );
  ANDN U79 ( .A(n37), .B(n34), .Z(n35) );
  NAND U80 ( .A(n38), .B(n39), .Z(n34) );
  OR U81 ( .A(n40), .B(n41), .Z(n39) );
  AND U82 ( .A(n42), .B(n43), .Z(n38) );
  OR U83 ( .A(n44), .B(n45), .Z(n43) );
  OR U84 ( .A(n46), .B(n47), .Z(n42) );
  NOR U85 ( .A(n48), .B(n49), .Z(n37) );
  ANDN U86 ( .A(n52), .B(n53), .Z(n51) );
  XOR U87 ( .A(\_MxM/Y0[5] ), .B(n54), .Z(n52) );
  XNOR U88 ( .A(n53), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U89 ( .A(n55), .B(n56), .Z(n53) );
  XNOR U90 ( .A(n54), .B(n57), .Z(n55) );
  AND U91 ( .A(n36), .B(n58), .Z(n57) );
  XOR U92 ( .A(n48), .B(n59), .Z(n58) );
  XOR U93 ( .A(n59), .B(n49), .Z(n48) );
  OR U94 ( .A(n60), .B(n61), .Z(n49) );
  IV U95 ( .A(n56), .Z(n59) );
  XNOR U96 ( .A(n47), .B(n46), .Z(n56) );
  OR U97 ( .A(n62), .B(n63), .Z(n46) );
  AND U98 ( .A(n64), .B(n65), .Z(n47) );
  XNOR U99 ( .A(n66), .B(n67), .Z(n65) );
  ANDN U100 ( .A(n68), .B(n69), .Z(n67) );
  XOR U101 ( .A(n66), .B(n70), .Z(n68) );
  XNOR U102 ( .A(n40), .B(n71), .Z(n64) );
  NAND U103 ( .A(n73), .B(n74), .Z(n41) );
  NANDN U104 ( .B(n75), .A(n76), .Z(n73) );
  NANDN U105 ( .B(n44), .A(n77), .Z(n72) );
  NANDN U106 ( .B(n45), .A(n78), .Z(n40) );
  IV U107 ( .A(n50), .Z(n54) );
  XNOR U108 ( .A(n80), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U109 ( .A(n82), .B(n83), .Z(n80) );
  XNOR U110 ( .A(n81), .B(n84), .Z(n82) );
  AND U111 ( .A(n36), .B(n85), .Z(n84) );
  XOR U112 ( .A(n60), .B(n86), .Z(n85) );
  XOR U113 ( .A(n86), .B(n61), .Z(n60) );
  OR U114 ( .A(n87), .B(n88), .Z(n61) );
  IV U115 ( .A(n83), .Z(n86) );
  XNOR U116 ( .A(n63), .B(n62), .Z(n83) );
  OR U117 ( .A(n89), .B(n90), .Z(n62) );
  XOR U118 ( .A(n70), .B(n69), .Z(n63) );
  XOR U119 ( .A(n66), .B(n91), .Z(n69) );
  AND U120 ( .A(n92), .B(n93), .Z(n91) );
  NANDN U121 ( .B(n44), .A(n94), .Z(n93) );
  OR U122 ( .A(n95), .B(n96), .Z(n92) );
  XOR U123 ( .A(n75), .B(n76), .Z(n70) );
  NANDN U124 ( .B(n45), .A(n99), .Z(n76) );
  XNOR U125 ( .A(n74), .B(n100), .Z(n75) );
  AND U126 ( .A(n78), .B(n77), .Z(n100) );
  ANDN U127 ( .A(n101), .B(n102), .Z(n74) );
  NANDN U128 ( .B(n103), .A(n104), .Z(n101) );
  IV U129 ( .A(n79), .Z(n81) );
  XNOR U130 ( .A(n106), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U131 ( .A(n108), .B(n109), .Z(n106) );
  XNOR U132 ( .A(n107), .B(n110), .Z(n108) );
  AND U133 ( .A(n36), .B(n111), .Z(n110) );
  XOR U134 ( .A(n87), .B(n112), .Z(n111) );
  XOR U135 ( .A(n112), .B(n88), .Z(n87) );
  OR U136 ( .A(n113), .B(n114), .Z(n88) );
  IV U137 ( .A(n109), .Z(n112) );
  XOR U138 ( .A(n98), .B(n97), .Z(n89) );
  XNOR U139 ( .A(n118), .B(n119), .Z(n97) );
  ANDN U140 ( .A(n122), .B(n123), .Z(n121) );
  XOR U141 ( .A(n120), .B(n124), .Z(n122) );
  XNOR U142 ( .A(n125), .B(n95), .Z(n118) );
  NAND U143 ( .A(n94), .B(n78), .Z(n95) );
  NANDN U144 ( .B(n44), .A(n127), .Z(n126) );
  XNOR U145 ( .A(n128), .B(n129), .Z(n96) );
  ANDN U146 ( .A(n130), .B(n131), .Z(n129) );
  XNOR U147 ( .A(n132), .B(n128), .Z(n130) );
  XOR U148 ( .A(n103), .B(n104), .Z(n98) );
  OR U149 ( .A(n133), .B(n45), .Z(n104) );
  AND U150 ( .A(n99), .B(n77), .Z(n134) );
  NAND U151 ( .A(n135), .B(n136), .Z(n102) );
  NANDN U152 ( .B(n137), .A(n138), .Z(n135) );
  IV U153 ( .A(n105), .Z(n107) );
  XNOR U154 ( .A(n140), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U155 ( .A(n141), .B(n142), .Z(n140) );
  XOR U156 ( .A(n139), .B(n143), .Z(n141) );
  AND U157 ( .A(n36), .B(n144), .Z(n143) );
  XOR U158 ( .A(n113), .B(n145), .Z(n144) );
  XOR U159 ( .A(n145), .B(n114), .Z(n113) );
  NANDN U160 ( .B(n146), .A(n147), .Z(n114) );
  IV U161 ( .A(n142), .Z(n145) );
  XOR U162 ( .A(n117), .B(n116), .Z(n142) );
  XNOR U163 ( .A(n115), .B(n148), .Z(n116) );
  AND U164 ( .A(n149), .B(n150), .Z(n148) );
  OR U165 ( .A(n151), .B(n152), .Z(n150) );
  AND U166 ( .A(n153), .B(n154), .Z(n149) );
  NANDN U167 ( .B(n44), .A(n155), .Z(n154) );
  NAND U168 ( .A(n156), .B(n157), .Z(n153) );
  XNOR U169 ( .A(n128), .B(n162), .Z(n131) );
  AND U170 ( .A(n78), .B(n127), .Z(n162) );
  XOR U171 ( .A(n163), .B(n164), .Z(n128) );
  ANDN U172 ( .A(n165), .B(n166), .Z(n164) );
  XNOR U173 ( .A(n167), .B(n163), .Z(n165) );
  XOR U174 ( .A(n168), .B(n132), .Z(n161) );
  NAND U175 ( .A(n94), .B(n99), .Z(n132) );
  IV U176 ( .A(n120), .Z(n168) );
  XOR U177 ( .A(n169), .B(n170), .Z(n120) );
  ANDN U178 ( .A(n171), .B(n172), .Z(n170) );
  XOR U179 ( .A(n169), .B(n173), .Z(n171) );
  XNOR U180 ( .A(n137), .B(n138), .Z(n124) );
  OR U181 ( .A(n174), .B(n45), .Z(n138) );
  XNOR U182 ( .A(n136), .B(n175), .Z(n137) );
  ANDN U183 ( .A(n77), .B(n133), .Z(n175) );
  ANDN U184 ( .A(n176), .B(n177), .Z(n136) );
  NANDN U185 ( .B(n178), .A(n179), .Z(n176) );
  XNOR U186 ( .A(n181), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U187 ( .A(n182), .B(n183), .Z(n181) );
  XNOR U188 ( .A(n184), .B(n180), .Z(n182) );
  NAND U189 ( .A(\_MxM/Y0[0] ), .B(n146), .Z(n180) );
  NAND U190 ( .A(n185), .B(n36), .Z(n184) );
  XOR U191 ( .A(e_input[7]), .B(g_input[7]), .Z(n36) );
  XNOR U192 ( .A(n147), .B(n183), .Z(n185) );
  XNOR U193 ( .A(n146), .B(n183), .Z(n147) );
  XNOR U194 ( .A(n160), .B(n159), .Z(n183) );
  XNOR U195 ( .A(n186), .B(n156), .Z(n159) );
  XNOR U196 ( .A(n187), .B(n151), .Z(n156) );
  NAND U197 ( .A(n78), .B(n155), .Z(n151) );
  NANDN U198 ( .B(n44), .A(n189), .Z(n188) );
  XNOR U199 ( .A(n157), .B(n158), .Z(n186) );
  XOR U200 ( .A(n193), .B(n194), .Z(n158) );
  AND U201 ( .A(n195), .B(n196), .Z(n194) );
  XNOR U202 ( .A(n193), .B(n197), .Z(n196) );
  XNOR U203 ( .A(n163), .B(n202), .Z(n166) );
  AND U204 ( .A(n99), .B(n127), .Z(n202) );
  XOR U205 ( .A(n203), .B(n204), .Z(n163) );
  ANDN U206 ( .A(n205), .B(n206), .Z(n204) );
  XNOR U207 ( .A(n207), .B(n203), .Z(n205) );
  XOR U208 ( .A(n208), .B(n167), .Z(n201) );
  NANDN U209 ( .B(n133), .A(n94), .Z(n167) );
  IV U210 ( .A(n169), .Z(n208) );
  XOR U211 ( .A(n209), .B(n210), .Z(n169) );
  ANDN U212 ( .A(n211), .B(n212), .Z(n210) );
  XOR U213 ( .A(n209), .B(n213), .Z(n211) );
  XNOR U214 ( .A(n178), .B(n179), .Z(n173) );
  NANDN U215 ( .B(n45), .A(n214), .Z(n179) );
  ANDN U216 ( .A(n77), .B(n174), .Z(n215) );
  NAND U217 ( .A(n216), .B(n217), .Z(n177) );
  NANDN U218 ( .B(n218), .A(n219), .Z(n216) );
  XNOR U219 ( .A(n197), .B(n195), .Z(n146) );
  XNOR U220 ( .A(n220), .B(n200), .Z(n195) );
  XNOR U221 ( .A(n191), .B(n192), .Z(n200) );
  NAND U222 ( .A(n99), .B(n155), .Z(n192) );
  XNOR U223 ( .A(n190), .B(n221), .Z(n191) );
  AND U224 ( .A(n189), .B(n78), .Z(n221) );
  XOR U225 ( .A(n222), .B(n223), .Z(n190) );
  AND U226 ( .A(n224), .B(n225), .Z(n223) );
  XNOR U227 ( .A(n226), .B(n222), .Z(n225) );
  XNOR U228 ( .A(n199), .B(n193), .Z(n220) );
  XOR U229 ( .A(n227), .B(n228), .Z(n193) );
  AND U230 ( .A(n230), .B(n231), .Z(n229) );
  NANDN U231 ( .B(n44), .A(n232), .Z(n231) );
  NANDN U232 ( .B(n233), .A(n234), .Z(n44) );
  AND U233 ( .A(n235), .B(g_input[7]), .Z(n234) );
  NANDN U234 ( .B(n236), .A(n237), .Z(n230) );
  XNOR U235 ( .A(n238), .B(n239), .Z(n198) );
  AND U236 ( .A(n240), .B(n241), .Z(n239) );
  XOR U237 ( .A(n237), .B(n242), .Z(n241) );
  XNOR U238 ( .A(n236), .B(n238), .Z(n242) );
  NAND U239 ( .A(n78), .B(n232), .Z(n236) );
  XNOR U240 ( .A(n246), .B(n243), .Z(n245) );
  XOR U241 ( .A(n224), .B(n247), .Z(n240) );
  XNOR U242 ( .A(n226), .B(n238), .Z(n247) );
  NANDN U243 ( .B(n133), .A(n155), .Z(n226) );
  XOR U244 ( .A(n222), .B(n248), .Z(n224) );
  AND U245 ( .A(n189), .B(n99), .Z(n248) );
  XNOR U246 ( .A(n252), .B(n249), .Z(n251) );
  XOR U247 ( .A(n253), .B(n254), .Z(n238) );
  AND U248 ( .A(n255), .B(n256), .Z(n254) );
  XOR U249 ( .A(n244), .B(n257), .Z(n256) );
  XNOR U250 ( .A(n246), .B(n253), .Z(n257) );
  NAND U251 ( .A(n99), .B(n232), .Z(n246) );
  XOR U252 ( .A(n243), .B(n258), .Z(n244) );
  AND U253 ( .A(n78), .B(e_input[0]), .Z(n258) );
  XNOR U254 ( .A(n235), .B(g_input[6]), .Z(n233) );
  NOR U255 ( .A(n259), .B(n260), .Z(n235) );
  XOR U256 ( .A(n261), .B(n262), .Z(n243) );
  AND U257 ( .A(n263), .B(n264), .Z(n262) );
  XNOR U258 ( .A(n265), .B(n261), .Z(n264) );
  XOR U259 ( .A(n250), .B(n266), .Z(n255) );
  XNOR U260 ( .A(n252), .B(n253), .Z(n266) );
  NANDN U261 ( .B(n174), .A(n155), .Z(n252) );
  XOR U262 ( .A(n249), .B(n267), .Z(n250) );
  ANDN U263 ( .A(n189), .B(n133), .Z(n267) );
  XOR U264 ( .A(n268), .B(n269), .Z(n249) );
  AND U265 ( .A(n270), .B(n271), .Z(n269) );
  XNOR U266 ( .A(n272), .B(n268), .Z(n271) );
  XOR U267 ( .A(n273), .B(n274), .Z(n253) );
  AND U268 ( .A(n275), .B(n276), .Z(n274) );
  XOR U269 ( .A(n263), .B(n277), .Z(n276) );
  XNOR U270 ( .A(n265), .B(n273), .Z(n277) );
  NANDN U271 ( .B(n133), .A(n232), .Z(n265) );
  XOR U272 ( .A(n261), .B(n278), .Z(n263) );
  AND U273 ( .A(n99), .B(e_input[0]), .Z(n278) );
  XNOR U274 ( .A(n279), .B(g_input[5]), .Z(n99) );
  NAND U275 ( .A(n280), .B(g_input[7]), .Z(n279) );
  XOR U276 ( .A(n260), .B(g_input[5]), .Z(n280) );
  XOR U277 ( .A(n259), .B(g_input[5]), .Z(n260) );
  NANDN U278 ( .B(n281), .A(n282), .Z(n259) );
  XOR U279 ( .A(n283), .B(n284), .Z(n261) );
  ANDN U280 ( .A(n285), .B(n286), .Z(n284) );
  XNOR U281 ( .A(n287), .B(n283), .Z(n285) );
  XOR U282 ( .A(n270), .B(n288), .Z(n275) );
  XNOR U283 ( .A(n272), .B(n273), .Z(n288) );
  NAND U284 ( .A(n155), .B(n214), .Z(n272) );
  XOR U285 ( .A(n268), .B(n289), .Z(n270) );
  ANDN U286 ( .A(n189), .B(n174), .Z(n289) );
  XOR U287 ( .A(n290), .B(n291), .Z(n268) );
  ANDN U288 ( .A(n292), .B(n293), .Z(n291) );
  XNOR U289 ( .A(n294), .B(n290), .Z(n292) );
  NAND U290 ( .A(n155), .B(n296), .Z(n294) );
  XNOR U291 ( .A(n290), .B(n297), .Z(n293) );
  AND U292 ( .A(n214), .B(n189), .Z(n297) );
  AND U293 ( .A(n298), .B(g_input[0]), .Z(n290) );
  NANDN U294 ( .B(n155), .A(n299), .Z(n298) );
  NAND U295 ( .A(n296), .B(n189), .Z(n299) );
  XNOR U296 ( .A(n300), .B(e_input[2]), .Z(n189) );
  NAND U297 ( .A(n301), .B(e_input[7]), .Z(n300) );
  XOR U298 ( .A(n302), .B(e_input[2]), .Z(n301) );
  XNOR U299 ( .A(n304), .B(n305), .Z(n228) );
  IV U300 ( .A(n286), .Z(n305) );
  XNOR U301 ( .A(n283), .B(n306), .Z(n286) );
  ANDN U302 ( .A(e_input[0]), .B(n133), .Z(n306) );
  XOR U303 ( .A(n307), .B(n308), .Z(n283) );
  AND U304 ( .A(n309), .B(n310), .Z(n308) );
  XOR U305 ( .A(n311), .B(n307), .Z(n310) );
  ANDN U306 ( .A(e_input[0]), .B(n174), .Z(n311) );
  XOR U307 ( .A(n312), .B(n307), .Z(n309) );
  AND U308 ( .A(n232), .B(n214), .Z(n312) );
  XOR U309 ( .A(n313), .B(n314), .Z(n307) );
  ANDN U310 ( .A(n315), .B(n316), .Z(n314) );
  XNOR U311 ( .A(n317), .B(n313), .Z(n315) );
  XOR U312 ( .A(n318), .B(n287), .Z(n304) );
  NANDN U313 ( .B(n174), .A(n232), .Z(n287) );
  IV U314 ( .A(n295), .Z(n318) );
  NAND U315 ( .A(n232), .B(n296), .Z(n317) );
  XNOR U316 ( .A(n313), .B(n319), .Z(n316) );
  AND U317 ( .A(n214), .B(e_input[0]), .Z(n319) );
  AND U318 ( .A(n320), .B(g_input[0]), .Z(n313) );
  NANDN U319 ( .B(n232), .A(n321), .Z(n320) );
  NAND U320 ( .A(n296), .B(e_input[0]), .Z(n321) );
  XNOR U321 ( .A(n322), .B(e_input[1]), .Z(n232) );
  NAND U322 ( .A(n323), .B(e_input[7]), .Z(n322) );
  XNOR U323 ( .A(e_input[1]), .B(n324), .Z(n323) );
  XNOR U324 ( .A(n203), .B(n326), .Z(n206) );
  ANDN U325 ( .A(n127), .B(n133), .Z(n326) );
  XOR U326 ( .A(n327), .B(g_input[4]), .Z(n133) );
  NAND U327 ( .A(n328), .B(g_input[7]), .Z(n327) );
  XOR U328 ( .A(n281), .B(g_input[4]), .Z(n328) );
  XNOR U329 ( .A(n282), .B(g_input[4]), .Z(n281) );
  NOR U330 ( .A(n329), .B(n330), .Z(n282) );
  XOR U331 ( .A(n331), .B(n332), .Z(n203) );
  AND U332 ( .A(n333), .B(n334), .Z(n332) );
  XOR U333 ( .A(n335), .B(n331), .Z(n334) );
  ANDN U334 ( .A(n127), .B(n174), .Z(n335) );
  XOR U335 ( .A(n336), .B(n331), .Z(n333) );
  AND U336 ( .A(n214), .B(n94), .Z(n336) );
  XOR U337 ( .A(n337), .B(n338), .Z(n331) );
  ANDN U338 ( .A(n339), .B(n340), .Z(n338) );
  XNOR U339 ( .A(n341), .B(n337), .Z(n339) );
  XOR U340 ( .A(n342), .B(n207), .Z(n325) );
  NANDN U341 ( .B(n174), .A(n94), .Z(n207) );
  NANDN U342 ( .B(n343), .A(n344), .Z(n329) );
  IV U343 ( .A(n209), .Z(n342) );
  XOR U344 ( .A(n345), .B(n341), .Z(n209) );
  NAND U345 ( .A(n94), .B(n296), .Z(n341) );
  IV U346 ( .A(n340), .Z(n345) );
  XNOR U347 ( .A(n337), .B(n346), .Z(n340) );
  AND U348 ( .A(n214), .B(n127), .Z(n346) );
  AND U349 ( .A(n347), .B(g_input[0]), .Z(n337) );
  NANDN U350 ( .B(n94), .A(n348), .Z(n347) );
  NAND U351 ( .A(n296), .B(n127), .Z(n348) );
  XNOR U352 ( .A(n349), .B(e_input[4]), .Z(n127) );
  NAND U353 ( .A(n350), .B(e_input[7]), .Z(n349) );
  XOR U354 ( .A(n351), .B(e_input[4]), .Z(n350) );
  XNOR U355 ( .A(n218), .B(n219), .Z(n213) );
  NANDN U356 ( .B(n45), .A(n296), .Z(n219) );
  XNOR U357 ( .A(n217), .B(n353), .Z(n218) );
  AND U358 ( .A(n214), .B(n77), .Z(n353) );
  XNOR U359 ( .A(n344), .B(g_input[2]), .Z(n343) );
  AND U360 ( .A(n355), .B(g_input[0]), .Z(n217) );
  NAND U361 ( .A(n356), .B(n45), .Z(n355) );
  NANDN U362 ( .B(n357), .A(n358), .Z(n45) );
  ANDN U363 ( .A(e_input[7]), .B(n359), .Z(n358) );
  NAND U364 ( .A(n296), .B(n77), .Z(n356) );
  XOR U365 ( .A(n359), .B(e_input[6]), .Z(n357) );
  OR U366 ( .A(n352), .B(n360), .Z(n359) );
  XOR U367 ( .A(n360), .B(e_input[5]), .Z(n352) );
  OR U368 ( .A(n351), .B(n361), .Z(n360) );
  XOR U369 ( .A(n361), .B(e_input[4]), .Z(n351) );
  OR U370 ( .A(n303), .B(n362), .Z(n361) );
  XOR U371 ( .A(n362), .B(e_input[3]), .Z(n303) );
  OR U372 ( .A(n302), .B(n363), .Z(n362) );
  XOR U373 ( .A(n363), .B(e_input[2]), .Z(n302) );
  NANDN U374 ( .B(e_input[0]), .A(n324), .Z(n363) );
  XNOR U375 ( .A(e_input[0]), .B(e_input[1]), .Z(n324) );
  XOR U376 ( .A(g_input[0]), .B(g_input[1]), .Z(n354) );
  AND U377 ( .A(n364), .B(n365), .Z(\_MxM/N31 ) );
  XOR U378 ( .A(\_MxM/n[13] ), .B(\_MxM/add_43/carry[13] ), .Z(n365) );
  AND U379 ( .A(\_MxM/N16 ), .B(n364), .Z(\_MxM/N30 ) );
  AND U380 ( .A(\_MxM/N15 ), .B(n364), .Z(\_MxM/N29 ) );
  AND U381 ( .A(\_MxM/N14 ), .B(n364), .Z(\_MxM/N28 ) );
  AND U382 ( .A(\_MxM/N13 ), .B(n364), .Z(\_MxM/N27 ) );
  AND U383 ( .A(\_MxM/N12 ), .B(n364), .Z(\_MxM/N26 ) );
  AND U384 ( .A(\_MxM/N11 ), .B(n364), .Z(\_MxM/N25 ) );
  AND U385 ( .A(\_MxM/N10 ), .B(n364), .Z(\_MxM/N24 ) );
  AND U386 ( .A(\_MxM/N9 ), .B(n364), .Z(\_MxM/N23 ) );
  AND U387 ( .A(\_MxM/N8 ), .B(n364), .Z(\_MxM/N22 ) );
  AND U388 ( .A(\_MxM/N7 ), .B(n364), .Z(\_MxM/N21 ) );
  AND U389 ( .A(\_MxM/N6 ), .B(n364), .Z(\_MxM/N20 ) );
  AND U390 ( .A(\_MxM/N5 ), .B(n364), .Z(\_MxM/N19 ) );
  NAND U391 ( .A(n366), .B(n367), .Z(n364) );
  AND U392 ( .A(n368), .B(n369), .Z(n367) );
  ANDN U393 ( .A(n22), .B(\_MxM/N18 ), .Z(n369) );
  NOR U394 ( .A(\_MxM/n[12] ), .B(\_MxM/n[11] ), .Z(n22) );
  AND U395 ( .A(\_MxM/n[10] ), .B(n370), .Z(n368) );
  NOR U396 ( .A(n24), .B(n25), .Z(n370) );
  OR U397 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n25) );
  OR U398 ( .A(\_MxM/n[5] ), .B(\_MxM/n[4] ), .Z(n24) );
  AND U399 ( .A(n371), .B(n372), .Z(n366) );
  AND U400 ( .A(\_MxM/n[2] ), .B(n373), .Z(n372) );
  AND U401 ( .A(\_MxM/n[1] ), .B(\_MxM/n[13] ), .Z(n373) );
  AND U402 ( .A(\_MxM/n[9] ), .B(n374), .Z(n371) );
  AND U403 ( .A(\_MxM/n[8] ), .B(\_MxM/n[3] ), .Z(n374) );
  IV U404 ( .A(\_MxM/n[0] ), .Z(\_MxM/N18 ) );
endmodule

