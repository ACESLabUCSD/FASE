
module MxM_TG_W8_N100 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n111 , \_MxM/n110 , \_MxM/n109 , \_MxM/n108 , \_MxM/n107 ,
         \_MxM/n106 , \_MxM/n105 , \_MxM/n104 , \_MxM/n103 , \_MxM/n102 ,
         \_MxM/n101 , \_MxM/n100 , \_MxM/n99 , \_MxM/n98 , \_MxM/n97 ,
         \_MxM/n96 , \_MxM/N18 , \_MxM/N17 , \_MxM/N16 , \_MxM/N15 ,
         \_MxM/N14 , \_MxM/N13 , \_MxM/N12 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 ,
         \_MxM/N7 , \_MxM/N6 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] ,
         \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/Y0[0] ,
         \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] , \_MxM/Y0[4] , \_MxM/Y0[5] ,
         \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/add_39/carry[6] ,
         \_MxM/add_39/carry[5] , \_MxM/add_39/carry[4] ,
         \_MxM/add_39/carry[3] , \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n96 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n97 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n98 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n99 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n100 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n101 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n102 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n103 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n104 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n105 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n106 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n107 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n108 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n109 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n110 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n111 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N14 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N13 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N12 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N10 ) );
  MUX U1 ( .IN0(g_input[3]), .IN1(n375), .SEL(g_input[7]), .F(n1) );
  IV U2 ( .A(n1), .Z(n224) );
  XNOR U3 ( .A(n385), .B(n386), .Z(n256) );
  MUX U4 ( .IN0(g_input[6]), .IN1(n281), .SEL(g_input[7]), .F(n130) );
  MUX U5 ( .IN0(n150), .IN1(n2), .SEL(n149), .F(n118) );
  IV U6 ( .A(n148), .Z(n2) );
  MUX U7 ( .IN0(n208), .IN1(n3), .SEL(n209), .F(n167) );
  IV U8 ( .A(n210), .Z(n3) );
  MUX U9 ( .IN0(n4), .IN1(n131), .SEL(n50), .F(n99) );
  IV U10 ( .A(\_MxM/Y0[4] ), .Z(n4) );
  MUX U11 ( .IN0(n5), .IN1(n274), .SEL(n275), .F(n322) );
  IV U12 ( .A(n344), .Z(n5) );
  MUX U13 ( .IN0(n311), .IN1(n327), .SEL(n313), .F(n291) );
  XOR U14 ( .A(n154), .B(n185), .Z(n155) );
  MUX U15 ( .IN0(e_input[2]), .IN1(n350), .SEL(e_input[7]), .F(n238) );
  XNOR U16 ( .A(n372), .B(n253), .Z(n259) );
  NAND U17 ( .A(n147), .B(n177), .Z(n176) );
  MUX U18 ( .IN0(n6), .IN1(n169), .SEL(n168), .F(n141) );
  IV U19 ( .A(n167), .Z(n6) );
  XNOR U20 ( .A(n99), .B(n100), .Z(n81) );
  MUX U21 ( .IN0(n7), .IN1(n190), .SEL(n44), .F(n157) );
  IV U22 ( .A(\_MxM/Y0[2] ), .Z(n7) );
  MUX U23 ( .IN0(e_input[1]), .IN1(n8), .SEL(e_input[7]), .F(n280) );
  IV U24 ( .A(n371), .Z(n8) );
  XOR U25 ( .A(n227), .B(n262), .Z(n228) );
  XOR U26 ( .A(n170), .B(n148), .Z(n149) );
  MUX U27 ( .IN0(n241), .IN1(n9), .SEL(n240), .F(n202) );
  IV U28 ( .A(n239), .Z(n9) );
  MUX U29 ( .IN0(n242), .IN1(n10), .SEL(n243), .F(n208) );
  IV U30 ( .A(n244), .Z(n10) );
  XNOR U31 ( .A(n175), .B(n174), .Z(n169) );
  XOR U32 ( .A(n99), .B(n109), .Z(n107) );
  NOR U33 ( .A(g_input[0]), .B(n402), .Z(n391) );
  XNOR U34 ( .A(n365), .B(n366), .Z(n344) );
  MUX U35 ( .IN0(g_input[4]), .IN1(n330), .SEL(g_input[7]), .F(n11) );
  IV U36 ( .A(n11), .Z(n184) );
  XNOR U37 ( .A(n211), .B(n182), .Z(n174) );
  NAND U38 ( .A(n202), .B(n237), .Z(n236) );
  XNOR U39 ( .A(n260), .B(n259), .Z(n244) );
  XNOR U40 ( .A(n223), .B(n222), .Z(n210) );
  MUX U41 ( .IN0(\_MxM/Y0[6] ), .IN1(n81), .SEL(n76), .F(n70) );
  XOR U42 ( .A(n157), .B(n162), .Z(n160) );
  MUX U43 ( .IN0(g_input[2]), .IN1(n390), .SEL(g_input[7]), .F(n261) );
  XOR U44 ( .A(n354), .B(n335), .Z(n275) );
  XNOR U45 ( .A(n248), .B(n216), .Z(n222) );
  MUX U46 ( .IN0(n247), .IN1(n245), .SEL(n246), .F(n12) );
  IV U47 ( .A(n12), .Z(n207) );
  AND U48 ( .A(n124), .B(n90), .Z(n123) );
  XNOR U49 ( .A(n140), .B(n141), .Z(n161) );
  MUX U50 ( .IN0(n230), .IN1(n13), .SEL(n41), .F(n190) );
  IV U51 ( .A(\_MxM/Y0[1] ), .Z(n13) );
  MUX U52 ( .IN0(\_MxM/Y0[7] ), .IN1(n70), .SEL(n71), .F(n14) );
  IV U53 ( .A(n14), .Z(n67) );
  NAND U54 ( .A(\_MxM/Y0[4] ), .B(rst), .Z(n51) );
  NAND U55 ( .A(n15), .B(n16), .Z(\_MxM/n99 ) );
  NANDN U56 ( .B(n17), .A(o[3]), .Z(n16) );
  AND U57 ( .A(n18), .B(n19), .Z(n15) );
  NAND U58 ( .A(n20), .B(o[3]), .Z(n19) );
  NAND U59 ( .A(n21), .B(n22), .Z(n18) );
  NAND U60 ( .A(n23), .B(n24), .Z(\_MxM/n98 ) );
  NANDN U61 ( .B(n17), .A(o[2]), .Z(n24) );
  AND U62 ( .A(n25), .B(n26), .Z(n23) );
  NAND U63 ( .A(n20), .B(o[2]), .Z(n26) );
  NANDN U64 ( .B(n27), .A(n22), .Z(n25) );
  NAND U65 ( .A(n28), .B(n29), .Z(\_MxM/n97 ) );
  NANDN U66 ( .B(n17), .A(o[1]), .Z(n29) );
  AND U67 ( .A(n30), .B(n31), .Z(n28) );
  NAND U68 ( .A(n20), .B(o[1]), .Z(n31) );
  NANDN U69 ( .B(n32), .A(n22), .Z(n30) );
  NAND U70 ( .A(n33), .B(n34), .Z(\_MxM/n96 ) );
  NANDN U71 ( .B(n17), .A(o[0]), .Z(n34) );
  AND U72 ( .A(n35), .B(n36), .Z(n33) );
  NAND U73 ( .A(n20), .B(o[0]), .Z(n36) );
  NANDN U74 ( .B(n37), .A(n22), .Z(n35) );
  NAND U75 ( .A(n38), .B(n39), .Z(\_MxM/n111 ) );
  OR U76 ( .A(n37), .B(n40), .Z(n39) );
  XNOR U77 ( .A(n41), .B(\_MxM/Y0[1] ), .Z(n37) );
  NANDN U78 ( .B(n17), .A(\_MxM/Y0[0] ), .Z(n38) );
  NAND U79 ( .A(n42), .B(n43), .Z(\_MxM/n110 ) );
  OR U80 ( .A(n32), .B(n40), .Z(n43) );
  XOR U81 ( .A(n44), .B(\_MxM/Y0[2] ), .Z(n32) );
  NANDN U82 ( .B(n17), .A(\_MxM/Y0[1] ), .Z(n42) );
  NAND U83 ( .A(n45), .B(n46), .Z(\_MxM/n109 ) );
  OR U84 ( .A(n27), .B(n40), .Z(n46) );
  XOR U85 ( .A(n47), .B(\_MxM/Y0[3] ), .Z(n27) );
  NANDN U86 ( .B(n17), .A(\_MxM/Y0[2] ), .Z(n45) );
  NAND U87 ( .A(n48), .B(n49), .Z(\_MxM/n108 ) );
  NANDN U88 ( .B(n40), .A(n21), .Z(n49) );
  XNOR U89 ( .A(n50), .B(\_MxM/Y0[4] ), .Z(n21) );
  NANDN U90 ( .B(n17), .A(\_MxM/Y0[3] ), .Z(n48) );
  NAND U91 ( .A(n51), .B(n52), .Z(\_MxM/n107 ) );
  NANDN U92 ( .B(n40), .A(n53), .Z(n52) );
  NAND U93 ( .A(n54), .B(n55), .Z(\_MxM/n106 ) );
  NANDN U94 ( .B(n40), .A(n56), .Z(n55) );
  NANDN U95 ( .B(n17), .A(\_MxM/Y0[5] ), .Z(n54) );
  NAND U96 ( .A(n57), .B(n58), .Z(\_MxM/n105 ) );
  OR U97 ( .A(n59), .B(n40), .Z(n58) );
  NANDN U98 ( .B(n17), .A(\_MxM/Y0[6] ), .Z(n57) );
  NAND U99 ( .A(n60), .B(n61), .Z(\_MxM/n104 ) );
  OR U100 ( .A(n40), .B(n62), .Z(n61) );
  NANDN U101 ( .B(rst), .A(n20), .Z(n40) );
  NANDN U102 ( .B(n17), .A(\_MxM/Y0[7] ), .Z(n60) );
  NAND U103 ( .A(n63), .B(n64), .Z(\_MxM/n103 ) );
  NANDN U104 ( .B(n17), .A(o[7]), .Z(n64) );
  AND U105 ( .A(n65), .B(n66), .Z(n63) );
  NAND U106 ( .A(n20), .B(o[7]), .Z(n66) );
  NANDN U107 ( .B(n62), .A(n22), .Z(n65) );
  XOR U108 ( .A(n67), .B(n68), .Z(n62) );
  XNOR U109 ( .A(\_MxM/Y0[7] ), .B(n69), .Z(n68) );
  NAND U110 ( .A(n72), .B(n73), .Z(\_MxM/n102 ) );
  NANDN U111 ( .B(n17), .A(o[6]), .Z(n73) );
  AND U112 ( .A(n74), .B(n75), .Z(n72) );
  NAND U113 ( .A(n20), .B(o[6]), .Z(n75) );
  NANDN U114 ( .B(n59), .A(n22), .Z(n74) );
  XOR U115 ( .A(n71), .B(\_MxM/Y0[7] ), .Z(n59) );
  XOR U116 ( .A(n70), .B(n69), .Z(n71) );
  NAND U117 ( .A(n77), .B(n78), .Z(\_MxM/n101 ) );
  NANDN U118 ( .B(n17), .A(o[5]), .Z(n78) );
  AND U119 ( .A(n79), .B(n80), .Z(n77) );
  NAND U120 ( .A(n20), .B(o[5]), .Z(n80) );
  NAND U121 ( .A(n56), .B(n22), .Z(n79) );
  XNOR U122 ( .A(n76), .B(\_MxM/Y0[6] ), .Z(n56) );
  XOR U123 ( .A(n81), .B(n82), .Z(n76) );
  ANDN U124 ( .A(n69), .B(n83), .Z(n82) );
  NANDN U125 ( .B(n84), .A(n85), .Z(n69) );
  ANDN U126 ( .A(n86), .B(n83), .Z(n84) );
  NAND U127 ( .A(n87), .B(n88), .Z(n83) );
  OR U128 ( .A(n89), .B(n90), .Z(n88) );
  AND U129 ( .A(n91), .B(n92), .Z(n87) );
  OR U130 ( .A(n93), .B(n94), .Z(n92) );
  OR U131 ( .A(n95), .B(n96), .Z(n91) );
  NOR U132 ( .A(n97), .B(n98), .Z(n86) );
  ANDN U133 ( .A(n101), .B(n102), .Z(n100) );
  XNOR U134 ( .A(\_MxM/Y0[5] ), .B(n99), .Z(n101) );
  NAND U135 ( .A(n103), .B(n104), .Z(\_MxM/n100 ) );
  NANDN U136 ( .B(n17), .A(o[4]), .Z(n104) );
  IV U137 ( .A(rst), .Z(n17) );
  AND U138 ( .A(n105), .B(n106), .Z(n103) );
  NAND U139 ( .A(n20), .B(o[4]), .Z(n106) );
  NAND U140 ( .A(n22), .B(n53), .Z(n105) );
  XNOR U141 ( .A(n102), .B(\_MxM/Y0[5] ), .Z(n53) );
  XNOR U142 ( .A(n107), .B(n108), .Z(n102) );
  AND U143 ( .A(n85), .B(n110), .Z(n109) );
  XOR U144 ( .A(n97), .B(n111), .Z(n110) );
  XOR U145 ( .A(n111), .B(n98), .Z(n97) );
  OR U146 ( .A(n112), .B(n113), .Z(n98) );
  IV U147 ( .A(n108), .Z(n111) );
  XNOR U148 ( .A(n96), .B(n95), .Z(n108) );
  OR U149 ( .A(n114), .B(n115), .Z(n95) );
  AND U150 ( .A(n116), .B(n117), .Z(n96) );
  XNOR U151 ( .A(n118), .B(n119), .Z(n117) );
  ANDN U152 ( .A(n120), .B(n121), .Z(n119) );
  XOR U153 ( .A(n118), .B(n122), .Z(n120) );
  XNOR U154 ( .A(n89), .B(n123), .Z(n116) );
  NAND U155 ( .A(n125), .B(n126), .Z(n90) );
  NANDN U156 ( .B(n127), .A(n128), .Z(n125) );
  NANDN U157 ( .B(n93), .A(n129), .Z(n124) );
  NANDN U158 ( .B(n94), .A(n130), .Z(n89) );
  XNOR U159 ( .A(n132), .B(n133), .Z(n50) );
  XNOR U160 ( .A(n134), .B(n135), .Z(n132) );
  AND U161 ( .A(n85), .B(n136), .Z(n135) );
  XOR U162 ( .A(n112), .B(n137), .Z(n136) );
  XOR U163 ( .A(n137), .B(n113), .Z(n112) );
  OR U164 ( .A(n138), .B(n139), .Z(n113) );
  IV U165 ( .A(n133), .Z(n137) );
  XNOR U166 ( .A(n115), .B(n114), .Z(n133) );
  OR U167 ( .A(n140), .B(n141), .Z(n114) );
  XOR U168 ( .A(n122), .B(n121), .Z(n115) );
  XOR U169 ( .A(n118), .B(n142), .Z(n121) );
  AND U170 ( .A(n143), .B(n144), .Z(n142) );
  NANDN U171 ( .B(n93), .A(n145), .Z(n144) );
  OR U172 ( .A(n146), .B(n147), .Z(n143) );
  XOR U173 ( .A(n127), .B(n128), .Z(n122) );
  NANDN U174 ( .B(n94), .A(n151), .Z(n128) );
  XNOR U175 ( .A(n126), .B(n152), .Z(n127) );
  AND U176 ( .A(n130), .B(n129), .Z(n152) );
  ANDN U177 ( .A(n153), .B(n154), .Z(n126) );
  NANDN U178 ( .B(n155), .A(n156), .Z(n153) );
  IV U179 ( .A(n131), .Z(n134) );
  XOR U180 ( .A(n157), .B(n158), .Z(n131) );
  ANDN U181 ( .A(n159), .B(n47), .Z(n158) );
  XNOR U182 ( .A(n160), .B(n161), .Z(n47) );
  AND U183 ( .A(n85), .B(n163), .Z(n162) );
  XOR U184 ( .A(n138), .B(n164), .Z(n163) );
  XOR U185 ( .A(n164), .B(n139), .Z(n138) );
  OR U186 ( .A(n165), .B(n166), .Z(n139) );
  IV U187 ( .A(n161), .Z(n164) );
  XOR U188 ( .A(n150), .B(n149), .Z(n140) );
  XOR U189 ( .A(n171), .B(n172), .Z(n148) );
  ANDN U190 ( .A(n173), .B(n174), .Z(n172) );
  XOR U191 ( .A(n171), .B(n175), .Z(n173) );
  XNOR U192 ( .A(n176), .B(n146), .Z(n170) );
  NAND U193 ( .A(n145), .B(n130), .Z(n146) );
  NANDN U194 ( .B(n93), .A(n178), .Z(n177) );
  XNOR U195 ( .A(n179), .B(n180), .Z(n147) );
  ANDN U196 ( .A(n181), .B(n182), .Z(n180) );
  XNOR U197 ( .A(n183), .B(n179), .Z(n181) );
  XOR U198 ( .A(n155), .B(n156), .Z(n150) );
  OR U199 ( .A(n184), .B(n94), .Z(n156) );
  AND U200 ( .A(n151), .B(n129), .Z(n185) );
  NAND U201 ( .A(n186), .B(n187), .Z(n154) );
  NANDN U202 ( .B(n188), .A(n189), .Z(n186) );
  XNOR U203 ( .A(\_MxM/Y0[3] ), .B(n157), .Z(n159) );
  XNOR U204 ( .A(n191), .B(n192), .Z(n44) );
  XOR U205 ( .A(n190), .B(n193), .Z(n191) );
  AND U206 ( .A(n85), .B(n194), .Z(n193) );
  XOR U207 ( .A(n165), .B(n195), .Z(n194) );
  XOR U208 ( .A(n195), .B(n166), .Z(n165) );
  NANDN U209 ( .B(n196), .A(n197), .Z(n166) );
  IV U210 ( .A(n192), .Z(n195) );
  XOR U211 ( .A(n169), .B(n168), .Z(n192) );
  XNOR U212 ( .A(n167), .B(n198), .Z(n168) );
  AND U213 ( .A(n199), .B(n200), .Z(n198) );
  OR U214 ( .A(n201), .B(n202), .Z(n200) );
  AND U215 ( .A(n203), .B(n204), .Z(n199) );
  NANDN U216 ( .B(n93), .A(n205), .Z(n204) );
  NAND U217 ( .A(n206), .B(n207), .Z(n203) );
  XNOR U218 ( .A(n179), .B(n212), .Z(n182) );
  AND U219 ( .A(n130), .B(n178), .Z(n212) );
  XOR U220 ( .A(n213), .B(n214), .Z(n179) );
  ANDN U221 ( .A(n215), .B(n216), .Z(n214) );
  XNOR U222 ( .A(n217), .B(n213), .Z(n215) );
  XOR U223 ( .A(n218), .B(n183), .Z(n211) );
  NAND U224 ( .A(n145), .B(n151), .Z(n183) );
  IV U225 ( .A(n171), .Z(n218) );
  XOR U226 ( .A(n219), .B(n220), .Z(n171) );
  ANDN U227 ( .A(n221), .B(n222), .Z(n220) );
  XOR U228 ( .A(n219), .B(n223), .Z(n221) );
  XNOR U229 ( .A(n188), .B(n189), .Z(n175) );
  OR U230 ( .A(n224), .B(n94), .Z(n189) );
  XNOR U231 ( .A(n187), .B(n225), .Z(n188) );
  ANDN U232 ( .A(n129), .B(n184), .Z(n225) );
  ANDN U233 ( .A(n226), .B(n227), .Z(n187) );
  NANDN U234 ( .B(n228), .A(n229), .Z(n226) );
  XOR U235 ( .A(n231), .B(n232), .Z(n41) );
  XNOR U236 ( .A(n233), .B(n230), .Z(n231) );
  NAND U237 ( .A(n234), .B(n85), .Z(n233) );
  XOR U238 ( .A(e_input[7]), .B(g_input[7]), .Z(n85) );
  XNOR U239 ( .A(n196), .B(n232), .Z(n234) );
  XOR U240 ( .A(n197), .B(n232), .Z(n196) );
  XOR U241 ( .A(n210), .B(n209), .Z(n232) );
  XNOR U242 ( .A(n235), .B(n206), .Z(n209) );
  XNOR U243 ( .A(n236), .B(n201), .Z(n206) );
  NAND U244 ( .A(n130), .B(n205), .Z(n201) );
  NANDN U245 ( .B(n93), .A(n238), .Z(n237) );
  XNOR U246 ( .A(n207), .B(n208), .Z(n235) );
  XNOR U247 ( .A(n213), .B(n249), .Z(n216) );
  AND U248 ( .A(n151), .B(n178), .Z(n249) );
  XOR U249 ( .A(n250), .B(n251), .Z(n213) );
  ANDN U250 ( .A(n252), .B(n253), .Z(n251) );
  XNOR U251 ( .A(n254), .B(n250), .Z(n252) );
  XOR U252 ( .A(n255), .B(n217), .Z(n248) );
  NANDN U253 ( .B(n184), .A(n145), .Z(n217) );
  IV U254 ( .A(n219), .Z(n255) );
  XOR U255 ( .A(n256), .B(n257), .Z(n219) );
  ANDN U256 ( .A(n258), .B(n259), .Z(n257) );
  XOR U257 ( .A(n256), .B(n260), .Z(n258) );
  XNOR U258 ( .A(n228), .B(n229), .Z(n223) );
  NANDN U259 ( .B(n94), .A(n261), .Z(n229) );
  ANDN U260 ( .A(n129), .B(n224), .Z(n262) );
  NAND U261 ( .A(n263), .B(n264), .Z(n227) );
  NANDN U262 ( .B(n265), .A(n266), .Z(n263) );
  NANDN U263 ( .B(n197), .A(\_MxM/Y0[0] ), .Z(n230) );
  XOR U264 ( .A(n244), .B(n243), .Z(n197) );
  XNOR U265 ( .A(n267), .B(n247), .Z(n243) );
  XNOR U266 ( .A(n240), .B(n241), .Z(n247) );
  NAND U267 ( .A(n151), .B(n205), .Z(n241) );
  XNOR U268 ( .A(n239), .B(n268), .Z(n240) );
  AND U269 ( .A(n238), .B(n130), .Z(n268) );
  XOR U270 ( .A(n269), .B(n270), .Z(n239) );
  AND U271 ( .A(n271), .B(n272), .Z(n270) );
  XNOR U272 ( .A(n273), .B(n269), .Z(n272) );
  XNOR U273 ( .A(n246), .B(n242), .Z(n267) );
  XOR U274 ( .A(n274), .B(n275), .Z(n242) );
  XOR U275 ( .A(n276), .B(n277), .Z(n246) );
  AND U276 ( .A(n278), .B(n279), .Z(n277) );
  NANDN U277 ( .B(n93), .A(n280), .Z(n279) );
  NANDN U278 ( .B(n281), .A(n282), .Z(n93) );
  AND U279 ( .A(n283), .B(g_input[7]), .Z(n282) );
  NANDN U280 ( .B(n284), .A(n285), .Z(n278) );
  IV U281 ( .A(n245), .Z(n276) );
  XNOR U282 ( .A(n286), .B(n287), .Z(n245) );
  AND U283 ( .A(n288), .B(n289), .Z(n287) );
  XOR U284 ( .A(n285), .B(n290), .Z(n289) );
  XNOR U285 ( .A(n284), .B(n286), .Z(n290) );
  NAND U286 ( .A(n130), .B(n280), .Z(n284) );
  XOR U287 ( .A(n291), .B(n292), .Z(n285) );
  AND U288 ( .A(n293), .B(n294), .Z(n292) );
  XNOR U289 ( .A(n295), .B(n291), .Z(n294) );
  XOR U290 ( .A(n271), .B(n296), .Z(n288) );
  XNOR U291 ( .A(n273), .B(n286), .Z(n296) );
  NANDN U292 ( .B(n184), .A(n205), .Z(n273) );
  XOR U293 ( .A(n269), .B(n297), .Z(n271) );
  AND U294 ( .A(n238), .B(n151), .Z(n297) );
  XOR U295 ( .A(n298), .B(n299), .Z(n269) );
  AND U296 ( .A(n300), .B(n301), .Z(n299) );
  XNOR U297 ( .A(n302), .B(n298), .Z(n301) );
  XOR U298 ( .A(n303), .B(n304), .Z(n286) );
  AND U299 ( .A(n305), .B(n306), .Z(n304) );
  XOR U300 ( .A(n293), .B(n307), .Z(n306) );
  XNOR U301 ( .A(n295), .B(n303), .Z(n307) );
  NAND U302 ( .A(n151), .B(n280), .Z(n295) );
  XOR U303 ( .A(n291), .B(n308), .Z(n293) );
  AND U304 ( .A(n130), .B(e_input[0]), .Z(n308) );
  XNOR U305 ( .A(n283), .B(g_input[6]), .Z(n281) );
  NOR U306 ( .A(n309), .B(n310), .Z(n283) );
  XNOR U307 ( .A(n314), .B(n311), .Z(n313) );
  XOR U308 ( .A(n300), .B(n315), .Z(n305) );
  XNOR U309 ( .A(n302), .B(n303), .Z(n315) );
  NANDN U310 ( .B(n224), .A(n205), .Z(n302) );
  XOR U311 ( .A(n298), .B(n316), .Z(n300) );
  ANDN U312 ( .A(n238), .B(n184), .Z(n316) );
  XOR U313 ( .A(n317), .B(n318), .Z(n298) );
  AND U314 ( .A(n319), .B(n320), .Z(n318) );
  XNOR U315 ( .A(n321), .B(n317), .Z(n320) );
  XOR U316 ( .A(n322), .B(n323), .Z(n303) );
  AND U317 ( .A(n324), .B(n325), .Z(n323) );
  XOR U318 ( .A(n312), .B(n326), .Z(n325) );
  XNOR U319 ( .A(n314), .B(n322), .Z(n326) );
  NANDN U320 ( .B(n184), .A(n280), .Z(n314) );
  XOR U321 ( .A(n311), .B(n327), .Z(n312) );
  AND U322 ( .A(n151), .B(e_input[0]), .Z(n327) );
  XNOR U323 ( .A(n328), .B(g_input[5]), .Z(n151) );
  NAND U324 ( .A(n329), .B(g_input[7]), .Z(n328) );
  XOR U325 ( .A(n310), .B(g_input[5]), .Z(n329) );
  XOR U326 ( .A(n309), .B(g_input[5]), .Z(n310) );
  NANDN U327 ( .B(n330), .A(n331), .Z(n309) );
  XOR U328 ( .A(n332), .B(n333), .Z(n311) );
  ANDN U329 ( .A(n334), .B(n335), .Z(n333) );
  XNOR U330 ( .A(n336), .B(n332), .Z(n334) );
  XOR U331 ( .A(n319), .B(n337), .Z(n324) );
  XNOR U332 ( .A(n321), .B(n322), .Z(n337) );
  NAND U333 ( .A(n205), .B(n261), .Z(n321) );
  XOR U334 ( .A(n317), .B(n338), .Z(n319) );
  ANDN U335 ( .A(n238), .B(n224), .Z(n338) );
  XOR U336 ( .A(n339), .B(n340), .Z(n317) );
  ANDN U337 ( .A(n341), .B(n342), .Z(n340) );
  XNOR U338 ( .A(n343), .B(n339), .Z(n341) );
  XNOR U339 ( .A(n345), .B(n343), .Z(n274) );
  NAND U340 ( .A(n205), .B(n346), .Z(n343) );
  IV U341 ( .A(n342), .Z(n345) );
  XNOR U342 ( .A(n339), .B(n347), .Z(n342) );
  AND U343 ( .A(n261), .B(n238), .Z(n347) );
  AND U344 ( .A(n348), .B(g_input[0]), .Z(n339) );
  NANDN U345 ( .B(n205), .A(n349), .Z(n348) );
  NAND U346 ( .A(n346), .B(n238), .Z(n349) );
  XNOR U347 ( .A(n351), .B(e_input[3]), .Z(n205) );
  NAND U348 ( .A(n352), .B(e_input[7]), .Z(n351) );
  XOR U349 ( .A(n353), .B(e_input[3]), .Z(n352) );
  XNOR U350 ( .A(n332), .B(n355), .Z(n335) );
  ANDN U351 ( .A(e_input[0]), .B(n184), .Z(n355) );
  XOR U352 ( .A(n356), .B(n357), .Z(n332) );
  AND U353 ( .A(n358), .B(n359), .Z(n357) );
  XOR U354 ( .A(n360), .B(n356), .Z(n359) );
  ANDN U355 ( .A(e_input[0]), .B(n224), .Z(n360) );
  XOR U356 ( .A(n361), .B(n356), .Z(n358) );
  AND U357 ( .A(n280), .B(n261), .Z(n361) );
  XOR U358 ( .A(n362), .B(n363), .Z(n356) );
  ANDN U359 ( .A(n364), .B(n365), .Z(n363) );
  XNOR U360 ( .A(n366), .B(n362), .Z(n364) );
  XOR U361 ( .A(n367), .B(n336), .Z(n354) );
  NANDN U362 ( .B(n224), .A(n280), .Z(n336) );
  IV U363 ( .A(n344), .Z(n367) );
  NAND U364 ( .A(n280), .B(n346), .Z(n366) );
  XNOR U365 ( .A(n362), .B(n368), .Z(n365) );
  AND U366 ( .A(n261), .B(e_input[0]), .Z(n368) );
  AND U367 ( .A(n369), .B(g_input[0]), .Z(n362) );
  NANDN U368 ( .B(n280), .A(n370), .Z(n369) );
  NAND U369 ( .A(n346), .B(e_input[0]), .Z(n370) );
  XNOR U370 ( .A(n250), .B(n373), .Z(n253) );
  ANDN U371 ( .A(n178), .B(n184), .Z(n373) );
  XNOR U372 ( .A(n331), .B(g_input[4]), .Z(n330) );
  NOR U373 ( .A(n374), .B(n375), .Z(n331) );
  XOR U374 ( .A(n376), .B(n377), .Z(n250) );
  AND U375 ( .A(n378), .B(n379), .Z(n377) );
  XOR U376 ( .A(n380), .B(n376), .Z(n379) );
  ANDN U377 ( .A(n178), .B(n224), .Z(n380) );
  XOR U378 ( .A(n381), .B(n376), .Z(n378) );
  AND U379 ( .A(n261), .B(n145), .Z(n381) );
  XOR U380 ( .A(n382), .B(n383), .Z(n376) );
  ANDN U381 ( .A(n384), .B(n385), .Z(n383) );
  XNOR U382 ( .A(n386), .B(n382), .Z(n384) );
  XOR U383 ( .A(n387), .B(n254), .Z(n372) );
  NANDN U384 ( .B(n224), .A(n145), .Z(n254) );
  XOR U385 ( .A(n389), .B(n388), .Z(n375) );
  IV U386 ( .A(g_input[3]), .Z(n388) );
  IV U387 ( .A(n374), .Z(n389) );
  NANDN U388 ( .B(n390), .A(n391), .Z(n374) );
  IV U389 ( .A(n256), .Z(n387) );
  NAND U390 ( .A(n145), .B(n346), .Z(n386) );
  XNOR U391 ( .A(n382), .B(n392), .Z(n385) );
  AND U392 ( .A(n261), .B(n178), .Z(n392) );
  AND U393 ( .A(n393), .B(g_input[0]), .Z(n382) );
  NANDN U394 ( .B(n145), .A(n394), .Z(n393) );
  NAND U395 ( .A(n346), .B(n178), .Z(n394) );
  XNOR U396 ( .A(n395), .B(e_input[4]), .Z(n178) );
  NAND U397 ( .A(n396), .B(e_input[7]), .Z(n395) );
  XOR U398 ( .A(n397), .B(e_input[4]), .Z(n396) );
  XNOR U399 ( .A(n398), .B(e_input[5]), .Z(n145) );
  NAND U400 ( .A(n399), .B(e_input[7]), .Z(n398) );
  XOR U401 ( .A(n400), .B(e_input[5]), .Z(n399) );
  XNOR U402 ( .A(n265), .B(n266), .Z(n260) );
  NANDN U403 ( .B(n94), .A(n346), .Z(n266) );
  XNOR U404 ( .A(n264), .B(n401), .Z(n265) );
  AND U405 ( .A(n261), .B(n129), .Z(n401) );
  XNOR U406 ( .A(n391), .B(g_input[2]), .Z(n390) );
  AND U407 ( .A(n403), .B(g_input[0]), .Z(n264) );
  NAND U408 ( .A(n404), .B(n94), .Z(n403) );
  NANDN U409 ( .B(n405), .A(n406), .Z(n94) );
  ANDN U410 ( .A(e_input[7]), .B(n407), .Z(n406) );
  NAND U411 ( .A(n346), .B(n129), .Z(n404) );
  XNOR U412 ( .A(n408), .B(e_input[6]), .Z(n129) );
  NAND U413 ( .A(n409), .B(e_input[7]), .Z(n408) );
  XOR U414 ( .A(n405), .B(e_input[6]), .Z(n409) );
  XOR U415 ( .A(n407), .B(e_input[6]), .Z(n405) );
  OR U416 ( .A(n400), .B(n410), .Z(n407) );
  XOR U417 ( .A(n410), .B(e_input[5]), .Z(n400) );
  OR U418 ( .A(n397), .B(n411), .Z(n410) );
  XOR U419 ( .A(n411), .B(e_input[4]), .Z(n397) );
  OR U420 ( .A(n353), .B(n412), .Z(n411) );
  XOR U421 ( .A(n412), .B(e_input[3]), .Z(n353) );
  OR U422 ( .A(n350), .B(n413), .Z(n412) );
  XOR U423 ( .A(n413), .B(e_input[2]), .Z(n350) );
  NANDN U424 ( .B(e_input[0]), .A(n371), .Z(n413) );
  XNOR U425 ( .A(e_input[0]), .B(e_input[1]), .Z(n371) );
  XNOR U426 ( .A(n414), .B(g_input[1]), .Z(n346) );
  NAND U427 ( .A(n415), .B(g_input[7]), .Z(n414) );
  XOR U428 ( .A(g_input[1]), .B(n402), .Z(n415) );
  XOR U429 ( .A(g_input[0]), .B(g_input[1]), .Z(n402) );
  NOR U430 ( .A(rst), .B(n20), .Z(n22) );
  NAND U431 ( .A(n416), .B(n417), .Z(n20) );
  ANDN U432 ( .A(n418), .B(\_MxM/n[2] ), .Z(n417) );
  NOR U433 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n418) );
  ANDN U434 ( .A(n419), .B(n420), .Z(n416) );
  ANDN U435 ( .A(\_MxM/N12 ), .B(\_MxM/n[1] ), .Z(n419) );
  AND U436 ( .A(n421), .B(n422), .Z(\_MxM/N18 ) );
  XOR U437 ( .A(\_MxM/n[6] ), .B(\_MxM/add_39/carry[6] ), .Z(n422) );
  AND U438 ( .A(\_MxM/N10 ), .B(n421), .Z(\_MxM/N17 ) );
  AND U439 ( .A(\_MxM/N9 ), .B(n421), .Z(\_MxM/N16 ) );
  AND U440 ( .A(\_MxM/N8 ), .B(n421), .Z(\_MxM/N15 ) );
  AND U441 ( .A(\_MxM/N7 ), .B(n421), .Z(\_MxM/N14 ) );
  AND U442 ( .A(\_MxM/N6 ), .B(n421), .Z(\_MxM/N13 ) );
  NAND U443 ( .A(n423), .B(n424), .Z(n421) );
  ANDN U444 ( .A(n425), .B(n420), .Z(n424) );
  OR U445 ( .A(\_MxM/n[3] ), .B(\_MxM/n[4] ), .Z(n420) );
  NOR U446 ( .A(\_MxM/N12 ), .B(\_MxM/n[2] ), .Z(n425) );
  AND U447 ( .A(\_MxM/n[6] ), .B(n426), .Z(n423) );
  AND U448 ( .A(\_MxM/n[5] ), .B(\_MxM/n[1] ), .Z(n426) );
  IV U449 ( .A(\_MxM/n[0] ), .Z(\_MxM/N12 ) );
endmodule

