
module MxM_TG_W8_N1000 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n57 , \_MxM/n54 , \_MxM/n51 , \_MxM/n48 , \_MxM/n45 ,
         \_MxM/n42 , \_MxM/n39 , \_MxM/n36 , \_MxM/N23 , \_MxM/N22 ,
         \_MxM/N21 , \_MxM/N20 , \_MxM/N19 , \_MxM/N18 , \_MxM/N17 ,
         \_MxM/N16 , \_MxM/N15 , \_MxM/N14 , \_MxM/N12 , \_MxM/N11 ,
         \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/N7 , \_MxM/N6 , \_MxM/N5 ,
         \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] ,
         \_MxM/n[5] , \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] ,
         \_MxM/Y1[0] , \_MxM/Y1[1] , \_MxM/Y1[2] , \_MxM/Y1[3] , \_MxM/Y1[4] ,
         \_MxM/Y1[5] , \_MxM/Y1[6] , \_MxM/Y1[7] , \_MxM/Y0[7] , \_MxM/Y0[6] ,
         \_MxM/Y0[5] , \_MxM/Y0[4] , \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] ,
         \_MxM/Y0[0] , \_MxM/add_43/carry[9] , \_MxM/add_43/carry[8] ,
         \_MxM/add_43/carry[7] , \_MxM/add_43/carry[6] ,
         \_MxM/add_43/carry[5] , \_MxM/add_43/carry[4] ,
         \_MxM/add_43/carry[3] , \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368;

  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n36 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n39 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n42 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n45 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n48 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n51 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n54 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n57 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N14 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_43/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_43/carry[6] ), .COUT(\_MxM/add_43/carry[7] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_43/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_43/carry[7] ), .COUT(\_MxM/add_43/carry[8] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_43/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_43/carry[8] ), .COUT(\_MxM/add_43/carry[9] ), .SUM(\_MxM/N12 ) );
  MUX U1 ( .IN0(n1), .IN1(n223), .SEL(n224), .F(n269) );
  IV U2 ( .A(n291), .Z(n1) );
  MUX U3 ( .IN0(n239), .IN1(n254), .SEL(n241), .F(n233) );
  XOR U4 ( .A(n173), .B(n211), .Z(n174) );
  MUX U5 ( .IN0(e_input[5]), .IN1(n348), .SEL(e_input[7]), .F(n90) );
  XNOR U6 ( .A(n116), .B(n117), .Z(n115) );
  NAND U7 ( .A(n148), .B(n184), .Z(n183) );
  MUX U8 ( .IN0(n2), .IN1(n101), .SEL(n102), .F(n75) );
  IV U9 ( .A(\_MxM/Y0[3] ), .Z(n2) );
  XOR U10 ( .A(n325), .B(g_input[3]), .Z(n326) );
  XNOR U11 ( .A(n194), .B(n225), .Z(n195) );
  MUX U12 ( .IN0(e_input[3]), .IN1(n299), .SEL(e_input[7]), .F(n151) );
  MUX U13 ( .IN0(e_input[6]), .IN1(n353), .SEL(e_input[7]), .F(n73) );
  XNOR U14 ( .A(n157), .B(n127), .Z(n119) );
  MUX U15 ( .IN0(n154), .IN1(n3), .SEL(n155), .F(n111) );
  IV U16 ( .A(n156), .Z(n3) );
  MUX U17 ( .IN0(n4), .IN1(n75), .SEL(n76), .F(n46) );
  IV U18 ( .A(\_MxM/Y0[4] ), .Z(n4) );
  XNOR U19 ( .A(n312), .B(n313), .Z(n291) );
  MUX U20 ( .IN0(n245), .IN1(n263), .SEL(n247), .F(n218) );
  XOR U21 ( .A(n98), .B(n130), .Z(n99) );
  MUX U22 ( .IN0(n196), .IN1(n194), .SEL(n195), .F(n5) );
  IV U23 ( .A(n5), .Z(n153) );
  XNOR U24 ( .A(n209), .B(n208), .Z(n193) );
  NAND U25 ( .A(n92), .B(n122), .Z(n121) );
  XNOR U26 ( .A(n169), .B(n168), .Z(n156) );
  XNOR U27 ( .A(n120), .B(n119), .Z(n113) );
  XNOR U28 ( .A(n46), .B(n47), .Z(n28) );
  NOR U29 ( .A(g_input[0]), .B(n350), .Z(n340) );
  XOR U30 ( .A(n289), .B(n290), .Z(n223) );
  XNOR U31 ( .A(n321), .B(n202), .Z(n208) );
  MUX U32 ( .IN0(n94), .IN1(n115), .SEL(n93), .F(n62) );
  MUX U33 ( .IN0(g_input[6]), .IN1(n229), .SEL(g_input[7]), .F(n74) );
  MUX U34 ( .IN0(n6), .IN1(n113), .SEL(n112), .F(n86) );
  IV U35 ( .A(n111), .Z(n6) );
  MUX U36 ( .IN0(n7), .IN1(n135), .SEL(n136), .F(n101) );
  IV U37 ( .A(\_MxM/Y0[2] ), .Z(n7) );
  MUX U38 ( .IN0(\_MxM/Y0[6] ), .IN1(n28), .SEL(n27), .F(n25) );
  MUX U39 ( .IN0(g_input[1]), .IN1(n350), .SEL(g_input[7]), .F(n292) );
  MUX U40 ( .IN0(g_input[2]), .IN1(n339), .SEL(g_input[7]), .F(n210) );
  MUX U41 ( .IN0(g_input[3]), .IN1(n326), .SEL(g_input[7]), .F(n8) );
  IV U42 ( .A(n8), .Z(n170) );
  XNOR U43 ( .A(n197), .B(n162), .Z(n168) );
  MUX U44 ( .IN0(n188), .IN1(n9), .SEL(n187), .F(n148) );
  IV U45 ( .A(n186), .Z(n9) );
  AND U46 ( .A(n68), .B(n37), .Z(n67) );
  MUX U47 ( .IN0(n10), .IN1(n176), .SEL(n177), .F(n135) );
  IV U48 ( .A(\_MxM/Y0[1] ), .Z(n10) );
  XNOR U49 ( .A(n85), .B(n86), .Z(n105) );
  MUX U50 ( .IN0(\_MxM/Y0[7] ), .IN1(n25), .SEL(n26), .F(n11) );
  IV U51 ( .A(n11), .Z(n22) );
  MUX U52 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n12), .F(\_MxM/n57 ) );
  MUX U53 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n12), .F(\_MxM/n54 ) );
  MUX U54 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n12), .F(\_MxM/n51 ) );
  MUX U55 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n12), .F(\_MxM/n48 ) );
  MUX U56 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n12), .F(\_MxM/n45 ) );
  MUX U57 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n12), .F(\_MxM/n42 ) );
  IV U58 ( .A(n13), .Z(n12) );
  MUX U59 ( .IN0(o[6]), .IN1(\_MxM/Y1[6] ), .SEL(n13), .F(\_MxM/n39 ) );
  MUX U60 ( .IN0(o[7]), .IN1(\_MxM/Y1[7] ), .SEL(n13), .F(\_MxM/n36 ) );
  AND U61 ( .A(n14), .B(n15), .Z(n13) );
  AND U62 ( .A(n16), .B(n17), .Z(n15) );
  ANDN U63 ( .A(n18), .B(\_MxM/n[7] ), .Z(n17) );
  NOR U64 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n18) );
  NOR U65 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n16) );
  AND U66 ( .A(n19), .B(n20), .Z(n14) );
  NOR U67 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n20) );
  NOR U68 ( .A(\_MxM/n[0] ), .B(n21), .Z(n19) );
  XNOR U69 ( .A(n22), .B(n23), .Z(\_MxM/Y1[7] ) );
  XNOR U70 ( .A(\_MxM/Y0[7] ), .B(n24), .Z(n23) );
  XNOR U71 ( .A(n26), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XOR U72 ( .A(n25), .B(n24), .Z(n26) );
  XNOR U73 ( .A(n27), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XOR U74 ( .A(n28), .B(n29), .Z(n27) );
  ANDN U75 ( .A(n24), .B(n30), .Z(n29) );
  NANDN U76 ( .B(n31), .A(n32), .Z(n24) );
  ANDN U77 ( .A(n33), .B(n30), .Z(n31) );
  NAND U78 ( .A(n34), .B(n35), .Z(n30) );
  OR U79 ( .A(n36), .B(n37), .Z(n35) );
  AND U80 ( .A(n38), .B(n39), .Z(n34) );
  OR U81 ( .A(n40), .B(n41), .Z(n39) );
  OR U82 ( .A(n42), .B(n43), .Z(n38) );
  NOR U83 ( .A(n44), .B(n45), .Z(n33) );
  ANDN U84 ( .A(n48), .B(n49), .Z(n47) );
  XOR U85 ( .A(\_MxM/Y0[5] ), .B(n50), .Z(n48) );
  XNOR U86 ( .A(n49), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U87 ( .A(n51), .B(n52), .Z(n49) );
  XNOR U88 ( .A(n50), .B(n53), .Z(n51) );
  AND U89 ( .A(n32), .B(n54), .Z(n53) );
  XOR U90 ( .A(n44), .B(n55), .Z(n54) );
  XOR U91 ( .A(n55), .B(n45), .Z(n44) );
  OR U92 ( .A(n56), .B(n57), .Z(n45) );
  IV U93 ( .A(n52), .Z(n55) );
  XNOR U94 ( .A(n43), .B(n42), .Z(n52) );
  OR U95 ( .A(n58), .B(n59), .Z(n42) );
  AND U96 ( .A(n60), .B(n61), .Z(n43) );
  XNOR U97 ( .A(n62), .B(n63), .Z(n61) );
  ANDN U98 ( .A(n64), .B(n65), .Z(n63) );
  XOR U99 ( .A(n62), .B(n66), .Z(n64) );
  XNOR U100 ( .A(n36), .B(n67), .Z(n60) );
  NAND U101 ( .A(n69), .B(n70), .Z(n37) );
  NANDN U102 ( .B(n71), .A(n72), .Z(n69) );
  NANDN U103 ( .B(n40), .A(n73), .Z(n68) );
  NANDN U104 ( .B(n41), .A(n74), .Z(n36) );
  IV U105 ( .A(n46), .Z(n50) );
  XNOR U106 ( .A(n76), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U107 ( .A(n78), .B(n79), .Z(n76) );
  XNOR U108 ( .A(n77), .B(n80), .Z(n78) );
  AND U109 ( .A(n32), .B(n81), .Z(n80) );
  XOR U110 ( .A(n56), .B(n82), .Z(n81) );
  XOR U111 ( .A(n82), .B(n57), .Z(n56) );
  OR U112 ( .A(n83), .B(n84), .Z(n57) );
  IV U113 ( .A(n79), .Z(n82) );
  XNOR U114 ( .A(n59), .B(n58), .Z(n79) );
  OR U115 ( .A(n85), .B(n86), .Z(n58) );
  XOR U116 ( .A(n66), .B(n65), .Z(n59) );
  XOR U117 ( .A(n62), .B(n87), .Z(n65) );
  AND U118 ( .A(n88), .B(n89), .Z(n87) );
  NANDN U119 ( .B(n40), .A(n90), .Z(n89) );
  OR U120 ( .A(n91), .B(n92), .Z(n88) );
  XOR U121 ( .A(n71), .B(n72), .Z(n66) );
  NANDN U122 ( .B(n41), .A(n95), .Z(n72) );
  XNOR U123 ( .A(n70), .B(n96), .Z(n71) );
  AND U124 ( .A(n74), .B(n73), .Z(n96) );
  ANDN U125 ( .A(n97), .B(n98), .Z(n70) );
  NANDN U126 ( .B(n99), .A(n100), .Z(n97) );
  IV U127 ( .A(n75), .Z(n77) );
  XNOR U128 ( .A(n102), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U129 ( .A(n104), .B(n105), .Z(n102) );
  XNOR U130 ( .A(n103), .B(n106), .Z(n104) );
  AND U131 ( .A(n32), .B(n107), .Z(n106) );
  XOR U132 ( .A(n83), .B(n108), .Z(n107) );
  XOR U133 ( .A(n108), .B(n84), .Z(n83) );
  OR U134 ( .A(n109), .B(n110), .Z(n84) );
  IV U135 ( .A(n105), .Z(n108) );
  XOR U136 ( .A(n94), .B(n93), .Z(n85) );
  XNOR U137 ( .A(n114), .B(n115), .Z(n93) );
  ANDN U138 ( .A(n118), .B(n119), .Z(n117) );
  XOR U139 ( .A(n116), .B(n120), .Z(n118) );
  XNOR U140 ( .A(n121), .B(n91), .Z(n114) );
  NAND U141 ( .A(n90), .B(n74), .Z(n91) );
  NANDN U142 ( .B(n40), .A(n123), .Z(n122) );
  XNOR U143 ( .A(n124), .B(n125), .Z(n92) );
  ANDN U144 ( .A(n126), .B(n127), .Z(n125) );
  XNOR U145 ( .A(n128), .B(n124), .Z(n126) );
  XOR U146 ( .A(n99), .B(n100), .Z(n94) );
  OR U147 ( .A(n129), .B(n41), .Z(n100) );
  AND U148 ( .A(n95), .B(n73), .Z(n130) );
  NAND U149 ( .A(n131), .B(n132), .Z(n98) );
  NANDN U150 ( .B(n133), .A(n134), .Z(n131) );
  IV U151 ( .A(n101), .Z(n103) );
  XNOR U152 ( .A(n136), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U153 ( .A(n137), .B(n138), .Z(n136) );
  XOR U154 ( .A(n135), .B(n139), .Z(n137) );
  AND U155 ( .A(n32), .B(n140), .Z(n139) );
  XOR U156 ( .A(n109), .B(n141), .Z(n140) );
  XOR U157 ( .A(n141), .B(n110), .Z(n109) );
  NANDN U158 ( .B(n142), .A(n143), .Z(n110) );
  IV U159 ( .A(n138), .Z(n141) );
  XOR U160 ( .A(n113), .B(n112), .Z(n138) );
  XNOR U161 ( .A(n111), .B(n144), .Z(n112) );
  AND U162 ( .A(n145), .B(n146), .Z(n144) );
  OR U163 ( .A(n147), .B(n148), .Z(n146) );
  AND U164 ( .A(n149), .B(n150), .Z(n145) );
  NANDN U165 ( .B(n40), .A(n151), .Z(n150) );
  NAND U166 ( .A(n152), .B(n153), .Z(n149) );
  XNOR U167 ( .A(n124), .B(n158), .Z(n127) );
  AND U168 ( .A(n74), .B(n123), .Z(n158) );
  XOR U169 ( .A(n159), .B(n160), .Z(n124) );
  ANDN U170 ( .A(n161), .B(n162), .Z(n160) );
  XNOR U171 ( .A(n163), .B(n159), .Z(n161) );
  XOR U172 ( .A(n164), .B(n128), .Z(n157) );
  NAND U173 ( .A(n90), .B(n95), .Z(n128) );
  IV U174 ( .A(n116), .Z(n164) );
  XOR U175 ( .A(n165), .B(n166), .Z(n116) );
  ANDN U176 ( .A(n167), .B(n168), .Z(n166) );
  XOR U177 ( .A(n165), .B(n169), .Z(n167) );
  XNOR U178 ( .A(n133), .B(n134), .Z(n120) );
  OR U179 ( .A(n170), .B(n41), .Z(n134) );
  XNOR U180 ( .A(n132), .B(n171), .Z(n133) );
  ANDN U181 ( .A(n73), .B(n129), .Z(n171) );
  ANDN U182 ( .A(n172), .B(n173), .Z(n132) );
  NANDN U183 ( .B(n174), .A(n175), .Z(n172) );
  XNOR U184 ( .A(n177), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U185 ( .A(n178), .B(n179), .Z(n177) );
  XNOR U186 ( .A(n180), .B(n176), .Z(n178) );
  NAND U187 ( .A(\_MxM/Y0[0] ), .B(n142), .Z(n176) );
  NAND U188 ( .A(n181), .B(n32), .Z(n180) );
  XOR U189 ( .A(e_input[7]), .B(g_input[7]), .Z(n32) );
  XNOR U190 ( .A(n143), .B(n179), .Z(n181) );
  XNOR U191 ( .A(n142), .B(n179), .Z(n143) );
  XNOR U192 ( .A(n156), .B(n155), .Z(n179) );
  XNOR U193 ( .A(n182), .B(n152), .Z(n155) );
  XNOR U194 ( .A(n183), .B(n147), .Z(n152) );
  NAND U195 ( .A(n74), .B(n151), .Z(n147) );
  NANDN U196 ( .B(n40), .A(n185), .Z(n184) );
  XNOR U197 ( .A(n153), .B(n154), .Z(n182) );
  XOR U198 ( .A(n189), .B(n190), .Z(n154) );
  AND U199 ( .A(n191), .B(n192), .Z(n190) );
  XNOR U200 ( .A(n189), .B(n193), .Z(n192) );
  XNOR U201 ( .A(n159), .B(n198), .Z(n162) );
  AND U202 ( .A(n95), .B(n123), .Z(n198) );
  XOR U203 ( .A(n199), .B(n200), .Z(n159) );
  ANDN U204 ( .A(n201), .B(n202), .Z(n200) );
  XNOR U205 ( .A(n203), .B(n199), .Z(n201) );
  XOR U206 ( .A(n204), .B(n163), .Z(n197) );
  NANDN U207 ( .B(n129), .A(n90), .Z(n163) );
  IV U208 ( .A(n165), .Z(n204) );
  XOR U209 ( .A(n205), .B(n206), .Z(n165) );
  ANDN U210 ( .A(n207), .B(n208), .Z(n206) );
  XOR U211 ( .A(n205), .B(n209), .Z(n207) );
  XNOR U212 ( .A(n174), .B(n175), .Z(n169) );
  NANDN U213 ( .B(n41), .A(n210), .Z(n175) );
  ANDN U214 ( .A(n73), .B(n170), .Z(n211) );
  NAND U215 ( .A(n212), .B(n213), .Z(n173) );
  NANDN U216 ( .B(n214), .A(n215), .Z(n212) );
  XNOR U217 ( .A(n193), .B(n191), .Z(n142) );
  XNOR U218 ( .A(n216), .B(n196), .Z(n191) );
  XNOR U219 ( .A(n187), .B(n188), .Z(n196) );
  NAND U220 ( .A(n95), .B(n151), .Z(n188) );
  XNOR U221 ( .A(n186), .B(n217), .Z(n187) );
  AND U222 ( .A(n185), .B(n74), .Z(n217) );
  XOR U223 ( .A(n218), .B(n219), .Z(n186) );
  AND U224 ( .A(n220), .B(n221), .Z(n219) );
  XNOR U225 ( .A(n222), .B(n218), .Z(n221) );
  XNOR U226 ( .A(n195), .B(n189), .Z(n216) );
  XOR U227 ( .A(n223), .B(n224), .Z(n189) );
  AND U228 ( .A(n226), .B(n227), .Z(n225) );
  NANDN U229 ( .B(n40), .A(n228), .Z(n227) );
  NANDN U230 ( .B(n229), .A(n230), .Z(n40) );
  AND U231 ( .A(n231), .B(g_input[7]), .Z(n230) );
  NANDN U232 ( .B(n232), .A(n233), .Z(n226) );
  XNOR U233 ( .A(n234), .B(n235), .Z(n194) );
  AND U234 ( .A(n236), .B(n237), .Z(n235) );
  XOR U235 ( .A(n233), .B(n238), .Z(n237) );
  XNOR U236 ( .A(n232), .B(n234), .Z(n238) );
  NAND U237 ( .A(n74), .B(n228), .Z(n232) );
  XNOR U238 ( .A(n242), .B(n239), .Z(n241) );
  XOR U239 ( .A(n220), .B(n243), .Z(n236) );
  XNOR U240 ( .A(n222), .B(n234), .Z(n243) );
  NANDN U241 ( .B(n129), .A(n151), .Z(n222) );
  XOR U242 ( .A(n218), .B(n244), .Z(n220) );
  AND U243 ( .A(n185), .B(n95), .Z(n244) );
  XNOR U244 ( .A(n248), .B(n245), .Z(n247) );
  XOR U245 ( .A(n249), .B(n250), .Z(n234) );
  AND U246 ( .A(n251), .B(n252), .Z(n250) );
  XOR U247 ( .A(n240), .B(n253), .Z(n252) );
  XNOR U248 ( .A(n242), .B(n249), .Z(n253) );
  NAND U249 ( .A(n95), .B(n228), .Z(n242) );
  XOR U250 ( .A(n239), .B(n254), .Z(n240) );
  AND U251 ( .A(n74), .B(e_input[0]), .Z(n254) );
  XNOR U252 ( .A(n231), .B(g_input[6]), .Z(n229) );
  NOR U253 ( .A(n255), .B(n256), .Z(n231) );
  XOR U254 ( .A(n257), .B(n258), .Z(n239) );
  AND U255 ( .A(n259), .B(n260), .Z(n258) );
  XNOR U256 ( .A(n261), .B(n257), .Z(n260) );
  XOR U257 ( .A(n246), .B(n262), .Z(n251) );
  XNOR U258 ( .A(n248), .B(n249), .Z(n262) );
  NANDN U259 ( .B(n170), .A(n151), .Z(n248) );
  XOR U260 ( .A(n245), .B(n263), .Z(n246) );
  ANDN U261 ( .A(n185), .B(n129), .Z(n263) );
  XOR U262 ( .A(n264), .B(n265), .Z(n245) );
  AND U263 ( .A(n266), .B(n267), .Z(n265) );
  XNOR U264 ( .A(n268), .B(n264), .Z(n267) );
  XOR U265 ( .A(n269), .B(n270), .Z(n249) );
  AND U266 ( .A(n271), .B(n272), .Z(n270) );
  XOR U267 ( .A(n259), .B(n273), .Z(n272) );
  XNOR U268 ( .A(n261), .B(n269), .Z(n273) );
  NANDN U269 ( .B(n129), .A(n228), .Z(n261) );
  XOR U270 ( .A(n257), .B(n274), .Z(n259) );
  AND U271 ( .A(n95), .B(e_input[0]), .Z(n274) );
  XNOR U272 ( .A(n275), .B(g_input[5]), .Z(n95) );
  NAND U273 ( .A(n276), .B(g_input[7]), .Z(n275) );
  XOR U274 ( .A(n256), .B(g_input[5]), .Z(n276) );
  XOR U275 ( .A(n255), .B(g_input[5]), .Z(n256) );
  NANDN U276 ( .B(n277), .A(n278), .Z(n255) );
  XOR U277 ( .A(n279), .B(n280), .Z(n257) );
  ANDN U278 ( .A(n281), .B(n282), .Z(n280) );
  XNOR U279 ( .A(n283), .B(n279), .Z(n281) );
  XOR U280 ( .A(n266), .B(n284), .Z(n271) );
  XNOR U281 ( .A(n268), .B(n269), .Z(n284) );
  NAND U282 ( .A(n151), .B(n210), .Z(n268) );
  XOR U283 ( .A(n264), .B(n285), .Z(n266) );
  ANDN U284 ( .A(n185), .B(n170), .Z(n285) );
  XOR U285 ( .A(n286), .B(n287), .Z(n264) );
  ANDN U286 ( .A(n288), .B(n289), .Z(n287) );
  XNOR U287 ( .A(n290), .B(n286), .Z(n288) );
  NAND U288 ( .A(n151), .B(n292), .Z(n290) );
  XNOR U289 ( .A(n286), .B(n293), .Z(n289) );
  AND U290 ( .A(n210), .B(n185), .Z(n293) );
  AND U291 ( .A(n294), .B(g_input[0]), .Z(n286) );
  NANDN U292 ( .B(n151), .A(n295), .Z(n294) );
  NAND U293 ( .A(n292), .B(n185), .Z(n295) );
  XNOR U294 ( .A(n296), .B(e_input[2]), .Z(n185) );
  NAND U295 ( .A(n297), .B(e_input[7]), .Z(n296) );
  XOR U296 ( .A(n298), .B(e_input[2]), .Z(n297) );
  XNOR U297 ( .A(n300), .B(n301), .Z(n224) );
  IV U298 ( .A(n282), .Z(n301) );
  XNOR U299 ( .A(n279), .B(n302), .Z(n282) );
  ANDN U300 ( .A(e_input[0]), .B(n129), .Z(n302) );
  XOR U301 ( .A(n303), .B(n304), .Z(n279) );
  AND U302 ( .A(n305), .B(n306), .Z(n304) );
  XOR U303 ( .A(n307), .B(n303), .Z(n306) );
  ANDN U304 ( .A(e_input[0]), .B(n170), .Z(n307) );
  XOR U305 ( .A(n308), .B(n303), .Z(n305) );
  AND U306 ( .A(n228), .B(n210), .Z(n308) );
  XOR U307 ( .A(n309), .B(n310), .Z(n303) );
  ANDN U308 ( .A(n311), .B(n312), .Z(n310) );
  XNOR U309 ( .A(n313), .B(n309), .Z(n311) );
  XOR U310 ( .A(n314), .B(n283), .Z(n300) );
  NANDN U311 ( .B(n170), .A(n228), .Z(n283) );
  IV U312 ( .A(n291), .Z(n314) );
  NAND U313 ( .A(n228), .B(n292), .Z(n313) );
  XNOR U314 ( .A(n309), .B(n315), .Z(n312) );
  AND U315 ( .A(n210), .B(e_input[0]), .Z(n315) );
  AND U316 ( .A(n316), .B(g_input[0]), .Z(n309) );
  NANDN U317 ( .B(n228), .A(n317), .Z(n316) );
  NAND U318 ( .A(n292), .B(e_input[0]), .Z(n317) );
  XNOR U319 ( .A(n318), .B(e_input[1]), .Z(n228) );
  NAND U320 ( .A(n319), .B(e_input[7]), .Z(n318) );
  XNOR U321 ( .A(e_input[1]), .B(n320), .Z(n319) );
  XNOR U322 ( .A(n199), .B(n322), .Z(n202) );
  ANDN U323 ( .A(n123), .B(n129), .Z(n322) );
  XOR U324 ( .A(n323), .B(g_input[4]), .Z(n129) );
  NAND U325 ( .A(n324), .B(g_input[7]), .Z(n323) );
  XOR U326 ( .A(n277), .B(g_input[4]), .Z(n324) );
  XNOR U327 ( .A(n278), .B(g_input[4]), .Z(n277) );
  NOR U328 ( .A(n325), .B(n326), .Z(n278) );
  XOR U329 ( .A(n327), .B(n328), .Z(n199) );
  AND U330 ( .A(n329), .B(n330), .Z(n328) );
  XOR U331 ( .A(n331), .B(n327), .Z(n330) );
  ANDN U332 ( .A(n123), .B(n170), .Z(n331) );
  XOR U333 ( .A(n332), .B(n327), .Z(n329) );
  AND U334 ( .A(n210), .B(n90), .Z(n332) );
  XOR U335 ( .A(n333), .B(n334), .Z(n327) );
  ANDN U336 ( .A(n335), .B(n336), .Z(n334) );
  XNOR U337 ( .A(n337), .B(n333), .Z(n335) );
  XOR U338 ( .A(n338), .B(n203), .Z(n321) );
  NANDN U339 ( .B(n170), .A(n90), .Z(n203) );
  NANDN U340 ( .B(n339), .A(n340), .Z(n325) );
  IV U341 ( .A(n205), .Z(n338) );
  XOR U342 ( .A(n341), .B(n337), .Z(n205) );
  NAND U343 ( .A(n90), .B(n292), .Z(n337) );
  IV U344 ( .A(n336), .Z(n341) );
  XNOR U345 ( .A(n333), .B(n342), .Z(n336) );
  AND U346 ( .A(n210), .B(n123), .Z(n342) );
  AND U347 ( .A(n343), .B(g_input[0]), .Z(n333) );
  NANDN U348 ( .B(n90), .A(n344), .Z(n343) );
  NAND U349 ( .A(n292), .B(n123), .Z(n344) );
  XNOR U350 ( .A(n345), .B(e_input[4]), .Z(n123) );
  NAND U351 ( .A(n346), .B(e_input[7]), .Z(n345) );
  XOR U352 ( .A(n347), .B(e_input[4]), .Z(n346) );
  XNOR U353 ( .A(n214), .B(n215), .Z(n209) );
  NANDN U354 ( .B(n41), .A(n292), .Z(n215) );
  XNOR U355 ( .A(n213), .B(n349), .Z(n214) );
  AND U356 ( .A(n210), .B(n73), .Z(n349) );
  XNOR U357 ( .A(n340), .B(g_input[2]), .Z(n339) );
  AND U358 ( .A(n351), .B(g_input[0]), .Z(n213) );
  NAND U359 ( .A(n352), .B(n41), .Z(n351) );
  NANDN U360 ( .B(n353), .A(n354), .Z(n41) );
  ANDN U361 ( .A(e_input[7]), .B(n355), .Z(n354) );
  NAND U362 ( .A(n292), .B(n73), .Z(n352) );
  XOR U363 ( .A(n355), .B(e_input[6]), .Z(n353) );
  OR U364 ( .A(n348), .B(n356), .Z(n355) );
  XOR U365 ( .A(n356), .B(e_input[5]), .Z(n348) );
  OR U366 ( .A(n347), .B(n357), .Z(n356) );
  XOR U367 ( .A(n357), .B(e_input[4]), .Z(n347) );
  OR U368 ( .A(n299), .B(n358), .Z(n357) );
  XOR U369 ( .A(n358), .B(e_input[3]), .Z(n299) );
  OR U370 ( .A(n298), .B(n359), .Z(n358) );
  XOR U371 ( .A(n359), .B(e_input[2]), .Z(n298) );
  NANDN U372 ( .B(e_input[0]), .A(n320), .Z(n359) );
  XNOR U373 ( .A(e_input[0]), .B(e_input[1]), .Z(n320) );
  XOR U374 ( .A(g_input[0]), .B(g_input[1]), .Z(n350) );
  AND U375 ( .A(n360), .B(n361), .Z(\_MxM/N23 ) );
  XOR U376 ( .A(\_MxM/n[9] ), .B(\_MxM/add_43/carry[9] ), .Z(n361) );
  AND U377 ( .A(\_MxM/N12 ), .B(n360), .Z(\_MxM/N22 ) );
  AND U378 ( .A(\_MxM/N11 ), .B(n360), .Z(\_MxM/N21 ) );
  AND U379 ( .A(\_MxM/N10 ), .B(n360), .Z(\_MxM/N20 ) );
  AND U380 ( .A(\_MxM/N9 ), .B(n360), .Z(\_MxM/N19 ) );
  AND U381 ( .A(\_MxM/N8 ), .B(n360), .Z(\_MxM/N18 ) );
  AND U382 ( .A(\_MxM/N7 ), .B(n360), .Z(\_MxM/N17 ) );
  AND U383 ( .A(\_MxM/N6 ), .B(n360), .Z(\_MxM/N16 ) );
  AND U384 ( .A(\_MxM/N5 ), .B(n360), .Z(\_MxM/N15 ) );
  NAND U385 ( .A(n362), .B(n363), .Z(n360) );
  AND U386 ( .A(n364), .B(n365), .Z(n363) );
  AND U387 ( .A(\_MxM/n[1] ), .B(n366), .Z(n365) );
  NOR U388 ( .A(\_MxM/N14 ), .B(n21), .Z(n366) );
  OR U389 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n21) );
  AND U390 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n364) );
  AND U391 ( .A(n367), .B(n368), .Z(n362) );
  AND U392 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n368) );
  AND U393 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n367) );
  IV U394 ( .A(\_MxM/n[0] ), .Z(\_MxM/N14 ) );
endmodule

