
module MAC_TG_N16 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236;
  wire   [15:0] o_reg;

  DFF \o_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[0])
         );
  DFF \o_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[1])
         );
  DFF \o_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[2])
         );
  DFF \o_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[3])
         );
  DFF \o_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[4])
         );
  DFF \o_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[5])
         );
  DFF \o_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[6])
         );
  DFF \o_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[7])
         );
  DFF \o_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[8])
         );
  DFF \o_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[9])
         );
  DFF \o_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[10]) );
  DFF \o_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[11]) );
  DFF \o_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[12]) );
  DFF \o_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[13]) );
  DFF \o_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[14]) );
  DFF \o_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[15]) );
  MUX U19 ( .IN0(n1026), .IN1(n17), .SEL(n1027), .F(n1013) );
  IV U20 ( .A(n1028), .Z(n17) );
  MUX U21 ( .IN0(n883), .IN1(n885), .SEL(n884), .F(n861) );
  XNOR U22 ( .A(n997), .B(n988), .Z(n846) );
  MUX U23 ( .IN0(n981), .IN1(n992), .SEL(n982), .F(n969) );
  MUX U24 ( .IN0(n785), .IN1(n18), .SEL(n786), .F(n763) );
  IV U25 ( .A(n787), .Z(n18) );
  XNOR U26 ( .A(n759), .B(n760), .Z(n769) );
  XNOR U27 ( .A(n945), .B(n936), .Z(n754) );
  XNOR U28 ( .A(n738), .B(n739), .Z(n734) );
  MUX U29 ( .IN0(n276), .IN1(n19), .SEL(n277), .F(n239) );
  IV U30 ( .A(n278), .Z(n19) );
  MUX U31 ( .IN0(n324), .IN1(n360), .SEL(n325), .F(n284) );
  MUX U32 ( .IN0(n387), .IN1(n437), .SEL(n388), .F(n335) );
  MUX U33 ( .IN0(n398), .IN1(n20), .SEL(n399), .F(n344) );
  IV U34 ( .A(n400), .Z(n20) );
  MUX U35 ( .IN0(n656), .IN1(n21), .SEL(n657), .F(n590) );
  IV U36 ( .A(n658), .Z(n21) );
  MUX U37 ( .IN0(n307), .IN1(n22), .SEL(n308), .F(n269) );
  IV U38 ( .A(n309), .Z(n22) );
  MUX U39 ( .IN0(n357), .IN1(n23), .SEL(n358), .F(n318) );
  IV U40 ( .A(n359), .Z(n23) );
  MUX U41 ( .IN0(n506), .IN1(n24), .SEL(n507), .F(n451) );
  IV U42 ( .A(n508), .Z(n24) );
  MUX U43 ( .IN0(n579), .IN1(n25), .SEL(n580), .F(n517) );
  IV U44 ( .A(n581), .Z(n25) );
  MUX U45 ( .IN0(n474), .IN1(n26), .SEL(n475), .F(n422) );
  IV U46 ( .A(n476), .Z(n26) );
  MUX U47 ( .IN0(n442), .IN1(n27), .SEL(n443), .F(n391) );
  IV U48 ( .A(n444), .Z(n27) );
  MUX U49 ( .IN0(n1116), .IN1(n28), .SEL(n724), .F(n627) );
  IV U50 ( .A(n723), .Z(n28) );
  MUX U51 ( .IN0(n29), .IN1(n162), .SEL(n163), .F(n144) );
  IV U52 ( .A(n164), .Z(n29) );
  MUX U53 ( .IN0(n604), .IN1(n30), .SEL(n605), .F(n543) );
  IV U54 ( .A(n606), .Z(n30) );
  MUX U55 ( .IN0(n221), .IN1(o_reg[10]), .SEL(n94), .F(n182) );
  MUX U56 ( .IN0(n383), .IN1(o_reg[6]), .SEL(n98), .F(n331) );
  MUX U57 ( .IN0(n1007), .IN1(n1018), .SEL(n1008), .F(n993) );
  MUX U58 ( .IN0(n849), .IN1(n872), .SEL(n850), .F(n827) );
  MUX U59 ( .IN0(n1013), .IN1(n31), .SEL(n1014), .F(n999) );
  IV U60 ( .A(n1015), .Z(n31) );
  MUX U61 ( .IN0(n32), .IN1(n911), .SEL(n741), .F(n886) );
  IV U62 ( .A(n740), .Z(n32) );
  XNOR U63 ( .A(n877), .B(n858), .Z(n862) );
  MUX U64 ( .IN0(n1088), .IN1(n1093), .SEL(n1089), .F(n1073) );
  MUX U65 ( .IN0(n1083), .IN1(n33), .SEL(n1084), .F(n1067) );
  IV U66 ( .A(n1085), .Z(n33) );
  MUX U67 ( .IN0(n1181), .IN1(n34), .SEL(n1182), .F(n1165) );
  IV U68 ( .A(n1183), .Z(n34) );
  MUX U69 ( .IN0(n991), .IN1(n844), .SEL(n846), .F(n979) );
  XNOR U70 ( .A(n807), .B(n786), .Z(n791) );
  XNOR U71 ( .A(n943), .B(n944), .Z(n774) );
  MUX U72 ( .IN0(n361), .IN1(n416), .SEL(n362), .F(n324) );
  MUX U73 ( .IN0(n353), .IN1(n35), .SEL(n354), .F(n312) );
  IV U74 ( .A(n355), .Z(n35) );
  MUX U75 ( .IN0(n344), .IN1(n36), .SEL(n345), .F(n303) );
  IV U76 ( .A(n346), .Z(n36) );
  MUX U77 ( .IN0(n575), .IN1(n37), .SEL(n576), .F(n511) );
  IV U78 ( .A(n577), .Z(n37) );
  MUX U79 ( .IN0(n600), .IN1(n665), .SEL(n601), .F(n539) );
  MUX U80 ( .IN0(n590), .IN1(n38), .SEL(n591), .F(n529) );
  IV U81 ( .A(n592), .Z(n38) );
  MUX U82 ( .IN0(n935), .IN1(n39), .SEL(n936), .F(n716) );
  IV U83 ( .A(n937), .Z(n39) );
  MUX U84 ( .IN0(n166), .IN1(n40), .SEL(n167), .F(n146) );
  IV U85 ( .A(n168), .Z(n40) );
  MUX U86 ( .IN0(n243), .IN1(n41), .SEL(n244), .F(n209) );
  IV U87 ( .A(n245), .Z(n41) );
  MUX U88 ( .IN0(n402), .IN1(n42), .SEL(n403), .F(n348) );
  IV U89 ( .A(n404), .Z(n42) );
  MUX U90 ( .IN0(n462), .IN1(n43), .SEL(n463), .F(n411) );
  IV U91 ( .A(n464), .Z(n43) );
  MUX U92 ( .IN0(n636), .IN1(n44), .SEL(n637), .F(n570) );
  IV U93 ( .A(n638), .Z(n44) );
  MUX U94 ( .IN0(n1214), .IN1(n45), .SEL(n1121), .F(n645) );
  IV U95 ( .A(n1120), .Z(n45) );
  XNOR U96 ( .A(n726), .B(n692), .Z(n696) );
  MUX U97 ( .IN0(n233), .IN1(n266), .SEL(n235), .F(n190) );
  MUX U98 ( .IN0(n299), .IN1(n46), .SEL(n300), .F(n261) );
  IV U99 ( .A(n301), .Z(n46) );
  MUX U100 ( .IN0(n497), .IN1(n47), .SEL(n498), .F(n442) );
  IV U101 ( .A(n499), .Z(n47) );
  MUX U102 ( .IN0(n48), .IN1(n616), .SEL(n617), .F(n548) );
  IV U103 ( .A(n618), .Z(n48) );
  MUX U104 ( .IN0(n422), .IN1(n49), .SEL(n423), .F(n368) );
  IV U105 ( .A(n424), .Z(n49) );
  MUX U106 ( .IN0(n431), .IN1(n50), .SEL(n432), .F(n378) );
  IV U107 ( .A(n433), .Z(n50) );
  MUX U108 ( .IN0(n670), .IN1(n51), .SEL(n671), .F(n604) );
  IV U109 ( .A(n672), .Z(n51) );
  MUX U110 ( .IN0(n159), .IN1(o_reg[12]), .SEL(n160), .F(n140) );
  MUX U111 ( .IN0(n291), .IN1(o_reg[8]), .SEL(n96), .F(n253) );
  MUX U112 ( .IN0(n489), .IN1(o_reg[4]), .SEL(n100), .F(n434) );
  MUX U113 ( .IN0(n895), .IN1(n929), .SEL(n896), .F(n873) );
  MUX U114 ( .IN0(n879), .IN1(n52), .SEL(n880), .F(n855) );
  IV U115 ( .A(n881), .Z(n52) );
  MUX U116 ( .IN0(n1017), .IN1(n890), .SEL(n892), .F(n1003) );
  MUX U117 ( .IN0(n993), .IN1(n1006), .SEL(n994), .F(n981) );
  MUX U118 ( .IN0(n999), .IN1(n53), .SEL(n1000), .F(n987) );
  IV U119 ( .A(n1001), .Z(n53) );
  MUX U120 ( .IN0(n837), .IN1(n839), .SEL(n838), .F(n813) );
  MUX U121 ( .IN0(n1092), .IN1(n932), .SEL(n933), .F(n1077) );
  MUX U122 ( .IN0(n1067), .IN1(n1082), .SEL(n1069), .F(n1051) );
  MUX U123 ( .IN0(n1200), .IN1(n1205), .SEL(n1201), .F(n1196) );
  XNOR U124 ( .A(n973), .B(n962), .Z(n800) );
  XNOR U125 ( .A(n781), .B(n782), .Z(n793) );
  MUX U126 ( .IN0(n763), .IN1(n54), .SEL(n764), .F(n728) );
  IV U127 ( .A(n765), .Z(n54) );
  MUX U128 ( .IN0(n941), .IN1(n954), .SEL(n942), .F(n744) );
  MUX U129 ( .IN0(n1132), .IN1(n1154), .SEL(n1134), .F(n1112) );
  MUX U130 ( .IN0(n466), .IN1(n522), .SEL(n467), .F(n417) );
  MUX U131 ( .IN0(n447), .IN1(n55), .SEL(n448), .F(n398) );
  IV U132 ( .A(n449), .Z(n55) );
  MUX U133 ( .IN0(n641), .IN1(n56), .SEL(n642), .F(n575) );
  IV U134 ( .A(n643), .Z(n56) );
  MUX U135 ( .IN0(n1126), .IN1(n57), .SEL(n1127), .F(n632) );
  IV U136 ( .A(n1128), .Z(n57) );
  MUX U137 ( .IN0(n280), .IN1(n58), .SEL(n281), .F(n243) );
  IV U138 ( .A(n282), .Z(n58) );
  MUX U139 ( .IN0(n539), .IN1(n599), .SEL(n540), .F(n478) );
  MUX U140 ( .IN0(n348), .IN1(n59), .SEL(n349), .F(n307) );
  IV U141 ( .A(n350), .Z(n59) );
  MUX U142 ( .IN0(n570), .IN1(n60), .SEL(n571), .F(n506) );
  IV U143 ( .A(n572), .Z(n60) );
  XNOR U144 ( .A(n934), .B(n716), .Z(n719) );
  MUX U145 ( .IN0(n695), .IN1(n61), .SEL(n696), .F(n660) );
  IV U146 ( .A(n697), .Z(n61) );
  MUX U147 ( .IN0(n148), .IN1(n62), .SEL(n149), .F(n131) );
  IV U148 ( .A(n150), .Z(n62) );
  XNOR U149 ( .A(n456), .B(n408), .Z(n414) );
  XNOR U150 ( .A(n528), .B(n472), .Z(n475) );
  MUX U151 ( .IN0(n627), .IN1(n63), .SEL(n628), .F(n559) );
  IV U152 ( .A(n629), .Z(n63) );
  XNOR U153 ( .A(n162), .B(n194), .Z(n187) );
  MUX U154 ( .IN0(n64), .IN1(n548), .SEL(n549), .F(n483) );
  IV U155 ( .A(n550), .Z(n64) );
  XOR U156 ( .A(n723), .B(n724), .Z(n705) );
  MUX U157 ( .IN0(n140), .IN1(o_reg[13]), .SEL(n141), .F(n126) );
  MUX U158 ( .IN0(n253), .IN1(o_reg[9]), .SEL(n95), .F(n221) );
  MUX U159 ( .IN0(n65), .IN1(n328), .SEL(n329), .F(n290) );
  IV U160 ( .A(n330), .Z(n65) );
  MUX U161 ( .IN0(o_reg[3]), .IN1(n551), .SEL(n101), .F(n489) );
  XNOR U162 ( .A(n1011), .B(n1000), .Z(n870) );
  MUX U163 ( .IN0(n827), .IN1(n848), .SEL(n828), .F(n803) );
  MUX U164 ( .IN0(n861), .IN1(n863), .SEL(n862), .F(n837) );
  MUX U165 ( .IN0(n833), .IN1(n66), .SEL(n834), .F(n809) );
  IV U166 ( .A(n835), .Z(n66) );
  XNOR U167 ( .A(n983), .B(n984), .Z(n844) );
  MUX U168 ( .IN0(n1073), .IN1(n1087), .SEL(n1075), .F(n1057) );
  MUX U169 ( .IN0(n1102), .IN1(n1107), .SEL(n1103), .F(n1098) );
  MUX U170 ( .IN0(n1190), .IN1(n1122), .SEL(n1123), .F(n1175) );
  MUX U171 ( .IN0(n1171), .IN1(n1185), .SEL(n1173), .F(n1155) );
  MUX U172 ( .IN0(n975), .IN1(n67), .SEL(n976), .F(n961) );
  IV U173 ( .A(n977), .Z(n67) );
  XNOR U174 ( .A(n971), .B(n972), .Z(n822) );
  MUX U175 ( .IN0(n921), .IN1(n926), .SEL(n922), .F(n917) );
  MUX U176 ( .IN0(n1221), .IN1(n1229), .SEL(n1222), .F(n1217) );
  MUX U177 ( .IN0(n736), .IN1(n756), .SEL(n737), .F(n699) );
  MUX U178 ( .IN0(n728), .IN1(n68), .SEL(n729), .F(n691) );
  IV U179 ( .A(n730), .Z(n68) );
  MUX U180 ( .IN0(n767), .IN1(n769), .SEL(n768), .F(n732) );
  MUX U181 ( .IN0(n239), .IN1(n69), .SEL(n240), .F(n203) );
  IV U182 ( .A(n241), .Z(n69) );
  MUX U183 ( .IN0(n295), .IN1(n334), .SEL(n296), .F(n257) );
  MUX U184 ( .IN0(n417), .IN1(n465), .SEL(n418), .F(n361) );
  MUX U185 ( .IN0(n493), .IN1(n554), .SEL(n494), .F(n438) );
  MUX U186 ( .IN0(n649), .IN1(n1232), .SEL(n650), .F(n583) );
  MUX U187 ( .IN0(n632), .IN1(n70), .SEL(n633), .F(n564) );
  IV U188 ( .A(n634), .Z(n70) );
  MUX U189 ( .IN0(n939), .IN1(n752), .SEL(n754), .F(n718) );
  MUX U190 ( .IN0(n303), .IN1(n71), .SEL(n304), .F(n267) );
  IV U191 ( .A(n305), .Z(n71) );
  MUX U192 ( .IN0(n708), .IN1(n743), .SEL(n709), .F(n674) );
  MUX U193 ( .IN0(n1130), .IN1(n72), .SEL(n1119), .F(n636) );
  IV U194 ( .A(n1118), .Z(n72) );
  MUX U195 ( .IN0(n478), .IN1(n538), .SEL(n479), .F(n425) );
  XNOR U196 ( .A(n351), .B(n315), .Z(n321) );
  MUX U197 ( .IN0(n339), .IN1(n73), .SEL(n340), .F(n299) );
  IV U198 ( .A(n341), .Z(n73) );
  XNOR U199 ( .A(n500), .B(n448), .Z(n453) );
  XNOR U200 ( .A(n509), .B(n459), .Z(n463) );
  MUX U201 ( .IN0(n559), .IN1(n74), .SEL(n560), .F(n497) );
  IV U202 ( .A(n561), .Z(n74) );
  XNOR U203 ( .A(n588), .B(n530), .Z(n536) );
  MUX U204 ( .IN0(n678), .IN1(n75), .SEL(n679), .F(n616) );
  IV U205 ( .A(n680), .Z(n75) );
  XNOR U206 ( .A(n1208), .B(n642), .Z(n646) );
  MUX U207 ( .IN0(n152), .IN1(n175), .SEL(n153), .F(n134) );
  MUX U208 ( .IN0(n703), .IN1(n76), .SEL(n704), .F(n670) );
  IV U209 ( .A(n705), .Z(n76) );
  XOR U210 ( .A(n143), .B(n144), .Z(n158) );
  XOR U211 ( .A(n200), .B(n199), .Z(n220) );
  XOR U212 ( .A(n232), .B(n231), .Z(n252) );
  MUX U213 ( .IN0(o_reg[7]), .IN1(n331), .SEL(n97), .F(n291) );
  XOR U214 ( .A(n378), .B(n371), .Z(n421) );
  MUX U215 ( .IN0(n81), .IN1(o_reg[2]), .SEL(n102), .F(n551) );
  MUX U216 ( .IN0(o_reg[14]), .IN1(n126), .SEL(n127), .F(n103) );
  MUX U217 ( .IN0(n902), .IN1(n77), .SEL(n903), .F(n879) );
  IV U218 ( .A(n904), .Z(n77) );
  MUX U219 ( .IN0(n873), .IN1(n894), .SEL(n874), .F(n849) );
  XNOR U220 ( .A(n1024), .B(n1014), .Z(n892) );
  XNOR U221 ( .A(n995), .B(n996), .Z(n868) );
  MUX U222 ( .IN0(n987), .IN1(n78), .SEL(n988), .F(n975) );
  IV U223 ( .A(n989), .Z(n78) );
  XNOR U224 ( .A(n853), .B(n834), .Z(n838) );
  MUX U225 ( .IN0(n969), .IN1(n980), .SEL(n970), .F(n955) );
  MUX U226 ( .IN0(n1165), .IN1(n1180), .SEL(n1167), .F(n1149) );
  MUX U227 ( .IN0(n779), .IN1(n802), .SEL(n780), .F(n757) );
  MUX U228 ( .IN0(n1057), .IN1(n1072), .SEL(n1059), .F(n1034) );
  MUX U229 ( .IN0(n1051), .IN1(n1066), .SEL(n1053), .F(n1040) );
  MUX U230 ( .IN0(n1155), .IN1(n1170), .SEL(n1157), .F(n1132) );
  XNOR U231 ( .A(n959), .B(n948), .Z(n776) );
  XNOR U232 ( .A(n1104), .B(n1105), .Z(n1092) );
  XNOR U233 ( .A(n1202), .B(n1203), .Z(n1190) );
  XNOR U234 ( .A(n783), .B(n764), .Z(n768) );
  XNOR U235 ( .A(n923), .B(n924), .Z(n906) );
  MUX U236 ( .IN0(n335), .IN1(n386), .SEL(n336), .F(n295) );
  MUX U237 ( .IN0(n523), .IN1(n582), .SEL(n524), .F(n466) );
  MUX U238 ( .IN0(n555), .IN1(n622), .SEL(n556), .F(n493) );
  MUX U239 ( .IN0(n666), .IN1(n698), .SEL(n667), .F(n600) );
  XNOR U240 ( .A(n746), .B(n747), .Z(n752) );
  MUX U241 ( .IN0(n215), .IN1(n246), .SEL(n216), .F(n176) );
  MUX U242 ( .IN0(n529), .IN1(n79), .SEL(n530), .F(n472) );
  IV U243 ( .A(n531), .Z(n79) );
  XNOR U244 ( .A(n1215), .B(n1211), .Z(n1121) );
  XNOR U245 ( .A(n1136), .B(n1127), .Z(n1119) );
  XNOR U246 ( .A(n237), .B(n206), .Z(n212) );
  XNOR U247 ( .A(n396), .B(n345), .Z(n349) );
  XNOR U248 ( .A(n405), .B(n354), .Z(n358) );
  XNOR U249 ( .A(n573), .B(n514), .Z(n520) );
  XNOR U250 ( .A(n562), .B(n503), .Z(n507) );
  XNOR U251 ( .A(n689), .B(n657), .Z(n663) );
  MUX U252 ( .IN0(n131), .IN1(n80), .SEL(n132), .F(n120) );
  IV U253 ( .A(n133), .Z(n80) );
  XOR U254 ( .A(n150), .B(n149), .Z(n143) );
  XOR U255 ( .A(n245), .B(n244), .Z(n232) );
  XNOR U256 ( .A(n548), .B(n614), .Z(n607) );
  XOR U257 ( .A(n581), .B(n580), .Z(n561) );
  XOR U258 ( .A(n647), .B(n646), .Z(n629) );
  XOR U259 ( .A(n265), .B(n264), .Z(n289) );
  XNOR U260 ( .A(n328), .B(n376), .Z(n365) );
  MUX U261 ( .IN0(n434), .IN1(o_reg[5]), .SEL(n99), .F(n383) );
  MUX U262 ( .IN0(n685), .IN1(o_reg[1]), .SEL(n686), .F(n81) );
  IV U263 ( .A(n81), .Z(n619) );
  XNOR U264 ( .A(n126), .B(n112), .Z(n128) );
  XOR U265 ( .A(n182), .B(n181), .Z(n186) );
  XNOR U266 ( .A(n1009), .B(n1010), .Z(n890) );
  XNOR U267 ( .A(n851), .B(n852), .Z(n863) );
  XNOR U268 ( .A(n829), .B(n830), .Z(n839) );
  XNOR U269 ( .A(n805), .B(n806), .Z(n817) );
  MUX U270 ( .IN0(n809), .IN1(n82), .SEL(n810), .F(n785) );
  IV U271 ( .A(n811), .Z(n82) );
  MUX U272 ( .IN0(n979), .IN1(n822), .SEL(n824), .F(n965) );
  MUX U273 ( .IN0(n1098), .IN1(n1101), .SEL(n1099), .F(n1083) );
  MUX U274 ( .IN0(n955), .IN1(n968), .SEL(n956), .F(n941) );
  MUX U275 ( .IN0(n1196), .IN1(n1199), .SEL(n1197), .F(n1181) );
  MUX U276 ( .IN0(n757), .IN1(n778), .SEL(n758), .F(n736) );
  MUX U277 ( .IN0(n961), .IN1(n83), .SEL(n962), .F(n947) );
  IV U278 ( .A(n963), .Z(n83) );
  MUX U279 ( .IN0(n1040), .IN1(n1050), .SEL(n1042), .F(n1026) );
  MUX U280 ( .IN0(n1217), .IN1(n1220), .SEL(n1218), .F(n1210) );
  MUX U281 ( .IN0(n1138), .IN1(n1148), .SEL(n1140), .F(n1126) );
  XNOR U282 ( .A(n1090), .B(n1091), .Z(n932) );
  MUX U283 ( .IN0(n247), .IN1(n283), .SEL(n248), .F(n215) );
  MUX U284 ( .IN0(n407), .IN1(n84), .SEL(n408), .F(n353) );
  IV U285 ( .A(n409), .Z(n84) );
  MUX U286 ( .IN0(n623), .IN1(n1111), .SEL(n624), .F(n555) );
  MUX U287 ( .IN0(n85), .IN1(n1233), .SEL(n1226), .F(n649) );
  IV U288 ( .A(n1227), .Z(n85) );
  XNOR U289 ( .A(n1188), .B(n1189), .Z(n1122) );
  XNOR U290 ( .A(n761), .B(n729), .Z(n733) );
  XNOR U291 ( .A(n915), .B(n903), .Z(n909) );
  XNOR U292 ( .A(n1022), .B(n1023), .Z(n913) );
  MUX U293 ( .IN0(n257), .IN1(n294), .SEL(n258), .F(n224) );
  MUX U294 ( .IN0(n718), .IN1(n86), .SEL(n719), .F(n681) );
  IV U295 ( .A(n720), .Z(n86) );
  XNOR U296 ( .A(n165), .B(n146), .Z(n149) );
  XNOR U297 ( .A(n274), .B(n240), .Z(n244) );
  XNOR U298 ( .A(n302), .B(n267), .Z(n271) );
  XNOR U299 ( .A(n445), .B(n399), .Z(n403) );
  MUX U300 ( .IN0(n674), .IN1(n707), .SEL(n675), .F(n614) );
  XNOR U301 ( .A(n639), .B(n576), .Z(n580) );
  XNOR U302 ( .A(n630), .B(n567), .Z(n571) );
  XNOR U303 ( .A(n654), .B(n591), .Z(n597) );
  XOR U304 ( .A(n697), .B(n696), .Z(n714) );
  XOR U305 ( .A(n174), .B(n173), .Z(n164) );
  XOR U306 ( .A(n282), .B(n281), .Z(n265) );
  MUX U307 ( .IN0(n425), .IN1(n477), .SEL(n426), .F(n376) );
  XOR U308 ( .A(n359), .B(n358), .Z(n341) );
  XOR U309 ( .A(n415), .B(n414), .Z(n395) );
  XOR U310 ( .A(n464), .B(n463), .Z(n444) );
  XOR U311 ( .A(n521), .B(n520), .Z(n499) );
  XOR U312 ( .A(n664), .B(n663), .Z(n680) );
  MUX U313 ( .IN0(n134), .IN1(n151), .SEL(n135), .F(n118) );
  XOR U314 ( .A(n301), .B(n300), .Z(n330) );
  XOR U315 ( .A(n431), .B(n429), .Z(n470) );
  XOR U316 ( .A(n629), .B(n628), .Z(n672) );
  XNOR U317 ( .A(n142), .B(n138), .Z(n141) );
  XOR U318 ( .A(n221), .B(n219), .Z(n222) );
  XNOR U319 ( .A(n875), .B(n876), .Z(n885) );
  MUX U320 ( .IN0(n1186), .IN1(n1191), .SEL(n1187), .F(n1171) );
  MUX U321 ( .IN0(n803), .IN1(n826), .SEL(n804), .F(n779) );
  XNOR U322 ( .A(n985), .B(n976), .Z(n824) );
  XNOR U323 ( .A(n831), .B(n810), .Z(n815) );
  MUX U324 ( .IN0(n1149), .IN1(n1164), .SEL(n1151), .F(n1138) );
  XNOR U325 ( .A(n957), .B(n958), .Z(n798) );
  MUX U326 ( .IN0(n917), .IN1(n920), .SEL(n918), .F(n902) );
  MUX U327 ( .IN0(n1034), .IN1(n1056), .SEL(n1036), .F(n1019) );
  XNOR U328 ( .A(n1096), .B(n1084), .Z(n933) );
  MUX U329 ( .IN0(n458), .IN1(n87), .SEL(n459), .F(n407) );
  IV U330 ( .A(n460), .Z(n87) );
  MUX U331 ( .IN0(n438), .IN1(n492), .SEL(n439), .F(n387) );
  MUX U332 ( .IN0(n502), .IN1(n88), .SEL(n503), .F(n447) );
  IV U333 ( .A(n504), .Z(n88) );
  MUX U334 ( .IN0(n583), .IN1(n648), .SEL(n584), .F(n523) );
  MUX U335 ( .IN0(n744), .IN1(n940), .SEL(n745), .F(n708) );
  MUX U336 ( .IN0(n1210), .IN1(n89), .SEL(n1211), .F(n641) );
  IV U337 ( .A(n1212), .Z(n89) );
  MUX U338 ( .IN0(n1112), .IN1(n1131), .SEL(n1113), .F(n623) );
  XNOR U339 ( .A(n1194), .B(n1182), .Z(n1123) );
  MUX U340 ( .IN0(n699), .IN1(n735), .SEL(n700), .F(n666) );
  MUX U341 ( .IN0(n732), .IN1(n734), .SEL(n733), .F(n695) );
  MUX U342 ( .IN0(n691), .IN1(n90), .SEL(n692), .F(n656) );
  IV U343 ( .A(n693), .Z(n90) );
  MUX U344 ( .IN0(n947), .IN1(n91), .SEL(n948), .F(n935) );
  IV U345 ( .A(n949), .Z(n91) );
  XNOR U346 ( .A(n1038), .B(n1027), .Z(n914) );
  MUX U347 ( .IN0(n645), .IN1(n92), .SEL(n646), .F(n579) );
  IV U348 ( .A(n647), .Z(n92) );
  XOR U349 ( .A(n910), .B(n909), .Z(n740) );
  MUX U350 ( .IN0(n176), .IN1(n214), .SEL(n177), .F(n152) );
  MUX U351 ( .IN0(n224), .IN1(n256), .SEL(n225), .F(n194) );
  XNOR U352 ( .A(n201), .B(n167), .Z(n173) );
  XNOR U353 ( .A(n310), .B(n277), .Z(n281) );
  XNOR U354 ( .A(n342), .B(n304), .Z(n308) );
  MUX U355 ( .IN0(n681), .IN1(n715), .SEL(n683), .F(n610) );
  XNOR U356 ( .A(n1124), .B(n633), .Z(n637) );
  XOR U357 ( .A(n1120), .B(n1121), .Z(n723) );
  MUX U358 ( .IN0(n712), .IN1(n93), .SEL(n713), .F(n678) );
  IV U359 ( .A(n714), .Z(n93) );
  XOR U360 ( .A(n133), .B(n132), .Z(n130) );
  XOR U361 ( .A(n213), .B(n212), .Z(n200) );
  XOR U362 ( .A(n322), .B(n321), .Z(n301) );
  XOR U363 ( .A(n424), .B(n423), .Z(n430) );
  XOR U364 ( .A(n476), .B(n475), .Z(n482) );
  XOR U365 ( .A(n537), .B(n536), .Z(n550) );
  XOR U366 ( .A(n598), .B(n597), .Z(n618) );
  XOR U367 ( .A(n341), .B(n340), .Z(n382) );
  XOR U368 ( .A(n395), .B(n394), .Z(n433) );
  XOR U369 ( .A(n444), .B(n443), .Z(n488) );
  XOR U370 ( .A(n499), .B(n498), .Z(n547) );
  XOR U371 ( .A(n561), .B(n560), .Z(n606) );
  XOR U372 ( .A(n159), .B(n157), .Z(n161) );
  XOR U373 ( .A(n253), .B(n251), .Z(n254) );
  XNOR U374 ( .A(n687), .B(n671), .Z(n686) );
  MUX U375 ( .IN0(o_reg[15]), .IN1(n103), .SEL(n104), .F(o[15]) );
  XOR U376 ( .A(o_reg[10]), .B(n94), .Z(o[9]) );
  XOR U377 ( .A(o_reg[9]), .B(n95), .Z(o[8]) );
  XOR U378 ( .A(o_reg[8]), .B(n96), .Z(o[7]) );
  XNOR U379 ( .A(n97), .B(o_reg[7]), .Z(o[6]) );
  XOR U380 ( .A(o_reg[6]), .B(n98), .Z(o[5]) );
  XOR U381 ( .A(o_reg[5]), .B(n99), .Z(o[4]) );
  XOR U382 ( .A(o_reg[4]), .B(n100), .Z(o[3]) );
  XNOR U383 ( .A(n101), .B(o_reg[3]), .Z(o[2]) );
  XOR U384 ( .A(o_reg[2]), .B(n102), .Z(o[1]) );
  XNOR U385 ( .A(o_reg[15]), .B(n104), .Z(o[14]) );
  XOR U386 ( .A(n105), .B(n106), .Z(n104) );
  XNOR U387 ( .A(n107), .B(n108), .Z(n106) );
  XOR U388 ( .A(n109), .B(n110), .Z(n108) );
  ANDN U389 ( .A(n111), .B(n112), .Z(n110) );
  AND U390 ( .A(n113), .B(n114), .Z(n109) );
  AND U391 ( .A(n115), .B(n116), .Z(n114) );
  NAND U392 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U393 ( .B(n119), .A(n120), .Z(n115) );
  AND U394 ( .A(n121), .B(n122), .Z(n113) );
  NAND U395 ( .A(n123), .B(n124), .Z(n122) );
  NAND U396 ( .A(n125), .B(n112), .Z(n121) );
  XNOR U397 ( .A(n103), .B(n118), .Z(n105) );
  XNOR U398 ( .A(o_reg[14]), .B(n127), .Z(o[13]) );
  XNOR U399 ( .A(n128), .B(n125), .Z(n127) );
  XOR U400 ( .A(n124), .B(n123), .Z(n125) );
  IV U401 ( .A(n111), .Z(n123) );
  OR U402 ( .A(n129), .B(n130), .Z(n111) );
  XOR U403 ( .A(n119), .B(n107), .Z(n124) );
  IV U404 ( .A(n120), .Z(n107) );
  XNOR U405 ( .A(n118), .B(n117), .Z(n119) );
  NAND U406 ( .A(g_input[15]), .B(e_input[15]), .Z(n117) );
  XNOR U407 ( .A(n137), .B(n134), .Z(n135) );
  ANDN U408 ( .A(n138), .B(n139), .Z(n112) );
  XOR U409 ( .A(o_reg[13]), .B(n141), .Z(o[12]) );
  XOR U410 ( .A(n130), .B(n129), .Z(n138) );
  NANDN U411 ( .B(n143), .A(n144), .Z(n129) );
  XOR U412 ( .A(n131), .B(n145), .Z(n132) );
  ANDN U413 ( .A(n146), .B(n147), .Z(n145) );
  XNOR U414 ( .A(n136), .B(n137), .Z(n133) );
  NAND U415 ( .A(e_input[15]), .B(g_input[14]), .Z(n137) );
  XNOR U416 ( .A(n134), .B(n151), .Z(n136) );
  AND U417 ( .A(g_input[15]), .B(e_input[14]), .Z(n151) );
  XNOR U418 ( .A(n155), .B(n152), .Z(n153) );
  XNOR U419 ( .A(n156), .B(n139), .Z(n142) );
  OR U420 ( .A(n157), .B(n158), .Z(n139) );
  IV U421 ( .A(n140), .Z(n156) );
  XOR U422 ( .A(o_reg[12]), .B(n160), .Z(o[11]) );
  XOR U423 ( .A(n161), .B(n158), .Z(n160) );
  XNOR U424 ( .A(n169), .B(n147), .Z(n165) );
  NAND U425 ( .A(e_input[13]), .B(g_input[15]), .Z(n147) );
  IV U426 ( .A(n148), .Z(n169) );
  XOR U427 ( .A(n170), .B(n171), .Z(n148) );
  AND U428 ( .A(n172), .B(n173), .Z(n171) );
  XNOR U429 ( .A(n170), .B(n174), .Z(n172) );
  XNOR U430 ( .A(n154), .B(n155), .Z(n150) );
  NAND U431 ( .A(e_input[15]), .B(g_input[13]), .Z(n155) );
  XNOR U432 ( .A(n152), .B(n175), .Z(n154) );
  AND U433 ( .A(g_input[14]), .B(e_input[14]), .Z(n175) );
  XNOR U434 ( .A(n179), .B(n176), .Z(n177) );
  OR U435 ( .A(n180), .B(n181), .Z(n157) );
  XOR U436 ( .A(n182), .B(n183), .Z(n159) );
  ANDN U437 ( .A(n184), .B(n185), .Z(n183) );
  XOR U438 ( .A(o_reg[11]), .B(n182), .Z(n184) );
  XNOR U439 ( .A(n185), .B(o_reg[11]), .Z(o[10]) );
  XNOR U440 ( .A(n186), .B(n180), .Z(n185) );
  XNOR U441 ( .A(n164), .B(n163), .Z(n180) );
  XNOR U442 ( .A(n187), .B(n188), .Z(n163) );
  XOR U443 ( .A(n189), .B(n190), .Z(n188) );
  AND U444 ( .A(n191), .B(n192), .Z(n189) );
  NAND U445 ( .A(n193), .B(n194), .Z(n192) );
  NANDN U446 ( .B(n195), .A(n190), .Z(n191) );
  XOR U447 ( .A(n196), .B(n197), .Z(n162) );
  AND U448 ( .A(n198), .B(n199), .Z(n197) );
  XNOR U449 ( .A(n196), .B(n200), .Z(n198) );
  XOR U450 ( .A(n166), .B(n202), .Z(n167) );
  AND U451 ( .A(g_input[15]), .B(e_input[12]), .Z(n202) );
  XOR U452 ( .A(n203), .B(n204), .Z(n166) );
  AND U453 ( .A(n205), .B(n206), .Z(n204) );
  XNOR U454 ( .A(n207), .B(n203), .Z(n205) );
  XNOR U455 ( .A(n208), .B(n168), .Z(n201) );
  NAND U456 ( .A(e_input[13]), .B(g_input[14]), .Z(n168) );
  IV U457 ( .A(n170), .Z(n208) );
  XOR U458 ( .A(n209), .B(n210), .Z(n170) );
  AND U459 ( .A(n211), .B(n212), .Z(n210) );
  XNOR U460 ( .A(n209), .B(n213), .Z(n211) );
  XNOR U461 ( .A(n178), .B(n179), .Z(n174) );
  NAND U462 ( .A(e_input[15]), .B(g_input[12]), .Z(n179) );
  XNOR U463 ( .A(n176), .B(n214), .Z(n178) );
  AND U464 ( .A(g_input[13]), .B(e_input[14]), .Z(n214) );
  XNOR U465 ( .A(n218), .B(n215), .Z(n216) );
  OR U466 ( .A(n219), .B(n220), .Z(n181) );
  XOR U467 ( .A(n222), .B(n220), .Z(n94) );
  XNOR U468 ( .A(n223), .B(n195), .Z(n199) );
  XNOR U469 ( .A(n194), .B(n193), .Z(n195) );
  NAND U470 ( .A(g_input[15]), .B(e_input[11]), .Z(n193) );
  XNOR U471 ( .A(n227), .B(n224), .Z(n225) );
  XNOR U472 ( .A(n190), .B(n196), .Z(n223) );
  XOR U473 ( .A(n228), .B(n229), .Z(n196) );
  AND U474 ( .A(n230), .B(n231), .Z(n229) );
  XNOR U475 ( .A(n228), .B(n232), .Z(n230) );
  XNOR U476 ( .A(n233), .B(n236), .Z(n235) );
  XOR U477 ( .A(n203), .B(n238), .Z(n206) );
  AND U478 ( .A(g_input[14]), .B(e_input[12]), .Z(n238) );
  XNOR U479 ( .A(n242), .B(n207), .Z(n237) );
  NAND U480 ( .A(e_input[13]), .B(g_input[13]), .Z(n207) );
  IV U481 ( .A(n209), .Z(n242) );
  XNOR U482 ( .A(n217), .B(n218), .Z(n213) );
  NAND U483 ( .A(e_input[15]), .B(g_input[11]), .Z(n218) );
  XNOR U484 ( .A(n215), .B(n246), .Z(n217) );
  AND U485 ( .A(g_input[12]), .B(e_input[14]), .Z(n246) );
  XNOR U486 ( .A(n250), .B(n247), .Z(n248) );
  OR U487 ( .A(n251), .B(n252), .Z(n219) );
  XOR U488 ( .A(n254), .B(n252), .Z(n95) );
  XOR U489 ( .A(n255), .B(n236), .Z(n231) );
  XNOR U490 ( .A(n226), .B(n227), .Z(n236) );
  NAND U491 ( .A(e_input[11]), .B(g_input[14]), .Z(n227) );
  XNOR U492 ( .A(n224), .B(n256), .Z(n226) );
  AND U493 ( .A(g_input[15]), .B(e_input[10]), .Z(n256) );
  XNOR U494 ( .A(n260), .B(n257), .Z(n258) );
  XNOR U495 ( .A(n234), .B(n228), .Z(n255) );
  XOR U496 ( .A(n261), .B(n262), .Z(n228) );
  AND U497 ( .A(n263), .B(n264), .Z(n262) );
  XNOR U498 ( .A(n261), .B(n265), .Z(n263) );
  XOR U499 ( .A(n233), .B(n266), .Z(n234) );
  ANDN U500 ( .A(n267), .B(n268), .Z(n266) );
  XOR U501 ( .A(n269), .B(n270), .Z(n233) );
  AND U502 ( .A(n271), .B(n272), .Z(n270) );
  XNOR U503 ( .A(n269), .B(n273), .Z(n272) );
  XOR U504 ( .A(n239), .B(n275), .Z(n240) );
  AND U505 ( .A(g_input[13]), .B(e_input[12]), .Z(n275) );
  XNOR U506 ( .A(n279), .B(n241), .Z(n274) );
  NAND U507 ( .A(e_input[13]), .B(g_input[12]), .Z(n241) );
  IV U508 ( .A(n243), .Z(n279) );
  XNOR U509 ( .A(n249), .B(n250), .Z(n245) );
  NAND U510 ( .A(e_input[15]), .B(g_input[10]), .Z(n250) );
  XNOR U511 ( .A(n247), .B(n283), .Z(n249) );
  AND U512 ( .A(g_input[11]), .B(e_input[14]), .Z(n283) );
  XOR U513 ( .A(n284), .B(n285), .Z(n247) );
  ANDN U514 ( .A(n286), .B(n287), .Z(n285) );
  XNOR U515 ( .A(n288), .B(n284), .Z(n286) );
  NANDN U516 ( .B(n289), .A(n290), .Z(n251) );
  XOR U517 ( .A(n292), .B(n289), .Z(n96) );
  XOR U518 ( .A(n293), .B(n273), .Z(n264) );
  XNOR U519 ( .A(n259), .B(n260), .Z(n273) );
  NAND U520 ( .A(e_input[11]), .B(g_input[13]), .Z(n260) );
  XNOR U521 ( .A(n257), .B(n294), .Z(n259) );
  AND U522 ( .A(g_input[14]), .B(e_input[10]), .Z(n294) );
  XNOR U523 ( .A(n298), .B(n295), .Z(n296) );
  XNOR U524 ( .A(n271), .B(n261), .Z(n293) );
  XNOR U525 ( .A(n306), .B(n268), .Z(n302) );
  NAND U526 ( .A(e_input[9]), .B(g_input[15]), .Z(n268) );
  IV U527 ( .A(n269), .Z(n306) );
  XOR U528 ( .A(n276), .B(n311), .Z(n277) );
  AND U529 ( .A(g_input[12]), .B(e_input[12]), .Z(n311) );
  XOR U530 ( .A(n312), .B(n313), .Z(n276) );
  AND U531 ( .A(n314), .B(n315), .Z(n313) );
  XNOR U532 ( .A(n316), .B(n312), .Z(n314) );
  XNOR U533 ( .A(n317), .B(n278), .Z(n310) );
  NAND U534 ( .A(e_input[13]), .B(g_input[11]), .Z(n278) );
  IV U535 ( .A(n280), .Z(n317) );
  XOR U536 ( .A(n318), .B(n319), .Z(n280) );
  AND U537 ( .A(n320), .B(n321), .Z(n319) );
  XNOR U538 ( .A(n318), .B(n322), .Z(n320) );
  XNOR U539 ( .A(n287), .B(n288), .Z(n282) );
  NAND U540 ( .A(e_input[15]), .B(g_input[9]), .Z(n288) );
  XNOR U541 ( .A(n284), .B(n323), .Z(n287) );
  AND U542 ( .A(g_input[10]), .B(e_input[14]), .Z(n323) );
  XNOR U543 ( .A(n327), .B(n324), .Z(n325) );
  XNOR U544 ( .A(n290), .B(n291), .Z(n292) );
  XOR U545 ( .A(n332), .B(n330), .Z(n97) );
  XOR U546 ( .A(n333), .B(n309), .Z(n300) );
  XNOR U547 ( .A(n297), .B(n298), .Z(n309) );
  NAND U548 ( .A(e_input[11]), .B(g_input[12]), .Z(n298) );
  XNOR U549 ( .A(n295), .B(n334), .Z(n297) );
  AND U550 ( .A(g_input[13]), .B(e_input[10]), .Z(n334) );
  XNOR U551 ( .A(n338), .B(n335), .Z(n336) );
  XNOR U552 ( .A(n308), .B(n299), .Z(n333) );
  XOR U553 ( .A(n303), .B(n343), .Z(n304) );
  AND U554 ( .A(g_input[15]), .B(e_input[8]), .Z(n343) );
  XNOR U555 ( .A(n347), .B(n305), .Z(n342) );
  NAND U556 ( .A(e_input[9]), .B(g_input[14]), .Z(n305) );
  IV U557 ( .A(n307), .Z(n347) );
  XOR U558 ( .A(n312), .B(n352), .Z(n315) );
  AND U559 ( .A(g_input[11]), .B(e_input[12]), .Z(n352) );
  XNOR U560 ( .A(n356), .B(n316), .Z(n351) );
  NAND U561 ( .A(e_input[13]), .B(g_input[10]), .Z(n316) );
  IV U562 ( .A(n318), .Z(n356) );
  XNOR U563 ( .A(n326), .B(n327), .Z(n322) );
  NAND U564 ( .A(e_input[15]), .B(g_input[8]), .Z(n327) );
  XNOR U565 ( .A(n324), .B(n360), .Z(n326) );
  AND U566 ( .A(g_input[9]), .B(e_input[14]), .Z(n360) );
  XNOR U567 ( .A(n364), .B(n361), .Z(n362) );
  XNOR U568 ( .A(n329), .B(n331), .Z(n332) );
  XNOR U569 ( .A(n365), .B(n366), .Z(n329) );
  XOR U570 ( .A(n367), .B(n368), .Z(n366) );
  AND U571 ( .A(n369), .B(n370), .Z(n367) );
  OR U572 ( .A(n371), .B(n372), .Z(n370) );
  AND U573 ( .A(n373), .B(n374), .Z(n369) );
  NAND U574 ( .A(n375), .B(n376), .Z(n374) );
  NANDN U575 ( .B(n377), .A(n368), .Z(n373) );
  XOR U576 ( .A(n378), .B(n379), .Z(n328) );
  ANDN U577 ( .A(n380), .B(n381), .Z(n379) );
  XNOR U578 ( .A(n378), .B(n382), .Z(n380) );
  XOR U579 ( .A(n384), .B(n382), .Z(n98) );
  XOR U580 ( .A(n385), .B(n350), .Z(n340) );
  XNOR U581 ( .A(n337), .B(n338), .Z(n350) );
  NAND U582 ( .A(e_input[11]), .B(g_input[11]), .Z(n338) );
  XNOR U583 ( .A(n335), .B(n386), .Z(n337) );
  AND U584 ( .A(g_input[12]), .B(e_input[10]), .Z(n386) );
  XNOR U585 ( .A(n390), .B(n387), .Z(n388) );
  XNOR U586 ( .A(n349), .B(n339), .Z(n385) );
  XOR U587 ( .A(n391), .B(n392), .Z(n339) );
  AND U588 ( .A(n393), .B(n394), .Z(n392) );
  XNOR U589 ( .A(n391), .B(n395), .Z(n393) );
  XOR U590 ( .A(n344), .B(n397), .Z(n345) );
  AND U591 ( .A(g_input[14]), .B(e_input[8]), .Z(n397) );
  XNOR U592 ( .A(n401), .B(n346), .Z(n396) );
  NAND U593 ( .A(e_input[9]), .B(g_input[13]), .Z(n346) );
  IV U594 ( .A(n348), .Z(n401) );
  XOR U595 ( .A(n353), .B(n406), .Z(n354) );
  AND U596 ( .A(g_input[10]), .B(e_input[12]), .Z(n406) );
  XNOR U597 ( .A(n410), .B(n355), .Z(n405) );
  NAND U598 ( .A(e_input[13]), .B(g_input[9]), .Z(n355) );
  IV U599 ( .A(n357), .Z(n410) );
  XOR U600 ( .A(n411), .B(n412), .Z(n357) );
  AND U601 ( .A(n413), .B(n414), .Z(n412) );
  XNOR U602 ( .A(n411), .B(n415), .Z(n413) );
  XNOR U603 ( .A(n363), .B(n364), .Z(n359) );
  NAND U604 ( .A(e_input[15]), .B(g_input[7]), .Z(n364) );
  XNOR U605 ( .A(n361), .B(n416), .Z(n363) );
  AND U606 ( .A(g_input[8]), .B(e_input[14]), .Z(n416) );
  XNOR U607 ( .A(n420), .B(n417), .Z(n418) );
  XOR U608 ( .A(n381), .B(n383), .Z(n384) );
  XNOR U609 ( .A(n421), .B(n372), .Z(n381) );
  XNOR U610 ( .A(n377), .B(n368), .Z(n372) );
  XNOR U611 ( .A(n376), .B(n375), .Z(n377) );
  NAND U612 ( .A(e_input[7]), .B(g_input[15]), .Z(n375) );
  XNOR U613 ( .A(n428), .B(n425), .Z(n426) );
  OR U614 ( .A(n429), .B(n430), .Z(n371) );
  XOR U615 ( .A(n435), .B(n433), .Z(n99) );
  XOR U616 ( .A(n436), .B(n404), .Z(n394) );
  XNOR U617 ( .A(n389), .B(n390), .Z(n404) );
  NAND U618 ( .A(e_input[11]), .B(g_input[10]), .Z(n390) );
  XNOR U619 ( .A(n387), .B(n437), .Z(n389) );
  AND U620 ( .A(g_input[11]), .B(e_input[10]), .Z(n437) );
  XNOR U621 ( .A(n441), .B(n438), .Z(n439) );
  XNOR U622 ( .A(n403), .B(n391), .Z(n436) );
  XOR U623 ( .A(n398), .B(n446), .Z(n399) );
  AND U624 ( .A(g_input[13]), .B(e_input[8]), .Z(n446) );
  XNOR U625 ( .A(n450), .B(n400), .Z(n445) );
  NAND U626 ( .A(e_input[9]), .B(g_input[12]), .Z(n400) );
  IV U627 ( .A(n402), .Z(n450) );
  XOR U628 ( .A(n451), .B(n452), .Z(n402) );
  AND U629 ( .A(n453), .B(n454), .Z(n452) );
  XNOR U630 ( .A(n451), .B(n455), .Z(n454) );
  XOR U631 ( .A(n407), .B(n457), .Z(n408) );
  AND U632 ( .A(g_input[9]), .B(e_input[12]), .Z(n457) );
  XNOR U633 ( .A(n461), .B(n409), .Z(n456) );
  NAND U634 ( .A(e_input[13]), .B(g_input[8]), .Z(n409) );
  IV U635 ( .A(n411), .Z(n461) );
  XNOR U636 ( .A(n419), .B(n420), .Z(n415) );
  NAND U637 ( .A(e_input[15]), .B(g_input[6]), .Z(n420) );
  XNOR U638 ( .A(n417), .B(n465), .Z(n419) );
  AND U639 ( .A(g_input[7]), .B(e_input[14]), .Z(n465) );
  XNOR U640 ( .A(n469), .B(n466), .Z(n467) );
  XNOR U641 ( .A(n432), .B(n434), .Z(n435) );
  XOR U642 ( .A(n470), .B(n430), .Z(n432) );
  XOR U643 ( .A(n422), .B(n471), .Z(n423) );
  ANDN U644 ( .A(n472), .B(n473), .Z(n471) );
  XNOR U645 ( .A(n427), .B(n428), .Z(n424) );
  NAND U646 ( .A(g_input[14]), .B(e_input[7]), .Z(n428) );
  XNOR U647 ( .A(n425), .B(n477), .Z(n427) );
  AND U648 ( .A(e_input[6]), .B(g_input[15]), .Z(n477) );
  XNOR U649 ( .A(n481), .B(n478), .Z(n479) );
  NANDN U650 ( .B(n482), .A(n483), .Z(n429) );
  XOR U651 ( .A(n484), .B(n485), .Z(n431) );
  AND U652 ( .A(n486), .B(n487), .Z(n485) );
  XNOR U653 ( .A(n484), .B(n488), .Z(n487) );
  XOR U654 ( .A(n490), .B(n488), .Z(n100) );
  XOR U655 ( .A(n491), .B(n455), .Z(n443) );
  XNOR U656 ( .A(n440), .B(n441), .Z(n455) );
  NAND U657 ( .A(e_input[11]), .B(g_input[9]), .Z(n441) );
  XNOR U658 ( .A(n438), .B(n492), .Z(n440) );
  AND U659 ( .A(g_input[10]), .B(e_input[10]), .Z(n492) );
  XNOR U660 ( .A(n496), .B(n493), .Z(n494) );
  XNOR U661 ( .A(n453), .B(n442), .Z(n491) );
  XOR U662 ( .A(n447), .B(n501), .Z(n448) );
  AND U663 ( .A(g_input[12]), .B(e_input[8]), .Z(n501) );
  XNOR U664 ( .A(n505), .B(n449), .Z(n500) );
  NAND U665 ( .A(e_input[9]), .B(g_input[11]), .Z(n449) );
  IV U666 ( .A(n451), .Z(n505) );
  XOR U667 ( .A(n458), .B(n510), .Z(n459) );
  AND U668 ( .A(g_input[8]), .B(e_input[12]), .Z(n510) );
  XOR U669 ( .A(n511), .B(n512), .Z(n458) );
  AND U670 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U671 ( .A(n515), .B(n511), .Z(n513) );
  XNOR U672 ( .A(n516), .B(n460), .Z(n509) );
  NAND U673 ( .A(e_input[13]), .B(g_input[7]), .Z(n460) );
  IV U674 ( .A(n462), .Z(n516) );
  XOR U675 ( .A(n517), .B(n518), .Z(n462) );
  AND U676 ( .A(n519), .B(n520), .Z(n518) );
  XNOR U677 ( .A(n517), .B(n521), .Z(n519) );
  XNOR U678 ( .A(n468), .B(n469), .Z(n464) );
  NAND U679 ( .A(e_input[15]), .B(g_input[5]), .Z(n469) );
  XNOR U680 ( .A(n466), .B(n522), .Z(n468) );
  AND U681 ( .A(g_input[6]), .B(e_input[14]), .Z(n522) );
  XNOR U682 ( .A(n526), .B(n523), .Z(n524) );
  XNOR U683 ( .A(n486), .B(n489), .Z(n490) );
  XOR U684 ( .A(n527), .B(n482), .Z(n486) );
  XNOR U685 ( .A(n532), .B(n473), .Z(n528) );
  NAND U686 ( .A(g_input[15]), .B(e_input[5]), .Z(n473) );
  IV U687 ( .A(n474), .Z(n532) );
  XOR U688 ( .A(n533), .B(n534), .Z(n474) );
  AND U689 ( .A(n535), .B(n536), .Z(n534) );
  XNOR U690 ( .A(n533), .B(n537), .Z(n535) );
  XNOR U691 ( .A(n480), .B(n481), .Z(n476) );
  NAND U692 ( .A(g_input[13]), .B(e_input[7]), .Z(n481) );
  XNOR U693 ( .A(n478), .B(n538), .Z(n480) );
  AND U694 ( .A(e_input[6]), .B(g_input[14]), .Z(n538) );
  XNOR U695 ( .A(n542), .B(n539), .Z(n540) );
  XNOR U696 ( .A(n483), .B(n484), .Z(n527) );
  XOR U697 ( .A(n543), .B(n544), .Z(n484) );
  ANDN U698 ( .A(n545), .B(n546), .Z(n544) );
  XNOR U699 ( .A(n543), .B(n547), .Z(n545) );
  XOR U700 ( .A(n552), .B(n547), .Z(n101) );
  XOR U701 ( .A(n553), .B(n508), .Z(n498) );
  XNOR U702 ( .A(n495), .B(n496), .Z(n508) );
  NAND U703 ( .A(e_input[11]), .B(g_input[8]), .Z(n496) );
  XNOR U704 ( .A(n493), .B(n554), .Z(n495) );
  AND U705 ( .A(g_input[9]), .B(e_input[10]), .Z(n554) );
  XNOR U706 ( .A(n558), .B(n555), .Z(n556) );
  XNOR U707 ( .A(n507), .B(n497), .Z(n553) );
  XOR U708 ( .A(n502), .B(n563), .Z(n503) );
  AND U709 ( .A(g_input[11]), .B(e_input[8]), .Z(n563) );
  XOR U710 ( .A(n564), .B(n565), .Z(n502) );
  AND U711 ( .A(n566), .B(n567), .Z(n565) );
  XNOR U712 ( .A(n568), .B(n564), .Z(n566) );
  XNOR U713 ( .A(n569), .B(n504), .Z(n562) );
  NAND U714 ( .A(e_input[9]), .B(g_input[10]), .Z(n504) );
  IV U715 ( .A(n506), .Z(n569) );
  XOR U716 ( .A(n511), .B(n574), .Z(n514) );
  AND U717 ( .A(g_input[7]), .B(e_input[12]), .Z(n574) );
  XNOR U718 ( .A(n578), .B(n515), .Z(n573) );
  NAND U719 ( .A(e_input[13]), .B(g_input[6]), .Z(n515) );
  IV U720 ( .A(n517), .Z(n578) );
  XNOR U721 ( .A(n525), .B(n526), .Z(n521) );
  NAND U722 ( .A(e_input[15]), .B(g_input[4]), .Z(n526) );
  XNOR U723 ( .A(n523), .B(n582), .Z(n525) );
  AND U724 ( .A(g_input[5]), .B(e_input[14]), .Z(n582) );
  XNOR U725 ( .A(n586), .B(n583), .Z(n584) );
  XNOR U726 ( .A(n546), .B(n551), .Z(n552) );
  XOR U727 ( .A(n587), .B(n550), .Z(n546) );
  XOR U728 ( .A(n529), .B(n589), .Z(n530) );
  AND U729 ( .A(e_input[4]), .B(g_input[15]), .Z(n589) );
  XNOR U730 ( .A(n593), .B(n531), .Z(n588) );
  NAND U731 ( .A(g_input[14]), .B(e_input[5]), .Z(n531) );
  IV U732 ( .A(n533), .Z(n593) );
  XOR U733 ( .A(n594), .B(n595), .Z(n533) );
  AND U734 ( .A(n596), .B(n597), .Z(n595) );
  XNOR U735 ( .A(n594), .B(n598), .Z(n596) );
  XNOR U736 ( .A(n541), .B(n542), .Z(n537) );
  NAND U737 ( .A(g_input[12]), .B(e_input[7]), .Z(n542) );
  XNOR U738 ( .A(n539), .B(n599), .Z(n541) );
  AND U739 ( .A(e_input[6]), .B(g_input[13]), .Z(n599) );
  XNOR U740 ( .A(n603), .B(n600), .Z(n601) );
  XNOR U741 ( .A(n549), .B(n543), .Z(n587) );
  XNOR U742 ( .A(n607), .B(n608), .Z(n549) );
  XOR U743 ( .A(n609), .B(n610), .Z(n608) );
  AND U744 ( .A(n611), .B(n612), .Z(n609) );
  NAND U745 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U746 ( .B(n615), .A(n610), .Z(n611) );
  XOR U747 ( .A(n620), .B(n606), .Z(n102) );
  XOR U748 ( .A(n621), .B(n572), .Z(n560) );
  XNOR U749 ( .A(n557), .B(n558), .Z(n572) );
  NAND U750 ( .A(e_input[11]), .B(g_input[7]), .Z(n558) );
  XNOR U751 ( .A(n555), .B(n622), .Z(n557) );
  AND U752 ( .A(g_input[8]), .B(e_input[10]), .Z(n622) );
  XNOR U753 ( .A(n626), .B(n623), .Z(n624) );
  XNOR U754 ( .A(n571), .B(n559), .Z(n621) );
  XOR U755 ( .A(n564), .B(n631), .Z(n567) );
  AND U756 ( .A(g_input[10]), .B(e_input[8]), .Z(n631) );
  XNOR U757 ( .A(n635), .B(n568), .Z(n630) );
  NAND U758 ( .A(e_input[9]), .B(g_input[9]), .Z(n568) );
  IV U759 ( .A(n570), .Z(n635) );
  XOR U760 ( .A(n575), .B(n640), .Z(n576) );
  AND U761 ( .A(g_input[6]), .B(e_input[12]), .Z(n640) );
  XNOR U762 ( .A(n644), .B(n577), .Z(n639) );
  NAND U763 ( .A(e_input[13]), .B(g_input[5]), .Z(n577) );
  IV U764 ( .A(n579), .Z(n644) );
  XNOR U765 ( .A(n585), .B(n586), .Z(n581) );
  NAND U766 ( .A(e_input[15]), .B(g_input[3]), .Z(n586) );
  XNOR U767 ( .A(n583), .B(n648), .Z(n585) );
  AND U768 ( .A(g_input[4]), .B(e_input[14]), .Z(n648) );
  XNOR U769 ( .A(n652), .B(n649), .Z(n650) );
  XOR U770 ( .A(n605), .B(n619), .Z(n620) );
  XOR U771 ( .A(n653), .B(n618), .Z(n605) );
  XOR U772 ( .A(n590), .B(n655), .Z(n591) );
  AND U773 ( .A(e_input[4]), .B(g_input[14]), .Z(n655) );
  XNOR U774 ( .A(n659), .B(n592), .Z(n654) );
  NAND U775 ( .A(g_input[13]), .B(e_input[5]), .Z(n592) );
  IV U776 ( .A(n594), .Z(n659) );
  XOR U777 ( .A(n660), .B(n661), .Z(n594) );
  AND U778 ( .A(n662), .B(n663), .Z(n661) );
  XNOR U779 ( .A(n660), .B(n664), .Z(n662) );
  XNOR U780 ( .A(n602), .B(n603), .Z(n598) );
  NAND U781 ( .A(g_input[11]), .B(e_input[7]), .Z(n603) );
  XNOR U782 ( .A(n600), .B(n665), .Z(n602) );
  AND U783 ( .A(e_input[6]), .B(g_input[12]), .Z(n665) );
  XNOR U784 ( .A(n669), .B(n666), .Z(n667) );
  XOR U785 ( .A(n617), .B(n604), .Z(n653) );
  XOR U786 ( .A(n673), .B(n615), .Z(n617) );
  XNOR U787 ( .A(n614), .B(n613), .Z(n615) );
  NAND U788 ( .A(e_input[3]), .B(g_input[15]), .Z(n613) );
  XNOR U789 ( .A(n677), .B(n674), .Z(n675) );
  XNOR U790 ( .A(n610), .B(n616), .Z(n673) );
  XNOR U791 ( .A(n681), .B(n684), .Z(n683) );
  XOR U792 ( .A(o_reg[1]), .B(n686), .Z(o[0]) );
  XOR U793 ( .A(n688), .B(n680), .Z(n671) );
  XOR U794 ( .A(n656), .B(n690), .Z(n657) );
  AND U795 ( .A(e_input[4]), .B(g_input[13]), .Z(n690) );
  XNOR U796 ( .A(n694), .B(n658), .Z(n689) );
  NAND U797 ( .A(g_input[12]), .B(e_input[5]), .Z(n658) );
  IV U798 ( .A(n660), .Z(n694) );
  XNOR U799 ( .A(n668), .B(n669), .Z(n664) );
  NAND U800 ( .A(g_input[10]), .B(e_input[7]), .Z(n669) );
  XNOR U801 ( .A(n666), .B(n698), .Z(n668) );
  AND U802 ( .A(e_input[6]), .B(g_input[11]), .Z(n698) );
  XNOR U803 ( .A(n702), .B(n699), .Z(n700) );
  XNOR U804 ( .A(n679), .B(n670), .Z(n688) );
  XOR U805 ( .A(n706), .B(n684), .Z(n679) );
  XNOR U806 ( .A(n676), .B(n677), .Z(n684) );
  NAND U807 ( .A(g_input[14]), .B(e_input[3]), .Z(n677) );
  XNOR U808 ( .A(n674), .B(n707), .Z(n676) );
  AND U809 ( .A(e_input[2]), .B(g_input[15]), .Z(n707) );
  XNOR U810 ( .A(n711), .B(n708), .Z(n709) );
  XNOR U811 ( .A(n682), .B(n678), .Z(n706) );
  XOR U812 ( .A(n681), .B(n715), .Z(n682) );
  ANDN U813 ( .A(n716), .B(n717), .Z(n715) );
  XNOR U814 ( .A(n672), .B(n721), .Z(n687) );
  IV U815 ( .A(n685), .Z(n721) );
  AND U816 ( .A(n722), .B(o_reg[0]), .Z(n685) );
  XNOR U817 ( .A(n704), .B(n705), .Z(n722) );
  XOR U818 ( .A(n725), .B(n714), .Z(n704) );
  XOR U819 ( .A(n691), .B(n727), .Z(n692) );
  AND U820 ( .A(e_input[4]), .B(g_input[12]), .Z(n727) );
  XNOR U821 ( .A(n731), .B(n693), .Z(n726) );
  NAND U822 ( .A(g_input[11]), .B(e_input[5]), .Z(n693) );
  IV U823 ( .A(n695), .Z(n731) );
  XNOR U824 ( .A(n701), .B(n702), .Z(n697) );
  NAND U825 ( .A(g_input[9]), .B(e_input[7]), .Z(n702) );
  XNOR U826 ( .A(n699), .B(n735), .Z(n701) );
  AND U827 ( .A(e_input[6]), .B(g_input[10]), .Z(n735) );
  XNOR U828 ( .A(n739), .B(n736), .Z(n737) );
  XNOR U829 ( .A(n713), .B(n703), .Z(n725) );
  XOR U830 ( .A(n740), .B(n741), .Z(n703) );
  XOR U831 ( .A(n742), .B(n720), .Z(n713) );
  XNOR U832 ( .A(n710), .B(n711), .Z(n720) );
  NAND U833 ( .A(g_input[13]), .B(e_input[3]), .Z(n711) );
  XNOR U834 ( .A(n708), .B(n743), .Z(n710) );
  AND U835 ( .A(e_input[2]), .B(g_input[14]), .Z(n743) );
  XNOR U836 ( .A(n747), .B(n744), .Z(n745) );
  XNOR U837 ( .A(n719), .B(n712), .Z(n742) );
  XOR U838 ( .A(n748), .B(n749), .Z(n712) );
  AND U839 ( .A(n750), .B(n751), .Z(n749) );
  XOR U840 ( .A(n752), .B(n753), .Z(n751) );
  XOR U841 ( .A(n748), .B(n754), .Z(n753) );
  XOR U842 ( .A(n733), .B(n755), .Z(n750) );
  XOR U843 ( .A(n748), .B(n734), .Z(n755) );
  NAND U844 ( .A(e_input[7]), .B(g_input[8]), .Z(n739) );
  XOR U845 ( .A(n736), .B(n756), .Z(n738) );
  AND U846 ( .A(e_input[6]), .B(g_input[9]), .Z(n756) );
  XNOR U847 ( .A(n760), .B(n757), .Z(n758) );
  XOR U848 ( .A(n728), .B(n762), .Z(n729) );
  AND U849 ( .A(e_input[4]), .B(g_input[11]), .Z(n762) );
  XNOR U850 ( .A(n766), .B(n730), .Z(n761) );
  NAND U851 ( .A(g_input[10]), .B(e_input[5]), .Z(n730) );
  IV U852 ( .A(n732), .Z(n766) );
  XOR U853 ( .A(n770), .B(n771), .Z(n748) );
  AND U854 ( .A(n772), .B(n773), .Z(n771) );
  XOR U855 ( .A(n774), .B(n775), .Z(n773) );
  XOR U856 ( .A(n770), .B(n776), .Z(n775) );
  XOR U857 ( .A(n768), .B(n777), .Z(n772) );
  XOR U858 ( .A(n770), .B(n769), .Z(n777) );
  NAND U859 ( .A(e_input[7]), .B(g_input[7]), .Z(n760) );
  XOR U860 ( .A(n757), .B(n778), .Z(n759) );
  AND U861 ( .A(g_input[8]), .B(e_input[6]), .Z(n778) );
  XNOR U862 ( .A(n782), .B(n779), .Z(n780) );
  XOR U863 ( .A(n763), .B(n784), .Z(n764) );
  AND U864 ( .A(e_input[4]), .B(g_input[10]), .Z(n784) );
  XNOR U865 ( .A(n788), .B(n765), .Z(n783) );
  NAND U866 ( .A(g_input[9]), .B(e_input[5]), .Z(n765) );
  IV U867 ( .A(n767), .Z(n788) );
  XOR U868 ( .A(n789), .B(n790), .Z(n767) );
  AND U869 ( .A(n791), .B(n792), .Z(n790) );
  XOR U870 ( .A(n793), .B(n789), .Z(n792) );
  XOR U871 ( .A(n794), .B(n795), .Z(n770) );
  AND U872 ( .A(n796), .B(n797), .Z(n795) );
  XOR U873 ( .A(n798), .B(n799), .Z(n797) );
  XOR U874 ( .A(n794), .B(n800), .Z(n799) );
  XOR U875 ( .A(n791), .B(n801), .Z(n796) );
  XOR U876 ( .A(n794), .B(n793), .Z(n801) );
  NAND U877 ( .A(e_input[7]), .B(g_input[6]), .Z(n782) );
  XOR U878 ( .A(n779), .B(n802), .Z(n781) );
  AND U879 ( .A(g_input[7]), .B(e_input[6]), .Z(n802) );
  XNOR U880 ( .A(n806), .B(n803), .Z(n804) );
  XOR U881 ( .A(n785), .B(n808), .Z(n786) );
  AND U882 ( .A(e_input[4]), .B(g_input[9]), .Z(n808) );
  XNOR U883 ( .A(n812), .B(n787), .Z(n807) );
  NAND U884 ( .A(e_input[5]), .B(g_input[8]), .Z(n787) );
  IV U885 ( .A(n789), .Z(n812) );
  XOR U886 ( .A(n813), .B(n814), .Z(n789) );
  AND U887 ( .A(n815), .B(n816), .Z(n814) );
  XOR U888 ( .A(n817), .B(n813), .Z(n816) );
  XOR U889 ( .A(n818), .B(n819), .Z(n794) );
  AND U890 ( .A(n820), .B(n821), .Z(n819) );
  XOR U891 ( .A(n822), .B(n823), .Z(n821) );
  XOR U892 ( .A(n818), .B(n824), .Z(n823) );
  XOR U893 ( .A(n815), .B(n825), .Z(n820) );
  XOR U894 ( .A(n818), .B(n817), .Z(n825) );
  NAND U895 ( .A(e_input[7]), .B(g_input[5]), .Z(n806) );
  XOR U896 ( .A(n803), .B(n826), .Z(n805) );
  AND U897 ( .A(g_input[6]), .B(e_input[6]), .Z(n826) );
  XNOR U898 ( .A(n830), .B(n827), .Z(n828) );
  XOR U899 ( .A(n809), .B(n832), .Z(n810) );
  AND U900 ( .A(g_input[8]), .B(e_input[4]), .Z(n832) );
  XNOR U901 ( .A(n836), .B(n811), .Z(n831) );
  NAND U902 ( .A(e_input[5]), .B(g_input[7]), .Z(n811) );
  IV U903 ( .A(n813), .Z(n836) );
  XOR U904 ( .A(n840), .B(n841), .Z(n818) );
  AND U905 ( .A(n842), .B(n843), .Z(n841) );
  XOR U906 ( .A(n844), .B(n845), .Z(n843) );
  XOR U907 ( .A(n840), .B(n846), .Z(n845) );
  XOR U908 ( .A(n838), .B(n847), .Z(n842) );
  XOR U909 ( .A(n840), .B(n839), .Z(n847) );
  NAND U910 ( .A(e_input[7]), .B(g_input[4]), .Z(n830) );
  XOR U911 ( .A(n827), .B(n848), .Z(n829) );
  AND U912 ( .A(g_input[5]), .B(e_input[6]), .Z(n848) );
  XNOR U913 ( .A(n852), .B(n849), .Z(n850) );
  XOR U914 ( .A(n833), .B(n854), .Z(n834) );
  AND U915 ( .A(g_input[7]), .B(e_input[4]), .Z(n854) );
  XOR U916 ( .A(n855), .B(n856), .Z(n833) );
  AND U917 ( .A(n857), .B(n858), .Z(n856) );
  XNOR U918 ( .A(n859), .B(n855), .Z(n857) );
  XNOR U919 ( .A(n860), .B(n835), .Z(n853) );
  NAND U920 ( .A(e_input[5]), .B(g_input[6]), .Z(n835) );
  IV U921 ( .A(n837), .Z(n860) );
  XOR U922 ( .A(n864), .B(n865), .Z(n840) );
  AND U923 ( .A(n866), .B(n867), .Z(n865) );
  XOR U924 ( .A(n868), .B(n869), .Z(n867) );
  XOR U925 ( .A(n864), .B(n870), .Z(n869) );
  XOR U926 ( .A(n862), .B(n871), .Z(n866) );
  XOR U927 ( .A(n864), .B(n863), .Z(n871) );
  NAND U928 ( .A(e_input[7]), .B(g_input[3]), .Z(n852) );
  XOR U929 ( .A(n849), .B(n872), .Z(n851) );
  AND U930 ( .A(g_input[4]), .B(e_input[6]), .Z(n872) );
  XNOR U931 ( .A(n876), .B(n873), .Z(n874) );
  XOR U932 ( .A(n855), .B(n878), .Z(n858) );
  AND U933 ( .A(g_input[6]), .B(e_input[4]), .Z(n878) );
  XNOR U934 ( .A(n882), .B(n859), .Z(n877) );
  NAND U935 ( .A(e_input[5]), .B(g_input[5]), .Z(n859) );
  IV U936 ( .A(n861), .Z(n882) );
  XOR U937 ( .A(n886), .B(n887), .Z(n864) );
  AND U938 ( .A(n888), .B(n889), .Z(n887) );
  XOR U939 ( .A(n890), .B(n891), .Z(n889) );
  XOR U940 ( .A(n886), .B(n892), .Z(n891) );
  XOR U941 ( .A(n884), .B(n893), .Z(n888) );
  XOR U942 ( .A(n886), .B(n885), .Z(n893) );
  NAND U943 ( .A(e_input[7]), .B(g_input[2]), .Z(n876) );
  XOR U944 ( .A(n873), .B(n894), .Z(n875) );
  AND U945 ( .A(g_input[3]), .B(e_input[6]), .Z(n894) );
  XNOR U946 ( .A(n898), .B(n895), .Z(n896) );
  XOR U947 ( .A(n899), .B(n900), .Z(n884) );
  IV U948 ( .A(n880), .Z(n900) );
  XOR U949 ( .A(n879), .B(n901), .Z(n880) );
  AND U950 ( .A(g_input[5]), .B(e_input[4]), .Z(n901) );
  XNOR U951 ( .A(n905), .B(n881), .Z(n899) );
  NAND U952 ( .A(e_input[5]), .B(g_input[4]), .Z(n881) );
  IV U953 ( .A(n883), .Z(n905) );
  XOR U954 ( .A(n906), .B(n907), .Z(n883) );
  AND U955 ( .A(n908), .B(n909), .Z(n907) );
  XNOR U956 ( .A(n906), .B(n910), .Z(n908) );
  XOR U957 ( .A(n912), .B(n913), .Z(n741) );
  XNOR U958 ( .A(n914), .B(n911), .Z(n912) );
  XOR U959 ( .A(n902), .B(n916), .Z(n903) );
  AND U960 ( .A(g_input[4]), .B(e_input[4]), .Z(n916) );
  XOR U961 ( .A(n919), .B(n917), .Z(n918) );
  AND U962 ( .A(g_input[3]), .B(e_input[4]), .Z(n919) );
  AND U963 ( .A(g_input[2]), .B(e_input[5]), .Z(n920) );
  XNOR U964 ( .A(n924), .B(n921), .Z(n922) );
  XNOR U965 ( .A(n925), .B(n904), .Z(n915) );
  NAND U966 ( .A(e_input[5]), .B(g_input[3]), .Z(n904) );
  IV U967 ( .A(n906), .Z(n925) );
  NAND U968 ( .A(e_input[5]), .B(g_input[1]), .Z(n924) );
  XOR U969 ( .A(n921), .B(n926), .Z(n923) );
  AND U970 ( .A(g_input[2]), .B(e_input[4]), .Z(n926) );
  AND U971 ( .A(n927), .B(g_input[0]), .Z(n921) );
  NANDN U972 ( .B(e_input[5]), .A(n928), .Z(n927) );
  NAND U973 ( .A(g_input[1]), .B(e_input[4]), .Z(n928) );
  XNOR U974 ( .A(n897), .B(n898), .Z(n910) );
  NAND U975 ( .A(e_input[7]), .B(g_input[1]), .Z(n898) );
  XNOR U976 ( .A(n895), .B(n929), .Z(n897) );
  AND U977 ( .A(g_input[2]), .B(e_input[6]), .Z(n929) );
  AND U978 ( .A(n930), .B(g_input[0]), .Z(n895) );
  NANDN U979 ( .B(e_input[7]), .A(n931), .Z(n930) );
  NAND U980 ( .A(g_input[1]), .B(e_input[6]), .Z(n931) );
  XOR U981 ( .A(n932), .B(n933), .Z(n911) );
  XNOR U982 ( .A(n938), .B(n717), .Z(n934) );
  NAND U983 ( .A(g_input[15]), .B(e_input[1]), .Z(n717) );
  IV U984 ( .A(n718), .Z(n938) );
  NAND U985 ( .A(g_input[12]), .B(e_input[3]), .Z(n747) );
  XOR U986 ( .A(n744), .B(n940), .Z(n746) );
  AND U987 ( .A(e_input[2]), .B(g_input[13]), .Z(n940) );
  XNOR U988 ( .A(n944), .B(n941), .Z(n942) );
  XOR U989 ( .A(n935), .B(n946), .Z(n936) );
  AND U990 ( .A(e_input[0]), .B(g_input[15]), .Z(n946) );
  XNOR U991 ( .A(n950), .B(n937), .Z(n945) );
  NAND U992 ( .A(g_input[14]), .B(e_input[1]), .Z(n937) );
  IV U993 ( .A(n939), .Z(n950) );
  XOR U994 ( .A(n951), .B(n952), .Z(n939) );
  AND U995 ( .A(n776), .B(n953), .Z(n952) );
  XOR U996 ( .A(n951), .B(n774), .Z(n953) );
  NAND U997 ( .A(g_input[11]), .B(e_input[3]), .Z(n944) );
  XOR U998 ( .A(n941), .B(n954), .Z(n943) );
  AND U999 ( .A(e_input[2]), .B(g_input[12]), .Z(n954) );
  XNOR U1000 ( .A(n958), .B(n955), .Z(n956) );
  XOR U1001 ( .A(n947), .B(n960), .Z(n948) );
  AND U1002 ( .A(e_input[0]), .B(g_input[14]), .Z(n960) );
  XNOR U1003 ( .A(n964), .B(n949), .Z(n959) );
  NAND U1004 ( .A(g_input[13]), .B(e_input[1]), .Z(n949) );
  IV U1005 ( .A(n951), .Z(n964) );
  XOR U1006 ( .A(n965), .B(n966), .Z(n951) );
  AND U1007 ( .A(n800), .B(n967), .Z(n966) );
  XOR U1008 ( .A(n965), .B(n798), .Z(n967) );
  NAND U1009 ( .A(g_input[10]), .B(e_input[3]), .Z(n958) );
  XOR U1010 ( .A(n955), .B(n968), .Z(n957) );
  AND U1011 ( .A(e_input[2]), .B(g_input[11]), .Z(n968) );
  XNOR U1012 ( .A(n972), .B(n969), .Z(n970) );
  XOR U1013 ( .A(n961), .B(n974), .Z(n962) );
  AND U1014 ( .A(e_input[0]), .B(g_input[13]), .Z(n974) );
  XNOR U1015 ( .A(n978), .B(n963), .Z(n973) );
  NAND U1016 ( .A(g_input[12]), .B(e_input[1]), .Z(n963) );
  IV U1017 ( .A(n965), .Z(n978) );
  NAND U1018 ( .A(g_input[9]), .B(e_input[3]), .Z(n972) );
  XOR U1019 ( .A(n969), .B(n980), .Z(n971) );
  AND U1020 ( .A(e_input[2]), .B(g_input[10]), .Z(n980) );
  XNOR U1021 ( .A(n984), .B(n981), .Z(n982) );
  XOR U1022 ( .A(n975), .B(n986), .Z(n976) );
  AND U1023 ( .A(e_input[0]), .B(g_input[12]), .Z(n986) );
  XNOR U1024 ( .A(n990), .B(n977), .Z(n985) );
  NAND U1025 ( .A(g_input[11]), .B(e_input[1]), .Z(n977) );
  IV U1026 ( .A(n979), .Z(n990) );
  NAND U1027 ( .A(g_input[8]), .B(e_input[3]), .Z(n984) );
  XOR U1028 ( .A(n981), .B(n992), .Z(n983) );
  AND U1029 ( .A(e_input[2]), .B(g_input[9]), .Z(n992) );
  XNOR U1030 ( .A(n996), .B(n993), .Z(n994) );
  XOR U1031 ( .A(n987), .B(n998), .Z(n988) );
  AND U1032 ( .A(e_input[0]), .B(g_input[11]), .Z(n998) );
  XNOR U1033 ( .A(n1002), .B(n989), .Z(n997) );
  NAND U1034 ( .A(g_input[10]), .B(e_input[1]), .Z(n989) );
  IV U1035 ( .A(n991), .Z(n1002) );
  XOR U1036 ( .A(n1003), .B(n1004), .Z(n991) );
  AND U1037 ( .A(n870), .B(n1005), .Z(n1004) );
  XOR U1038 ( .A(n1003), .B(n868), .Z(n1005) );
  NAND U1039 ( .A(g_input[7]), .B(e_input[3]), .Z(n996) );
  XOR U1040 ( .A(n993), .B(n1006), .Z(n995) );
  AND U1041 ( .A(e_input[2]), .B(g_input[8]), .Z(n1006) );
  XNOR U1042 ( .A(n1010), .B(n1007), .Z(n1008) );
  XOR U1043 ( .A(n999), .B(n1012), .Z(n1000) );
  AND U1044 ( .A(e_input[0]), .B(g_input[10]), .Z(n1012) );
  XNOR U1045 ( .A(n1016), .B(n1001), .Z(n1011) );
  NAND U1046 ( .A(g_input[9]), .B(e_input[1]), .Z(n1001) );
  IV U1047 ( .A(n1003), .Z(n1016) );
  NAND U1048 ( .A(g_input[6]), .B(e_input[3]), .Z(n1010) );
  XOR U1049 ( .A(n1007), .B(n1018), .Z(n1009) );
  AND U1050 ( .A(e_input[2]), .B(g_input[7]), .Z(n1018) );
  XOR U1051 ( .A(n1019), .B(n1020), .Z(n1007) );
  AND U1052 ( .A(n1021), .B(n1022), .Z(n1020) );
  XNOR U1053 ( .A(n1023), .B(n1019), .Z(n1021) );
  XOR U1054 ( .A(n1013), .B(n1025), .Z(n1014) );
  AND U1055 ( .A(e_input[0]), .B(g_input[9]), .Z(n1025) );
  XNOR U1056 ( .A(n1029), .B(n1015), .Z(n1024) );
  NAND U1057 ( .A(g_input[8]), .B(e_input[1]), .Z(n1015) );
  IV U1058 ( .A(n1017), .Z(n1029) );
  XOR U1059 ( .A(n1030), .B(n1031), .Z(n1017) );
  AND U1060 ( .A(n914), .B(n1032), .Z(n1031) );
  XOR U1061 ( .A(n1030), .B(n913), .Z(n1032) );
  NAND U1062 ( .A(g_input[5]), .B(e_input[3]), .Z(n1023) );
  XOR U1063 ( .A(n1019), .B(n1033), .Z(n1022) );
  AND U1064 ( .A(e_input[2]), .B(g_input[6]), .Z(n1033) );
  XNOR U1065 ( .A(n1037), .B(n1034), .Z(n1036) );
  XOR U1066 ( .A(n1026), .B(n1039), .Z(n1027) );
  AND U1067 ( .A(e_input[0]), .B(g_input[8]), .Z(n1039) );
  XNOR U1068 ( .A(n1043), .B(n1040), .Z(n1042) );
  XNOR U1069 ( .A(n1044), .B(n1028), .Z(n1038) );
  NAND U1070 ( .A(g_input[7]), .B(e_input[1]), .Z(n1028) );
  IV U1071 ( .A(n1030), .Z(n1044) );
  XOR U1072 ( .A(n1045), .B(n1046), .Z(n1030) );
  AND U1073 ( .A(n1047), .B(n1048), .Z(n1046) );
  XOR U1074 ( .A(n1041), .B(n1049), .Z(n1048) );
  XNOR U1075 ( .A(n1043), .B(n1045), .Z(n1049) );
  NAND U1076 ( .A(g_input[6]), .B(e_input[1]), .Z(n1043) );
  XOR U1077 ( .A(n1040), .B(n1050), .Z(n1041) );
  AND U1078 ( .A(e_input[0]), .B(g_input[7]), .Z(n1050) );
  XNOR U1079 ( .A(n1054), .B(n1051), .Z(n1053) );
  XOR U1080 ( .A(n1035), .B(n1055), .Z(n1047) );
  XNOR U1081 ( .A(n1037), .B(n1045), .Z(n1055) );
  NAND U1082 ( .A(e_input[3]), .B(g_input[4]), .Z(n1037) );
  XOR U1083 ( .A(n1034), .B(n1056), .Z(n1035) );
  AND U1084 ( .A(e_input[2]), .B(g_input[5]), .Z(n1056) );
  XNOR U1085 ( .A(n1060), .B(n1057), .Z(n1059) );
  XOR U1086 ( .A(n1061), .B(n1062), .Z(n1045) );
  AND U1087 ( .A(n1063), .B(n1064), .Z(n1062) );
  XOR U1088 ( .A(n1052), .B(n1065), .Z(n1064) );
  XNOR U1089 ( .A(n1054), .B(n1061), .Z(n1065) );
  NAND U1090 ( .A(g_input[5]), .B(e_input[1]), .Z(n1054) );
  XOR U1091 ( .A(n1051), .B(n1066), .Z(n1052) );
  AND U1092 ( .A(e_input[0]), .B(g_input[6]), .Z(n1066) );
  XNOR U1093 ( .A(n1070), .B(n1067), .Z(n1069) );
  XOR U1094 ( .A(n1058), .B(n1071), .Z(n1063) );
  XNOR U1095 ( .A(n1060), .B(n1061), .Z(n1071) );
  NAND U1096 ( .A(e_input[3]), .B(g_input[3]), .Z(n1060) );
  XOR U1097 ( .A(n1057), .B(n1072), .Z(n1058) );
  AND U1098 ( .A(g_input[4]), .B(e_input[2]), .Z(n1072) );
  XNOR U1099 ( .A(n1076), .B(n1073), .Z(n1075) );
  XOR U1100 ( .A(n1077), .B(n1078), .Z(n1061) );
  AND U1101 ( .A(n1079), .B(n1080), .Z(n1078) );
  XOR U1102 ( .A(n1068), .B(n1081), .Z(n1080) );
  XNOR U1103 ( .A(n1070), .B(n1077), .Z(n1081) );
  NAND U1104 ( .A(g_input[4]), .B(e_input[1]), .Z(n1070) );
  XOR U1105 ( .A(n1067), .B(n1082), .Z(n1068) );
  AND U1106 ( .A(e_input[0]), .B(g_input[5]), .Z(n1082) );
  XOR U1107 ( .A(n1074), .B(n1086), .Z(n1079) );
  XNOR U1108 ( .A(n1076), .B(n1077), .Z(n1086) );
  NAND U1109 ( .A(e_input[3]), .B(g_input[2]), .Z(n1076) );
  XOR U1110 ( .A(n1073), .B(n1087), .Z(n1074) );
  AND U1111 ( .A(g_input[3]), .B(e_input[2]), .Z(n1087) );
  XNOR U1112 ( .A(n1091), .B(n1088), .Z(n1089) );
  NAND U1113 ( .A(e_input[3]), .B(g_input[1]), .Z(n1091) );
  XOR U1114 ( .A(n1088), .B(n1093), .Z(n1090) );
  AND U1115 ( .A(g_input[2]), .B(e_input[2]), .Z(n1093) );
  AND U1116 ( .A(n1094), .B(g_input[0]), .Z(n1088) );
  NANDN U1117 ( .B(e_input[3]), .A(n1095), .Z(n1094) );
  NAND U1118 ( .A(g_input[1]), .B(e_input[2]), .Z(n1095) );
  XOR U1119 ( .A(n1083), .B(n1097), .Z(n1084) );
  AND U1120 ( .A(e_input[0]), .B(g_input[4]), .Z(n1097) );
  XOR U1121 ( .A(n1100), .B(n1098), .Z(n1099) );
  AND U1122 ( .A(e_input[0]), .B(g_input[3]), .Z(n1100) );
  AND U1123 ( .A(e_input[1]), .B(g_input[2]), .Z(n1101) );
  XNOR U1124 ( .A(n1105), .B(n1102), .Z(n1103) );
  XNOR U1125 ( .A(n1106), .B(n1085), .Z(n1096) );
  NAND U1126 ( .A(g_input[3]), .B(e_input[1]), .Z(n1085) );
  IV U1127 ( .A(n1092), .Z(n1106) );
  NAND U1128 ( .A(g_input[1]), .B(e_input[1]), .Z(n1105) );
  XOR U1129 ( .A(n1102), .B(n1107), .Z(n1104) );
  AND U1130 ( .A(e_input[0]), .B(g_input[2]), .Z(n1107) );
  AND U1131 ( .A(n1108), .B(g_input[0]), .Z(n1102) );
  NANDN U1132 ( .B(e_input[1]), .A(n1109), .Z(n1108) );
  NAND U1133 ( .A(g_input[1]), .B(e_input[0]), .Z(n1109) );
  XOR U1134 ( .A(n1110), .B(n638), .Z(n628) );
  XNOR U1135 ( .A(n625), .B(n626), .Z(n638) );
  NAND U1136 ( .A(e_input[11]), .B(g_input[6]), .Z(n626) );
  XNOR U1137 ( .A(n623), .B(n1111), .Z(n625) );
  AND U1138 ( .A(g_input[7]), .B(e_input[10]), .Z(n1111) );
  XNOR U1139 ( .A(n1115), .B(n1112), .Z(n1113) );
  XNOR U1140 ( .A(n637), .B(n627), .Z(n1110) );
  XOR U1141 ( .A(n1117), .B(n1118), .Z(n724) );
  XNOR U1142 ( .A(n1119), .B(n1116), .Z(n1117) );
  XOR U1143 ( .A(n1122), .B(n1123), .Z(n1116) );
  XOR U1144 ( .A(n632), .B(n1125), .Z(n633) );
  AND U1145 ( .A(g_input[9]), .B(e_input[8]), .Z(n1125) );
  XNOR U1146 ( .A(n1129), .B(n634), .Z(n1124) );
  NAND U1147 ( .A(e_input[9]), .B(g_input[8]), .Z(n634) );
  IV U1148 ( .A(n636), .Z(n1129) );
  XNOR U1149 ( .A(n1114), .B(n1115), .Z(n1118) );
  NAND U1150 ( .A(e_input[11]), .B(g_input[5]), .Z(n1115) );
  XNOR U1151 ( .A(n1112), .B(n1131), .Z(n1114) );
  AND U1152 ( .A(g_input[6]), .B(e_input[10]), .Z(n1131) );
  XNOR U1153 ( .A(n1135), .B(n1132), .Z(n1134) );
  XOR U1154 ( .A(n1126), .B(n1137), .Z(n1127) );
  AND U1155 ( .A(g_input[8]), .B(e_input[8]), .Z(n1137) );
  XNOR U1156 ( .A(n1141), .B(n1138), .Z(n1140) );
  XNOR U1157 ( .A(n1142), .B(n1128), .Z(n1136) );
  NAND U1158 ( .A(e_input[9]), .B(g_input[7]), .Z(n1128) );
  IV U1159 ( .A(n1130), .Z(n1142) );
  XOR U1160 ( .A(n1143), .B(n1144), .Z(n1130) );
  AND U1161 ( .A(n1145), .B(n1146), .Z(n1144) );
  XOR U1162 ( .A(n1139), .B(n1147), .Z(n1146) );
  XNOR U1163 ( .A(n1141), .B(n1143), .Z(n1147) );
  NAND U1164 ( .A(e_input[9]), .B(g_input[6]), .Z(n1141) );
  XOR U1165 ( .A(n1138), .B(n1148), .Z(n1139) );
  AND U1166 ( .A(g_input[7]), .B(e_input[8]), .Z(n1148) );
  XNOR U1167 ( .A(n1152), .B(n1149), .Z(n1151) );
  XOR U1168 ( .A(n1133), .B(n1153), .Z(n1145) );
  XNOR U1169 ( .A(n1135), .B(n1143), .Z(n1153) );
  NAND U1170 ( .A(e_input[11]), .B(g_input[4]), .Z(n1135) );
  XOR U1171 ( .A(n1132), .B(n1154), .Z(n1133) );
  AND U1172 ( .A(g_input[5]), .B(e_input[10]), .Z(n1154) );
  XNOR U1173 ( .A(n1158), .B(n1155), .Z(n1157) );
  XOR U1174 ( .A(n1159), .B(n1160), .Z(n1143) );
  AND U1175 ( .A(n1161), .B(n1162), .Z(n1160) );
  XOR U1176 ( .A(n1150), .B(n1163), .Z(n1162) );
  XNOR U1177 ( .A(n1152), .B(n1159), .Z(n1163) );
  NAND U1178 ( .A(e_input[9]), .B(g_input[5]), .Z(n1152) );
  XOR U1179 ( .A(n1149), .B(n1164), .Z(n1150) );
  AND U1180 ( .A(g_input[6]), .B(e_input[8]), .Z(n1164) );
  XNOR U1181 ( .A(n1168), .B(n1165), .Z(n1167) );
  XOR U1182 ( .A(n1156), .B(n1169), .Z(n1161) );
  XNOR U1183 ( .A(n1158), .B(n1159), .Z(n1169) );
  NAND U1184 ( .A(e_input[11]), .B(g_input[3]), .Z(n1158) );
  XOR U1185 ( .A(n1155), .B(n1170), .Z(n1156) );
  AND U1186 ( .A(g_input[4]), .B(e_input[10]), .Z(n1170) );
  XNOR U1187 ( .A(n1174), .B(n1171), .Z(n1173) );
  XOR U1188 ( .A(n1175), .B(n1176), .Z(n1159) );
  AND U1189 ( .A(n1177), .B(n1178), .Z(n1176) );
  XOR U1190 ( .A(n1166), .B(n1179), .Z(n1178) );
  XNOR U1191 ( .A(n1168), .B(n1175), .Z(n1179) );
  NAND U1192 ( .A(e_input[9]), .B(g_input[4]), .Z(n1168) );
  XOR U1193 ( .A(n1165), .B(n1180), .Z(n1166) );
  AND U1194 ( .A(g_input[5]), .B(e_input[8]), .Z(n1180) );
  XOR U1195 ( .A(n1172), .B(n1184), .Z(n1177) );
  XNOR U1196 ( .A(n1174), .B(n1175), .Z(n1184) );
  NAND U1197 ( .A(e_input[11]), .B(g_input[2]), .Z(n1174) );
  XOR U1198 ( .A(n1171), .B(n1185), .Z(n1172) );
  AND U1199 ( .A(g_input[3]), .B(e_input[10]), .Z(n1185) );
  XNOR U1200 ( .A(n1189), .B(n1186), .Z(n1187) );
  NAND U1201 ( .A(e_input[11]), .B(g_input[1]), .Z(n1189) );
  XOR U1202 ( .A(n1186), .B(n1191), .Z(n1188) );
  AND U1203 ( .A(g_input[2]), .B(e_input[10]), .Z(n1191) );
  AND U1204 ( .A(n1192), .B(g_input[0]), .Z(n1186) );
  NANDN U1205 ( .B(e_input[11]), .A(n1193), .Z(n1192) );
  NAND U1206 ( .A(g_input[1]), .B(e_input[10]), .Z(n1193) );
  XOR U1207 ( .A(n1181), .B(n1195), .Z(n1182) );
  AND U1208 ( .A(g_input[4]), .B(e_input[8]), .Z(n1195) );
  XOR U1209 ( .A(n1198), .B(n1196), .Z(n1197) );
  AND U1210 ( .A(g_input[3]), .B(e_input[8]), .Z(n1198) );
  AND U1211 ( .A(g_input[2]), .B(e_input[9]), .Z(n1199) );
  XNOR U1212 ( .A(n1203), .B(n1200), .Z(n1201) );
  XNOR U1213 ( .A(n1204), .B(n1183), .Z(n1194) );
  NAND U1214 ( .A(e_input[9]), .B(g_input[3]), .Z(n1183) );
  IV U1215 ( .A(n1190), .Z(n1204) );
  NAND U1216 ( .A(e_input[9]), .B(g_input[1]), .Z(n1203) );
  XOR U1217 ( .A(n1200), .B(n1205), .Z(n1202) );
  AND U1218 ( .A(g_input[2]), .B(e_input[8]), .Z(n1205) );
  AND U1219 ( .A(n1206), .B(g_input[0]), .Z(n1200) );
  NANDN U1220 ( .B(e_input[9]), .A(n1207), .Z(n1206) );
  NAND U1221 ( .A(g_input[1]), .B(e_input[8]), .Z(n1207) );
  XOR U1222 ( .A(n641), .B(n1209), .Z(n642) );
  AND U1223 ( .A(g_input[5]), .B(e_input[12]), .Z(n1209) );
  XNOR U1224 ( .A(n1213), .B(n643), .Z(n1208) );
  NAND U1225 ( .A(e_input[13]), .B(g_input[4]), .Z(n643) );
  IV U1226 ( .A(n645), .Z(n1213) );
  XOR U1227 ( .A(n1210), .B(n1216), .Z(n1211) );
  AND U1228 ( .A(g_input[4]), .B(e_input[12]), .Z(n1216) );
  XOR U1229 ( .A(n1219), .B(n1217), .Z(n1218) );
  AND U1230 ( .A(g_input[3]), .B(e_input[12]), .Z(n1219) );
  AND U1231 ( .A(g_input[2]), .B(e_input[13]), .Z(n1220) );
  XNOR U1232 ( .A(n1224), .B(n1221), .Z(n1222) );
  XNOR U1233 ( .A(n1225), .B(n1212), .Z(n1215) );
  NAND U1234 ( .A(e_input[13]), .B(g_input[3]), .Z(n1212) );
  IV U1235 ( .A(n1214), .Z(n1225) );
  XNOR U1236 ( .A(n1226), .B(n1227), .Z(n1120) );
  XOR U1237 ( .A(n1228), .B(n1224), .Z(n1214) );
  NAND U1238 ( .A(e_input[13]), .B(g_input[1]), .Z(n1224) );
  IV U1239 ( .A(n1223), .Z(n1228) );
  XOR U1240 ( .A(n1221), .B(n1229), .Z(n1223) );
  AND U1241 ( .A(g_input[2]), .B(e_input[12]), .Z(n1229) );
  AND U1242 ( .A(n1230), .B(g_input[0]), .Z(n1221) );
  NANDN U1243 ( .B(e_input[13]), .A(n1231), .Z(n1230) );
  NAND U1244 ( .A(g_input[1]), .B(e_input[12]), .Z(n1231) );
  XNOR U1245 ( .A(n651), .B(n652), .Z(n647) );
  NAND U1246 ( .A(e_input[15]), .B(g_input[2]), .Z(n652) );
  XNOR U1247 ( .A(n649), .B(n1232), .Z(n651) );
  AND U1248 ( .A(g_input[3]), .B(e_input[14]), .Z(n1232) );
  XNOR U1249 ( .A(n1233), .B(n1234), .Z(n1226) );
  AND U1250 ( .A(g_input[2]), .B(e_input[14]), .Z(n1234) );
  NAND U1251 ( .A(e_input[15]), .B(g_input[1]), .Z(n1227) );
  AND U1252 ( .A(n1235), .B(g_input[0]), .Z(n1233) );
  NANDN U1253 ( .B(e_input[15]), .A(n1236), .Z(n1235) );
  NAND U1254 ( .A(g_input[1]), .B(e_input[14]), .Z(n1236) );
endmodule

