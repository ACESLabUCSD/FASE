
module MxM_W8_N10000 ( clk, rst, A, X, Y );
  input [7:0] A;
  input [7:0] X;
  output [7:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, \add_25/carry[13] ,
         \add_25/carry[12] , \add_25/carry[11] , \add_25/carry[10] ,
         \add_25/carry[9] , \add_25/carry[8] , \add_25/carry[7] ,
         \add_25/carry[6] , \add_25/carry[5] , \add_25/carry[4] ,
         \add_25/carry[3] , \add_25/carry[2] , n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599;
  wire   [7:0] Y0;
  wire   [13:0] n;

  DFF \n_reg[0]  ( .D(n166), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n165), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n164), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n163), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n162), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n161), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n160), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \n_reg[7]  ( .D(n159), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[7]) );
  DFF \n_reg[8]  ( .D(n158), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[8]) );
  DFF \n_reg[9]  ( .D(n157), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[9]) );
  DFF \n_reg[10]  ( .D(n156), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[10]) );
  DFF \n_reg[11]  ( .D(n155), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[11]) );
  DFF \n_reg[12]  ( .D(n154), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[12]) );
  DFF \n_reg[13]  ( .D(n153), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[13]) );
  DFF \Y0_reg[0]  ( .D(n152), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n151), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n150), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n149), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n148), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n147), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n146), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n145), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y_reg[7]  ( .D(n144), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n143), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n142), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n141), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n140), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n139), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n138), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n137), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  HADDER \add_25/U1_1_6  ( .IN0(n[6]), .IN1(\add_25/carry[6] ), .COUT(
        \add_25/carry[7] ), .SUM(N13) );
  HADDER \add_25/U1_1_7  ( .IN0(n[7]), .IN1(\add_25/carry[7] ), .COUT(
        \add_25/carry[8] ), .SUM(N14) );
  HADDER \add_25/U1_1_8  ( .IN0(n[8]), .IN1(\add_25/carry[8] ), .COUT(
        \add_25/carry[9] ), .SUM(N15) );
  HADDER \add_25/U1_1_9  ( .IN0(n[9]), .IN1(\add_25/carry[9] ), .COUT(
        \add_25/carry[10] ), .SUM(N16) );
  HADDER \add_25/U1_1_10  ( .IN0(n[10]), .IN1(\add_25/carry[10] ), .COUT(
        \add_25/carry[11] ), .SUM(N17) );
  HADDER \add_25/U1_1_11  ( .IN0(n[11]), .IN1(\add_25/carry[11] ), .COUT(
        \add_25/carry[12] ), .SUM(N18) );
  HADDER \add_25/U1_1_12  ( .IN0(n[12]), .IN1(\add_25/carry[12] ), .COUT(
        \add_25/carry[13] ), .SUM(N19) );
  MUX U169 ( .IN0(n492), .IN1(n508), .SEL(n494), .F(n473) );
  MUX U170 ( .IN0(A[3]), .IN1(n557), .SEL(A[7]), .F(n167) );
  IV U171 ( .A(n167), .Z(n402) );
  MUX U172 ( .IN0(n442), .IN1(n440), .SEL(n441), .F(n397) );
  NAND U173 ( .A(n315), .B(n349), .Z(n348) );
  MUX U174 ( .IN0(n425), .IN1(n168), .SEL(n424), .F(n380) );
  IV U175 ( .A(n423), .Z(n168) );
  MUX U176 ( .IN0(n169), .IN1(n325), .SEL(n326), .F(n293) );
  IV U177 ( .A(Y0[3]), .Z(n169) );
  XOR U178 ( .A(n556), .B(A[3]), .Z(n557) );
  XNOR U179 ( .A(n544), .B(n545), .Z(n523) );
  MUX U180 ( .IN0(X[6]), .IN1(n582), .SEL(X[7]), .F(n291) );
  MUX U181 ( .IN0(X[3]), .IN1(n532), .SEL(X[7]), .F(n383) );
  MUX U182 ( .IN0(n386), .IN1(n170), .SEL(n387), .F(n338) );
  IV U183 ( .A(n388), .Z(n170) );
  XNOR U184 ( .A(n389), .B(n354), .Z(n346) );
  MUX U185 ( .IN0(n171), .IN1(n408), .SEL(n409), .F(n363) );
  IV U186 ( .A(Y0[1]), .Z(n171) );
  XOR U187 ( .A(n261), .B(n271), .Z(n269) );
  MUX U188 ( .IN0(n172), .IN1(n562), .SEL(n563), .F(n558) );
  IV U189 ( .A(n564), .Z(n172) );
  MUX U190 ( .IN0(A[4]), .IN1(n509), .SEL(A[7]), .F(n173) );
  IV U191 ( .A(n173), .Z(n356) );
  MUX U192 ( .IN0(A[5]), .IN1(n491), .SEL(A[7]), .F(n319) );
  XOR U193 ( .A(n405), .B(n444), .Z(n406) );
  MUX U194 ( .IN0(A[6]), .IN1(n463), .SEL(A[7]), .F(n292) );
  MUX U195 ( .IN0(n426), .IN1(n174), .SEL(n427), .F(n386) );
  IV U196 ( .A(n428), .Z(n174) );
  XNOR U197 ( .A(n308), .B(n309), .Z(n332) );
  XOR U198 ( .A(n293), .B(n303), .Z(n301) );
  NOR U199 ( .A(A[0]), .B(n579), .Z(n567) );
  MUX U200 ( .IN0(n175), .IN1(n456), .SEL(n457), .F(n503) );
  IV U201 ( .A(n523), .Z(n175) );
  MUX U202 ( .IN0(n558), .IN1(n561), .SEL(n559), .F(n434) );
  MUX U203 ( .IN0(n473), .IN1(n489), .SEL(n475), .F(n467) );
  MUX U204 ( .IN0(n318), .IN1(n342), .SEL(n317), .F(n280) );
  NAND U205 ( .A(n380), .B(n421), .Z(n420) );
  XNOR U206 ( .A(n442), .B(n441), .Z(n428) );
  XNOR U207 ( .A(n347), .B(n346), .Z(n340) );
  XNOR U208 ( .A(n401), .B(n400), .Z(n388) );
  MUX U209 ( .IN0(Y0[6]), .IN1(n243), .SEL(n238), .F(n231) );
  XOR U210 ( .A(n325), .B(n333), .Z(n331) );
  MUX U211 ( .IN0(A[2]), .IN1(n566), .SEL(A[7]), .F(n443) );
  XOR U212 ( .A(n533), .B(n514), .Z(n457) );
  XNOR U213 ( .A(n432), .B(n394), .Z(n400) );
  MUX U214 ( .IN0(n431), .IN1(n429), .SEL(n430), .F(n176) );
  IV U215 ( .A(n176), .Z(n385) );
  AND U216 ( .A(n286), .B(n252), .Z(n285) );
  MUX U217 ( .IN0(n177), .IN1(n340), .SEL(n339), .F(n309) );
  IV U218 ( .A(n338), .Z(n177) );
  MUX U219 ( .IN0(n178), .IN1(n363), .SEL(n364), .F(n325) );
  IV U220 ( .A(Y0[2]), .Z(n178) );
  MUX U221 ( .IN0(Y0[7]), .IN1(n231), .SEL(n232), .F(n179) );
  IV U222 ( .A(n179), .Z(n228) );
  XOR U223 ( .A(n409), .B(Y0[1]), .Z(n197) );
  ANDN U224 ( .A(n180), .B(n[0]), .Z(n166) );
  AND U225 ( .A(N8), .B(n180), .Z(n165) );
  AND U226 ( .A(N9), .B(n180), .Z(n164) );
  AND U227 ( .A(N10), .B(n180), .Z(n163) );
  AND U228 ( .A(N11), .B(n180), .Z(n162) );
  AND U229 ( .A(N12), .B(n180), .Z(n161) );
  AND U230 ( .A(N13), .B(n180), .Z(n160) );
  AND U231 ( .A(N14), .B(n180), .Z(n159) );
  AND U232 ( .A(N15), .B(n180), .Z(n158) );
  AND U233 ( .A(N16), .B(n180), .Z(n157) );
  AND U234 ( .A(N17), .B(n180), .Z(n156) );
  AND U235 ( .A(N18), .B(n180), .Z(n155) );
  AND U236 ( .A(N19), .B(n180), .Z(n154) );
  AND U237 ( .A(n180), .B(n181), .Z(n153) );
  XOR U238 ( .A(n[13]), .B(\add_25/carry[13] ), .Z(n181) );
  ANDN U239 ( .A(n182), .B(rst), .Z(n180) );
  NAND U240 ( .A(n183), .B(n184), .Z(n182) );
  AND U241 ( .A(n185), .B(n186), .Z(n184) );
  ANDN U242 ( .A(n187), .B(n188), .Z(n186) );
  NOR U243 ( .A(n189), .B(n190), .Z(n187) );
  AND U244 ( .A(n191), .B(n[13]), .Z(n185) );
  AND U245 ( .A(n[10]), .B(n[0]), .Z(n191) );
  AND U246 ( .A(n192), .B(n193), .Z(n183) );
  AND U247 ( .A(n[3]), .B(n194), .Z(n193) );
  AND U248 ( .A(n[2]), .B(n[1]), .Z(n194) );
  AND U249 ( .A(n[9]), .B(n[8]), .Z(n192) );
  NAND U250 ( .A(n195), .B(n196), .Z(n152) );
  OR U251 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U252 ( .B(n199), .A(Y0[0]), .Z(n195) );
  NAND U253 ( .A(n200), .B(n201), .Z(n151) );
  NANDN U254 ( .B(n198), .A(n202), .Z(n201) );
  NANDN U255 ( .B(n203), .A(rst), .Z(n200) );
  NAND U256 ( .A(n204), .B(n205), .Z(n150) );
  NANDN U257 ( .B(n198), .A(n206), .Z(n205) );
  NANDN U258 ( .B(n199), .A(Y0[2]), .Z(n204) );
  NAND U259 ( .A(n207), .B(n208), .Z(n149) );
  NANDN U260 ( .B(n198), .A(n209), .Z(n208) );
  NANDN U261 ( .B(n199), .A(Y0[3]), .Z(n207) );
  NAND U262 ( .A(n210), .B(n211), .Z(n148) );
  NANDN U263 ( .B(n198), .A(n212), .Z(n211) );
  NANDN U264 ( .B(n199), .A(Y0[4]), .Z(n210) );
  NAND U265 ( .A(n213), .B(n214), .Z(n147) );
  NANDN U266 ( .B(n198), .A(n215), .Z(n214) );
  NANDN U267 ( .B(n199), .A(Y0[5]), .Z(n213) );
  NAND U268 ( .A(n216), .B(n217), .Z(n146) );
  OR U269 ( .A(n218), .B(n198), .Z(n217) );
  NANDN U270 ( .B(n199), .A(Y0[6]), .Z(n216) );
  NAND U271 ( .A(n219), .B(n220), .Z(n145) );
  OR U272 ( .A(n198), .B(n221), .Z(n220) );
  NANDN U273 ( .B(n222), .A(n199), .Z(n198) );
  NANDN U274 ( .B(n199), .A(Y0[7]), .Z(n219) );
  NAND U275 ( .A(n223), .B(n224), .Z(n144) );
  NANDN U276 ( .B(n199), .A(Y[7]), .Z(n224) );
  AND U277 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U278 ( .B(n222), .A(Y[7]), .Z(n226) );
  OR U279 ( .A(n221), .B(n227), .Z(n225) );
  XOR U280 ( .A(n228), .B(n229), .Z(n221) );
  XNOR U281 ( .A(Y0[7]), .B(n230), .Z(n229) );
  NAND U282 ( .A(n233), .B(n234), .Z(n143) );
  NANDN U283 ( .B(n199), .A(Y[6]), .Z(n234) );
  AND U284 ( .A(n235), .B(n236), .Z(n233) );
  NANDN U285 ( .B(n222), .A(Y[6]), .Z(n236) );
  OR U286 ( .A(n218), .B(n227), .Z(n235) );
  XOR U287 ( .A(n232), .B(Y0[7]), .Z(n218) );
  XOR U288 ( .A(n231), .B(n230), .Z(n232) );
  NAND U289 ( .A(n239), .B(n240), .Z(n142) );
  NANDN U290 ( .B(n199), .A(Y[5]), .Z(n240) );
  AND U291 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U292 ( .B(n222), .A(Y[5]), .Z(n242) );
  NANDN U293 ( .B(n227), .A(n215), .Z(n241) );
  XNOR U294 ( .A(n238), .B(Y0[6]), .Z(n215) );
  XOR U295 ( .A(n243), .B(n244), .Z(n238) );
  ANDN U296 ( .A(n230), .B(n245), .Z(n244) );
  NANDN U297 ( .B(n246), .A(n247), .Z(n230) );
  ANDN U298 ( .A(n248), .B(n245), .Z(n246) );
  NAND U299 ( .A(n249), .B(n250), .Z(n245) );
  OR U300 ( .A(n251), .B(n252), .Z(n250) );
  AND U301 ( .A(n253), .B(n254), .Z(n249) );
  OR U302 ( .A(n255), .B(n256), .Z(n254) );
  OR U303 ( .A(n257), .B(n258), .Z(n253) );
  NOR U304 ( .A(n259), .B(n260), .Z(n248) );
  IV U305 ( .A(n237), .Z(n243) );
  XOR U306 ( .A(n261), .B(n262), .Z(n237) );
  ANDN U307 ( .A(n263), .B(n264), .Z(n262) );
  XNOR U308 ( .A(Y0[5]), .B(n261), .Z(n263) );
  NAND U309 ( .A(n265), .B(n266), .Z(n141) );
  NANDN U310 ( .B(n199), .A(Y[4]), .Z(n266) );
  AND U311 ( .A(n267), .B(n268), .Z(n265) );
  NANDN U312 ( .B(n222), .A(Y[4]), .Z(n268) );
  NANDN U313 ( .B(n227), .A(n212), .Z(n267) );
  XNOR U314 ( .A(n264), .B(Y0[5]), .Z(n212) );
  XNOR U315 ( .A(n269), .B(n270), .Z(n264) );
  AND U316 ( .A(n247), .B(n272), .Z(n271) );
  XOR U317 ( .A(n259), .B(n273), .Z(n272) );
  XOR U318 ( .A(n273), .B(n260), .Z(n259) );
  OR U319 ( .A(n274), .B(n275), .Z(n260) );
  IV U320 ( .A(n270), .Z(n273) );
  XNOR U321 ( .A(n258), .B(n257), .Z(n270) );
  OR U322 ( .A(n276), .B(n277), .Z(n257) );
  AND U323 ( .A(n278), .B(n279), .Z(n258) );
  XNOR U324 ( .A(n280), .B(n281), .Z(n279) );
  ANDN U325 ( .A(n282), .B(n283), .Z(n281) );
  XOR U326 ( .A(n280), .B(n284), .Z(n282) );
  XNOR U327 ( .A(n251), .B(n285), .Z(n278) );
  NAND U328 ( .A(n287), .B(n288), .Z(n252) );
  NANDN U329 ( .B(n289), .A(n290), .Z(n287) );
  NANDN U330 ( .B(n255), .A(n291), .Z(n286) );
  NANDN U331 ( .B(n256), .A(n292), .Z(n251) );
  XOR U332 ( .A(n293), .B(n294), .Z(n261) );
  ANDN U333 ( .A(n295), .B(n296), .Z(n294) );
  XNOR U334 ( .A(Y0[4]), .B(n293), .Z(n295) );
  NAND U335 ( .A(n297), .B(n298), .Z(n140) );
  NANDN U336 ( .B(n199), .A(Y[3]), .Z(n298) );
  AND U337 ( .A(n299), .B(n300), .Z(n297) );
  NANDN U338 ( .B(n222), .A(Y[3]), .Z(n300) );
  NANDN U339 ( .B(n227), .A(n209), .Z(n299) );
  XNOR U340 ( .A(n296), .B(Y0[4]), .Z(n209) );
  XNOR U341 ( .A(n301), .B(n302), .Z(n296) );
  AND U342 ( .A(n247), .B(n304), .Z(n303) );
  XOR U343 ( .A(n274), .B(n305), .Z(n304) );
  XOR U344 ( .A(n305), .B(n275), .Z(n274) );
  OR U345 ( .A(n306), .B(n307), .Z(n275) );
  IV U346 ( .A(n302), .Z(n305) );
  XNOR U347 ( .A(n277), .B(n276), .Z(n302) );
  OR U348 ( .A(n308), .B(n309), .Z(n276) );
  XOR U349 ( .A(n284), .B(n283), .Z(n277) );
  XOR U350 ( .A(n280), .B(n310), .Z(n283) );
  AND U351 ( .A(n311), .B(n312), .Z(n310) );
  NANDN U352 ( .B(n255), .A(n313), .Z(n312) );
  OR U353 ( .A(n314), .B(n315), .Z(n311) );
  XOR U354 ( .A(n289), .B(n290), .Z(n284) );
  NANDN U355 ( .B(n256), .A(n319), .Z(n290) );
  XNOR U356 ( .A(n288), .B(n320), .Z(n289) );
  AND U357 ( .A(n292), .B(n291), .Z(n320) );
  ANDN U358 ( .A(n321), .B(n322), .Z(n288) );
  NANDN U359 ( .B(n323), .A(n324), .Z(n321) );
  NAND U360 ( .A(n327), .B(n328), .Z(n139) );
  NANDN U361 ( .B(n199), .A(Y[2]), .Z(n328) );
  AND U362 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U363 ( .B(n222), .A(Y[2]), .Z(n330) );
  NANDN U364 ( .B(n227), .A(n206), .Z(n329) );
  XNOR U365 ( .A(n326), .B(Y0[3]), .Z(n206) );
  XNOR U366 ( .A(n331), .B(n332), .Z(n326) );
  AND U367 ( .A(n247), .B(n334), .Z(n333) );
  XOR U368 ( .A(n306), .B(n335), .Z(n334) );
  XOR U369 ( .A(n335), .B(n307), .Z(n306) );
  OR U370 ( .A(n336), .B(n337), .Z(n307) );
  IV U371 ( .A(n332), .Z(n335) );
  XOR U372 ( .A(n318), .B(n317), .Z(n308) );
  XNOR U373 ( .A(n341), .B(n342), .Z(n317) );
  IV U374 ( .A(n316), .Z(n342) );
  XOR U375 ( .A(n343), .B(n344), .Z(n316) );
  ANDN U376 ( .A(n345), .B(n346), .Z(n344) );
  XOR U377 ( .A(n343), .B(n347), .Z(n345) );
  XNOR U378 ( .A(n348), .B(n314), .Z(n341) );
  NAND U379 ( .A(n313), .B(n292), .Z(n314) );
  NANDN U380 ( .B(n255), .A(n350), .Z(n349) );
  XNOR U381 ( .A(n351), .B(n352), .Z(n315) );
  ANDN U382 ( .A(n353), .B(n354), .Z(n352) );
  XNOR U383 ( .A(n355), .B(n351), .Z(n353) );
  XOR U384 ( .A(n323), .B(n324), .Z(n318) );
  OR U385 ( .A(n356), .B(n256), .Z(n324) );
  XNOR U386 ( .A(n357), .B(n358), .Z(n323) );
  AND U387 ( .A(n319), .B(n291), .Z(n358) );
  IV U388 ( .A(n322), .Z(n357) );
  NAND U389 ( .A(n359), .B(n360), .Z(n322) );
  NANDN U390 ( .B(n361), .A(n362), .Z(n359) );
  NAND U391 ( .A(n365), .B(n366), .Z(n138) );
  NANDN U392 ( .B(n199), .A(Y[1]), .Z(n366) );
  AND U393 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U394 ( .B(n222), .A(Y[1]), .Z(n368) );
  NANDN U395 ( .B(n227), .A(n202), .Z(n367) );
  XNOR U396 ( .A(n364), .B(Y0[2]), .Z(n202) );
  XNOR U397 ( .A(n369), .B(n370), .Z(n364) );
  XOR U398 ( .A(n363), .B(n371), .Z(n369) );
  AND U399 ( .A(n247), .B(n372), .Z(n371) );
  XOR U400 ( .A(n336), .B(n373), .Z(n372) );
  XOR U401 ( .A(n373), .B(n337), .Z(n336) );
  NANDN U402 ( .B(n374), .A(n375), .Z(n337) );
  IV U403 ( .A(n370), .Z(n373) );
  XOR U404 ( .A(n340), .B(n339), .Z(n370) );
  XNOR U405 ( .A(n338), .B(n376), .Z(n339) );
  AND U406 ( .A(n377), .B(n378), .Z(n376) );
  OR U407 ( .A(n379), .B(n380), .Z(n378) );
  AND U408 ( .A(n381), .B(n382), .Z(n377) );
  NANDN U409 ( .B(n255), .A(n383), .Z(n382) );
  NAND U410 ( .A(n384), .B(n385), .Z(n381) );
  XNOR U411 ( .A(n351), .B(n390), .Z(n354) );
  AND U412 ( .A(n292), .B(n350), .Z(n390) );
  XOR U413 ( .A(n391), .B(n392), .Z(n351) );
  ANDN U414 ( .A(n393), .B(n394), .Z(n392) );
  XNOR U415 ( .A(n395), .B(n391), .Z(n393) );
  XOR U416 ( .A(n396), .B(n355), .Z(n389) );
  NAND U417 ( .A(n313), .B(n319), .Z(n355) );
  IV U418 ( .A(n343), .Z(n396) );
  XOR U419 ( .A(n397), .B(n398), .Z(n343) );
  ANDN U420 ( .A(n399), .B(n400), .Z(n398) );
  XOR U421 ( .A(n397), .B(n401), .Z(n399) );
  XNOR U422 ( .A(n361), .B(n362), .Z(n347) );
  OR U423 ( .A(n402), .B(n256), .Z(n362) );
  XNOR U424 ( .A(n360), .B(n403), .Z(n361) );
  ANDN U425 ( .A(n291), .B(n356), .Z(n403) );
  ANDN U426 ( .A(n404), .B(n405), .Z(n360) );
  NANDN U427 ( .B(n406), .A(n407), .Z(n404) );
  NAND U428 ( .A(n410), .B(n411), .Z(n137) );
  NANDN U429 ( .B(n199), .A(Y[0]), .Z(n411) );
  AND U430 ( .A(n412), .B(n413), .Z(n410) );
  NANDN U431 ( .B(n222), .A(Y[0]), .Z(n413) );
  IV U432 ( .A(n414), .Z(n222) );
  OR U433 ( .A(n227), .B(n197), .Z(n412) );
  IV U434 ( .A(Y0[1]), .Z(n203) );
  XOR U435 ( .A(n415), .B(n416), .Z(n409) );
  XNOR U436 ( .A(n417), .B(n408), .Z(n415) );
  NAND U437 ( .A(Y0[0]), .B(n374), .Z(n408) );
  NAND U438 ( .A(n418), .B(n247), .Z(n417) );
  XOR U439 ( .A(A[7]), .B(X[7]), .Z(n247) );
  XNOR U440 ( .A(n375), .B(n416), .Z(n418) );
  XNOR U441 ( .A(n374), .B(n416), .Z(n375) );
  XNOR U442 ( .A(n388), .B(n387), .Z(n416) );
  XNOR U443 ( .A(n419), .B(n384), .Z(n387) );
  XNOR U444 ( .A(n420), .B(n379), .Z(n384) );
  NAND U445 ( .A(n292), .B(n383), .Z(n379) );
  NANDN U446 ( .B(n255), .A(n422), .Z(n421) );
  XNOR U447 ( .A(n385), .B(n386), .Z(n419) );
  XNOR U448 ( .A(n391), .B(n433), .Z(n394) );
  AND U449 ( .A(n319), .B(n350), .Z(n433) );
  XOR U450 ( .A(n434), .B(n435), .Z(n391) );
  ANDN U451 ( .A(n436), .B(n437), .Z(n435) );
  XNOR U452 ( .A(n438), .B(n434), .Z(n436) );
  XOR U453 ( .A(n439), .B(n395), .Z(n432) );
  NANDN U454 ( .B(n356), .A(n313), .Z(n395) );
  IV U455 ( .A(n397), .Z(n439) );
  XNOR U456 ( .A(n406), .B(n407), .Z(n401) );
  NANDN U457 ( .B(n256), .A(n443), .Z(n407) );
  ANDN U458 ( .A(n291), .B(n402), .Z(n444) );
  NAND U459 ( .A(n445), .B(n446), .Z(n405) );
  NANDN U460 ( .B(n447), .A(n448), .Z(n445) );
  XNOR U461 ( .A(n428), .B(n427), .Z(n374) );
  XNOR U462 ( .A(n449), .B(n431), .Z(n427) );
  XNOR U463 ( .A(n424), .B(n425), .Z(n431) );
  NAND U464 ( .A(n319), .B(n383), .Z(n425) );
  XNOR U465 ( .A(n423), .B(n450), .Z(n424) );
  AND U466 ( .A(n422), .B(n292), .Z(n450) );
  XOR U467 ( .A(n451), .B(n452), .Z(n423) );
  AND U468 ( .A(n453), .B(n454), .Z(n452) );
  XNOR U469 ( .A(n455), .B(n451), .Z(n454) );
  XNOR U470 ( .A(n430), .B(n426), .Z(n449) );
  XOR U471 ( .A(n456), .B(n457), .Z(n426) );
  XOR U472 ( .A(n458), .B(n459), .Z(n430) );
  AND U473 ( .A(n460), .B(n461), .Z(n459) );
  NANDN U474 ( .B(n255), .A(n462), .Z(n461) );
  NANDN U475 ( .B(n463), .A(n464), .Z(n255) );
  AND U476 ( .A(n465), .B(A[7]), .Z(n464) );
  NANDN U477 ( .B(n466), .A(n467), .Z(n460) );
  IV U478 ( .A(n429), .Z(n458) );
  XNOR U479 ( .A(n468), .B(n469), .Z(n429) );
  AND U480 ( .A(n470), .B(n471), .Z(n469) );
  XOR U481 ( .A(n467), .B(n472), .Z(n471) );
  XNOR U482 ( .A(n466), .B(n468), .Z(n472) );
  NAND U483 ( .A(n292), .B(n462), .Z(n466) );
  XNOR U484 ( .A(n476), .B(n473), .Z(n475) );
  XOR U485 ( .A(n453), .B(n477), .Z(n470) );
  XNOR U486 ( .A(n455), .B(n468), .Z(n477) );
  NANDN U487 ( .B(n356), .A(n383), .Z(n455) );
  XOR U488 ( .A(n451), .B(n478), .Z(n453) );
  AND U489 ( .A(n422), .B(n319), .Z(n478) );
  XOR U490 ( .A(n479), .B(n480), .Z(n451) );
  AND U491 ( .A(n481), .B(n482), .Z(n480) );
  XNOR U492 ( .A(n483), .B(n479), .Z(n482) );
  XOR U493 ( .A(n484), .B(n485), .Z(n468) );
  AND U494 ( .A(n486), .B(n487), .Z(n485) );
  XOR U495 ( .A(n474), .B(n488), .Z(n487) );
  XNOR U496 ( .A(n476), .B(n484), .Z(n488) );
  NAND U497 ( .A(n319), .B(n462), .Z(n476) );
  XOR U498 ( .A(n473), .B(n489), .Z(n474) );
  AND U499 ( .A(n292), .B(X[0]), .Z(n489) );
  XNOR U500 ( .A(n465), .B(A[6]), .Z(n463) );
  NOR U501 ( .A(n490), .B(n491), .Z(n465) );
  XNOR U502 ( .A(n495), .B(n492), .Z(n494) );
  XOR U503 ( .A(n481), .B(n496), .Z(n486) );
  XNOR U504 ( .A(n483), .B(n484), .Z(n496) );
  NANDN U505 ( .B(n402), .A(n383), .Z(n483) );
  XOR U506 ( .A(n479), .B(n497), .Z(n481) );
  ANDN U507 ( .A(n422), .B(n356), .Z(n497) );
  XOR U508 ( .A(n498), .B(n499), .Z(n479) );
  AND U509 ( .A(n500), .B(n501), .Z(n499) );
  XNOR U510 ( .A(n502), .B(n498), .Z(n501) );
  XOR U511 ( .A(n503), .B(n504), .Z(n484) );
  AND U512 ( .A(n505), .B(n506), .Z(n504) );
  XOR U513 ( .A(n493), .B(n507), .Z(n506) );
  XNOR U514 ( .A(n495), .B(n503), .Z(n507) );
  NANDN U515 ( .B(n356), .A(n462), .Z(n495) );
  XOR U516 ( .A(n492), .B(n508), .Z(n493) );
  AND U517 ( .A(n319), .B(X[0]), .Z(n508) );
  XOR U518 ( .A(n490), .B(A[5]), .Z(n491) );
  NANDN U519 ( .B(n509), .A(n510), .Z(n490) );
  XOR U520 ( .A(n511), .B(n512), .Z(n492) );
  ANDN U521 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U522 ( .A(n515), .B(n511), .Z(n513) );
  XOR U523 ( .A(n500), .B(n516), .Z(n505) );
  XNOR U524 ( .A(n502), .B(n503), .Z(n516) );
  NAND U525 ( .A(n383), .B(n443), .Z(n502) );
  XOR U526 ( .A(n498), .B(n517), .Z(n500) );
  ANDN U527 ( .A(n422), .B(n402), .Z(n517) );
  XOR U528 ( .A(n518), .B(n519), .Z(n498) );
  ANDN U529 ( .A(n520), .B(n521), .Z(n519) );
  XNOR U530 ( .A(n522), .B(n518), .Z(n520) );
  XNOR U531 ( .A(n524), .B(n522), .Z(n456) );
  NAND U532 ( .A(n383), .B(n525), .Z(n522) );
  IV U533 ( .A(n521), .Z(n524) );
  XNOR U534 ( .A(n518), .B(n526), .Z(n521) );
  AND U535 ( .A(n443), .B(n422), .Z(n526) );
  AND U536 ( .A(n527), .B(A[0]), .Z(n518) );
  NANDN U537 ( .B(n383), .A(n528), .Z(n527) );
  NAND U538 ( .A(n525), .B(n422), .Z(n528) );
  XNOR U539 ( .A(n529), .B(X[2]), .Z(n422) );
  NAND U540 ( .A(n530), .B(X[7]), .Z(n529) );
  XOR U541 ( .A(n531), .B(X[2]), .Z(n530) );
  XNOR U542 ( .A(n511), .B(n534), .Z(n514) );
  ANDN U543 ( .A(X[0]), .B(n356), .Z(n534) );
  XOR U544 ( .A(n535), .B(n536), .Z(n511) );
  AND U545 ( .A(n537), .B(n538), .Z(n536) );
  XOR U546 ( .A(n539), .B(n535), .Z(n538) );
  ANDN U547 ( .A(X[0]), .B(n402), .Z(n539) );
  XOR U548 ( .A(n540), .B(n535), .Z(n537) );
  AND U549 ( .A(n462), .B(n443), .Z(n540) );
  XOR U550 ( .A(n541), .B(n542), .Z(n535) );
  ANDN U551 ( .A(n543), .B(n544), .Z(n542) );
  XNOR U552 ( .A(n545), .B(n541), .Z(n543) );
  XOR U553 ( .A(n546), .B(n515), .Z(n533) );
  NANDN U554 ( .B(n402), .A(n462), .Z(n515) );
  IV U555 ( .A(n523), .Z(n546) );
  NAND U556 ( .A(n462), .B(n525), .Z(n545) );
  XNOR U557 ( .A(n541), .B(n547), .Z(n544) );
  AND U558 ( .A(n443), .B(X[0]), .Z(n547) );
  AND U559 ( .A(n548), .B(A[0]), .Z(n541) );
  NANDN U560 ( .B(n462), .A(n549), .Z(n548) );
  NAND U561 ( .A(n525), .B(X[0]), .Z(n549) );
  XNOR U562 ( .A(n550), .B(X[1]), .Z(n462) );
  NAND U563 ( .A(n551), .B(X[7]), .Z(n550) );
  XNOR U564 ( .A(X[1]), .B(n552), .Z(n551) );
  XOR U565 ( .A(n553), .B(n554), .Z(n441) );
  IV U566 ( .A(n437), .Z(n554) );
  XNOR U567 ( .A(n434), .B(n555), .Z(n437) );
  ANDN U568 ( .A(n350), .B(n356), .Z(n555) );
  XNOR U569 ( .A(n510), .B(A[4]), .Z(n509) );
  NOR U570 ( .A(n556), .B(n557), .Z(n510) );
  XOR U571 ( .A(n560), .B(n558), .Z(n559) );
  ANDN U572 ( .A(n350), .B(n402), .Z(n560) );
  AND U573 ( .A(n443), .B(n313), .Z(n561) );
  XOR U574 ( .A(n565), .B(n438), .Z(n553) );
  NANDN U575 ( .B(n402), .A(n313), .Z(n438) );
  NANDN U576 ( .B(n566), .A(n567), .Z(n556) );
  IV U577 ( .A(n440), .Z(n565) );
  XOR U578 ( .A(n568), .B(n564), .Z(n440) );
  NAND U579 ( .A(n313), .B(n525), .Z(n564) );
  IV U580 ( .A(n563), .Z(n568) );
  XNOR U581 ( .A(n562), .B(n569), .Z(n563) );
  AND U582 ( .A(n443), .B(n350), .Z(n569) );
  AND U583 ( .A(n570), .B(A[0]), .Z(n562) );
  NANDN U584 ( .B(n313), .A(n571), .Z(n570) );
  NAND U585 ( .A(n525), .B(n350), .Z(n571) );
  XNOR U586 ( .A(n572), .B(X[4]), .Z(n350) );
  NAND U587 ( .A(n573), .B(X[7]), .Z(n572) );
  XOR U588 ( .A(n574), .B(X[4]), .Z(n573) );
  XNOR U589 ( .A(n575), .B(X[5]), .Z(n313) );
  NAND U590 ( .A(n576), .B(X[7]), .Z(n575) );
  XOR U591 ( .A(n577), .B(X[5]), .Z(n576) );
  XNOR U592 ( .A(n447), .B(n448), .Z(n442) );
  NANDN U593 ( .B(n256), .A(n525), .Z(n448) );
  XNOR U594 ( .A(n446), .B(n578), .Z(n447) );
  AND U595 ( .A(n443), .B(n291), .Z(n578) );
  XNOR U596 ( .A(n567), .B(A[2]), .Z(n566) );
  AND U597 ( .A(n580), .B(A[0]), .Z(n446) );
  NAND U598 ( .A(n581), .B(n256), .Z(n580) );
  NANDN U599 ( .B(n582), .A(n583), .Z(n256) );
  ANDN U600 ( .A(X[7]), .B(n584), .Z(n583) );
  NAND U601 ( .A(n525), .B(n291), .Z(n581) );
  XOR U602 ( .A(n584), .B(X[6]), .Z(n582) );
  OR U603 ( .A(n577), .B(n585), .Z(n584) );
  XOR U604 ( .A(n585), .B(X[5]), .Z(n577) );
  OR U605 ( .A(n574), .B(n586), .Z(n585) );
  XOR U606 ( .A(n586), .B(X[4]), .Z(n574) );
  OR U607 ( .A(n532), .B(n587), .Z(n586) );
  XOR U608 ( .A(n587), .B(X[3]), .Z(n532) );
  OR U609 ( .A(n531), .B(n588), .Z(n587) );
  XOR U610 ( .A(n588), .B(X[2]), .Z(n531) );
  NANDN U611 ( .B(X[0]), .A(n552), .Z(n588) );
  XNOR U612 ( .A(X[0]), .B(X[1]), .Z(n552) );
  XNOR U613 ( .A(n589), .B(A[1]), .Z(n525) );
  NAND U614 ( .A(n590), .B(A[7]), .Z(n589) );
  XOR U615 ( .A(A[1]), .B(n579), .Z(n590) );
  XOR U616 ( .A(A[0]), .B(A[1]), .Z(n579) );
  NANDN U617 ( .B(n414), .A(n199), .Z(n227) );
  IV U618 ( .A(rst), .Z(n199) );
  NAND U619 ( .A(n591), .B(n592), .Z(n414) );
  AND U620 ( .A(n593), .B(n594), .Z(n592) );
  ANDN U621 ( .A(n595), .B(n[3]), .Z(n594) );
  NOR U622 ( .A(n[8]), .B(n[9]), .Z(n595) );
  ANDN U623 ( .A(n596), .B(n[13]), .Z(n593) );
  NOR U624 ( .A(n[1]), .B(n[2]), .Z(n596) );
  AND U625 ( .A(n597), .B(n598), .Z(n591) );
  ANDN U626 ( .A(n599), .B(n190), .Z(n598) );
  OR U627 ( .A(n[6]), .B(n[7]), .Z(n190) );
  NOR U628 ( .A(n[0]), .B(n[10]), .Z(n599) );
  NOR U629 ( .A(n188), .B(n189), .Z(n597) );
  OR U630 ( .A(n[4]), .B(n[5]), .Z(n189) );
  OR U631 ( .A(n[12]), .B(n[11]), .Z(n188) );
endmodule

