
module MxM_TG_W8_N10000 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n166 , \_MxM/n165 , \_MxM/n164 , \_MxM/n163 , \_MxM/n162 ,
         \_MxM/n161 , \_MxM/n160 , \_MxM/n159 , \_MxM/n158 , \_MxM/n157 ,
         \_MxM/n156 , \_MxM/n155 , \_MxM/n154 , \_MxM/n153 , \_MxM/n152 ,
         \_MxM/n151 , \_MxM/n150 , \_MxM/n149 , \_MxM/n148 , \_MxM/n147 ,
         \_MxM/n146 , \_MxM/n145 , \_MxM/n144 , \_MxM/n143 , \_MxM/n142 ,
         \_MxM/n141 , \_MxM/n140 , \_MxM/n139 , \_MxM/n138 , \_MxM/n137 ,
         \_MxM/N19 , \_MxM/N18 , \_MxM/N17 , \_MxM/N16 , \_MxM/N15 ,
         \_MxM/N14 , \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 ,
         \_MxM/N8 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] ,
         \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] ,
         \_MxM/n[9] , \_MxM/n[10] , \_MxM/n[11] , \_MxM/n[12] , \_MxM/n[13] ,
         \_MxM/Y0[0] , \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] , \_MxM/Y0[4] ,
         \_MxM/Y0[5] , \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/add_39/carry[13] ,
         \_MxM/add_39/carry[12] , \_MxM/add_39/carry[11] ,
         \_MxM/add_39/carry[10] , \_MxM/add_39/carry[9] ,
         \_MxM/add_39/carry[8] , \_MxM/add_39/carry[7] ,
         \_MxM/add_39/carry[6] , \_MxM/add_39/carry[5] ,
         \_MxM/add_39/carry[4] , \_MxM/add_39/carry[3] ,
         \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n137 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n138 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n139 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n140 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n141 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n142 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n143 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n144 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n145 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n146 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n147 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n148 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n149 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n150 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n151 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n152 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[13]  ( .D(\_MxM/n153 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[13] ) );
  DFF \_MxM/n_reg[12]  ( .D(\_MxM/n154 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[12] ) );
  DFF \_MxM/n_reg[11]  ( .D(\_MxM/n155 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[11] ) );
  DFF \_MxM/n_reg[10]  ( .D(\_MxM/n156 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[10] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/n157 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/n158 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/n159 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n160 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n161 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n162 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n163 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n164 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n165 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n166 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N14 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N15 ) );
  HADDER \_MxM/add_39/U1_1_9  ( .IN0(\_MxM/n[9] ), .IN1(\_MxM/add_39/carry[9] ), .COUT(\_MxM/add_39/carry[10] ), .SUM(\_MxM/N16 ) );
  HADDER \_MxM/add_39/U1_1_10  ( .IN0(\_MxM/n[10] ), .IN1(
        \_MxM/add_39/carry[10] ), .COUT(\_MxM/add_39/carry[11] ), .SUM(
        \_MxM/N17 ) );
  HADDER \_MxM/add_39/U1_1_11  ( .IN0(\_MxM/n[11] ), .IN1(
        \_MxM/add_39/carry[11] ), .COUT(\_MxM/add_39/carry[12] ), .SUM(
        \_MxM/N18 ) );
  HADDER \_MxM/add_39/U1_1_12  ( .IN0(\_MxM/n[12] ), .IN1(
        \_MxM/add_39/carry[12] ), .COUT(\_MxM/add_39/carry[13] ), .SUM(
        \_MxM/N19 ) );
  MUX U1 ( .IN0(n326), .IN1(n342), .SEL(n328), .F(n307) );
  MUX U2 ( .IN0(g_input[3]), .IN1(n391), .SEL(g_input[7]), .F(n1) );
  IV U3 ( .A(n1), .Z(n236) );
  MUX U4 ( .IN0(n276), .IN1(n274), .SEL(n275), .F(n231) );
  NAND U5 ( .A(n149), .B(n183), .Z(n182) );
  MUX U6 ( .IN0(n259), .IN1(n2), .SEL(n258), .F(n214) );
  IV U7 ( .A(n257), .Z(n2) );
  MUX U8 ( .IN0(n3), .IN1(n159), .SEL(n160), .F(n127) );
  IV U9 ( .A(\_MxM/Y0[3] ), .Z(n3) );
  XOR U10 ( .A(n390), .B(g_input[3]), .Z(n391) );
  XNOR U11 ( .A(n378), .B(n379), .Z(n357) );
  MUX U12 ( .IN0(e_input[6]), .IN1(n416), .SEL(e_input[7]), .F(n125) );
  MUX U13 ( .IN0(e_input[3]), .IN1(n366), .SEL(e_input[7]), .F(n217) );
  MUX U14 ( .IN0(n220), .IN1(n4), .SEL(n221), .F(n172) );
  IV U15 ( .A(n222), .Z(n4) );
  XNOR U16 ( .A(n223), .B(n188), .Z(n180) );
  MUX U17 ( .IN0(n5), .IN1(n242), .SEL(n243), .F(n197) );
  IV U18 ( .A(\_MxM/Y0[1] ), .Z(n5) );
  XOR U19 ( .A(n95), .B(n105), .Z(n103) );
  MUX U20 ( .IN0(n6), .IN1(n396), .SEL(n397), .F(n392) );
  IV U21 ( .A(n398), .Z(n6) );
  MUX U22 ( .IN0(g_input[4]), .IN1(n343), .SEL(g_input[7]), .F(n7) );
  IV U23 ( .A(n7), .Z(n190) );
  MUX U24 ( .IN0(g_input[5]), .IN1(n325), .SEL(g_input[7]), .F(n153) );
  XOR U25 ( .A(n239), .B(n278), .Z(n240) );
  MUX U26 ( .IN0(g_input[6]), .IN1(n297), .SEL(g_input[7]), .F(n126) );
  MUX U27 ( .IN0(n260), .IN1(n8), .SEL(n261), .F(n220) );
  IV U28 ( .A(n262), .Z(n8) );
  XNOR U29 ( .A(n142), .B(n143), .Z(n166) );
  XOR U30 ( .A(n127), .B(n137), .Z(n135) );
  NOR U31 ( .A(g_input[0]), .B(n413), .Z(n401) );
  MUX U32 ( .IN0(n9), .IN1(n290), .SEL(n291), .F(n337) );
  IV U33 ( .A(n357), .Z(n9) );
  MUX U34 ( .IN0(n392), .IN1(n395), .SEL(n393), .F(n268) );
  MUX U35 ( .IN0(n307), .IN1(n323), .SEL(n309), .F(n301) );
  MUX U36 ( .IN0(n152), .IN1(n176), .SEL(n151), .F(n114) );
  NAND U37 ( .A(n214), .B(n255), .Z(n254) );
  XNOR U38 ( .A(n276), .B(n275), .Z(n262) );
  XNOR U39 ( .A(n181), .B(n180), .Z(n174) );
  XNOR U40 ( .A(n235), .B(n234), .Z(n222) );
  MUX U41 ( .IN0(\_MxM/Y0[6] ), .IN1(n77), .SEL(n72), .F(n65) );
  XOR U42 ( .A(n159), .B(n167), .Z(n165) );
  MUX U43 ( .IN0(g_input[2]), .IN1(n400), .SEL(g_input[7]), .F(n277) );
  XOR U44 ( .A(n367), .B(n348), .Z(n291) );
  XNOR U45 ( .A(n266), .B(n228), .Z(n234) );
  MUX U46 ( .IN0(n265), .IN1(n263), .SEL(n264), .F(n10) );
  IV U47 ( .A(n10), .Z(n219) );
  AND U48 ( .A(n120), .B(n86), .Z(n119) );
  MUX U49 ( .IN0(n11), .IN1(n174), .SEL(n173), .F(n143) );
  IV U50 ( .A(n172), .Z(n11) );
  MUX U51 ( .IN0(n12), .IN1(n197), .SEL(n198), .F(n159) );
  IV U52 ( .A(\_MxM/Y0[2] ), .Z(n12) );
  MUX U53 ( .IN0(\_MxM/Y0[7] ), .IN1(n65), .SEL(n66), .F(n13) );
  IV U54 ( .A(n13), .Z(n62) );
  XOR U55 ( .A(n243), .B(\_MxM/Y0[1] ), .Z(n31) );
  ANDN U56 ( .A(n14), .B(\_MxM/n[0] ), .Z(\_MxM/n166 ) );
  AND U57 ( .A(\_MxM/N8 ), .B(n14), .Z(\_MxM/n165 ) );
  AND U58 ( .A(\_MxM/N9 ), .B(n14), .Z(\_MxM/n164 ) );
  AND U59 ( .A(\_MxM/N10 ), .B(n14), .Z(\_MxM/n163 ) );
  AND U60 ( .A(\_MxM/N11 ), .B(n14), .Z(\_MxM/n162 ) );
  AND U61 ( .A(\_MxM/N12 ), .B(n14), .Z(\_MxM/n161 ) );
  AND U62 ( .A(\_MxM/N13 ), .B(n14), .Z(\_MxM/n160 ) );
  AND U63 ( .A(\_MxM/N14 ), .B(n14), .Z(\_MxM/n159 ) );
  AND U64 ( .A(\_MxM/N15 ), .B(n14), .Z(\_MxM/n158 ) );
  AND U65 ( .A(\_MxM/N16 ), .B(n14), .Z(\_MxM/n157 ) );
  AND U66 ( .A(\_MxM/N17 ), .B(n14), .Z(\_MxM/n156 ) );
  AND U67 ( .A(\_MxM/N18 ), .B(n14), .Z(\_MxM/n155 ) );
  AND U68 ( .A(\_MxM/N19 ), .B(n14), .Z(\_MxM/n154 ) );
  AND U69 ( .A(n14), .B(n15), .Z(\_MxM/n153 ) );
  XOR U70 ( .A(\_MxM/n[13] ), .B(\_MxM/add_39/carry[13] ), .Z(n15) );
  ANDN U71 ( .A(n16), .B(rst), .Z(n14) );
  NAND U72 ( .A(n17), .B(n18), .Z(n16) );
  AND U73 ( .A(n19), .B(n20), .Z(n18) );
  ANDN U74 ( .A(n21), .B(n22), .Z(n20) );
  NOR U75 ( .A(n23), .B(n24), .Z(n21) );
  AND U76 ( .A(n25), .B(\_MxM/n[13] ), .Z(n19) );
  AND U77 ( .A(\_MxM/n[10] ), .B(\_MxM/n[0] ), .Z(n25) );
  AND U78 ( .A(n26), .B(n27), .Z(n17) );
  AND U79 ( .A(\_MxM/n[3] ), .B(n28), .Z(n27) );
  AND U80 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n28) );
  AND U81 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n26) );
  NAND U82 ( .A(n29), .B(n30), .Z(\_MxM/n152 ) );
  OR U83 ( .A(n31), .B(n32), .Z(n30) );
  NANDN U84 ( .B(n33), .A(\_MxM/Y0[0] ), .Z(n29) );
  NAND U85 ( .A(n34), .B(n35), .Z(\_MxM/n151 ) );
  NANDN U86 ( .B(n32), .A(n36), .Z(n35) );
  NANDN U87 ( .B(n37), .A(rst), .Z(n34) );
  NAND U88 ( .A(n38), .B(n39), .Z(\_MxM/n150 ) );
  NANDN U89 ( .B(n32), .A(n40), .Z(n39) );
  NANDN U90 ( .B(n33), .A(\_MxM/Y0[2] ), .Z(n38) );
  NAND U91 ( .A(n41), .B(n42), .Z(\_MxM/n149 ) );
  NANDN U92 ( .B(n32), .A(n43), .Z(n42) );
  NANDN U93 ( .B(n33), .A(\_MxM/Y0[3] ), .Z(n41) );
  NAND U94 ( .A(n44), .B(n45), .Z(\_MxM/n148 ) );
  NANDN U95 ( .B(n32), .A(n46), .Z(n45) );
  NANDN U96 ( .B(n33), .A(\_MxM/Y0[4] ), .Z(n44) );
  NAND U97 ( .A(n47), .B(n48), .Z(\_MxM/n147 ) );
  NANDN U98 ( .B(n32), .A(n49), .Z(n48) );
  NANDN U99 ( .B(n33), .A(\_MxM/Y0[5] ), .Z(n47) );
  NAND U100 ( .A(n50), .B(n51), .Z(\_MxM/n146 ) );
  OR U101 ( .A(n52), .B(n32), .Z(n51) );
  NANDN U102 ( .B(n33), .A(\_MxM/Y0[6] ), .Z(n50) );
  NAND U103 ( .A(n53), .B(n54), .Z(\_MxM/n145 ) );
  OR U104 ( .A(n32), .B(n55), .Z(n54) );
  NANDN U105 ( .B(n56), .A(n33), .Z(n32) );
  NANDN U106 ( .B(n33), .A(\_MxM/Y0[7] ), .Z(n53) );
  NAND U107 ( .A(n57), .B(n58), .Z(\_MxM/n144 ) );
  NANDN U108 ( .B(n33), .A(o[7]), .Z(n58) );
  AND U109 ( .A(n59), .B(n60), .Z(n57) );
  NANDN U110 ( .B(n56), .A(o[7]), .Z(n60) );
  OR U111 ( .A(n55), .B(n61), .Z(n59) );
  XOR U112 ( .A(n62), .B(n63), .Z(n55) );
  XNOR U113 ( .A(\_MxM/Y0[7] ), .B(n64), .Z(n63) );
  NAND U114 ( .A(n67), .B(n68), .Z(\_MxM/n143 ) );
  NANDN U115 ( .B(n33), .A(o[6]), .Z(n68) );
  AND U116 ( .A(n69), .B(n70), .Z(n67) );
  NANDN U117 ( .B(n56), .A(o[6]), .Z(n70) );
  OR U118 ( .A(n52), .B(n61), .Z(n69) );
  XOR U119 ( .A(n66), .B(\_MxM/Y0[7] ), .Z(n52) );
  XOR U120 ( .A(n65), .B(n64), .Z(n66) );
  NAND U121 ( .A(n73), .B(n74), .Z(\_MxM/n142 ) );
  NANDN U122 ( .B(n33), .A(o[5]), .Z(n74) );
  AND U123 ( .A(n75), .B(n76), .Z(n73) );
  NANDN U124 ( .B(n56), .A(o[5]), .Z(n76) );
  NANDN U125 ( .B(n61), .A(n49), .Z(n75) );
  XNOR U126 ( .A(n72), .B(\_MxM/Y0[6] ), .Z(n49) );
  XOR U127 ( .A(n77), .B(n78), .Z(n72) );
  ANDN U128 ( .A(n64), .B(n79), .Z(n78) );
  NANDN U129 ( .B(n80), .A(n81), .Z(n64) );
  ANDN U130 ( .A(n82), .B(n79), .Z(n80) );
  NAND U131 ( .A(n83), .B(n84), .Z(n79) );
  OR U132 ( .A(n85), .B(n86), .Z(n84) );
  AND U133 ( .A(n87), .B(n88), .Z(n83) );
  OR U134 ( .A(n89), .B(n90), .Z(n88) );
  OR U135 ( .A(n91), .B(n92), .Z(n87) );
  NOR U136 ( .A(n93), .B(n94), .Z(n82) );
  IV U137 ( .A(n71), .Z(n77) );
  XOR U138 ( .A(n95), .B(n96), .Z(n71) );
  ANDN U139 ( .A(n97), .B(n98), .Z(n96) );
  XNOR U140 ( .A(\_MxM/Y0[5] ), .B(n95), .Z(n97) );
  NAND U141 ( .A(n99), .B(n100), .Z(\_MxM/n141 ) );
  NANDN U142 ( .B(n33), .A(o[4]), .Z(n100) );
  AND U143 ( .A(n101), .B(n102), .Z(n99) );
  NANDN U144 ( .B(n56), .A(o[4]), .Z(n102) );
  NANDN U145 ( .B(n61), .A(n46), .Z(n101) );
  XNOR U146 ( .A(n98), .B(\_MxM/Y0[5] ), .Z(n46) );
  XNOR U147 ( .A(n103), .B(n104), .Z(n98) );
  AND U148 ( .A(n81), .B(n106), .Z(n105) );
  XOR U149 ( .A(n93), .B(n107), .Z(n106) );
  XOR U150 ( .A(n107), .B(n94), .Z(n93) );
  OR U151 ( .A(n108), .B(n109), .Z(n94) );
  IV U152 ( .A(n104), .Z(n107) );
  XNOR U153 ( .A(n92), .B(n91), .Z(n104) );
  OR U154 ( .A(n110), .B(n111), .Z(n91) );
  AND U155 ( .A(n112), .B(n113), .Z(n92) );
  XNOR U156 ( .A(n114), .B(n115), .Z(n113) );
  ANDN U157 ( .A(n116), .B(n117), .Z(n115) );
  XOR U158 ( .A(n114), .B(n118), .Z(n116) );
  XNOR U159 ( .A(n85), .B(n119), .Z(n112) );
  NAND U160 ( .A(n121), .B(n122), .Z(n86) );
  NANDN U161 ( .B(n123), .A(n124), .Z(n121) );
  NANDN U162 ( .B(n89), .A(n125), .Z(n120) );
  NANDN U163 ( .B(n90), .A(n126), .Z(n85) );
  XOR U164 ( .A(n127), .B(n128), .Z(n95) );
  ANDN U165 ( .A(n129), .B(n130), .Z(n128) );
  XNOR U166 ( .A(\_MxM/Y0[4] ), .B(n127), .Z(n129) );
  NAND U167 ( .A(n131), .B(n132), .Z(\_MxM/n140 ) );
  NANDN U168 ( .B(n33), .A(o[3]), .Z(n132) );
  AND U169 ( .A(n133), .B(n134), .Z(n131) );
  NANDN U170 ( .B(n56), .A(o[3]), .Z(n134) );
  NANDN U171 ( .B(n61), .A(n43), .Z(n133) );
  XNOR U172 ( .A(n130), .B(\_MxM/Y0[4] ), .Z(n43) );
  XNOR U173 ( .A(n135), .B(n136), .Z(n130) );
  AND U174 ( .A(n81), .B(n138), .Z(n137) );
  XOR U175 ( .A(n108), .B(n139), .Z(n138) );
  XOR U176 ( .A(n139), .B(n109), .Z(n108) );
  OR U177 ( .A(n140), .B(n141), .Z(n109) );
  IV U178 ( .A(n136), .Z(n139) );
  XNOR U179 ( .A(n111), .B(n110), .Z(n136) );
  OR U180 ( .A(n142), .B(n143), .Z(n110) );
  XOR U181 ( .A(n118), .B(n117), .Z(n111) );
  XOR U182 ( .A(n114), .B(n144), .Z(n117) );
  AND U183 ( .A(n145), .B(n146), .Z(n144) );
  NANDN U184 ( .B(n89), .A(n147), .Z(n146) );
  OR U185 ( .A(n148), .B(n149), .Z(n145) );
  XOR U186 ( .A(n123), .B(n124), .Z(n118) );
  NANDN U187 ( .B(n90), .A(n153), .Z(n124) );
  XNOR U188 ( .A(n122), .B(n154), .Z(n123) );
  AND U189 ( .A(n126), .B(n125), .Z(n154) );
  ANDN U190 ( .A(n155), .B(n156), .Z(n122) );
  NANDN U191 ( .B(n157), .A(n158), .Z(n155) );
  NAND U192 ( .A(n161), .B(n162), .Z(\_MxM/n139 ) );
  NANDN U193 ( .B(n33), .A(o[2]), .Z(n162) );
  AND U194 ( .A(n163), .B(n164), .Z(n161) );
  NANDN U195 ( .B(n56), .A(o[2]), .Z(n164) );
  NANDN U196 ( .B(n61), .A(n40), .Z(n163) );
  XNOR U197 ( .A(n160), .B(\_MxM/Y0[3] ), .Z(n40) );
  XNOR U198 ( .A(n165), .B(n166), .Z(n160) );
  AND U199 ( .A(n81), .B(n168), .Z(n167) );
  XOR U200 ( .A(n140), .B(n169), .Z(n168) );
  XOR U201 ( .A(n169), .B(n141), .Z(n140) );
  OR U202 ( .A(n170), .B(n171), .Z(n141) );
  IV U203 ( .A(n166), .Z(n169) );
  XOR U204 ( .A(n152), .B(n151), .Z(n142) );
  XNOR U205 ( .A(n175), .B(n176), .Z(n151) );
  IV U206 ( .A(n150), .Z(n176) );
  XOR U207 ( .A(n177), .B(n178), .Z(n150) );
  ANDN U208 ( .A(n179), .B(n180), .Z(n178) );
  XOR U209 ( .A(n177), .B(n181), .Z(n179) );
  XNOR U210 ( .A(n182), .B(n148), .Z(n175) );
  NAND U211 ( .A(n147), .B(n126), .Z(n148) );
  NANDN U212 ( .B(n89), .A(n184), .Z(n183) );
  XNOR U213 ( .A(n185), .B(n186), .Z(n149) );
  ANDN U214 ( .A(n187), .B(n188), .Z(n186) );
  XNOR U215 ( .A(n189), .B(n185), .Z(n187) );
  XOR U216 ( .A(n157), .B(n158), .Z(n152) );
  OR U217 ( .A(n190), .B(n90), .Z(n158) );
  XNOR U218 ( .A(n191), .B(n192), .Z(n157) );
  AND U219 ( .A(n153), .B(n125), .Z(n192) );
  IV U220 ( .A(n156), .Z(n191) );
  NAND U221 ( .A(n193), .B(n194), .Z(n156) );
  NANDN U222 ( .B(n195), .A(n196), .Z(n193) );
  NAND U223 ( .A(n199), .B(n200), .Z(\_MxM/n138 ) );
  NANDN U224 ( .B(n33), .A(o[1]), .Z(n200) );
  AND U225 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U226 ( .B(n56), .A(o[1]), .Z(n202) );
  NANDN U227 ( .B(n61), .A(n36), .Z(n201) );
  XNOR U228 ( .A(n198), .B(\_MxM/Y0[2] ), .Z(n36) );
  XNOR U229 ( .A(n203), .B(n204), .Z(n198) );
  XOR U230 ( .A(n197), .B(n205), .Z(n203) );
  AND U231 ( .A(n81), .B(n206), .Z(n205) );
  XOR U232 ( .A(n170), .B(n207), .Z(n206) );
  XOR U233 ( .A(n207), .B(n171), .Z(n170) );
  NANDN U234 ( .B(n208), .A(n209), .Z(n171) );
  IV U235 ( .A(n204), .Z(n207) );
  XOR U236 ( .A(n174), .B(n173), .Z(n204) );
  XNOR U237 ( .A(n172), .B(n210), .Z(n173) );
  AND U238 ( .A(n211), .B(n212), .Z(n210) );
  OR U239 ( .A(n213), .B(n214), .Z(n212) );
  AND U240 ( .A(n215), .B(n216), .Z(n211) );
  NANDN U241 ( .B(n89), .A(n217), .Z(n216) );
  NAND U242 ( .A(n218), .B(n219), .Z(n215) );
  XNOR U243 ( .A(n185), .B(n224), .Z(n188) );
  AND U244 ( .A(n126), .B(n184), .Z(n224) );
  XOR U245 ( .A(n225), .B(n226), .Z(n185) );
  ANDN U246 ( .A(n227), .B(n228), .Z(n226) );
  XNOR U247 ( .A(n229), .B(n225), .Z(n227) );
  XOR U248 ( .A(n230), .B(n189), .Z(n223) );
  NAND U249 ( .A(n147), .B(n153), .Z(n189) );
  IV U250 ( .A(n177), .Z(n230) );
  XOR U251 ( .A(n231), .B(n232), .Z(n177) );
  ANDN U252 ( .A(n233), .B(n234), .Z(n232) );
  XOR U253 ( .A(n231), .B(n235), .Z(n233) );
  XNOR U254 ( .A(n195), .B(n196), .Z(n181) );
  OR U255 ( .A(n236), .B(n90), .Z(n196) );
  XNOR U256 ( .A(n194), .B(n237), .Z(n195) );
  ANDN U257 ( .A(n125), .B(n190), .Z(n237) );
  ANDN U258 ( .A(n238), .B(n239), .Z(n194) );
  NANDN U259 ( .B(n240), .A(n241), .Z(n238) );
  NAND U260 ( .A(n244), .B(n245), .Z(\_MxM/n137 ) );
  NANDN U261 ( .B(n33), .A(o[0]), .Z(n245) );
  AND U262 ( .A(n246), .B(n247), .Z(n244) );
  NANDN U263 ( .B(n56), .A(o[0]), .Z(n247) );
  IV U264 ( .A(n248), .Z(n56) );
  OR U265 ( .A(n61), .B(n31), .Z(n246) );
  IV U266 ( .A(\_MxM/Y0[1] ), .Z(n37) );
  XOR U267 ( .A(n249), .B(n250), .Z(n243) );
  XNOR U268 ( .A(n251), .B(n242), .Z(n249) );
  NAND U269 ( .A(\_MxM/Y0[0] ), .B(n208), .Z(n242) );
  NAND U270 ( .A(n252), .B(n81), .Z(n251) );
  XOR U271 ( .A(e_input[7]), .B(g_input[7]), .Z(n81) );
  XNOR U272 ( .A(n209), .B(n250), .Z(n252) );
  XNOR U273 ( .A(n208), .B(n250), .Z(n209) );
  XNOR U274 ( .A(n222), .B(n221), .Z(n250) );
  XNOR U275 ( .A(n253), .B(n218), .Z(n221) );
  XNOR U276 ( .A(n254), .B(n213), .Z(n218) );
  NAND U277 ( .A(n126), .B(n217), .Z(n213) );
  NANDN U278 ( .B(n89), .A(n256), .Z(n255) );
  XNOR U279 ( .A(n219), .B(n220), .Z(n253) );
  XNOR U280 ( .A(n225), .B(n267), .Z(n228) );
  AND U281 ( .A(n153), .B(n184), .Z(n267) );
  XOR U282 ( .A(n268), .B(n269), .Z(n225) );
  ANDN U283 ( .A(n270), .B(n271), .Z(n269) );
  XNOR U284 ( .A(n272), .B(n268), .Z(n270) );
  XOR U285 ( .A(n273), .B(n229), .Z(n266) );
  NANDN U286 ( .B(n190), .A(n147), .Z(n229) );
  IV U287 ( .A(n231), .Z(n273) );
  XNOR U288 ( .A(n240), .B(n241), .Z(n235) );
  NANDN U289 ( .B(n90), .A(n277), .Z(n241) );
  ANDN U290 ( .A(n125), .B(n236), .Z(n278) );
  NAND U291 ( .A(n279), .B(n280), .Z(n239) );
  NANDN U292 ( .B(n281), .A(n282), .Z(n279) );
  XNOR U293 ( .A(n262), .B(n261), .Z(n208) );
  XNOR U294 ( .A(n283), .B(n265), .Z(n261) );
  XNOR U295 ( .A(n258), .B(n259), .Z(n265) );
  NAND U296 ( .A(n153), .B(n217), .Z(n259) );
  XNOR U297 ( .A(n257), .B(n284), .Z(n258) );
  AND U298 ( .A(n256), .B(n126), .Z(n284) );
  XOR U299 ( .A(n285), .B(n286), .Z(n257) );
  AND U300 ( .A(n287), .B(n288), .Z(n286) );
  XNOR U301 ( .A(n289), .B(n285), .Z(n288) );
  XNOR U302 ( .A(n264), .B(n260), .Z(n283) );
  XOR U303 ( .A(n290), .B(n291), .Z(n260) );
  XOR U304 ( .A(n292), .B(n293), .Z(n264) );
  AND U305 ( .A(n294), .B(n295), .Z(n293) );
  NANDN U306 ( .B(n89), .A(n296), .Z(n295) );
  NANDN U307 ( .B(n297), .A(n298), .Z(n89) );
  AND U308 ( .A(n299), .B(g_input[7]), .Z(n298) );
  NANDN U309 ( .B(n300), .A(n301), .Z(n294) );
  IV U310 ( .A(n263), .Z(n292) );
  XNOR U311 ( .A(n302), .B(n303), .Z(n263) );
  AND U312 ( .A(n304), .B(n305), .Z(n303) );
  XOR U313 ( .A(n301), .B(n306), .Z(n305) );
  XNOR U314 ( .A(n300), .B(n302), .Z(n306) );
  NAND U315 ( .A(n126), .B(n296), .Z(n300) );
  XNOR U316 ( .A(n310), .B(n307), .Z(n309) );
  XOR U317 ( .A(n287), .B(n311), .Z(n304) );
  XNOR U318 ( .A(n289), .B(n302), .Z(n311) );
  NANDN U319 ( .B(n190), .A(n217), .Z(n289) );
  XOR U320 ( .A(n285), .B(n312), .Z(n287) );
  AND U321 ( .A(n256), .B(n153), .Z(n312) );
  XOR U322 ( .A(n313), .B(n314), .Z(n285) );
  AND U323 ( .A(n315), .B(n316), .Z(n314) );
  XNOR U324 ( .A(n317), .B(n313), .Z(n316) );
  XOR U325 ( .A(n318), .B(n319), .Z(n302) );
  AND U326 ( .A(n320), .B(n321), .Z(n319) );
  XOR U327 ( .A(n308), .B(n322), .Z(n321) );
  XNOR U328 ( .A(n310), .B(n318), .Z(n322) );
  NAND U329 ( .A(n153), .B(n296), .Z(n310) );
  XOR U330 ( .A(n307), .B(n323), .Z(n308) );
  AND U331 ( .A(n126), .B(e_input[0]), .Z(n323) );
  XNOR U332 ( .A(n299), .B(g_input[6]), .Z(n297) );
  NOR U333 ( .A(n324), .B(n325), .Z(n299) );
  XNOR U334 ( .A(n329), .B(n326), .Z(n328) );
  XOR U335 ( .A(n315), .B(n330), .Z(n320) );
  XNOR U336 ( .A(n317), .B(n318), .Z(n330) );
  NANDN U337 ( .B(n236), .A(n217), .Z(n317) );
  XOR U338 ( .A(n313), .B(n331), .Z(n315) );
  ANDN U339 ( .A(n256), .B(n190), .Z(n331) );
  XOR U340 ( .A(n332), .B(n333), .Z(n313) );
  AND U341 ( .A(n334), .B(n335), .Z(n333) );
  XNOR U342 ( .A(n336), .B(n332), .Z(n335) );
  XOR U343 ( .A(n337), .B(n338), .Z(n318) );
  AND U344 ( .A(n339), .B(n340), .Z(n338) );
  XOR U345 ( .A(n327), .B(n341), .Z(n340) );
  XNOR U346 ( .A(n329), .B(n337), .Z(n341) );
  NANDN U347 ( .B(n190), .A(n296), .Z(n329) );
  XOR U348 ( .A(n326), .B(n342), .Z(n327) );
  AND U349 ( .A(n153), .B(e_input[0]), .Z(n342) );
  XOR U350 ( .A(n324), .B(g_input[5]), .Z(n325) );
  NANDN U351 ( .B(n343), .A(n344), .Z(n324) );
  XOR U352 ( .A(n345), .B(n346), .Z(n326) );
  ANDN U353 ( .A(n347), .B(n348), .Z(n346) );
  XNOR U354 ( .A(n349), .B(n345), .Z(n347) );
  XOR U355 ( .A(n334), .B(n350), .Z(n339) );
  XNOR U356 ( .A(n336), .B(n337), .Z(n350) );
  NAND U357 ( .A(n217), .B(n277), .Z(n336) );
  XOR U358 ( .A(n332), .B(n351), .Z(n334) );
  ANDN U359 ( .A(n256), .B(n236), .Z(n351) );
  XOR U360 ( .A(n352), .B(n353), .Z(n332) );
  ANDN U361 ( .A(n354), .B(n355), .Z(n353) );
  XNOR U362 ( .A(n356), .B(n352), .Z(n354) );
  XNOR U363 ( .A(n358), .B(n356), .Z(n290) );
  NAND U364 ( .A(n217), .B(n359), .Z(n356) );
  IV U365 ( .A(n355), .Z(n358) );
  XNOR U366 ( .A(n352), .B(n360), .Z(n355) );
  AND U367 ( .A(n277), .B(n256), .Z(n360) );
  AND U368 ( .A(n361), .B(g_input[0]), .Z(n352) );
  NANDN U369 ( .B(n217), .A(n362), .Z(n361) );
  NAND U370 ( .A(n359), .B(n256), .Z(n362) );
  XNOR U371 ( .A(n363), .B(e_input[2]), .Z(n256) );
  NAND U372 ( .A(n364), .B(e_input[7]), .Z(n363) );
  XOR U373 ( .A(n365), .B(e_input[2]), .Z(n364) );
  XNOR U374 ( .A(n345), .B(n368), .Z(n348) );
  ANDN U375 ( .A(e_input[0]), .B(n190), .Z(n368) );
  XOR U376 ( .A(n369), .B(n370), .Z(n345) );
  AND U377 ( .A(n371), .B(n372), .Z(n370) );
  XOR U378 ( .A(n373), .B(n369), .Z(n372) );
  ANDN U379 ( .A(e_input[0]), .B(n236), .Z(n373) );
  XOR U380 ( .A(n374), .B(n369), .Z(n371) );
  AND U381 ( .A(n296), .B(n277), .Z(n374) );
  XOR U382 ( .A(n375), .B(n376), .Z(n369) );
  ANDN U383 ( .A(n377), .B(n378), .Z(n376) );
  XNOR U384 ( .A(n379), .B(n375), .Z(n377) );
  XOR U385 ( .A(n380), .B(n349), .Z(n367) );
  NANDN U386 ( .B(n236), .A(n296), .Z(n349) );
  IV U387 ( .A(n357), .Z(n380) );
  NAND U388 ( .A(n296), .B(n359), .Z(n379) );
  XNOR U389 ( .A(n375), .B(n381), .Z(n378) );
  AND U390 ( .A(n277), .B(e_input[0]), .Z(n381) );
  AND U391 ( .A(n382), .B(g_input[0]), .Z(n375) );
  NANDN U392 ( .B(n296), .A(n383), .Z(n382) );
  NAND U393 ( .A(n359), .B(e_input[0]), .Z(n383) );
  XNOR U394 ( .A(n384), .B(e_input[1]), .Z(n296) );
  NAND U395 ( .A(n385), .B(e_input[7]), .Z(n384) );
  XNOR U396 ( .A(e_input[1]), .B(n386), .Z(n385) );
  XOR U397 ( .A(n387), .B(n388), .Z(n275) );
  IV U398 ( .A(n271), .Z(n388) );
  XNOR U399 ( .A(n268), .B(n389), .Z(n271) );
  ANDN U400 ( .A(n184), .B(n190), .Z(n389) );
  XNOR U401 ( .A(n344), .B(g_input[4]), .Z(n343) );
  NOR U402 ( .A(n390), .B(n391), .Z(n344) );
  XOR U403 ( .A(n394), .B(n392), .Z(n393) );
  ANDN U404 ( .A(n184), .B(n236), .Z(n394) );
  AND U405 ( .A(n277), .B(n147), .Z(n395) );
  XOR U406 ( .A(n399), .B(n272), .Z(n387) );
  NANDN U407 ( .B(n236), .A(n147), .Z(n272) );
  NANDN U408 ( .B(n400), .A(n401), .Z(n390) );
  IV U409 ( .A(n274), .Z(n399) );
  XOR U410 ( .A(n402), .B(n398), .Z(n274) );
  NAND U411 ( .A(n147), .B(n359), .Z(n398) );
  IV U412 ( .A(n397), .Z(n402) );
  XNOR U413 ( .A(n396), .B(n403), .Z(n397) );
  AND U414 ( .A(n277), .B(n184), .Z(n403) );
  AND U415 ( .A(n404), .B(g_input[0]), .Z(n396) );
  NANDN U416 ( .B(n147), .A(n405), .Z(n404) );
  NAND U417 ( .A(n359), .B(n184), .Z(n405) );
  XNOR U418 ( .A(n406), .B(e_input[4]), .Z(n184) );
  NAND U419 ( .A(n407), .B(e_input[7]), .Z(n406) );
  XOR U420 ( .A(n408), .B(e_input[4]), .Z(n407) );
  XNOR U421 ( .A(n409), .B(e_input[5]), .Z(n147) );
  NAND U422 ( .A(n410), .B(e_input[7]), .Z(n409) );
  XOR U423 ( .A(n411), .B(e_input[5]), .Z(n410) );
  XNOR U424 ( .A(n281), .B(n282), .Z(n276) );
  NANDN U425 ( .B(n90), .A(n359), .Z(n282) );
  XNOR U426 ( .A(n280), .B(n412), .Z(n281) );
  AND U427 ( .A(n277), .B(n125), .Z(n412) );
  XNOR U428 ( .A(n401), .B(g_input[2]), .Z(n400) );
  AND U429 ( .A(n414), .B(g_input[0]), .Z(n280) );
  NAND U430 ( .A(n415), .B(n90), .Z(n414) );
  NANDN U431 ( .B(n416), .A(n417), .Z(n90) );
  ANDN U432 ( .A(e_input[7]), .B(n418), .Z(n417) );
  NAND U433 ( .A(n359), .B(n125), .Z(n415) );
  XOR U434 ( .A(n418), .B(e_input[6]), .Z(n416) );
  OR U435 ( .A(n411), .B(n419), .Z(n418) );
  XOR U436 ( .A(n419), .B(e_input[5]), .Z(n411) );
  OR U437 ( .A(n408), .B(n420), .Z(n419) );
  XOR U438 ( .A(n420), .B(e_input[4]), .Z(n408) );
  OR U439 ( .A(n366), .B(n421), .Z(n420) );
  XOR U440 ( .A(n421), .B(e_input[3]), .Z(n366) );
  OR U441 ( .A(n365), .B(n422), .Z(n421) );
  XOR U442 ( .A(n422), .B(e_input[2]), .Z(n365) );
  NANDN U443 ( .B(e_input[0]), .A(n386), .Z(n422) );
  XNOR U444 ( .A(e_input[0]), .B(e_input[1]), .Z(n386) );
  XNOR U445 ( .A(n423), .B(g_input[1]), .Z(n359) );
  NAND U446 ( .A(n424), .B(g_input[7]), .Z(n423) );
  XOR U447 ( .A(g_input[1]), .B(n413), .Z(n424) );
  XOR U448 ( .A(g_input[0]), .B(g_input[1]), .Z(n413) );
  NANDN U449 ( .B(n248), .A(n33), .Z(n61) );
  IV U450 ( .A(rst), .Z(n33) );
  NAND U451 ( .A(n425), .B(n426), .Z(n248) );
  AND U452 ( .A(n427), .B(n428), .Z(n426) );
  ANDN U453 ( .A(n429), .B(\_MxM/n[3] ), .Z(n428) );
  NOR U454 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n429) );
  ANDN U455 ( .A(n430), .B(\_MxM/n[13] ), .Z(n427) );
  NOR U456 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n430) );
  AND U457 ( .A(n431), .B(n432), .Z(n425) );
  ANDN U458 ( .A(n433), .B(n24), .Z(n432) );
  OR U459 ( .A(\_MxM/n[6] ), .B(\_MxM/n[7] ), .Z(n24) );
  NOR U460 ( .A(\_MxM/n[0] ), .B(\_MxM/n[10] ), .Z(n433) );
  NOR U461 ( .A(n22), .B(n23), .Z(n431) );
  OR U462 ( .A(\_MxM/n[4] ), .B(\_MxM/n[5] ), .Z(n23) );
  OR U463 ( .A(\_MxM/n[12] ), .B(\_MxM/n[11] ), .Z(n22) );
endmodule

