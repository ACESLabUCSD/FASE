
module MxM_W8_N1000 ( clk, rst, A, X, Y );
  input [7:0] A;
  input [7:0] X;
  output [7:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         \add_25/carry[9] , \add_25/carry[8] , \add_25/carry[7] ,
         \add_25/carry[6] , \add_25/carry[5] , \add_25/carry[4] ,
         \add_25/carry[3] , \add_25/carry[2] , n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575;
  wire   [7:0] Y0;
  wire   [9:0] n;

  DFF \n_reg[0]  ( .D(n148), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n147), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n146), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n145), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n144), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n143), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n142), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \n_reg[7]  ( .D(n141), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[7]) );
  DFF \n_reg[8]  ( .D(n140), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[8]) );
  DFF \n_reg[9]  ( .D(n139), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[9]) );
  DFF \Y0_reg[0]  ( .D(n138), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n137), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n136), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n135), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n134), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n133), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n132), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n131), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y_reg[7]  ( .D(n130), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n129), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n128), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n127), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n126), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n125), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n124), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n123), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  HADDER \add_25/U1_1_6  ( .IN0(n[6]), .IN1(\add_25/carry[6] ), .COUT(
        \add_25/carry[7] ), .SUM(N13) );
  HADDER \add_25/U1_1_7  ( .IN0(n[7]), .IN1(\add_25/carry[7] ), .COUT(
        \add_25/carry[8] ), .SUM(N14) );
  HADDER \add_25/U1_1_8  ( .IN0(n[8]), .IN1(\add_25/carry[8] ), .COUT(
        \add_25/carry[9] ), .SUM(N15) );
  MUX U151 ( .IN0(n470), .IN1(n486), .SEL(n472), .F(n451) );
  MUX U152 ( .IN0(A[3]), .IN1(n535), .SEL(A[7]), .F(n149) );
  IV U153 ( .A(n149), .Z(n380) );
  MUX U154 ( .IN0(n420), .IN1(n418), .SEL(n419), .F(n375) );
  NAND U155 ( .A(n293), .B(n327), .Z(n326) );
  MUX U156 ( .IN0(n403), .IN1(n150), .SEL(n402), .F(n358) );
  IV U157 ( .A(n401), .Z(n150) );
  MUX U158 ( .IN0(n151), .IN1(n303), .SEL(n304), .F(n271) );
  IV U159 ( .A(Y0[3]), .Z(n151) );
  XOR U160 ( .A(n534), .B(A[3]), .Z(n535) );
  XNOR U161 ( .A(n522), .B(n523), .Z(n501) );
  MUX U162 ( .IN0(X[6]), .IN1(n560), .SEL(X[7]), .F(n269) );
  MUX U163 ( .IN0(X[3]), .IN1(n510), .SEL(X[7]), .F(n361) );
  MUX U164 ( .IN0(n364), .IN1(n152), .SEL(n365), .F(n316) );
  IV U165 ( .A(n366), .Z(n152) );
  XNOR U166 ( .A(n367), .B(n332), .Z(n324) );
  MUX U167 ( .IN0(n153), .IN1(n386), .SEL(n387), .F(n341) );
  IV U168 ( .A(Y0[1]), .Z(n153) );
  XOR U169 ( .A(n239), .B(n249), .Z(n247) );
  MUX U170 ( .IN0(n154), .IN1(n540), .SEL(n541), .F(n536) );
  IV U171 ( .A(n542), .Z(n154) );
  MUX U172 ( .IN0(A[4]), .IN1(n487), .SEL(A[7]), .F(n155) );
  IV U173 ( .A(n155), .Z(n334) );
  MUX U174 ( .IN0(A[5]), .IN1(n469), .SEL(A[7]), .F(n297) );
  XOR U175 ( .A(n383), .B(n422), .Z(n384) );
  MUX U176 ( .IN0(A[6]), .IN1(n441), .SEL(A[7]), .F(n270) );
  MUX U177 ( .IN0(n404), .IN1(n156), .SEL(n405), .F(n364) );
  IV U178 ( .A(n406), .Z(n156) );
  XNOR U179 ( .A(n286), .B(n287), .Z(n310) );
  XOR U180 ( .A(n271), .B(n281), .Z(n279) );
  NOR U181 ( .A(A[0]), .B(n557), .Z(n545) );
  MUX U182 ( .IN0(n157), .IN1(n434), .SEL(n435), .F(n481) );
  IV U183 ( .A(n501), .Z(n157) );
  MUX U184 ( .IN0(n536), .IN1(n539), .SEL(n537), .F(n412) );
  MUX U185 ( .IN0(n451), .IN1(n467), .SEL(n453), .F(n445) );
  MUX U186 ( .IN0(n296), .IN1(n320), .SEL(n295), .F(n258) );
  NAND U187 ( .A(n358), .B(n399), .Z(n398) );
  XNOR U188 ( .A(n420), .B(n419), .Z(n406) );
  XNOR U189 ( .A(n325), .B(n324), .Z(n318) );
  XNOR U190 ( .A(n379), .B(n378), .Z(n366) );
  MUX U191 ( .IN0(Y0[6]), .IN1(n221), .SEL(n216), .F(n209) );
  XOR U192 ( .A(n303), .B(n311), .Z(n309) );
  MUX U193 ( .IN0(A[2]), .IN1(n544), .SEL(A[7]), .F(n421) );
  XOR U194 ( .A(n511), .B(n492), .Z(n435) );
  XNOR U195 ( .A(n410), .B(n372), .Z(n378) );
  MUX U196 ( .IN0(n409), .IN1(n407), .SEL(n408), .F(n158) );
  IV U197 ( .A(n158), .Z(n363) );
  AND U198 ( .A(n264), .B(n230), .Z(n263) );
  MUX U199 ( .IN0(n159), .IN1(n318), .SEL(n317), .F(n287) );
  IV U200 ( .A(n316), .Z(n159) );
  MUX U201 ( .IN0(n160), .IN1(n341), .SEL(n342), .F(n303) );
  IV U202 ( .A(Y0[2]), .Z(n160) );
  MUX U203 ( .IN0(Y0[7]), .IN1(n209), .SEL(n210), .F(n161) );
  IV U204 ( .A(n161), .Z(n206) );
  XOR U205 ( .A(n387), .B(Y0[1]), .Z(n175) );
  ANDN U206 ( .A(n162), .B(n[0]), .Z(n148) );
  AND U207 ( .A(N8), .B(n162), .Z(n147) );
  AND U208 ( .A(N9), .B(n162), .Z(n146) );
  AND U209 ( .A(N10), .B(n162), .Z(n145) );
  AND U210 ( .A(N11), .B(n162), .Z(n144) );
  AND U211 ( .A(N12), .B(n162), .Z(n143) );
  AND U212 ( .A(N13), .B(n162), .Z(n142) );
  AND U213 ( .A(N14), .B(n162), .Z(n141) );
  AND U214 ( .A(N15), .B(n162), .Z(n140) );
  AND U215 ( .A(n162), .B(n163), .Z(n139) );
  XOR U216 ( .A(n[9]), .B(\add_25/carry[9] ), .Z(n163) );
  ANDN U217 ( .A(n164), .B(rst), .Z(n162) );
  NAND U218 ( .A(n165), .B(n166), .Z(n164) );
  AND U219 ( .A(n167), .B(n168), .Z(n166) );
  AND U220 ( .A(n[1]), .B(n169), .Z(n168) );
  ANDN U221 ( .A(n[0]), .B(n170), .Z(n169) );
  AND U222 ( .A(n[5]), .B(n[2]), .Z(n167) );
  AND U223 ( .A(n171), .B(n172), .Z(n165) );
  AND U224 ( .A(n[7]), .B(n[6]), .Z(n172) );
  AND U225 ( .A(n[8]), .B(n[9]), .Z(n171) );
  NAND U226 ( .A(n173), .B(n174), .Z(n138) );
  OR U227 ( .A(n175), .B(n176), .Z(n174) );
  NANDN U228 ( .B(n177), .A(Y0[0]), .Z(n173) );
  NAND U229 ( .A(n178), .B(n179), .Z(n137) );
  NANDN U230 ( .B(n176), .A(n180), .Z(n179) );
  NANDN U231 ( .B(n181), .A(rst), .Z(n178) );
  NAND U232 ( .A(n182), .B(n183), .Z(n136) );
  NANDN U233 ( .B(n176), .A(n184), .Z(n183) );
  NANDN U234 ( .B(n177), .A(Y0[2]), .Z(n182) );
  NAND U235 ( .A(n185), .B(n186), .Z(n135) );
  NANDN U236 ( .B(n176), .A(n187), .Z(n186) );
  NANDN U237 ( .B(n177), .A(Y0[3]), .Z(n185) );
  NAND U238 ( .A(n188), .B(n189), .Z(n134) );
  NANDN U239 ( .B(n176), .A(n190), .Z(n189) );
  NANDN U240 ( .B(n177), .A(Y0[4]), .Z(n188) );
  NAND U241 ( .A(n191), .B(n192), .Z(n133) );
  NANDN U242 ( .B(n176), .A(n193), .Z(n192) );
  NANDN U243 ( .B(n177), .A(Y0[5]), .Z(n191) );
  NAND U244 ( .A(n194), .B(n195), .Z(n132) );
  OR U245 ( .A(n196), .B(n176), .Z(n195) );
  NANDN U246 ( .B(n177), .A(Y0[6]), .Z(n194) );
  NAND U247 ( .A(n197), .B(n198), .Z(n131) );
  OR U248 ( .A(n176), .B(n199), .Z(n198) );
  NANDN U249 ( .B(n200), .A(n177), .Z(n176) );
  NANDN U250 ( .B(n177), .A(Y0[7]), .Z(n197) );
  NAND U251 ( .A(n201), .B(n202), .Z(n130) );
  NANDN U252 ( .B(n177), .A(Y[7]), .Z(n202) );
  AND U253 ( .A(n203), .B(n204), .Z(n201) );
  NANDN U254 ( .B(n200), .A(Y[7]), .Z(n204) );
  OR U255 ( .A(n199), .B(n205), .Z(n203) );
  XOR U256 ( .A(n206), .B(n207), .Z(n199) );
  XNOR U257 ( .A(Y0[7]), .B(n208), .Z(n207) );
  NAND U258 ( .A(n211), .B(n212), .Z(n129) );
  NANDN U259 ( .B(n177), .A(Y[6]), .Z(n212) );
  AND U260 ( .A(n213), .B(n214), .Z(n211) );
  NANDN U261 ( .B(n200), .A(Y[6]), .Z(n214) );
  OR U262 ( .A(n196), .B(n205), .Z(n213) );
  XOR U263 ( .A(n210), .B(Y0[7]), .Z(n196) );
  XOR U264 ( .A(n209), .B(n208), .Z(n210) );
  NAND U265 ( .A(n217), .B(n218), .Z(n128) );
  NANDN U266 ( .B(n177), .A(Y[5]), .Z(n218) );
  AND U267 ( .A(n219), .B(n220), .Z(n217) );
  NANDN U268 ( .B(n200), .A(Y[5]), .Z(n220) );
  NANDN U269 ( .B(n205), .A(n193), .Z(n219) );
  XNOR U270 ( .A(n216), .B(Y0[6]), .Z(n193) );
  XOR U271 ( .A(n221), .B(n222), .Z(n216) );
  ANDN U272 ( .A(n208), .B(n223), .Z(n222) );
  NANDN U273 ( .B(n224), .A(n225), .Z(n208) );
  ANDN U274 ( .A(n226), .B(n223), .Z(n224) );
  NAND U275 ( .A(n227), .B(n228), .Z(n223) );
  OR U276 ( .A(n229), .B(n230), .Z(n228) );
  AND U277 ( .A(n231), .B(n232), .Z(n227) );
  OR U278 ( .A(n233), .B(n234), .Z(n232) );
  OR U279 ( .A(n235), .B(n236), .Z(n231) );
  NOR U280 ( .A(n237), .B(n238), .Z(n226) );
  IV U281 ( .A(n215), .Z(n221) );
  XOR U282 ( .A(n239), .B(n240), .Z(n215) );
  ANDN U283 ( .A(n241), .B(n242), .Z(n240) );
  XNOR U284 ( .A(Y0[5]), .B(n239), .Z(n241) );
  NAND U285 ( .A(n243), .B(n244), .Z(n127) );
  NANDN U286 ( .B(n177), .A(Y[4]), .Z(n244) );
  AND U287 ( .A(n245), .B(n246), .Z(n243) );
  NANDN U288 ( .B(n200), .A(Y[4]), .Z(n246) );
  NANDN U289 ( .B(n205), .A(n190), .Z(n245) );
  XNOR U290 ( .A(n242), .B(Y0[5]), .Z(n190) );
  XNOR U291 ( .A(n247), .B(n248), .Z(n242) );
  AND U292 ( .A(n225), .B(n250), .Z(n249) );
  XOR U293 ( .A(n237), .B(n251), .Z(n250) );
  XOR U294 ( .A(n251), .B(n238), .Z(n237) );
  OR U295 ( .A(n252), .B(n253), .Z(n238) );
  IV U296 ( .A(n248), .Z(n251) );
  XNOR U297 ( .A(n236), .B(n235), .Z(n248) );
  OR U298 ( .A(n254), .B(n255), .Z(n235) );
  AND U299 ( .A(n256), .B(n257), .Z(n236) );
  XNOR U300 ( .A(n258), .B(n259), .Z(n257) );
  ANDN U301 ( .A(n260), .B(n261), .Z(n259) );
  XOR U302 ( .A(n258), .B(n262), .Z(n260) );
  XNOR U303 ( .A(n229), .B(n263), .Z(n256) );
  NAND U304 ( .A(n265), .B(n266), .Z(n230) );
  NANDN U305 ( .B(n267), .A(n268), .Z(n265) );
  NANDN U306 ( .B(n233), .A(n269), .Z(n264) );
  NANDN U307 ( .B(n234), .A(n270), .Z(n229) );
  XOR U308 ( .A(n271), .B(n272), .Z(n239) );
  ANDN U309 ( .A(n273), .B(n274), .Z(n272) );
  XNOR U310 ( .A(Y0[4]), .B(n271), .Z(n273) );
  NAND U311 ( .A(n275), .B(n276), .Z(n126) );
  NANDN U312 ( .B(n177), .A(Y[3]), .Z(n276) );
  AND U313 ( .A(n277), .B(n278), .Z(n275) );
  NANDN U314 ( .B(n200), .A(Y[3]), .Z(n278) );
  NANDN U315 ( .B(n205), .A(n187), .Z(n277) );
  XNOR U316 ( .A(n274), .B(Y0[4]), .Z(n187) );
  XNOR U317 ( .A(n279), .B(n280), .Z(n274) );
  AND U318 ( .A(n225), .B(n282), .Z(n281) );
  XOR U319 ( .A(n252), .B(n283), .Z(n282) );
  XOR U320 ( .A(n283), .B(n253), .Z(n252) );
  OR U321 ( .A(n284), .B(n285), .Z(n253) );
  IV U322 ( .A(n280), .Z(n283) );
  XNOR U323 ( .A(n255), .B(n254), .Z(n280) );
  OR U324 ( .A(n286), .B(n287), .Z(n254) );
  XOR U325 ( .A(n262), .B(n261), .Z(n255) );
  XOR U326 ( .A(n258), .B(n288), .Z(n261) );
  AND U327 ( .A(n289), .B(n290), .Z(n288) );
  NANDN U328 ( .B(n233), .A(n291), .Z(n290) );
  OR U329 ( .A(n292), .B(n293), .Z(n289) );
  XOR U330 ( .A(n267), .B(n268), .Z(n262) );
  NANDN U331 ( .B(n234), .A(n297), .Z(n268) );
  XNOR U332 ( .A(n266), .B(n298), .Z(n267) );
  AND U333 ( .A(n270), .B(n269), .Z(n298) );
  ANDN U334 ( .A(n299), .B(n300), .Z(n266) );
  NANDN U335 ( .B(n301), .A(n302), .Z(n299) );
  NAND U336 ( .A(n305), .B(n306), .Z(n125) );
  NANDN U337 ( .B(n177), .A(Y[2]), .Z(n306) );
  AND U338 ( .A(n307), .B(n308), .Z(n305) );
  NANDN U339 ( .B(n200), .A(Y[2]), .Z(n308) );
  NANDN U340 ( .B(n205), .A(n184), .Z(n307) );
  XNOR U341 ( .A(n304), .B(Y0[3]), .Z(n184) );
  XNOR U342 ( .A(n309), .B(n310), .Z(n304) );
  AND U343 ( .A(n225), .B(n312), .Z(n311) );
  XOR U344 ( .A(n284), .B(n313), .Z(n312) );
  XOR U345 ( .A(n313), .B(n285), .Z(n284) );
  OR U346 ( .A(n314), .B(n315), .Z(n285) );
  IV U347 ( .A(n310), .Z(n313) );
  XOR U348 ( .A(n296), .B(n295), .Z(n286) );
  XNOR U349 ( .A(n319), .B(n320), .Z(n295) );
  IV U350 ( .A(n294), .Z(n320) );
  XOR U351 ( .A(n321), .B(n322), .Z(n294) );
  ANDN U352 ( .A(n323), .B(n324), .Z(n322) );
  XOR U353 ( .A(n321), .B(n325), .Z(n323) );
  XNOR U354 ( .A(n326), .B(n292), .Z(n319) );
  NAND U355 ( .A(n291), .B(n270), .Z(n292) );
  NANDN U356 ( .B(n233), .A(n328), .Z(n327) );
  XNOR U357 ( .A(n329), .B(n330), .Z(n293) );
  ANDN U358 ( .A(n331), .B(n332), .Z(n330) );
  XNOR U359 ( .A(n333), .B(n329), .Z(n331) );
  XOR U360 ( .A(n301), .B(n302), .Z(n296) );
  OR U361 ( .A(n334), .B(n234), .Z(n302) );
  XNOR U362 ( .A(n335), .B(n336), .Z(n301) );
  AND U363 ( .A(n297), .B(n269), .Z(n336) );
  IV U364 ( .A(n300), .Z(n335) );
  NAND U365 ( .A(n337), .B(n338), .Z(n300) );
  NANDN U366 ( .B(n339), .A(n340), .Z(n337) );
  NAND U367 ( .A(n343), .B(n344), .Z(n124) );
  NANDN U368 ( .B(n177), .A(Y[1]), .Z(n344) );
  AND U369 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U370 ( .B(n200), .A(Y[1]), .Z(n346) );
  NANDN U371 ( .B(n205), .A(n180), .Z(n345) );
  XNOR U372 ( .A(n342), .B(Y0[2]), .Z(n180) );
  XNOR U373 ( .A(n347), .B(n348), .Z(n342) );
  XOR U374 ( .A(n341), .B(n349), .Z(n347) );
  AND U375 ( .A(n225), .B(n350), .Z(n349) );
  XOR U376 ( .A(n314), .B(n351), .Z(n350) );
  XOR U377 ( .A(n351), .B(n315), .Z(n314) );
  NANDN U378 ( .B(n352), .A(n353), .Z(n315) );
  IV U379 ( .A(n348), .Z(n351) );
  XOR U380 ( .A(n318), .B(n317), .Z(n348) );
  XNOR U381 ( .A(n316), .B(n354), .Z(n317) );
  AND U382 ( .A(n355), .B(n356), .Z(n354) );
  OR U383 ( .A(n357), .B(n358), .Z(n356) );
  AND U384 ( .A(n359), .B(n360), .Z(n355) );
  NANDN U385 ( .B(n233), .A(n361), .Z(n360) );
  NAND U386 ( .A(n362), .B(n363), .Z(n359) );
  XNOR U387 ( .A(n329), .B(n368), .Z(n332) );
  AND U388 ( .A(n270), .B(n328), .Z(n368) );
  XOR U389 ( .A(n369), .B(n370), .Z(n329) );
  ANDN U390 ( .A(n371), .B(n372), .Z(n370) );
  XNOR U391 ( .A(n373), .B(n369), .Z(n371) );
  XOR U392 ( .A(n374), .B(n333), .Z(n367) );
  NAND U393 ( .A(n291), .B(n297), .Z(n333) );
  IV U394 ( .A(n321), .Z(n374) );
  XOR U395 ( .A(n375), .B(n376), .Z(n321) );
  ANDN U396 ( .A(n377), .B(n378), .Z(n376) );
  XOR U397 ( .A(n375), .B(n379), .Z(n377) );
  XNOR U398 ( .A(n339), .B(n340), .Z(n325) );
  OR U399 ( .A(n380), .B(n234), .Z(n340) );
  XNOR U400 ( .A(n338), .B(n381), .Z(n339) );
  ANDN U401 ( .A(n269), .B(n334), .Z(n381) );
  ANDN U402 ( .A(n382), .B(n383), .Z(n338) );
  NANDN U403 ( .B(n384), .A(n385), .Z(n382) );
  NAND U404 ( .A(n388), .B(n389), .Z(n123) );
  NANDN U405 ( .B(n177), .A(Y[0]), .Z(n389) );
  AND U406 ( .A(n390), .B(n391), .Z(n388) );
  NANDN U407 ( .B(n200), .A(Y[0]), .Z(n391) );
  IV U408 ( .A(n392), .Z(n200) );
  OR U409 ( .A(n205), .B(n175), .Z(n390) );
  IV U410 ( .A(Y0[1]), .Z(n181) );
  XOR U411 ( .A(n393), .B(n394), .Z(n387) );
  XNOR U412 ( .A(n395), .B(n386), .Z(n393) );
  NAND U413 ( .A(Y0[0]), .B(n352), .Z(n386) );
  NAND U414 ( .A(n396), .B(n225), .Z(n395) );
  XOR U415 ( .A(A[7]), .B(X[7]), .Z(n225) );
  XNOR U416 ( .A(n353), .B(n394), .Z(n396) );
  XNOR U417 ( .A(n352), .B(n394), .Z(n353) );
  XNOR U418 ( .A(n366), .B(n365), .Z(n394) );
  XNOR U419 ( .A(n397), .B(n362), .Z(n365) );
  XNOR U420 ( .A(n398), .B(n357), .Z(n362) );
  NAND U421 ( .A(n270), .B(n361), .Z(n357) );
  NANDN U422 ( .B(n233), .A(n400), .Z(n399) );
  XNOR U423 ( .A(n363), .B(n364), .Z(n397) );
  XNOR U424 ( .A(n369), .B(n411), .Z(n372) );
  AND U425 ( .A(n297), .B(n328), .Z(n411) );
  XOR U426 ( .A(n412), .B(n413), .Z(n369) );
  ANDN U427 ( .A(n414), .B(n415), .Z(n413) );
  XNOR U428 ( .A(n416), .B(n412), .Z(n414) );
  XOR U429 ( .A(n417), .B(n373), .Z(n410) );
  NANDN U430 ( .B(n334), .A(n291), .Z(n373) );
  IV U431 ( .A(n375), .Z(n417) );
  XNOR U432 ( .A(n384), .B(n385), .Z(n379) );
  NANDN U433 ( .B(n234), .A(n421), .Z(n385) );
  ANDN U434 ( .A(n269), .B(n380), .Z(n422) );
  NAND U435 ( .A(n423), .B(n424), .Z(n383) );
  NANDN U436 ( .B(n425), .A(n426), .Z(n423) );
  XNOR U437 ( .A(n406), .B(n405), .Z(n352) );
  XNOR U438 ( .A(n427), .B(n409), .Z(n405) );
  XNOR U439 ( .A(n402), .B(n403), .Z(n409) );
  NAND U440 ( .A(n297), .B(n361), .Z(n403) );
  XNOR U441 ( .A(n401), .B(n428), .Z(n402) );
  AND U442 ( .A(n400), .B(n270), .Z(n428) );
  XOR U443 ( .A(n429), .B(n430), .Z(n401) );
  AND U444 ( .A(n431), .B(n432), .Z(n430) );
  XNOR U445 ( .A(n433), .B(n429), .Z(n432) );
  XNOR U446 ( .A(n408), .B(n404), .Z(n427) );
  XOR U447 ( .A(n434), .B(n435), .Z(n404) );
  XOR U448 ( .A(n436), .B(n437), .Z(n408) );
  AND U449 ( .A(n438), .B(n439), .Z(n437) );
  NANDN U450 ( .B(n233), .A(n440), .Z(n439) );
  NANDN U451 ( .B(n441), .A(n442), .Z(n233) );
  AND U452 ( .A(n443), .B(A[7]), .Z(n442) );
  NANDN U453 ( .B(n444), .A(n445), .Z(n438) );
  IV U454 ( .A(n407), .Z(n436) );
  XNOR U455 ( .A(n446), .B(n447), .Z(n407) );
  AND U456 ( .A(n448), .B(n449), .Z(n447) );
  XOR U457 ( .A(n445), .B(n450), .Z(n449) );
  XNOR U458 ( .A(n444), .B(n446), .Z(n450) );
  NAND U459 ( .A(n270), .B(n440), .Z(n444) );
  XNOR U460 ( .A(n454), .B(n451), .Z(n453) );
  XOR U461 ( .A(n431), .B(n455), .Z(n448) );
  XNOR U462 ( .A(n433), .B(n446), .Z(n455) );
  NANDN U463 ( .B(n334), .A(n361), .Z(n433) );
  XOR U464 ( .A(n429), .B(n456), .Z(n431) );
  AND U465 ( .A(n400), .B(n297), .Z(n456) );
  XOR U466 ( .A(n457), .B(n458), .Z(n429) );
  AND U467 ( .A(n459), .B(n460), .Z(n458) );
  XNOR U468 ( .A(n461), .B(n457), .Z(n460) );
  XOR U469 ( .A(n462), .B(n463), .Z(n446) );
  AND U470 ( .A(n464), .B(n465), .Z(n463) );
  XOR U471 ( .A(n452), .B(n466), .Z(n465) );
  XNOR U472 ( .A(n454), .B(n462), .Z(n466) );
  NAND U473 ( .A(n297), .B(n440), .Z(n454) );
  XOR U474 ( .A(n451), .B(n467), .Z(n452) );
  AND U475 ( .A(n270), .B(X[0]), .Z(n467) );
  XNOR U476 ( .A(n443), .B(A[6]), .Z(n441) );
  NOR U477 ( .A(n468), .B(n469), .Z(n443) );
  XNOR U478 ( .A(n473), .B(n470), .Z(n472) );
  XOR U479 ( .A(n459), .B(n474), .Z(n464) );
  XNOR U480 ( .A(n461), .B(n462), .Z(n474) );
  NANDN U481 ( .B(n380), .A(n361), .Z(n461) );
  XOR U482 ( .A(n457), .B(n475), .Z(n459) );
  ANDN U483 ( .A(n400), .B(n334), .Z(n475) );
  XOR U484 ( .A(n476), .B(n477), .Z(n457) );
  AND U485 ( .A(n478), .B(n479), .Z(n477) );
  XNOR U486 ( .A(n480), .B(n476), .Z(n479) );
  XOR U487 ( .A(n481), .B(n482), .Z(n462) );
  AND U488 ( .A(n483), .B(n484), .Z(n482) );
  XOR U489 ( .A(n471), .B(n485), .Z(n484) );
  XNOR U490 ( .A(n473), .B(n481), .Z(n485) );
  NANDN U491 ( .B(n334), .A(n440), .Z(n473) );
  XOR U492 ( .A(n470), .B(n486), .Z(n471) );
  AND U493 ( .A(n297), .B(X[0]), .Z(n486) );
  XOR U494 ( .A(n468), .B(A[5]), .Z(n469) );
  NANDN U495 ( .B(n487), .A(n488), .Z(n468) );
  XOR U496 ( .A(n489), .B(n490), .Z(n470) );
  ANDN U497 ( .A(n491), .B(n492), .Z(n490) );
  XNOR U498 ( .A(n493), .B(n489), .Z(n491) );
  XOR U499 ( .A(n478), .B(n494), .Z(n483) );
  XNOR U500 ( .A(n480), .B(n481), .Z(n494) );
  NAND U501 ( .A(n361), .B(n421), .Z(n480) );
  XOR U502 ( .A(n476), .B(n495), .Z(n478) );
  ANDN U503 ( .A(n400), .B(n380), .Z(n495) );
  XOR U504 ( .A(n496), .B(n497), .Z(n476) );
  ANDN U505 ( .A(n498), .B(n499), .Z(n497) );
  XNOR U506 ( .A(n500), .B(n496), .Z(n498) );
  XNOR U507 ( .A(n502), .B(n500), .Z(n434) );
  NAND U508 ( .A(n361), .B(n503), .Z(n500) );
  IV U509 ( .A(n499), .Z(n502) );
  XNOR U510 ( .A(n496), .B(n504), .Z(n499) );
  AND U511 ( .A(n421), .B(n400), .Z(n504) );
  AND U512 ( .A(n505), .B(A[0]), .Z(n496) );
  NANDN U513 ( .B(n361), .A(n506), .Z(n505) );
  NAND U514 ( .A(n503), .B(n400), .Z(n506) );
  XNOR U515 ( .A(n507), .B(X[2]), .Z(n400) );
  NAND U516 ( .A(n508), .B(X[7]), .Z(n507) );
  XOR U517 ( .A(n509), .B(X[2]), .Z(n508) );
  XNOR U518 ( .A(n489), .B(n512), .Z(n492) );
  ANDN U519 ( .A(X[0]), .B(n334), .Z(n512) );
  XOR U520 ( .A(n513), .B(n514), .Z(n489) );
  AND U521 ( .A(n515), .B(n516), .Z(n514) );
  XOR U522 ( .A(n517), .B(n513), .Z(n516) );
  ANDN U523 ( .A(X[0]), .B(n380), .Z(n517) );
  XOR U524 ( .A(n518), .B(n513), .Z(n515) );
  AND U525 ( .A(n440), .B(n421), .Z(n518) );
  XOR U526 ( .A(n519), .B(n520), .Z(n513) );
  ANDN U527 ( .A(n521), .B(n522), .Z(n520) );
  XNOR U528 ( .A(n523), .B(n519), .Z(n521) );
  XOR U529 ( .A(n524), .B(n493), .Z(n511) );
  NANDN U530 ( .B(n380), .A(n440), .Z(n493) );
  IV U531 ( .A(n501), .Z(n524) );
  NAND U532 ( .A(n440), .B(n503), .Z(n523) );
  XNOR U533 ( .A(n519), .B(n525), .Z(n522) );
  AND U534 ( .A(n421), .B(X[0]), .Z(n525) );
  AND U535 ( .A(n526), .B(A[0]), .Z(n519) );
  NANDN U536 ( .B(n440), .A(n527), .Z(n526) );
  NAND U537 ( .A(n503), .B(X[0]), .Z(n527) );
  XNOR U538 ( .A(n528), .B(X[1]), .Z(n440) );
  NAND U539 ( .A(n529), .B(X[7]), .Z(n528) );
  XNOR U540 ( .A(X[1]), .B(n530), .Z(n529) );
  XOR U541 ( .A(n531), .B(n532), .Z(n419) );
  IV U542 ( .A(n415), .Z(n532) );
  XNOR U543 ( .A(n412), .B(n533), .Z(n415) );
  ANDN U544 ( .A(n328), .B(n334), .Z(n533) );
  XNOR U545 ( .A(n488), .B(A[4]), .Z(n487) );
  NOR U546 ( .A(n534), .B(n535), .Z(n488) );
  XOR U547 ( .A(n538), .B(n536), .Z(n537) );
  ANDN U548 ( .A(n328), .B(n380), .Z(n538) );
  AND U549 ( .A(n421), .B(n291), .Z(n539) );
  XOR U550 ( .A(n543), .B(n416), .Z(n531) );
  NANDN U551 ( .B(n380), .A(n291), .Z(n416) );
  NANDN U552 ( .B(n544), .A(n545), .Z(n534) );
  IV U553 ( .A(n418), .Z(n543) );
  XOR U554 ( .A(n546), .B(n542), .Z(n418) );
  NAND U555 ( .A(n291), .B(n503), .Z(n542) );
  IV U556 ( .A(n541), .Z(n546) );
  XNOR U557 ( .A(n540), .B(n547), .Z(n541) );
  AND U558 ( .A(n421), .B(n328), .Z(n547) );
  AND U559 ( .A(n548), .B(A[0]), .Z(n540) );
  NANDN U560 ( .B(n291), .A(n549), .Z(n548) );
  NAND U561 ( .A(n503), .B(n328), .Z(n549) );
  XNOR U562 ( .A(n550), .B(X[4]), .Z(n328) );
  NAND U563 ( .A(n551), .B(X[7]), .Z(n550) );
  XOR U564 ( .A(n552), .B(X[4]), .Z(n551) );
  XNOR U565 ( .A(n553), .B(X[5]), .Z(n291) );
  NAND U566 ( .A(n554), .B(X[7]), .Z(n553) );
  XOR U567 ( .A(n555), .B(X[5]), .Z(n554) );
  XNOR U568 ( .A(n425), .B(n426), .Z(n420) );
  NANDN U569 ( .B(n234), .A(n503), .Z(n426) );
  XNOR U570 ( .A(n424), .B(n556), .Z(n425) );
  AND U571 ( .A(n421), .B(n269), .Z(n556) );
  XNOR U572 ( .A(n545), .B(A[2]), .Z(n544) );
  AND U573 ( .A(n558), .B(A[0]), .Z(n424) );
  NAND U574 ( .A(n559), .B(n234), .Z(n558) );
  NANDN U575 ( .B(n560), .A(n561), .Z(n234) );
  ANDN U576 ( .A(X[7]), .B(n562), .Z(n561) );
  NAND U577 ( .A(n503), .B(n269), .Z(n559) );
  XOR U578 ( .A(n562), .B(X[6]), .Z(n560) );
  OR U579 ( .A(n555), .B(n563), .Z(n562) );
  XOR U580 ( .A(n563), .B(X[5]), .Z(n555) );
  OR U581 ( .A(n552), .B(n564), .Z(n563) );
  XOR U582 ( .A(n564), .B(X[4]), .Z(n552) );
  OR U583 ( .A(n510), .B(n565), .Z(n564) );
  XOR U584 ( .A(n565), .B(X[3]), .Z(n510) );
  OR U585 ( .A(n509), .B(n566), .Z(n565) );
  XOR U586 ( .A(n566), .B(X[2]), .Z(n509) );
  NANDN U587 ( .B(X[0]), .A(n530), .Z(n566) );
  XNOR U588 ( .A(X[0]), .B(X[1]), .Z(n530) );
  XNOR U589 ( .A(n567), .B(A[1]), .Z(n503) );
  NAND U590 ( .A(n568), .B(A[7]), .Z(n567) );
  XOR U591 ( .A(A[1]), .B(n557), .Z(n568) );
  XOR U592 ( .A(A[0]), .B(A[1]), .Z(n557) );
  NANDN U593 ( .B(n392), .A(n177), .Z(n205) );
  IV U594 ( .A(rst), .Z(n177) );
  NAND U595 ( .A(n569), .B(n570), .Z(n392) );
  AND U596 ( .A(n571), .B(n572), .Z(n570) );
  ANDN U597 ( .A(n573), .B(n[7]), .Z(n572) );
  NOR U598 ( .A(n[9]), .B(n[8]), .Z(n573) );
  NOR U599 ( .A(n[5]), .B(n[6]), .Z(n571) );
  AND U600 ( .A(n574), .B(n575), .Z(n569) );
  NOR U601 ( .A(n[1]), .B(n[2]), .Z(n575) );
  NOR U602 ( .A(n[0]), .B(n170), .Z(n574) );
  OR U603 ( .A(n[3]), .B(n[4]), .Z(n170) );
endmodule

