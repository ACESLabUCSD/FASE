
module MxM_TG_W8_N100 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n133 , \_MxM/n132 , \_MxM/n131 , \_MxM/n130 , \_MxM/n129 ,
         \_MxM/n128 , \_MxM/n127 , \_MxM/n126 , \_MxM/n125 , \_MxM/n124 ,
         \_MxM/n123 , \_MxM/n122 , \_MxM/n121 , \_MxM/n120 , \_MxM/n119 ,
         \_MxM/n118 , \_MxM/n117 , \_MxM/n116 , \_MxM/n115 , \_MxM/n114 ,
         \_MxM/n113 , \_MxM/n112 , \_MxM/n111 , \_MxM/N12 , \_MxM/N11 ,
         \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/Y0[0] , \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] , \_MxM/Y0[4] ,
         \_MxM/Y0[5] , \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/add_39/carry[6] ,
         \_MxM/add_39/carry[5] , \_MxM/add_39/carry[4] ,
         \_MxM/add_39/carry[3] , \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n111 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n112 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n113 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n114 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n115 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n116 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n117 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n118 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n119 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n120 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n121 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n122 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n123 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n124 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n125 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n126 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n127 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n128 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n129 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n130 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n131 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n132 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n133 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  MUX U1 ( .IN0(n319), .IN1(n335), .SEL(n321), .F(n300) );
  MUX U2 ( .IN0(g_input[3]), .IN1(n384), .SEL(g_input[7]), .F(n1) );
  IV U3 ( .A(n1), .Z(n229) );
  MUX U4 ( .IN0(n269), .IN1(n267), .SEL(n268), .F(n224) );
  NAND U5 ( .A(n142), .B(n176), .Z(n175) );
  MUX U6 ( .IN0(n252), .IN1(n2), .SEL(n251), .F(n207) );
  IV U7 ( .A(n250), .Z(n2) );
  MUX U8 ( .IN0(n3), .IN1(n152), .SEL(n153), .F(n120) );
  IV U9 ( .A(\_MxM/Y0[3] ), .Z(n3) );
  XOR U10 ( .A(n383), .B(g_input[3]), .Z(n384) );
  XNOR U11 ( .A(n371), .B(n372), .Z(n350) );
  MUX U12 ( .IN0(e_input[6]), .IN1(n409), .SEL(e_input[7]), .F(n118) );
  MUX U13 ( .IN0(e_input[3]), .IN1(n359), .SEL(e_input[7]), .F(n210) );
  MUX U14 ( .IN0(n213), .IN1(n4), .SEL(n214), .F(n165) );
  IV U15 ( .A(n215), .Z(n4) );
  XNOR U16 ( .A(n216), .B(n181), .Z(n173) );
  MUX U17 ( .IN0(n5), .IN1(n235), .SEL(n236), .F(n190) );
  IV U18 ( .A(\_MxM/Y0[1] ), .Z(n5) );
  XOR U19 ( .A(n88), .B(n98), .Z(n96) );
  MUX U20 ( .IN0(n6), .IN1(n389), .SEL(n390), .F(n385) );
  IV U21 ( .A(n391), .Z(n6) );
  MUX U22 ( .IN0(g_input[4]), .IN1(n336), .SEL(g_input[7]), .F(n7) );
  IV U23 ( .A(n7), .Z(n183) );
  MUX U24 ( .IN0(g_input[5]), .IN1(n318), .SEL(g_input[7]), .F(n146) );
  XOR U25 ( .A(n232), .B(n271), .Z(n233) );
  MUX U26 ( .IN0(g_input[6]), .IN1(n290), .SEL(g_input[7]), .F(n119) );
  MUX U27 ( .IN0(n253), .IN1(n8), .SEL(n254), .F(n213) );
  IV U28 ( .A(n255), .Z(n8) );
  XNOR U29 ( .A(n135), .B(n136), .Z(n159) );
  XOR U30 ( .A(n120), .B(n130), .Z(n128) );
  NOR U31 ( .A(g_input[0]), .B(n406), .Z(n394) );
  MUX U32 ( .IN0(n9), .IN1(n283), .SEL(n284), .F(n330) );
  IV U33 ( .A(n350), .Z(n9) );
  MUX U34 ( .IN0(n385), .IN1(n388), .SEL(n386), .F(n261) );
  MUX U35 ( .IN0(n300), .IN1(n316), .SEL(n302), .F(n294) );
  MUX U36 ( .IN0(n145), .IN1(n169), .SEL(n144), .F(n107) );
  NAND U37 ( .A(n207), .B(n248), .Z(n247) );
  XNOR U38 ( .A(n269), .B(n268), .Z(n255) );
  XNOR U39 ( .A(n174), .B(n173), .Z(n167) );
  XNOR U40 ( .A(n228), .B(n227), .Z(n215) );
  MUX U41 ( .IN0(\_MxM/Y0[6] ), .IN1(n70), .SEL(n65), .F(n58) );
  XOR U42 ( .A(n152), .B(n160), .Z(n158) );
  MUX U43 ( .IN0(g_input[2]), .IN1(n393), .SEL(g_input[7]), .F(n270) );
  XOR U44 ( .A(n360), .B(n341), .Z(n284) );
  XNOR U45 ( .A(n259), .B(n221), .Z(n227) );
  MUX U46 ( .IN0(n258), .IN1(n256), .SEL(n257), .F(n10) );
  IV U47 ( .A(n10), .Z(n212) );
  AND U48 ( .A(n113), .B(n79), .Z(n112) );
  MUX U49 ( .IN0(n11), .IN1(n167), .SEL(n166), .F(n136) );
  IV U50 ( .A(n165), .Z(n11) );
  MUX U51 ( .IN0(n12), .IN1(n190), .SEL(n191), .F(n152) );
  IV U52 ( .A(\_MxM/Y0[2] ), .Z(n12) );
  MUX U53 ( .IN0(\_MxM/Y0[7] ), .IN1(n58), .SEL(n59), .F(n13) );
  IV U54 ( .A(n13), .Z(n55) );
  XOR U55 ( .A(n236), .B(\_MxM/Y0[1] ), .Z(n24) );
  ANDN U56 ( .A(n14), .B(\_MxM/n[0] ), .Z(\_MxM/n133 ) );
  AND U57 ( .A(\_MxM/N8 ), .B(n14), .Z(\_MxM/n132 ) );
  AND U58 ( .A(\_MxM/N9 ), .B(n14), .Z(\_MxM/n131 ) );
  AND U59 ( .A(\_MxM/N10 ), .B(n14), .Z(\_MxM/n130 ) );
  AND U60 ( .A(\_MxM/N11 ), .B(n14), .Z(\_MxM/n129 ) );
  AND U61 ( .A(\_MxM/N12 ), .B(n14), .Z(\_MxM/n128 ) );
  AND U62 ( .A(n14), .B(n15), .Z(\_MxM/n127 ) );
  XOR U63 ( .A(\_MxM/n[6] ), .B(\_MxM/add_39/carry[6] ), .Z(n15) );
  ANDN U64 ( .A(n16), .B(rst), .Z(n14) );
  NAND U65 ( .A(n17), .B(n18), .Z(n16) );
  AND U66 ( .A(\_MxM/n[0] ), .B(n19), .Z(n18) );
  NOR U67 ( .A(n20), .B(\_MxM/n[2] ), .Z(n19) );
  AND U68 ( .A(n21), .B(\_MxM/n[6] ), .Z(n17) );
  AND U69 ( .A(\_MxM/n[5] ), .B(\_MxM/n[1] ), .Z(n21) );
  NAND U70 ( .A(n22), .B(n23), .Z(\_MxM/n126 ) );
  OR U71 ( .A(n24), .B(n25), .Z(n23) );
  NANDN U72 ( .B(n26), .A(\_MxM/Y0[0] ), .Z(n22) );
  NAND U73 ( .A(n27), .B(n28), .Z(\_MxM/n125 ) );
  NANDN U74 ( .B(n25), .A(n29), .Z(n28) );
  NANDN U75 ( .B(n30), .A(rst), .Z(n27) );
  NAND U76 ( .A(n31), .B(n32), .Z(\_MxM/n124 ) );
  NANDN U77 ( .B(n25), .A(n33), .Z(n32) );
  NANDN U78 ( .B(n26), .A(\_MxM/Y0[2] ), .Z(n31) );
  NAND U79 ( .A(n34), .B(n35), .Z(\_MxM/n123 ) );
  NANDN U80 ( .B(n25), .A(n36), .Z(n35) );
  NANDN U81 ( .B(n26), .A(\_MxM/Y0[3] ), .Z(n34) );
  NAND U82 ( .A(n37), .B(n38), .Z(\_MxM/n122 ) );
  NANDN U83 ( .B(n25), .A(n39), .Z(n38) );
  NANDN U84 ( .B(n26), .A(\_MxM/Y0[4] ), .Z(n37) );
  NAND U85 ( .A(n40), .B(n41), .Z(\_MxM/n121 ) );
  NANDN U86 ( .B(n25), .A(n42), .Z(n41) );
  NANDN U87 ( .B(n26), .A(\_MxM/Y0[5] ), .Z(n40) );
  NAND U88 ( .A(n43), .B(n44), .Z(\_MxM/n120 ) );
  OR U89 ( .A(n45), .B(n25), .Z(n44) );
  NANDN U90 ( .B(n26), .A(\_MxM/Y0[6] ), .Z(n43) );
  NAND U91 ( .A(n46), .B(n47), .Z(\_MxM/n119 ) );
  OR U92 ( .A(n25), .B(n48), .Z(n47) );
  NANDN U93 ( .B(n49), .A(n26), .Z(n25) );
  NANDN U94 ( .B(n26), .A(\_MxM/Y0[7] ), .Z(n46) );
  NAND U95 ( .A(n50), .B(n51), .Z(\_MxM/n118 ) );
  NANDN U96 ( .B(n26), .A(o[7]), .Z(n51) );
  AND U97 ( .A(n52), .B(n53), .Z(n50) );
  NANDN U98 ( .B(n49), .A(o[7]), .Z(n53) );
  OR U99 ( .A(n48), .B(n54), .Z(n52) );
  XOR U100 ( .A(n55), .B(n56), .Z(n48) );
  XNOR U101 ( .A(\_MxM/Y0[7] ), .B(n57), .Z(n56) );
  NAND U102 ( .A(n60), .B(n61), .Z(\_MxM/n117 ) );
  NANDN U103 ( .B(n26), .A(o[6]), .Z(n61) );
  AND U104 ( .A(n62), .B(n63), .Z(n60) );
  NANDN U105 ( .B(n49), .A(o[6]), .Z(n63) );
  OR U106 ( .A(n45), .B(n54), .Z(n62) );
  XOR U107 ( .A(n59), .B(\_MxM/Y0[7] ), .Z(n45) );
  XOR U108 ( .A(n58), .B(n57), .Z(n59) );
  NAND U109 ( .A(n66), .B(n67), .Z(\_MxM/n116 ) );
  NANDN U110 ( .B(n26), .A(o[5]), .Z(n67) );
  AND U111 ( .A(n68), .B(n69), .Z(n66) );
  NANDN U112 ( .B(n49), .A(o[5]), .Z(n69) );
  NANDN U113 ( .B(n54), .A(n42), .Z(n68) );
  XNOR U114 ( .A(n65), .B(\_MxM/Y0[6] ), .Z(n42) );
  XOR U115 ( .A(n70), .B(n71), .Z(n65) );
  ANDN U116 ( .A(n57), .B(n72), .Z(n71) );
  NANDN U117 ( .B(n73), .A(n74), .Z(n57) );
  ANDN U118 ( .A(n75), .B(n72), .Z(n73) );
  NAND U119 ( .A(n76), .B(n77), .Z(n72) );
  OR U120 ( .A(n78), .B(n79), .Z(n77) );
  AND U121 ( .A(n80), .B(n81), .Z(n76) );
  OR U122 ( .A(n82), .B(n83), .Z(n81) );
  OR U123 ( .A(n84), .B(n85), .Z(n80) );
  NOR U124 ( .A(n86), .B(n87), .Z(n75) );
  IV U125 ( .A(n64), .Z(n70) );
  XOR U126 ( .A(n88), .B(n89), .Z(n64) );
  ANDN U127 ( .A(n90), .B(n91), .Z(n89) );
  XNOR U128 ( .A(\_MxM/Y0[5] ), .B(n88), .Z(n90) );
  NAND U129 ( .A(n92), .B(n93), .Z(\_MxM/n115 ) );
  NANDN U130 ( .B(n26), .A(o[4]), .Z(n93) );
  AND U131 ( .A(n94), .B(n95), .Z(n92) );
  NANDN U132 ( .B(n49), .A(o[4]), .Z(n95) );
  NANDN U133 ( .B(n54), .A(n39), .Z(n94) );
  XNOR U134 ( .A(n91), .B(\_MxM/Y0[5] ), .Z(n39) );
  XNOR U135 ( .A(n96), .B(n97), .Z(n91) );
  AND U136 ( .A(n74), .B(n99), .Z(n98) );
  XOR U137 ( .A(n86), .B(n100), .Z(n99) );
  XOR U138 ( .A(n100), .B(n87), .Z(n86) );
  OR U139 ( .A(n101), .B(n102), .Z(n87) );
  IV U140 ( .A(n97), .Z(n100) );
  XNOR U141 ( .A(n85), .B(n84), .Z(n97) );
  OR U142 ( .A(n103), .B(n104), .Z(n84) );
  AND U143 ( .A(n105), .B(n106), .Z(n85) );
  XNOR U144 ( .A(n107), .B(n108), .Z(n106) );
  ANDN U145 ( .A(n109), .B(n110), .Z(n108) );
  XOR U146 ( .A(n107), .B(n111), .Z(n109) );
  XNOR U147 ( .A(n78), .B(n112), .Z(n105) );
  NAND U148 ( .A(n114), .B(n115), .Z(n79) );
  NANDN U149 ( .B(n116), .A(n117), .Z(n114) );
  NANDN U150 ( .B(n82), .A(n118), .Z(n113) );
  NANDN U151 ( .B(n83), .A(n119), .Z(n78) );
  XOR U152 ( .A(n120), .B(n121), .Z(n88) );
  ANDN U153 ( .A(n122), .B(n123), .Z(n121) );
  XNOR U154 ( .A(\_MxM/Y0[4] ), .B(n120), .Z(n122) );
  NAND U155 ( .A(n124), .B(n125), .Z(\_MxM/n114 ) );
  NANDN U156 ( .B(n26), .A(o[3]), .Z(n125) );
  AND U157 ( .A(n126), .B(n127), .Z(n124) );
  NANDN U158 ( .B(n49), .A(o[3]), .Z(n127) );
  NANDN U159 ( .B(n54), .A(n36), .Z(n126) );
  XNOR U160 ( .A(n123), .B(\_MxM/Y0[4] ), .Z(n36) );
  XNOR U161 ( .A(n128), .B(n129), .Z(n123) );
  AND U162 ( .A(n74), .B(n131), .Z(n130) );
  XOR U163 ( .A(n101), .B(n132), .Z(n131) );
  XOR U164 ( .A(n132), .B(n102), .Z(n101) );
  OR U165 ( .A(n133), .B(n134), .Z(n102) );
  IV U166 ( .A(n129), .Z(n132) );
  XNOR U167 ( .A(n104), .B(n103), .Z(n129) );
  OR U168 ( .A(n135), .B(n136), .Z(n103) );
  XOR U169 ( .A(n111), .B(n110), .Z(n104) );
  XOR U170 ( .A(n107), .B(n137), .Z(n110) );
  AND U171 ( .A(n138), .B(n139), .Z(n137) );
  NANDN U172 ( .B(n82), .A(n140), .Z(n139) );
  OR U173 ( .A(n141), .B(n142), .Z(n138) );
  XOR U174 ( .A(n116), .B(n117), .Z(n111) );
  NANDN U175 ( .B(n83), .A(n146), .Z(n117) );
  XNOR U176 ( .A(n115), .B(n147), .Z(n116) );
  AND U177 ( .A(n119), .B(n118), .Z(n147) );
  ANDN U178 ( .A(n148), .B(n149), .Z(n115) );
  NANDN U179 ( .B(n150), .A(n151), .Z(n148) );
  NAND U180 ( .A(n154), .B(n155), .Z(\_MxM/n113 ) );
  NANDN U181 ( .B(n26), .A(o[2]), .Z(n155) );
  AND U182 ( .A(n156), .B(n157), .Z(n154) );
  NANDN U183 ( .B(n49), .A(o[2]), .Z(n157) );
  NANDN U184 ( .B(n54), .A(n33), .Z(n156) );
  XNOR U185 ( .A(n153), .B(\_MxM/Y0[3] ), .Z(n33) );
  XNOR U186 ( .A(n158), .B(n159), .Z(n153) );
  AND U187 ( .A(n74), .B(n161), .Z(n160) );
  XOR U188 ( .A(n133), .B(n162), .Z(n161) );
  XOR U189 ( .A(n162), .B(n134), .Z(n133) );
  OR U190 ( .A(n163), .B(n164), .Z(n134) );
  IV U191 ( .A(n159), .Z(n162) );
  XOR U192 ( .A(n145), .B(n144), .Z(n135) );
  XNOR U193 ( .A(n168), .B(n169), .Z(n144) );
  IV U194 ( .A(n143), .Z(n169) );
  XOR U195 ( .A(n170), .B(n171), .Z(n143) );
  ANDN U196 ( .A(n172), .B(n173), .Z(n171) );
  XOR U197 ( .A(n170), .B(n174), .Z(n172) );
  XNOR U198 ( .A(n175), .B(n141), .Z(n168) );
  NAND U199 ( .A(n140), .B(n119), .Z(n141) );
  NANDN U200 ( .B(n82), .A(n177), .Z(n176) );
  XNOR U201 ( .A(n178), .B(n179), .Z(n142) );
  ANDN U202 ( .A(n180), .B(n181), .Z(n179) );
  XNOR U203 ( .A(n182), .B(n178), .Z(n180) );
  XOR U204 ( .A(n150), .B(n151), .Z(n145) );
  OR U205 ( .A(n183), .B(n83), .Z(n151) );
  XNOR U206 ( .A(n184), .B(n185), .Z(n150) );
  AND U207 ( .A(n146), .B(n118), .Z(n185) );
  IV U208 ( .A(n149), .Z(n184) );
  NAND U209 ( .A(n186), .B(n187), .Z(n149) );
  NANDN U210 ( .B(n188), .A(n189), .Z(n186) );
  NAND U211 ( .A(n192), .B(n193), .Z(\_MxM/n112 ) );
  NANDN U212 ( .B(n26), .A(o[1]), .Z(n193) );
  AND U213 ( .A(n194), .B(n195), .Z(n192) );
  NANDN U214 ( .B(n49), .A(o[1]), .Z(n195) );
  NANDN U215 ( .B(n54), .A(n29), .Z(n194) );
  XNOR U216 ( .A(n191), .B(\_MxM/Y0[2] ), .Z(n29) );
  XNOR U217 ( .A(n196), .B(n197), .Z(n191) );
  XOR U218 ( .A(n190), .B(n198), .Z(n196) );
  AND U219 ( .A(n74), .B(n199), .Z(n198) );
  XOR U220 ( .A(n163), .B(n200), .Z(n199) );
  XOR U221 ( .A(n200), .B(n164), .Z(n163) );
  NANDN U222 ( .B(n201), .A(n202), .Z(n164) );
  IV U223 ( .A(n197), .Z(n200) );
  XOR U224 ( .A(n167), .B(n166), .Z(n197) );
  XNOR U225 ( .A(n165), .B(n203), .Z(n166) );
  AND U226 ( .A(n204), .B(n205), .Z(n203) );
  OR U227 ( .A(n206), .B(n207), .Z(n205) );
  AND U228 ( .A(n208), .B(n209), .Z(n204) );
  NANDN U229 ( .B(n82), .A(n210), .Z(n209) );
  NAND U230 ( .A(n211), .B(n212), .Z(n208) );
  XNOR U231 ( .A(n178), .B(n217), .Z(n181) );
  AND U232 ( .A(n119), .B(n177), .Z(n217) );
  XOR U233 ( .A(n218), .B(n219), .Z(n178) );
  ANDN U234 ( .A(n220), .B(n221), .Z(n219) );
  XNOR U235 ( .A(n222), .B(n218), .Z(n220) );
  XOR U236 ( .A(n223), .B(n182), .Z(n216) );
  NAND U237 ( .A(n140), .B(n146), .Z(n182) );
  IV U238 ( .A(n170), .Z(n223) );
  XOR U239 ( .A(n224), .B(n225), .Z(n170) );
  ANDN U240 ( .A(n226), .B(n227), .Z(n225) );
  XOR U241 ( .A(n224), .B(n228), .Z(n226) );
  XNOR U242 ( .A(n188), .B(n189), .Z(n174) );
  OR U243 ( .A(n229), .B(n83), .Z(n189) );
  XNOR U244 ( .A(n187), .B(n230), .Z(n188) );
  ANDN U245 ( .A(n118), .B(n183), .Z(n230) );
  ANDN U246 ( .A(n231), .B(n232), .Z(n187) );
  NANDN U247 ( .B(n233), .A(n234), .Z(n231) );
  NAND U248 ( .A(n237), .B(n238), .Z(\_MxM/n111 ) );
  NANDN U249 ( .B(n26), .A(o[0]), .Z(n238) );
  AND U250 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U251 ( .B(n49), .A(o[0]), .Z(n240) );
  IV U252 ( .A(n241), .Z(n49) );
  OR U253 ( .A(n54), .B(n24), .Z(n239) );
  IV U254 ( .A(\_MxM/Y0[1] ), .Z(n30) );
  XOR U255 ( .A(n242), .B(n243), .Z(n236) );
  XNOR U256 ( .A(n244), .B(n235), .Z(n242) );
  NAND U257 ( .A(\_MxM/Y0[0] ), .B(n201), .Z(n235) );
  NAND U258 ( .A(n245), .B(n74), .Z(n244) );
  XOR U259 ( .A(e_input[7]), .B(g_input[7]), .Z(n74) );
  XNOR U260 ( .A(n202), .B(n243), .Z(n245) );
  XNOR U261 ( .A(n201), .B(n243), .Z(n202) );
  XNOR U262 ( .A(n215), .B(n214), .Z(n243) );
  XNOR U263 ( .A(n246), .B(n211), .Z(n214) );
  XNOR U264 ( .A(n247), .B(n206), .Z(n211) );
  NAND U265 ( .A(n119), .B(n210), .Z(n206) );
  NANDN U266 ( .B(n82), .A(n249), .Z(n248) );
  XNOR U267 ( .A(n212), .B(n213), .Z(n246) );
  XNOR U268 ( .A(n218), .B(n260), .Z(n221) );
  AND U269 ( .A(n146), .B(n177), .Z(n260) );
  XOR U270 ( .A(n261), .B(n262), .Z(n218) );
  ANDN U271 ( .A(n263), .B(n264), .Z(n262) );
  XNOR U272 ( .A(n265), .B(n261), .Z(n263) );
  XOR U273 ( .A(n266), .B(n222), .Z(n259) );
  NANDN U274 ( .B(n183), .A(n140), .Z(n222) );
  IV U275 ( .A(n224), .Z(n266) );
  XNOR U276 ( .A(n233), .B(n234), .Z(n228) );
  NANDN U277 ( .B(n83), .A(n270), .Z(n234) );
  ANDN U278 ( .A(n118), .B(n229), .Z(n271) );
  NAND U279 ( .A(n272), .B(n273), .Z(n232) );
  NANDN U280 ( .B(n274), .A(n275), .Z(n272) );
  XNOR U281 ( .A(n255), .B(n254), .Z(n201) );
  XNOR U282 ( .A(n276), .B(n258), .Z(n254) );
  XNOR U283 ( .A(n251), .B(n252), .Z(n258) );
  NAND U284 ( .A(n146), .B(n210), .Z(n252) );
  XNOR U285 ( .A(n250), .B(n277), .Z(n251) );
  AND U286 ( .A(n249), .B(n119), .Z(n277) );
  XOR U287 ( .A(n278), .B(n279), .Z(n250) );
  AND U288 ( .A(n280), .B(n281), .Z(n279) );
  XNOR U289 ( .A(n282), .B(n278), .Z(n281) );
  XNOR U290 ( .A(n257), .B(n253), .Z(n276) );
  XOR U291 ( .A(n283), .B(n284), .Z(n253) );
  XOR U292 ( .A(n285), .B(n286), .Z(n257) );
  AND U293 ( .A(n287), .B(n288), .Z(n286) );
  NANDN U294 ( .B(n82), .A(n289), .Z(n288) );
  NANDN U295 ( .B(n290), .A(n291), .Z(n82) );
  AND U296 ( .A(n292), .B(g_input[7]), .Z(n291) );
  NANDN U297 ( .B(n293), .A(n294), .Z(n287) );
  IV U298 ( .A(n256), .Z(n285) );
  XNOR U299 ( .A(n295), .B(n296), .Z(n256) );
  AND U300 ( .A(n297), .B(n298), .Z(n296) );
  XOR U301 ( .A(n294), .B(n299), .Z(n298) );
  XNOR U302 ( .A(n293), .B(n295), .Z(n299) );
  NAND U303 ( .A(n119), .B(n289), .Z(n293) );
  XNOR U304 ( .A(n303), .B(n300), .Z(n302) );
  XOR U305 ( .A(n280), .B(n304), .Z(n297) );
  XNOR U306 ( .A(n282), .B(n295), .Z(n304) );
  NANDN U307 ( .B(n183), .A(n210), .Z(n282) );
  XOR U308 ( .A(n278), .B(n305), .Z(n280) );
  AND U309 ( .A(n249), .B(n146), .Z(n305) );
  XOR U310 ( .A(n306), .B(n307), .Z(n278) );
  AND U311 ( .A(n308), .B(n309), .Z(n307) );
  XNOR U312 ( .A(n310), .B(n306), .Z(n309) );
  XOR U313 ( .A(n311), .B(n312), .Z(n295) );
  AND U314 ( .A(n313), .B(n314), .Z(n312) );
  XOR U315 ( .A(n301), .B(n315), .Z(n314) );
  XNOR U316 ( .A(n303), .B(n311), .Z(n315) );
  NAND U317 ( .A(n146), .B(n289), .Z(n303) );
  XOR U318 ( .A(n300), .B(n316), .Z(n301) );
  AND U319 ( .A(n119), .B(e_input[0]), .Z(n316) );
  XNOR U320 ( .A(n292), .B(g_input[6]), .Z(n290) );
  NOR U321 ( .A(n317), .B(n318), .Z(n292) );
  XNOR U322 ( .A(n322), .B(n319), .Z(n321) );
  XOR U323 ( .A(n308), .B(n323), .Z(n313) );
  XNOR U324 ( .A(n310), .B(n311), .Z(n323) );
  NANDN U325 ( .B(n229), .A(n210), .Z(n310) );
  XOR U326 ( .A(n306), .B(n324), .Z(n308) );
  ANDN U327 ( .A(n249), .B(n183), .Z(n324) );
  XOR U328 ( .A(n325), .B(n326), .Z(n306) );
  AND U329 ( .A(n327), .B(n328), .Z(n326) );
  XNOR U330 ( .A(n329), .B(n325), .Z(n328) );
  XOR U331 ( .A(n330), .B(n331), .Z(n311) );
  AND U332 ( .A(n332), .B(n333), .Z(n331) );
  XOR U333 ( .A(n320), .B(n334), .Z(n333) );
  XNOR U334 ( .A(n322), .B(n330), .Z(n334) );
  NANDN U335 ( .B(n183), .A(n289), .Z(n322) );
  XOR U336 ( .A(n319), .B(n335), .Z(n320) );
  AND U337 ( .A(n146), .B(e_input[0]), .Z(n335) );
  XOR U338 ( .A(n317), .B(g_input[5]), .Z(n318) );
  NANDN U339 ( .B(n336), .A(n337), .Z(n317) );
  XOR U340 ( .A(n338), .B(n339), .Z(n319) );
  ANDN U341 ( .A(n340), .B(n341), .Z(n339) );
  XNOR U342 ( .A(n342), .B(n338), .Z(n340) );
  XOR U343 ( .A(n327), .B(n343), .Z(n332) );
  XNOR U344 ( .A(n329), .B(n330), .Z(n343) );
  NAND U345 ( .A(n210), .B(n270), .Z(n329) );
  XOR U346 ( .A(n325), .B(n344), .Z(n327) );
  ANDN U347 ( .A(n249), .B(n229), .Z(n344) );
  XOR U348 ( .A(n345), .B(n346), .Z(n325) );
  ANDN U349 ( .A(n347), .B(n348), .Z(n346) );
  XNOR U350 ( .A(n349), .B(n345), .Z(n347) );
  XNOR U351 ( .A(n351), .B(n349), .Z(n283) );
  NAND U352 ( .A(n210), .B(n352), .Z(n349) );
  IV U353 ( .A(n348), .Z(n351) );
  XNOR U354 ( .A(n345), .B(n353), .Z(n348) );
  AND U355 ( .A(n270), .B(n249), .Z(n353) );
  AND U356 ( .A(n354), .B(g_input[0]), .Z(n345) );
  NANDN U357 ( .B(n210), .A(n355), .Z(n354) );
  NAND U358 ( .A(n352), .B(n249), .Z(n355) );
  XNOR U359 ( .A(n356), .B(e_input[2]), .Z(n249) );
  NAND U360 ( .A(n357), .B(e_input[7]), .Z(n356) );
  XOR U361 ( .A(n358), .B(e_input[2]), .Z(n357) );
  XNOR U362 ( .A(n338), .B(n361), .Z(n341) );
  ANDN U363 ( .A(e_input[0]), .B(n183), .Z(n361) );
  XOR U364 ( .A(n362), .B(n363), .Z(n338) );
  AND U365 ( .A(n364), .B(n365), .Z(n363) );
  XOR U366 ( .A(n366), .B(n362), .Z(n365) );
  ANDN U367 ( .A(e_input[0]), .B(n229), .Z(n366) );
  XOR U368 ( .A(n367), .B(n362), .Z(n364) );
  AND U369 ( .A(n289), .B(n270), .Z(n367) );
  XOR U370 ( .A(n368), .B(n369), .Z(n362) );
  ANDN U371 ( .A(n370), .B(n371), .Z(n369) );
  XNOR U372 ( .A(n372), .B(n368), .Z(n370) );
  XOR U373 ( .A(n373), .B(n342), .Z(n360) );
  NANDN U374 ( .B(n229), .A(n289), .Z(n342) );
  IV U375 ( .A(n350), .Z(n373) );
  NAND U376 ( .A(n289), .B(n352), .Z(n372) );
  XNOR U377 ( .A(n368), .B(n374), .Z(n371) );
  AND U378 ( .A(n270), .B(e_input[0]), .Z(n374) );
  AND U379 ( .A(n375), .B(g_input[0]), .Z(n368) );
  NANDN U380 ( .B(n289), .A(n376), .Z(n375) );
  NAND U381 ( .A(n352), .B(e_input[0]), .Z(n376) );
  XNOR U382 ( .A(n377), .B(e_input[1]), .Z(n289) );
  NAND U383 ( .A(n378), .B(e_input[7]), .Z(n377) );
  XNOR U384 ( .A(e_input[1]), .B(n379), .Z(n378) );
  XOR U385 ( .A(n380), .B(n381), .Z(n268) );
  IV U386 ( .A(n264), .Z(n381) );
  XNOR U387 ( .A(n261), .B(n382), .Z(n264) );
  ANDN U388 ( .A(n177), .B(n183), .Z(n382) );
  XNOR U389 ( .A(n337), .B(g_input[4]), .Z(n336) );
  NOR U390 ( .A(n383), .B(n384), .Z(n337) );
  XOR U391 ( .A(n387), .B(n385), .Z(n386) );
  ANDN U392 ( .A(n177), .B(n229), .Z(n387) );
  AND U393 ( .A(n270), .B(n140), .Z(n388) );
  XOR U394 ( .A(n392), .B(n265), .Z(n380) );
  NANDN U395 ( .B(n229), .A(n140), .Z(n265) );
  NANDN U396 ( .B(n393), .A(n394), .Z(n383) );
  IV U397 ( .A(n267), .Z(n392) );
  XOR U398 ( .A(n395), .B(n391), .Z(n267) );
  NAND U399 ( .A(n140), .B(n352), .Z(n391) );
  IV U400 ( .A(n390), .Z(n395) );
  XNOR U401 ( .A(n389), .B(n396), .Z(n390) );
  AND U402 ( .A(n270), .B(n177), .Z(n396) );
  AND U403 ( .A(n397), .B(g_input[0]), .Z(n389) );
  NANDN U404 ( .B(n140), .A(n398), .Z(n397) );
  NAND U405 ( .A(n352), .B(n177), .Z(n398) );
  XNOR U406 ( .A(n399), .B(e_input[4]), .Z(n177) );
  NAND U407 ( .A(n400), .B(e_input[7]), .Z(n399) );
  XOR U408 ( .A(n401), .B(e_input[4]), .Z(n400) );
  XNOR U409 ( .A(n402), .B(e_input[5]), .Z(n140) );
  NAND U410 ( .A(n403), .B(e_input[7]), .Z(n402) );
  XOR U411 ( .A(n404), .B(e_input[5]), .Z(n403) );
  XNOR U412 ( .A(n274), .B(n275), .Z(n269) );
  NANDN U413 ( .B(n83), .A(n352), .Z(n275) );
  XNOR U414 ( .A(n273), .B(n405), .Z(n274) );
  AND U415 ( .A(n270), .B(n118), .Z(n405) );
  XNOR U416 ( .A(n394), .B(g_input[2]), .Z(n393) );
  AND U417 ( .A(n407), .B(g_input[0]), .Z(n273) );
  NAND U418 ( .A(n408), .B(n83), .Z(n407) );
  NANDN U419 ( .B(n409), .A(n410), .Z(n83) );
  ANDN U420 ( .A(e_input[7]), .B(n411), .Z(n410) );
  NAND U421 ( .A(n352), .B(n118), .Z(n408) );
  XOR U422 ( .A(n411), .B(e_input[6]), .Z(n409) );
  OR U423 ( .A(n404), .B(n412), .Z(n411) );
  XOR U424 ( .A(n412), .B(e_input[5]), .Z(n404) );
  OR U425 ( .A(n401), .B(n413), .Z(n412) );
  XOR U426 ( .A(n413), .B(e_input[4]), .Z(n401) );
  OR U427 ( .A(n359), .B(n414), .Z(n413) );
  XOR U428 ( .A(n414), .B(e_input[3]), .Z(n359) );
  OR U429 ( .A(n358), .B(n415), .Z(n414) );
  XOR U430 ( .A(n415), .B(e_input[2]), .Z(n358) );
  NANDN U431 ( .B(e_input[0]), .A(n379), .Z(n415) );
  XNOR U432 ( .A(e_input[0]), .B(e_input[1]), .Z(n379) );
  XNOR U433 ( .A(n416), .B(g_input[1]), .Z(n352) );
  NAND U434 ( .A(n417), .B(g_input[7]), .Z(n416) );
  XOR U435 ( .A(g_input[1]), .B(n406), .Z(n417) );
  XOR U436 ( .A(g_input[0]), .B(g_input[1]), .Z(n406) );
  NANDN U437 ( .B(n241), .A(n26), .Z(n54) );
  IV U438 ( .A(rst), .Z(n26) );
  NAND U439 ( .A(n418), .B(n419), .Z(n241) );
  ANDN U440 ( .A(n420), .B(\_MxM/n[2] ), .Z(n419) );
  NOR U441 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n420) );
  ANDN U442 ( .A(n421), .B(n20), .Z(n418) );
  OR U443 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n20) );
  NOR U444 ( .A(\_MxM/n[0] ), .B(\_MxM/n[1] ), .Z(n421) );
endmodule

