
module MAC_TG_N16 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MAC/_MULT/X__[0] , \_MAC/_MULT/A__[0] , n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366;
  wire   [15:0] o_reg;
  assign \_MAC/_MULT/X__[0]  = e_input[0];
  assign \_MAC/_MULT/A__[0]  = g_input[0];

  DFF \o_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[0])
         );
  DFF \o_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[1])
         );
  DFF \o_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[2])
         );
  DFF \o_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[3])
         );
  DFF \o_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[4])
         );
  DFF \o_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[5])
         );
  DFF \o_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[6])
         );
  DFF \o_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[7])
         );
  DFF \o_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[8])
         );
  DFF \o_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[9])
         );
  DFF \o_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[10]) );
  DFF \o_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[11]) );
  DFF \o_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[12]) );
  DFF \o_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[13]) );
  DFF \o_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[14]) );
  DFF \o_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[15]) );
  MUX U19 ( .IN0(n1273), .IN1(n1291), .SEL(n1275), .F(n1254) );
  XOR U20 ( .A(n837), .B(n838), .Z(n849) );
  MUX U21 ( .IN0(n17), .IN1(n818), .SEL(n819), .F(n786) );
  IV U22 ( .A(n820), .Z(n17) );
  XOR U23 ( .A(n1040), .B(n1030), .Z(n831) );
  MUX U24 ( .IN0(n18), .IN1(n1025), .SEL(n1026), .F(n801) );
  IV U25 ( .A(n1027), .Z(n18) );
  MUX U26 ( .IN0(e_input[8]), .IN1(n1321), .SEL(e_input[15]), .F(n466) );
  MUX U27 ( .IN0(n19), .IN1(n770), .SEL(n771), .F(n679) );
  IV U28 ( .A(n772), .Z(n19) );
  XOR U29 ( .A(n1038), .B(n1039), .Z(n854) );
  MUX U30 ( .IN0(n988), .IN1(n991), .SEL(n989), .F(n973) );
  MUX U31 ( .IN0(n20), .IN1(n794), .SEL(n795), .F(n733) );
  IV U32 ( .A(n796), .Z(n20) );
  MUX U33 ( .IN0(n21), .IN1(n456), .SEL(n457), .F(n440) );
  IV U34 ( .A(n458), .Z(n21) );
  MUX U35 ( .IN0(e_input[9]), .IN1(n1322), .SEL(e_input[15]), .F(n446) );
  XNOR U36 ( .A(n1336), .B(n1337), .Z(n774) );
  MUX U37 ( .IN0(n1031), .IN1(n22), .SEL(n1030), .F(n1020) );
  IV U38 ( .A(n1029), .Z(n22) );
  XOR U39 ( .A(n1127), .B(n1116), .Z(n961) );
  MUX U40 ( .IN0(n1179), .IN1(n1195), .SEL(n1181), .F(n1162) );
  MUX U41 ( .IN0(n1254), .IN1(n1272), .SEL(n1256), .F(n1223) );
  MUX U42 ( .IN0(n23), .IN1(n813), .SEL(n814), .F(n794) );
  IV U43 ( .A(n815), .Z(n23) );
  MUX U44 ( .IN0(n24), .IN1(n500), .SEL(n501), .F(n480) );
  IV U45 ( .A(n502), .Z(n24) );
  MUX U46 ( .IN0(n25), .IN1(n381), .SEL(n382), .F(n364) );
  IV U47 ( .A(n383), .Z(n25) );
  MUX U48 ( .IN0(g_input[10]), .IN1(n1092), .SEL(g_input[15]), .F(n493) );
  MUX U49 ( .IN0(n578), .IN1(n26), .SEL(n576), .F(n189) );
  IV U50 ( .A(n643), .Z(n26) );
  MUX U51 ( .IN0(n1173), .IN1(n1188), .SEL(n1175), .F(n1156) );
  MUX U52 ( .IN0(n27), .IN1(n786), .SEL(n787), .F(n725) );
  IV U53 ( .A(n788), .Z(n27) );
  MUX U54 ( .IN0(n28), .IN1(n495), .SEL(n496), .F(n475) );
  IV U55 ( .A(n497), .Z(n28) );
  MUX U56 ( .IN0(n29), .IN1(n369), .SEL(n370), .F(n348) );
  IV U57 ( .A(n371), .Z(n29) );
  MUX U58 ( .IN0(g_input[7]), .IN1(n1232), .SEL(g_input[15]), .F(n551) );
  MUX U59 ( .IN0(n30), .IN1(n801), .SEL(n802), .F(n743) );
  IV U60 ( .A(n803), .Z(n30) );
  MUX U61 ( .IN0(n435), .IN1(n581), .SEL(n436), .F(n572) );
  MUX U62 ( .IN0(n469), .IN1(n31), .SEL(n468), .F(n448) );
  IV U63 ( .A(n467), .Z(n31) );
  XNOR U64 ( .A(n1323), .B(n771), .Z(n775) );
  MUX U65 ( .IN0(n132), .IN1(n126), .SEL(n124), .F(n32) );
  IV U66 ( .A(n32), .Z(n129) );
  MUX U67 ( .IN0(n981), .IN1(n979), .SEL(n980), .F(n952) );
  MUX U68 ( .IN0(n33), .IN1(n1213), .SEL(n1214), .F(n1209) );
  IV U69 ( .A(n1215), .Z(n33) );
  XOR U70 ( .A(n814), .B(n815), .Z(n824) );
  MUX U71 ( .IN0(n1223), .IN1(n1253), .SEL(n1225), .F(n753) );
  MUX U72 ( .IN0(n34), .IN1(n558), .SEL(n559), .F(n538) );
  IV U73 ( .A(n560), .Z(n34) );
  MUX U74 ( .IN0(g_input[11]), .IN1(n1078), .SEL(g_input[15]), .F(n388) );
  XOR U75 ( .A(n802), .B(n803), .Z(n808) );
  MUX U76 ( .IN0(n489), .IN1(n602), .SEL(n490), .F(n595) );
  MUX U77 ( .IN0(n366), .IN1(n35), .SEL(n365), .F(n343) );
  IV U78 ( .A(n364), .Z(n35) );
  NAND U79 ( .A(n189), .B(n641), .Z(n640) );
  MUX U80 ( .IN0(n148), .IN1(n134), .SEL(n124), .F(n36) );
  IV U81 ( .A(n36), .Z(n145) );
  XOR U82 ( .A(n1090), .B(n1080), .Z(n909) );
  MUX U83 ( .IN0(n1139), .IN1(n1161), .SEL(n1141), .F(n1122) );
  MUX U84 ( .IN0(g_input[1]), .IN1(n1349), .SEL(g_input[15]), .F(n998) );
  XOR U85 ( .A(n839), .B(n819), .Z(n823) );
  XOR U86 ( .A(n795), .B(n796), .Z(n792) );
  MUX U87 ( .IN0(n37), .IN1(n553), .SEL(n554), .F(n533) );
  IV U88 ( .A(n555), .Z(n37) );
  MUX U89 ( .IN0(n38), .IN1(n761), .SEL(n762), .F(n558) );
  IV U90 ( .A(n763), .Z(n38) );
  MUX U91 ( .IN0(g_input[2]), .IN1(n1339), .SEL(g_input[15]), .F(n777) );
  MUX U92 ( .IN0(g_input[12]), .IN1(n1058), .SEL(g_input[15]), .F(n367) );
  MUX U93 ( .IN0(n486), .IN1(n488), .SEL(n487), .F(n460) );
  MUX U94 ( .IN0(n507), .IN1(n609), .SEL(n508), .F(n602) );
  XNOR U95 ( .A(n575), .B(n576), .Z(n423) );
  MUX U96 ( .IN0(n176), .IN1(n151), .SEL(n124), .F(n39) );
  IV U97 ( .A(n39), .Z(n173) );
  MUX U98 ( .IN0(n40), .IN1(n1079), .SEL(n1080), .F(n1060) );
  IV U99 ( .A(n1081), .Z(n40) );
  MUX U100 ( .IN0(n41), .IN1(n725), .SEL(n726), .F(n381) );
  IV U101 ( .A(n727), .Z(n41) );
  XOR U102 ( .A(n1303), .B(n1288), .Z(n1228) );
  MUX U103 ( .IN0(e_input[11]), .IN1(n1302), .SEL(e_input[15]), .F(n419) );
  XOR U104 ( .A(n695), .B(n696), .Z(n600) );
  MUX U105 ( .IN0(e_input[6]), .IN1(n1007), .SEL(e_input[15]), .F(n327) );
  MUX U106 ( .IN0(n547), .IN1(n623), .SEL(n548), .F(n616) );
  MUX U107 ( .IN0(n745), .IN1(n42), .SEL(n744), .F(n397) );
  IV U108 ( .A(n743), .Z(n42) );
  XNOR U109 ( .A(n582), .B(n583), .Z(n436) );
  MUX U110 ( .IN0(n43), .IN1(n491), .SEL(n320), .F(n472) );
  IV U111 ( .A(n319), .Z(n43) );
  MUX U112 ( .IN0(n263), .IN1(n179), .SEL(n124), .F(n44) );
  IV U113 ( .A(n44), .Z(n198) );
  MUX U114 ( .IN0(n1156), .IN1(n1172), .SEL(n1158), .F(n1145) );
  MUX U115 ( .IN0(e_input[4]), .IN1(n1002), .SEL(e_input[15]), .F(n363) );
  MUX U116 ( .IN0(n45), .IN1(n733), .SEL(n734), .F(n390) );
  IV U117 ( .A(n735), .Z(n45) );
  MUX U118 ( .IN0(n46), .IN1(n440), .SEL(n441), .F(n429) );
  IV U119 ( .A(n442), .Z(n46) );
  MUX U120 ( .IN0(n524), .IN1(n526), .SEL(n525), .F(n504) );
  MUX U121 ( .IN0(n346), .IN1(n47), .SEL(n345), .F(n322) );
  IV U122 ( .A(n344), .Z(n47) );
  MUX U123 ( .IN0(n565), .IN1(n630), .SEL(n566), .F(n623) );
  XOR U124 ( .A(n744), .B(n745), .Z(n750) );
  XNOR U125 ( .A(n432), .B(n443), .Z(n433) );
  XNOR U126 ( .A(n589), .B(n590), .Z(n452) );
  MUX U127 ( .IN0(n48), .IN1(n509), .SEL(n336), .F(n491) );
  IV U128 ( .A(n335), .Z(n48) );
  XOR U129 ( .A(n199), .B(n202), .Z(n200) );
  MUX U130 ( .IN0(n1209), .IN1(n1212), .SEL(n1210), .F(n1189) );
  XOR U131 ( .A(n1026), .B(n1027), .Z(n829) );
  MUX U132 ( .IN0(n49), .IN1(n533), .SEL(n534), .F(n513) );
  IV U133 ( .A(n535), .Z(n49) );
  MUX U134 ( .IN0(n50), .IN1(n348), .SEL(n349), .F(n328) );
  IV U135 ( .A(n350), .Z(n50) );
  MUX U136 ( .IN0(e_input[5]), .IN1(n1003), .SEL(e_input[15]), .F(n341) );
  MUX U137 ( .IN0(n387), .IN1(n385), .SEL(n386), .F(n358) );
  MUX U138 ( .IN0(n639), .IN1(n637), .SEL(n638), .F(n630) );
  MUX U139 ( .IN0(n562), .IN1(n564), .SEL(n563), .F(n544) );
  XOR U140 ( .A(n195), .B(n684), .Z(n196) );
  XNOR U141 ( .A(n596), .B(n597), .Z(n471) );
  XOR U142 ( .A(n459), .B(n96), .Z(n449) );
  MUX U143 ( .IN0(n51), .IN1(n529), .SEL(n355), .F(n509) );
  IV U144 ( .A(n354), .Z(n51) );
  MUX U145 ( .IN0(n318), .IN1(n282), .SEL(n283), .F(n52) );
  IV U146 ( .A(n52), .Z(n302) );
  XOR U147 ( .A(n206), .B(n209), .Z(n207) );
  XOR U148 ( .A(n1072), .B(n1073), .Z(n907) );
  XOR U149 ( .A(n1028), .B(n1020), .Z(n810) );
  XNOR U150 ( .A(n995), .B(n996), .Z(n979) );
  MUX U151 ( .IN0(n53), .IN1(n475), .SEL(n476), .F(n456) );
  IV U152 ( .A(n477), .Z(n53) );
  MUX U153 ( .IN0(g_input[6]), .IN1(n1245), .SEL(g_input[15]), .F(n673) );
  MUX U154 ( .IN0(g_input[3]), .IN1(n1326), .SEL(g_input[15]), .F(n54) );
  IV U155 ( .A(n54), .Z(n712) );
  MUX U156 ( .IN0(g_input[5]), .IN1(n1265), .SEL(g_input[15]), .F(n678) );
  MUX U157 ( .IN0(g_input[4]), .IN1(n1283), .SEL(g_input[15]), .F(n55) );
  IV U158 ( .A(n55), .Z(n708) );
  MUX U159 ( .IN0(n790), .IN1(n56), .SEL(n791), .F(n729) );
  IV U160 ( .A(n792), .Z(n56) );
  MUX U161 ( .IN0(n504), .IN1(n506), .SEL(n505), .F(n486) );
  MUX U162 ( .IN0(n776), .IN1(n774), .SEL(n775), .F(n637) );
  XOR U163 ( .A(n1229), .B(n762), .Z(n766) );
  MUX U164 ( .IN0(g_input[13]), .IN1(n1043), .SEL(g_input[15]), .F(n192) );
  MUX U165 ( .IN0(n57), .IN1(n424), .SEL(n299), .F(n411) );
  IV U166 ( .A(n298), .Z(n57) );
  XNOR U167 ( .A(n603), .B(n604), .Z(n490) );
  MUX U168 ( .IN0(n58), .IN1(n549), .SEL(n377), .F(n529) );
  IV U169 ( .A(n376), .Z(n58) );
  NAND U170 ( .A(n343), .B(n362), .Z(n361) );
  MUX U171 ( .IN0(n334), .IN1(n280), .SEL(n281), .F(n318) );
  MUX U172 ( .IN0(n59), .IN1(n240), .SEL(n115), .F(n233) );
  IV U173 ( .A(o_reg[4]), .Z(n59) );
  XOR U174 ( .A(n213), .B(n216), .Z(n214) );
  MUX U175 ( .IN0(n60), .IN1(n1009), .SEL(n1010), .F(n1183) );
  IV U176 ( .A(n1201), .Z(n60) );
  MUX U177 ( .IN0(n61), .IN1(n1044), .SEL(n1045), .F(n1029) );
  IV U178 ( .A(n1046), .Z(n61) );
  XOR U179 ( .A(n1125), .B(n1126), .Z(n984) );
  MUX U180 ( .IN0(n451), .IN1(n588), .SEL(n452), .F(n581) );
  XOR U181 ( .A(n701), .B(n702), .Z(n614) );
  MUX U182 ( .IN0(n544), .IN1(n546), .SEL(n545), .F(n524) );
  XNOR U183 ( .A(n784), .B(n726), .Z(n730) );
  NAND U184 ( .A(n416), .B(n427), .Z(n426) );
  MUX U185 ( .IN0(e_input[7]), .IN1(n1008), .SEL(e_input[15]), .F(n309) );
  XOR U186 ( .A(n478), .B(n468), .Z(n461) );
  XNOR U187 ( .A(n610), .B(n611), .Z(n508) );
  MUX U188 ( .IN0(n405), .IN1(n62), .SEL(n404), .F(n372) );
  IV U189 ( .A(n403), .Z(n62) );
  MUX U190 ( .IN0(n63), .IN1(n567), .SEL(n568), .F(n549) );
  IV U191 ( .A(n569), .Z(n63) );
  MUX U192 ( .IN0(n64), .IN1(n278), .SEL(n279), .F(n334) );
  IV U193 ( .A(n353), .Z(n64) );
  MUX U194 ( .IN0(n65), .IN1(n247), .SEL(n116), .F(n240) );
  IV U195 ( .A(o_reg[3]), .Z(n65) );
  XOR U196 ( .A(n221), .B(n286), .Z(n112) );
  MUX U197 ( .IN0(n66), .IN1(n982), .SEL(n798), .F(n955) );
  IV U198 ( .A(n797), .Z(n66) );
  MUX U199 ( .IN0(n1145), .IN1(n1155), .SEL(n1147), .F(n1131) );
  MUX U200 ( .IN0(e_input[10]), .IN1(n1301), .SEL(e_input[15]), .F(n428) );
  XOR U201 ( .A(n689), .B(n690), .Z(n586) );
  MUX U202 ( .IN0(e_input[3]), .IN1(n1206), .SEL(e_input[15]), .F(n400) );
  MUX U203 ( .IN0(n67), .IN1(n453), .SEL(n410), .F(n437) );
  IV U204 ( .A(n409), .Z(n67) );
  MUX U205 ( .IN0(n68), .IN1(n328), .SEL(n329), .F(n317) );
  IV U206 ( .A(n330), .Z(n68) );
  XOR U207 ( .A(n498), .B(n483), .Z(n487) );
  XNOR U208 ( .A(n617), .B(n618), .Z(n528) );
  XOR U209 ( .A(n357), .B(n344), .Z(n345) );
  MUX U210 ( .IN0(n69), .IN1(n756), .SEL(n757), .F(n567) );
  IV U211 ( .A(n758), .Z(n69) );
  MUX U212 ( .IN0(n70), .IN1(n746), .SEL(n747), .F(n403) );
  IV U213 ( .A(n748), .Z(n70) );
  MUX U214 ( .IN0(n375), .IN1(n71), .SEL(n277), .F(n353) );
  IV U215 ( .A(n276), .Z(n71) );
  MUX U216 ( .IN0(o_reg[13]), .IN1(n130), .SEL(n131), .F(n127) );
  MUX U217 ( .IN0(n72), .IN1(n254), .SEL(n117), .F(n247) );
  IV U218 ( .A(o_reg[2]), .Z(n72) );
  XOR U219 ( .A(n226), .B(n229), .Z(n227) );
  MUX U220 ( .IN0(n1119), .IN1(n73), .SEL(n961), .F(n1100) );
  IV U221 ( .A(n959), .Z(n73) );
  MUX U222 ( .IN0(n873), .IN1(n74), .SEL(n874), .F(n847) );
  IV U223 ( .A(n875), .Z(n74) );
  MUX U224 ( .IN0(n1048), .IN1(n75), .SEL(n856), .F(n1033) );
  IV U225 ( .A(n854), .Z(n75) );
  MUX U226 ( .IN0(e_input[1]), .IN1(n76), .SEL(e_input[15]), .F(n1015) );
  IV U227 ( .A(n1220), .Z(n76) );
  MUX U228 ( .IN0(n77), .IN1(n390), .SEL(n391), .F(n369) );
  IV U229 ( .A(n392), .Z(n77) );
  XNOR U230 ( .A(n986), .B(n976), .Z(n980) );
  MUX U231 ( .IN0(n765), .IN1(n767), .SEL(n766), .F(n562) );
  MUX U232 ( .IN0(n731), .IN1(n729), .SEL(n730), .F(n385) );
  MUX U233 ( .IN0(e_input[14]), .IN1(n1352), .SEL(e_input[15]), .F(n162) );
  MUX U234 ( .IN0(n431), .IN1(n78), .SEL(n430), .F(n416) );
  IV U235 ( .A(n429), .Z(n78) );
  MUX U236 ( .IN0(n79), .IN1(n437), .SEL(n301), .F(n424) );
  IV U237 ( .A(n300), .Z(n79) );
  MUX U238 ( .IN0(n324), .IN1(n322), .SEL(n323), .F(n315) );
  XOR U239 ( .A(n516), .B(n501), .Z(n505) );
  XNOR U240 ( .A(n631), .B(n632), .Z(n566) );
  NAND U241 ( .A(n397), .B(n741), .Z(n740) );
  MUX U242 ( .IN0(n374), .IN1(n372), .SEL(n373), .F(n80) );
  IV U243 ( .A(n80), .Z(n352) );
  MUX U244 ( .IN0(n406), .IN1(n81), .SEL(n407), .F(n375) );
  IV U245 ( .A(n408), .Z(n81) );
  MUX U246 ( .IN0(n302), .IN1(n82), .SEL(n285), .F(n289) );
  IV U247 ( .A(n284), .Z(n82) );
  MUX U248 ( .IN0(o_reg[12]), .IN1(n146), .SEL(n147), .F(n130) );
  MUX U249 ( .IN0(n83), .IN1(n213), .SEL(n111), .F(n206) );
  IV U250 ( .A(o_reg[8]), .Z(n83) );
  XOR U251 ( .A(n233), .B(n236), .Z(n234) );
  MUX U252 ( .IN0(n927), .IN1(n84), .SEL(n928), .F(n900) );
  IV U253 ( .A(n929), .Z(n84) );
  MUX U254 ( .IN0(n1100), .IN1(n85), .SEL(n936), .F(n1083) );
  IV U255 ( .A(n934), .Z(n85) );
  XNOR U256 ( .A(n1214), .B(n1215), .Z(n1201) );
  MUX U257 ( .IN0(n822), .IN1(n86), .SEL(n823), .F(n790) );
  IV U258 ( .A(n824), .Z(n86) );
  MUX U259 ( .IN0(n87), .IN1(n753), .SEL(n754), .F(n553) );
  IV U260 ( .A(n755), .Z(n87) );
  MUX U261 ( .IN0(g_input[9]), .IN1(n1112), .SEL(g_input[15]), .F(n511) );
  MUX U262 ( .IN0(g_input[8]), .IN1(n1129), .SEL(g_input[15]), .F(n531) );
  MUX U263 ( .IN0(n1033), .IN1(n88), .SEL(n831), .F(n1021) );
  IV U264 ( .A(n829), .Z(n88) );
  MUX U265 ( .IN0(n450), .IN1(n96), .SEL(n449), .F(n432) );
  MUX U266 ( .IN0(n527), .IN1(n616), .SEL(n528), .F(n609) );
  XOR U267 ( .A(n715), .B(n778), .Z(n716) );
  XNOR U268 ( .A(n572), .B(n573), .Z(n571) );
  MUX U269 ( .IN0(n89), .IN1(n472), .SEL(n304), .F(n453) );
  IV U270 ( .A(n303), .Z(n89) );
  XOR U271 ( .A(n536), .B(n521), .Z(n525) );
  XOR U272 ( .A(n349), .B(n350), .Z(n346) );
  XNOR U273 ( .A(n379), .B(n365), .Z(n359) );
  XNOR U274 ( .A(n768), .B(n682), .Z(n638) );
  XNOR U275 ( .A(n776), .B(n775), .Z(n758) );
  XNOR U276 ( .A(n547), .B(n548), .Z(n354) );
  XNOR U277 ( .A(n372), .B(n393), .Z(n373) );
  XOR U278 ( .A(n321), .B(n311), .Z(n283) );
  MUX U279 ( .IN0(o_reg[11]), .IN1(n174), .SEL(n175), .F(n146) );
  MUX U280 ( .IN0(n90), .IN1(n220), .SEL(n112), .F(n213) );
  IV U281 ( .A(o_reg[7]), .Z(n90) );
  XOR U282 ( .A(n240), .B(n243), .Z(n241) );
  MUX U283 ( .IN0(n91), .IN1(n940), .SEL(n941), .F(n913) );
  IV U284 ( .A(n942), .Z(n91) );
  MUX U285 ( .IN0(n1083), .IN1(n92), .SEL(n909), .F(n1066) );
  IV U286 ( .A(n907), .Z(n92) );
  MUX U287 ( .IN0(n900), .IN1(n93), .SEL(n901), .F(n873) );
  IV U288 ( .A(n902), .Z(n93) );
  MUX U289 ( .IN0(n94), .IN1(n1227), .SEL(n1228), .F(n1277) );
  IV U290 ( .A(n1297), .Z(n94) );
  XOR U291 ( .A(n1325), .B(g_input[3]), .Z(n1326) );
  XOR U292 ( .A(n1199), .B(n1200), .Z(n1009) );
  MUX U293 ( .IN0(n95), .IN1(n513), .SEL(n514), .F(n495) );
  IV U294 ( .A(n515), .Z(n95) );
  XOR U295 ( .A(n816), .B(n787), .Z(n791) );
  XOR U296 ( .A(n1143), .B(n1134), .Z(n985) );
  MUX U297 ( .IN0(n470), .IN1(n595), .SEL(n471), .F(n588) );
  MUX U298 ( .IN0(n460), .IN1(n462), .SEL(n461), .F(n96) );
  XOR U299 ( .A(n707), .B(n709), .Z(n628) );
  MUX U300 ( .IN0(n360), .IN1(n358), .SEL(n359), .F(n344) );
  XNOR U301 ( .A(n1021), .B(n1022), .Z(n1011) );
  XNOR U302 ( .A(n981), .B(n980), .Z(n797) );
  XNOR U303 ( .A(n624), .B(n625), .Z(n548) );
  XOR U304 ( .A(n556), .B(n541), .Z(n545) );
  XNOR U305 ( .A(n731), .B(n730), .Z(n748) );
  MUX U306 ( .IN0(g_input[14]), .IN1(n1016), .SEL(g_input[15]), .F(n163) );
  MUX U307 ( .IN0(n191), .IN1(n571), .SEL(n190), .F(n168) );
  MUX U308 ( .IN0(n97), .IN1(n411), .SEL(n297), .F(n183) );
  IV U309 ( .A(n296), .Z(n97) );
  XNOR U310 ( .A(n489), .B(n490), .Z(n303) );
  XNOR U311 ( .A(n527), .B(n528), .Z(n335) );
  XNOR U312 ( .A(n565), .B(n566), .Z(n376) );
  XNOR U313 ( .A(n387), .B(n386), .Z(n405) );
  XNOR U314 ( .A(n758), .B(n757), .Z(n738) );
  XNOR U315 ( .A(n319), .B(n320), .Z(n282) );
  XNOR U316 ( .A(n334), .B(n333), .Z(n337) );
  XNOR U317 ( .A(n569), .B(n568), .Z(n408) );
  MUX U318 ( .IN0(o_reg[10]), .IN1(n98), .SEL(n109), .F(n174) );
  IV U319 ( .A(n199), .Z(n98) );
  MUX U320 ( .IN0(n99), .IN1(n226), .SEL(n113), .F(n220) );
  IV U321 ( .A(o_reg[6]), .Z(n99) );
  MUX U322 ( .IN0(o_reg[14]), .IN1(n127), .SEL(n128), .F(n120) );
  XOR U323 ( .A(n247), .B(n250), .Z(n248) );
  MUX U324 ( .IN0(n1137), .IN1(n100), .SEL(n985), .F(n1119) );
  IV U325 ( .A(n984), .Z(n100) );
  MUX U326 ( .IN0(n952), .IN1(n101), .SEL(n953), .F(n927) );
  IV U327 ( .A(n954), .Z(n101) );
  NOR U328 ( .A(\_MAC/_MULT/A__[0] ), .B(n1349), .Z(n1340) );
  MUX U329 ( .IN0(n1066), .IN1(n102), .SEL(n882), .F(n1048) );
  IV U330 ( .A(n880), .Z(n102) );
  MUX U331 ( .IN0(n847), .IN1(n103), .SEL(n848), .F(n822) );
  IV U332 ( .A(n849), .Z(n103) );
  XOR U333 ( .A(n1207), .B(n1192), .Z(n1010) );
  XOR U334 ( .A(n1295), .B(n1296), .Z(n1227) );
  MUX U335 ( .IN0(e_input[13]), .IN1(n1347), .SEL(e_input[15]), .F(n187) );
  MUX U336 ( .IN0(e_input[2]), .IN1(n1205), .SEL(e_input[15]), .F(n742) );
  MUX U337 ( .IN0(n434), .IN1(n432), .SEL(n433), .F(n104) );
  IV U338 ( .A(n104), .Z(n421) );
  XOR U339 ( .A(n329), .B(n330), .Z(n324) );
  XOR U340 ( .A(n759), .B(n559), .Z(n563) );
  XNOR U341 ( .A(n723), .B(n382), .Z(n386) );
  MUX U342 ( .IN0(n750), .IN1(n1011), .SEL(n749), .F(n402) );
  AND U343 ( .A(n157), .B(n138), .Z(n156) );
  XNOR U344 ( .A(n422), .B(n423), .Z(n296) );
  XNOR U345 ( .A(n435), .B(n436), .Z(n298) );
  XNOR U346 ( .A(n451), .B(n452), .Z(n300) );
  XNOR U347 ( .A(n470), .B(n471), .Z(n409) );
  XNOR U348 ( .A(n507), .B(n508), .Z(n319) );
  XNOR U349 ( .A(n360), .B(n359), .Z(n374) );
  XNOR U350 ( .A(n639), .B(n638), .Z(n569) );
  MUX U351 ( .IN0(n736), .IN1(n105), .SEL(n737), .F(n406) );
  IV U352 ( .A(n738), .Z(n105) );
  XNOR U353 ( .A(n303), .B(n304), .Z(n284) );
  XNOR U354 ( .A(n335), .B(n336), .Z(n280) );
  XNOR U355 ( .A(n354), .B(n355), .Z(n278) );
  XNOR U356 ( .A(n376), .B(n377), .Z(n276) );
  MUX U357 ( .IN0(n106), .IN1(n206), .SEL(n110), .F(n199) );
  IV U358 ( .A(o_reg[9]), .Z(n106) );
  MUX U359 ( .IN0(n107), .IN1(n233), .SEL(n114), .F(n226) );
  IV U360 ( .A(o_reg[5]), .Z(n107) );
  MUX U361 ( .IN0(n261), .IN1(n108), .SEL(n262), .F(n254) );
  IV U362 ( .A(o_reg[1]), .Z(n108) );
  MUX U363 ( .IN0(o_reg[15]), .IN1(n120), .SEL(n121), .F(n119) );
  XNOR U364 ( .A(n109), .B(o_reg[10]), .Z(o[9]) );
  XNOR U365 ( .A(n110), .B(o_reg[9]), .Z(o[8]) );
  XNOR U366 ( .A(n111), .B(o_reg[8]), .Z(o[7]) );
  XNOR U367 ( .A(n112), .B(o_reg[7]), .Z(o[6]) );
  XNOR U368 ( .A(n113), .B(o_reg[6]), .Z(o[5]) );
  XNOR U369 ( .A(n114), .B(o_reg[5]), .Z(o[4]) );
  XNOR U370 ( .A(n115), .B(o_reg[4]), .Z(o[3]) );
  XNOR U371 ( .A(n116), .B(o_reg[3]), .Z(o[2]) );
  XNOR U372 ( .A(n117), .B(o_reg[2]), .Z(o[1]) );
  XOR U373 ( .A(n118), .B(n119), .Z(o[15]) );
  XNOR U374 ( .A(o_reg[15]), .B(n122), .Z(n118) );
  XNOR U375 ( .A(o_reg[15]), .B(n121), .Z(o[14]) );
  XOR U376 ( .A(n120), .B(n122), .Z(n121) );
  NAND U377 ( .A(n123), .B(n124), .Z(n122) );
  NANDN U378 ( .B(n125), .A(n126), .Z(n123) );
  XNOR U379 ( .A(n128), .B(o_reg[14]), .Z(o[13]) );
  XNOR U380 ( .A(n129), .B(n127), .Z(n128) );
  XOR U381 ( .A(n132), .B(n125), .Z(n126) );
  NANDN U382 ( .B(n133), .A(n134), .Z(n125) );
  AND U383 ( .A(n135), .B(n136), .Z(n132) );
  OR U384 ( .A(n137), .B(n138), .Z(n136) );
  AND U385 ( .A(n139), .B(n140), .Z(n135) );
  OR U386 ( .A(n141), .B(n142), .Z(n140) );
  OR U387 ( .A(n143), .B(n144), .Z(n139) );
  XNOR U388 ( .A(n131), .B(o_reg[13]), .Z(o[12]) );
  XNOR U389 ( .A(n145), .B(n130), .Z(n131) );
  XNOR U390 ( .A(n149), .B(n133), .Z(n134) );
  NANDN U391 ( .B(n150), .A(n151), .Z(n133) );
  IV U392 ( .A(n148), .Z(n149) );
  XNOR U393 ( .A(n144), .B(n143), .Z(n148) );
  OR U394 ( .A(n152), .B(n153), .Z(n143) );
  AND U395 ( .A(n154), .B(n155), .Z(n144) );
  XNOR U396 ( .A(n137), .B(n156), .Z(n155) );
  NAND U397 ( .A(n158), .B(n159), .Z(n138) );
  NANDN U398 ( .B(n160), .A(n161), .Z(n158) );
  NANDN U399 ( .B(n141), .A(n162), .Z(n157) );
  NANDN U400 ( .B(n142), .A(n163), .Z(n137) );
  AND U401 ( .A(n164), .B(n165), .Z(n154) );
  OR U402 ( .A(n166), .B(n167), .Z(n165) );
  XNOR U403 ( .A(n168), .B(n169), .Z(n164) );
  ANDN U404 ( .A(n170), .B(n171), .Z(n169) );
  XOR U405 ( .A(n168), .B(n172), .Z(n170) );
  XNOR U406 ( .A(n147), .B(o_reg[12]), .Z(o[11]) );
  XNOR U407 ( .A(n173), .B(n146), .Z(n147) );
  XNOR U408 ( .A(n177), .B(n150), .Z(n151) );
  NANDN U409 ( .B(n178), .A(n179), .Z(n150) );
  IV U410 ( .A(n176), .Z(n177) );
  XNOR U411 ( .A(n153), .B(n152), .Z(n176) );
  NANDN U412 ( .B(n180), .A(n181), .Z(n152) );
  XNOR U413 ( .A(n167), .B(n166), .Z(n153) );
  NANDN U414 ( .B(n182), .A(n183), .Z(n166) );
  XOR U415 ( .A(n172), .B(n171), .Z(n167) );
  XOR U416 ( .A(n168), .B(n184), .Z(n171) );
  AND U417 ( .A(n185), .B(n186), .Z(n184) );
  NANDN U418 ( .B(n141), .A(n187), .Z(n186) );
  OR U419 ( .A(n188), .B(n189), .Z(n185) );
  XOR U420 ( .A(n160), .B(n161), .Z(n172) );
  NANDN U421 ( .B(n142), .A(n192), .Z(n161) );
  XNOR U422 ( .A(n159), .B(n193), .Z(n160) );
  AND U423 ( .A(n163), .B(n162), .Z(n193) );
  ANDN U424 ( .A(n194), .B(n195), .Z(n159) );
  NANDN U425 ( .B(n196), .A(n197), .Z(n194) );
  XNOR U426 ( .A(n175), .B(o_reg[11]), .Z(o[10]) );
  XNOR U427 ( .A(n198), .B(n174), .Z(n175) );
  XNOR U428 ( .A(n200), .B(n201), .Z(n109) );
  AND U429 ( .A(n124), .B(n203), .Z(n202) );
  XOR U430 ( .A(n204), .B(n205), .Z(n203) );
  XNOR U431 ( .A(n207), .B(n208), .Z(n110) );
  AND U432 ( .A(n124), .B(n210), .Z(n209) );
  XOR U433 ( .A(n211), .B(n212), .Z(n210) );
  XNOR U434 ( .A(n214), .B(n215), .Z(n111) );
  AND U435 ( .A(n124), .B(n217), .Z(n216) );
  XOR U436 ( .A(n218), .B(n219), .Z(n217) );
  XNOR U437 ( .A(n222), .B(n223), .Z(n221) );
  AND U438 ( .A(n124), .B(n224), .Z(n223) );
  XOR U439 ( .A(n225), .B(n286), .Z(n224) );
  IV U440 ( .A(n220), .Z(n222) );
  XNOR U441 ( .A(n227), .B(n228), .Z(n113) );
  AND U442 ( .A(n124), .B(n230), .Z(n229) );
  XOR U443 ( .A(n231), .B(n232), .Z(n230) );
  XNOR U444 ( .A(n234), .B(n235), .Z(n114) );
  AND U445 ( .A(n124), .B(n237), .Z(n236) );
  XOR U446 ( .A(n238), .B(n239), .Z(n237) );
  XNOR U447 ( .A(n241), .B(n242), .Z(n115) );
  AND U448 ( .A(n124), .B(n244), .Z(n243) );
  XOR U449 ( .A(n245), .B(n246), .Z(n244) );
  XNOR U450 ( .A(n248), .B(n249), .Z(n116) );
  AND U451 ( .A(n124), .B(n251), .Z(n250) );
  XOR U452 ( .A(n252), .B(n253), .Z(n251) );
  XNOR U453 ( .A(n255), .B(n256), .Z(n117) );
  XOR U454 ( .A(n254), .B(n257), .Z(n255) );
  AND U455 ( .A(n124), .B(n258), .Z(n257) );
  XOR U456 ( .A(n259), .B(n260), .Z(n258) );
  XNOR U457 ( .A(n264), .B(n178), .Z(n179) );
  OR U458 ( .A(n204), .B(n265), .Z(n178) );
  XOR U459 ( .A(n205), .B(n265), .Z(n204) );
  OR U460 ( .A(n211), .B(n266), .Z(n265) );
  XOR U461 ( .A(n212), .B(n266), .Z(n211) );
  OR U462 ( .A(n218), .B(n267), .Z(n266) );
  XOR U463 ( .A(n219), .B(n267), .Z(n218) );
  OR U464 ( .A(n225), .B(n268), .Z(n267) );
  XOR U465 ( .A(n286), .B(n268), .Z(n225) );
  OR U466 ( .A(n231), .B(n269), .Z(n268) );
  XOR U467 ( .A(n232), .B(n269), .Z(n231) );
  OR U468 ( .A(n238), .B(n270), .Z(n269) );
  XOR U469 ( .A(n239), .B(n270), .Z(n238) );
  OR U470 ( .A(n245), .B(n271), .Z(n270) );
  XOR U471 ( .A(n246), .B(n271), .Z(n245) );
  OR U472 ( .A(n252), .B(n272), .Z(n271) );
  XOR U473 ( .A(n253), .B(n272), .Z(n252) );
  OR U474 ( .A(n259), .B(n273), .Z(n272) );
  XOR U475 ( .A(n260), .B(n273), .Z(n259) );
  NANDN U476 ( .B(n274), .A(n275), .Z(n273) );
  IV U477 ( .A(n256), .Z(n260) );
  XOR U478 ( .A(n276), .B(n277), .Z(n256) );
  IV U479 ( .A(n249), .Z(n253) );
  XOR U480 ( .A(n278), .B(n279), .Z(n249) );
  IV U481 ( .A(n242), .Z(n246) );
  XOR U482 ( .A(n280), .B(n281), .Z(n242) );
  IV U483 ( .A(n235), .Z(n239) );
  XOR U484 ( .A(n282), .B(n283), .Z(n235) );
  IV U485 ( .A(n228), .Z(n232) );
  XOR U486 ( .A(n284), .B(n285), .Z(n228) );
  XNOR U487 ( .A(n288), .B(n289), .Z(n286) );
  IV U488 ( .A(n215), .Z(n219) );
  XNOR U489 ( .A(n290), .B(n291), .Z(n215) );
  IV U490 ( .A(n208), .Z(n212) );
  XNOR U491 ( .A(n292), .B(n293), .Z(n208) );
  IV U492 ( .A(n201), .Z(n205) );
  XNOR U493 ( .A(n294), .B(n295), .Z(n201) );
  IV U494 ( .A(n263), .Z(n264) );
  XOR U495 ( .A(n181), .B(n180), .Z(n263) );
  OR U496 ( .A(n295), .B(n294), .Z(n180) );
  XNOR U497 ( .A(n296), .B(n297), .Z(n294) );
  OR U498 ( .A(n293), .B(n292), .Z(n295) );
  XNOR U499 ( .A(n298), .B(n299), .Z(n292) );
  OR U500 ( .A(n291), .B(n290), .Z(n293) );
  XNOR U501 ( .A(n300), .B(n301), .Z(n290) );
  NANDN U502 ( .B(n288), .A(n289), .Z(n291) );
  XNOR U503 ( .A(n302), .B(n305), .Z(n285) );
  AND U504 ( .A(n287), .B(n306), .Z(n305) );
  AND U505 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U506 ( .B(n141), .A(n309), .Z(n308) );
  OR U507 ( .A(n310), .B(n311), .Z(n307) );
  AND U508 ( .A(n312), .B(n313), .Z(n287) );
  NANDN U509 ( .B(n314), .A(n315), .Z(n313) );
  NANDN U510 ( .B(n316), .A(n317), .Z(n312) );
  XOR U511 ( .A(n314), .B(n315), .Z(n311) );
  XOR U512 ( .A(n325), .B(n316), .Z(n314) );
  NAND U513 ( .A(n163), .B(n309), .Z(n316) );
  NANDN U514 ( .B(n317), .A(n326), .Z(n325) );
  NANDN U515 ( .B(n141), .A(n327), .Z(n326) );
  XOR U516 ( .A(n331), .B(n310), .Z(n321) );
  OR U517 ( .A(n332), .B(n333), .Z(n310) );
  IV U518 ( .A(n318), .Z(n331) );
  XOR U519 ( .A(n337), .B(n332), .Z(n281) );
  XOR U520 ( .A(n324), .B(n323), .Z(n332) );
  XOR U521 ( .A(n322), .B(n338), .Z(n323) );
  AND U522 ( .A(n339), .B(n340), .Z(n338) );
  NANDN U523 ( .B(n141), .A(n341), .Z(n340) );
  OR U524 ( .A(n342), .B(n343), .Z(n339) );
  NAND U525 ( .A(n192), .B(n309), .Z(n330) );
  XNOR U526 ( .A(n328), .B(n347), .Z(n329) );
  AND U527 ( .A(n327), .B(n163), .Z(n347) );
  NANDN U528 ( .B(n351), .A(n352), .Z(n333) );
  XOR U529 ( .A(n356), .B(n351), .Z(n279) );
  XOR U530 ( .A(n346), .B(n345), .Z(n351) );
  XNOR U531 ( .A(n361), .B(n342), .Z(n357) );
  NAND U532 ( .A(n163), .B(n341), .Z(n342) );
  NANDN U533 ( .B(n141), .A(n363), .Z(n362) );
  NAND U534 ( .A(n367), .B(n309), .Z(n350) );
  XNOR U535 ( .A(n348), .B(n368), .Z(n349) );
  AND U536 ( .A(n327), .B(n192), .Z(n368) );
  XNOR U537 ( .A(n352), .B(n353), .Z(n356) );
  XNOR U538 ( .A(n378), .B(n374), .Z(n277) );
  XNOR U539 ( .A(n364), .B(n380), .Z(n365) );
  AND U540 ( .A(n363), .B(n163), .Z(n380) );
  XOR U541 ( .A(n384), .B(n366), .Z(n379) );
  NAND U542 ( .A(n192), .B(n341), .Z(n366) );
  IV U543 ( .A(n358), .Z(n384) );
  XNOR U544 ( .A(n370), .B(n371), .Z(n360) );
  NAND U545 ( .A(n388), .B(n309), .Z(n371) );
  XNOR U546 ( .A(n369), .B(n389), .Z(n370) );
  AND U547 ( .A(n327), .B(n367), .Z(n389) );
  XNOR U548 ( .A(n373), .B(n375), .Z(n378) );
  AND U549 ( .A(n394), .B(n395), .Z(n393) );
  OR U550 ( .A(n396), .B(n397), .Z(n395) );
  AND U551 ( .A(n398), .B(n399), .Z(n394) );
  NANDN U552 ( .B(n141), .A(n400), .Z(n399) );
  NANDN U553 ( .B(n401), .A(n402), .Z(n398) );
  XNOR U554 ( .A(n409), .B(n410), .Z(n288) );
  XNOR U555 ( .A(n182), .B(n183), .Z(n181) );
  XOR U556 ( .A(n411), .B(n412), .Z(n297) );
  AND U557 ( .A(n413), .B(n414), .Z(n412) );
  OR U558 ( .A(n415), .B(n416), .Z(n414) );
  AND U559 ( .A(n417), .B(n418), .Z(n413) );
  NANDN U560 ( .B(n141), .A(n419), .Z(n418) );
  NAND U561 ( .A(n420), .B(n421), .Z(n417) );
  XOR U562 ( .A(n425), .B(n420), .Z(n299) );
  XNOR U563 ( .A(n426), .B(n415), .Z(n420) );
  NAND U564 ( .A(n419), .B(n163), .Z(n415) );
  NANDN U565 ( .B(n141), .A(n428), .Z(n427) );
  XNOR U566 ( .A(n421), .B(n424), .Z(n425) );
  XOR U567 ( .A(n438), .B(n434), .Z(n301) );
  XNOR U568 ( .A(n430), .B(n431), .Z(n434) );
  NAND U569 ( .A(n419), .B(n192), .Z(n431) );
  XNOR U570 ( .A(n429), .B(n439), .Z(n430) );
  AND U571 ( .A(n163), .B(n428), .Z(n439) );
  XNOR U572 ( .A(n433), .B(n437), .Z(n438) );
  AND U573 ( .A(n444), .B(n445), .Z(n443) );
  NANDN U574 ( .B(n141), .A(n446), .Z(n445) );
  OR U575 ( .A(n447), .B(n448), .Z(n444) );
  XOR U576 ( .A(n454), .B(n450), .Z(n410) );
  XNOR U577 ( .A(n441), .B(n442), .Z(n450) );
  NAND U578 ( .A(n419), .B(n367), .Z(n442) );
  XNOR U579 ( .A(n440), .B(n455), .Z(n441) );
  AND U580 ( .A(n192), .B(n428), .Z(n455) );
  XNOR U581 ( .A(n449), .B(n453), .Z(n454) );
  XNOR U582 ( .A(n463), .B(n447), .Z(n459) );
  NAND U583 ( .A(n446), .B(n163), .Z(n447) );
  NANDN U584 ( .B(n464), .A(n465), .Z(n463) );
  NANDN U585 ( .B(n141), .A(n466), .Z(n465) );
  IV U586 ( .A(n448), .Z(n464) );
  XNOR U587 ( .A(n473), .B(n462), .Z(n304) );
  XNOR U588 ( .A(n457), .B(n458), .Z(n462) );
  NAND U589 ( .A(n419), .B(n388), .Z(n458) );
  XNOR U590 ( .A(n456), .B(n474), .Z(n457) );
  AND U591 ( .A(n367), .B(n428), .Z(n474) );
  XNOR U592 ( .A(n461), .B(n472), .Z(n473) );
  XNOR U593 ( .A(n467), .B(n479), .Z(n468) );
  AND U594 ( .A(n163), .B(n466), .Z(n479) );
  XOR U595 ( .A(n480), .B(n481), .Z(n467) );
  ANDN U596 ( .A(n482), .B(n483), .Z(n481) );
  XNOR U597 ( .A(n484), .B(n480), .Z(n482) );
  XOR U598 ( .A(n485), .B(n469), .Z(n478) );
  NAND U599 ( .A(n446), .B(n192), .Z(n469) );
  IV U600 ( .A(n460), .Z(n485) );
  XNOR U601 ( .A(n492), .B(n488), .Z(n320) );
  XNOR U602 ( .A(n476), .B(n477), .Z(n488) );
  NAND U603 ( .A(n419), .B(n493), .Z(n477) );
  XNOR U604 ( .A(n475), .B(n494), .Z(n476) );
  AND U605 ( .A(n388), .B(n428), .Z(n494) );
  XNOR U606 ( .A(n487), .B(n491), .Z(n492) );
  XNOR U607 ( .A(n480), .B(n499), .Z(n483) );
  AND U608 ( .A(n192), .B(n466), .Z(n499) );
  XOR U609 ( .A(n503), .B(n484), .Z(n498) );
  NAND U610 ( .A(n446), .B(n367), .Z(n484) );
  IV U611 ( .A(n486), .Z(n503) );
  XNOR U612 ( .A(n510), .B(n506), .Z(n336) );
  XNOR U613 ( .A(n496), .B(n497), .Z(n506) );
  NAND U614 ( .A(n419), .B(n511), .Z(n497) );
  XNOR U615 ( .A(n495), .B(n512), .Z(n496) );
  AND U616 ( .A(n493), .B(n428), .Z(n512) );
  XNOR U617 ( .A(n505), .B(n509), .Z(n510) );
  XNOR U618 ( .A(n500), .B(n517), .Z(n501) );
  AND U619 ( .A(n367), .B(n466), .Z(n517) );
  XOR U620 ( .A(n518), .B(n519), .Z(n500) );
  ANDN U621 ( .A(n520), .B(n521), .Z(n519) );
  XNOR U622 ( .A(n522), .B(n518), .Z(n520) );
  XOR U623 ( .A(n523), .B(n502), .Z(n516) );
  NAND U624 ( .A(n446), .B(n388), .Z(n502) );
  IV U625 ( .A(n504), .Z(n523) );
  XNOR U626 ( .A(n530), .B(n526), .Z(n355) );
  XNOR U627 ( .A(n514), .B(n515), .Z(n526) );
  NAND U628 ( .A(n419), .B(n531), .Z(n515) );
  XNOR U629 ( .A(n513), .B(n532), .Z(n514) );
  AND U630 ( .A(n511), .B(n428), .Z(n532) );
  XNOR U631 ( .A(n525), .B(n529), .Z(n530) );
  XNOR U632 ( .A(n518), .B(n537), .Z(n521) );
  AND U633 ( .A(n388), .B(n466), .Z(n537) );
  XOR U634 ( .A(n538), .B(n539), .Z(n518) );
  ANDN U635 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U636 ( .A(n542), .B(n538), .Z(n540) );
  XOR U637 ( .A(n543), .B(n522), .Z(n536) );
  NAND U638 ( .A(n446), .B(n493), .Z(n522) );
  IV U639 ( .A(n524), .Z(n543) );
  XNOR U640 ( .A(n550), .B(n546), .Z(n377) );
  XNOR U641 ( .A(n534), .B(n535), .Z(n546) );
  NAND U642 ( .A(n419), .B(n551), .Z(n535) );
  XNOR U643 ( .A(n533), .B(n552), .Z(n534) );
  AND U644 ( .A(n531), .B(n428), .Z(n552) );
  XNOR U645 ( .A(n545), .B(n549), .Z(n550) );
  XNOR U646 ( .A(n538), .B(n557), .Z(n541) );
  AND U647 ( .A(n493), .B(n466), .Z(n557) );
  XOR U648 ( .A(n561), .B(n542), .Z(n556) );
  NAND U649 ( .A(n446), .B(n511), .Z(n542) );
  IV U650 ( .A(n544), .Z(n561) );
  XOR U651 ( .A(n191), .B(n190), .Z(n182) );
  XNOR U652 ( .A(n570), .B(n571), .Z(n190) );
  ANDN U653 ( .A(n574), .B(n423), .Z(n573) );
  XOR U654 ( .A(n577), .B(n578), .Z(n575) );
  IV U655 ( .A(n572), .Z(n577) );
  XOR U656 ( .A(n572), .B(n422), .Z(n574) );
  XNOR U657 ( .A(n579), .B(n580), .Z(n422) );
  XOR U658 ( .A(n584), .B(n585), .Z(n582) );
  IV U659 ( .A(n581), .Z(n584) );
  XNOR U660 ( .A(n586), .B(n587), .Z(n435) );
  XOR U661 ( .A(n591), .B(n592), .Z(n589) );
  IV U662 ( .A(n588), .Z(n591) );
  XNOR U663 ( .A(n593), .B(n594), .Z(n451) );
  XOR U664 ( .A(n598), .B(n599), .Z(n596) );
  IV U665 ( .A(n595), .Z(n598) );
  XNOR U666 ( .A(n600), .B(n601), .Z(n470) );
  XOR U667 ( .A(n605), .B(n606), .Z(n603) );
  IV U668 ( .A(n602), .Z(n605) );
  XNOR U669 ( .A(n607), .B(n608), .Z(n489) );
  XOR U670 ( .A(n612), .B(n613), .Z(n610) );
  IV U671 ( .A(n609), .Z(n612) );
  XNOR U672 ( .A(n614), .B(n615), .Z(n507) );
  XOR U673 ( .A(n619), .B(n620), .Z(n617) );
  IV U674 ( .A(n616), .Z(n619) );
  XNOR U675 ( .A(n621), .B(n622), .Z(n527) );
  XOR U676 ( .A(n626), .B(n627), .Z(n624) );
  IV U677 ( .A(n623), .Z(n626) );
  XNOR U678 ( .A(n628), .B(n629), .Z(n547) );
  XOR U679 ( .A(n633), .B(n634), .Z(n631) );
  IV U680 ( .A(n630), .Z(n633) );
  XNOR U681 ( .A(n635), .B(n636), .Z(n565) );
  XNOR U682 ( .A(n640), .B(n188), .Z(n570) );
  NAND U683 ( .A(n187), .B(n163), .Z(n188) );
  NANDN U684 ( .B(n141), .A(n642), .Z(n641) );
  XNOR U685 ( .A(n643), .B(n644), .Z(n576) );
  AND U686 ( .A(n163), .B(n642), .Z(n644) );
  NAND U687 ( .A(n187), .B(n192), .Z(n578) );
  XOR U688 ( .A(n645), .B(n646), .Z(n643) );
  ANDN U689 ( .A(n647), .B(n583), .Z(n646) );
  XNOR U690 ( .A(n645), .B(n648), .Z(n583) );
  AND U691 ( .A(n192), .B(n642), .Z(n648) );
  XNOR U692 ( .A(n585), .B(n645), .Z(n647) );
  NAND U693 ( .A(n187), .B(n367), .Z(n585) );
  XOR U694 ( .A(n649), .B(n650), .Z(n645) );
  ANDN U695 ( .A(n651), .B(n590), .Z(n650) );
  XNOR U696 ( .A(n649), .B(n652), .Z(n590) );
  AND U697 ( .A(n367), .B(n642), .Z(n652) );
  XNOR U698 ( .A(n592), .B(n649), .Z(n651) );
  NAND U699 ( .A(n187), .B(n388), .Z(n592) );
  XOR U700 ( .A(n653), .B(n654), .Z(n649) );
  ANDN U701 ( .A(n655), .B(n597), .Z(n654) );
  XNOR U702 ( .A(n653), .B(n656), .Z(n597) );
  AND U703 ( .A(n388), .B(n642), .Z(n656) );
  XNOR U704 ( .A(n599), .B(n653), .Z(n655) );
  NAND U705 ( .A(n187), .B(n493), .Z(n599) );
  XOR U706 ( .A(n657), .B(n658), .Z(n653) );
  ANDN U707 ( .A(n659), .B(n604), .Z(n658) );
  XNOR U708 ( .A(n657), .B(n660), .Z(n604) );
  AND U709 ( .A(n493), .B(n642), .Z(n660) );
  XNOR U710 ( .A(n606), .B(n657), .Z(n659) );
  NAND U711 ( .A(n187), .B(n511), .Z(n606) );
  XOR U712 ( .A(n661), .B(n662), .Z(n657) );
  ANDN U713 ( .A(n663), .B(n611), .Z(n662) );
  XNOR U714 ( .A(n661), .B(n664), .Z(n611) );
  AND U715 ( .A(n511), .B(n642), .Z(n664) );
  XNOR U716 ( .A(n613), .B(n661), .Z(n663) );
  NAND U717 ( .A(n187), .B(n531), .Z(n613) );
  XOR U718 ( .A(n665), .B(n666), .Z(n661) );
  ANDN U719 ( .A(n667), .B(n618), .Z(n666) );
  XNOR U720 ( .A(n665), .B(n668), .Z(n618) );
  AND U721 ( .A(n531), .B(n642), .Z(n668) );
  XNOR U722 ( .A(n620), .B(n665), .Z(n667) );
  NAND U723 ( .A(n187), .B(n551), .Z(n620) );
  XOR U724 ( .A(n669), .B(n670), .Z(n665) );
  ANDN U725 ( .A(n671), .B(n625), .Z(n670) );
  XNOR U726 ( .A(n669), .B(n672), .Z(n625) );
  AND U727 ( .A(n551), .B(n642), .Z(n672) );
  XNOR U728 ( .A(n627), .B(n669), .Z(n671) );
  NAND U729 ( .A(n187), .B(n673), .Z(n627) );
  XOR U730 ( .A(n674), .B(n675), .Z(n669) );
  ANDN U731 ( .A(n676), .B(n632), .Z(n675) );
  XNOR U732 ( .A(n674), .B(n677), .Z(n632) );
  AND U733 ( .A(n673), .B(n642), .Z(n677) );
  XNOR U734 ( .A(n634), .B(n674), .Z(n676) );
  NAND U735 ( .A(n187), .B(n678), .Z(n634) );
  XOR U736 ( .A(n679), .B(n680), .Z(n674) );
  ANDN U737 ( .A(n681), .B(n682), .Z(n680) );
  XNOR U738 ( .A(n683), .B(n679), .Z(n681) );
  XOR U739 ( .A(n196), .B(n197), .Z(n191) );
  NANDN U740 ( .B(n142), .A(n367), .Z(n197) );
  AND U741 ( .A(n192), .B(n162), .Z(n684) );
  NAND U742 ( .A(n685), .B(n686), .Z(n195) );
  NANDN U743 ( .B(n579), .A(n580), .Z(n685) );
  NANDN U744 ( .B(n142), .A(n388), .Z(n580) );
  XNOR U745 ( .A(n686), .B(n687), .Z(n579) );
  AND U746 ( .A(n367), .B(n162), .Z(n687) );
  ANDN U747 ( .A(n688), .B(n689), .Z(n686) );
  NANDN U748 ( .B(n586), .A(n587), .Z(n688) );
  NANDN U749 ( .B(n142), .A(n493), .Z(n587) );
  AND U750 ( .A(n388), .B(n162), .Z(n690) );
  NAND U751 ( .A(n691), .B(n692), .Z(n689) );
  NANDN U752 ( .B(n593), .A(n594), .Z(n691) );
  NANDN U753 ( .B(n142), .A(n511), .Z(n594) );
  XNOR U754 ( .A(n692), .B(n693), .Z(n593) );
  AND U755 ( .A(n493), .B(n162), .Z(n693) );
  ANDN U756 ( .A(n694), .B(n695), .Z(n692) );
  NANDN U757 ( .B(n600), .A(n601), .Z(n694) );
  NANDN U758 ( .B(n142), .A(n531), .Z(n601) );
  AND U759 ( .A(n511), .B(n162), .Z(n696) );
  NAND U760 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U761 ( .B(n607), .A(n608), .Z(n697) );
  NANDN U762 ( .B(n142), .A(n551), .Z(n608) );
  XNOR U763 ( .A(n698), .B(n699), .Z(n607) );
  AND U764 ( .A(n531), .B(n162), .Z(n699) );
  ANDN U765 ( .A(n700), .B(n701), .Z(n698) );
  NANDN U766 ( .B(n614), .A(n615), .Z(n700) );
  NANDN U767 ( .B(n142), .A(n673), .Z(n615) );
  AND U768 ( .A(n551), .B(n162), .Z(n702) );
  NAND U769 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U770 ( .B(n621), .A(n622), .Z(n703) );
  NANDN U771 ( .B(n142), .A(n678), .Z(n622) );
  XNOR U772 ( .A(n704), .B(n705), .Z(n621) );
  AND U773 ( .A(n673), .B(n162), .Z(n705) );
  ANDN U774 ( .A(n706), .B(n707), .Z(n704) );
  NANDN U775 ( .B(n628), .A(n629), .Z(n706) );
  OR U776 ( .A(n708), .B(n142), .Z(n629) );
  AND U777 ( .A(n678), .B(n162), .Z(n709) );
  NAND U778 ( .A(n710), .B(n711), .Z(n707) );
  NANDN U779 ( .B(n635), .A(n636), .Z(n710) );
  OR U780 ( .A(n712), .B(n142), .Z(n636) );
  XNOR U781 ( .A(n711), .B(n713), .Z(n635) );
  ANDN U782 ( .A(n162), .B(n708), .Z(n713) );
  ANDN U783 ( .A(n714), .B(n715), .Z(n711) );
  NANDN U784 ( .B(n716), .A(n717), .Z(n714) );
  XOR U785 ( .A(n262), .B(o_reg[1]), .Z(o[0]) );
  XOR U786 ( .A(n718), .B(n719), .Z(n262) );
  XNOR U787 ( .A(n720), .B(n261), .Z(n718) );
  NANDN U788 ( .B(n275), .A(o_reg[0]), .Z(n261) );
  NAND U789 ( .A(n721), .B(n124), .Z(n720) );
  XOR U790 ( .A(e_input[15]), .B(g_input[15]), .Z(n124) );
  XNOR U791 ( .A(n274), .B(n719), .Z(n721) );
  XOR U792 ( .A(n275), .B(n719), .Z(n274) );
  XOR U793 ( .A(n408), .B(n407), .Z(n719) );
  XNOR U794 ( .A(n722), .B(n405), .Z(n407) );
  XNOR U795 ( .A(n381), .B(n724), .Z(n382) );
  AND U796 ( .A(n363), .B(n192), .Z(n724) );
  XOR U797 ( .A(n728), .B(n383), .Z(n723) );
  NAND U798 ( .A(n367), .B(n341), .Z(n383) );
  IV U799 ( .A(n385), .Z(n728) );
  XNOR U800 ( .A(n391), .B(n392), .Z(n387) );
  NAND U801 ( .A(n493), .B(n309), .Z(n392) );
  XNOR U802 ( .A(n390), .B(n732), .Z(n391) );
  AND U803 ( .A(n327), .B(n388), .Z(n732) );
  XNOR U804 ( .A(n404), .B(n406), .Z(n722) );
  XNOR U805 ( .A(n739), .B(n401), .Z(n404) );
  XOR U806 ( .A(n740), .B(n396), .Z(n401) );
  NAND U807 ( .A(n163), .B(n400), .Z(n396) );
  NANDN U808 ( .B(n141), .A(n742), .Z(n741) );
  XNOR U809 ( .A(n402), .B(n403), .Z(n739) );
  XNOR U810 ( .A(n751), .B(n564), .Z(n568) );
  XNOR U811 ( .A(n554), .B(n555), .Z(n564) );
  NAND U812 ( .A(n419), .B(n673), .Z(n555) );
  XNOR U813 ( .A(n553), .B(n752), .Z(n554) );
  AND U814 ( .A(n551), .B(n428), .Z(n752) );
  XNOR U815 ( .A(n563), .B(n567), .Z(n751) );
  XNOR U816 ( .A(n558), .B(n760), .Z(n559) );
  AND U817 ( .A(n511), .B(n466), .Z(n760) );
  XOR U818 ( .A(n764), .B(n560), .Z(n759) );
  NAND U819 ( .A(n446), .B(n531), .Z(n560) );
  IV U820 ( .A(n562), .Z(n764) );
  XNOR U821 ( .A(n679), .B(n769), .Z(n682) );
  AND U822 ( .A(n678), .B(n642), .Z(n769) );
  XOR U823 ( .A(n773), .B(n683), .Z(n768) );
  NANDN U824 ( .B(n708), .A(n187), .Z(n683) );
  IV U825 ( .A(n637), .Z(n773) );
  XNOR U826 ( .A(n716), .B(n717), .Z(n639) );
  NANDN U827 ( .B(n142), .A(n777), .Z(n717) );
  ANDN U828 ( .A(n162), .B(n712), .Z(n778) );
  NAND U829 ( .A(n779), .B(n780), .Z(n715) );
  NANDN U830 ( .B(n781), .A(n782), .Z(n779) );
  XOR U831 ( .A(n738), .B(n737), .Z(n275) );
  XNOR U832 ( .A(n783), .B(n748), .Z(n737) );
  XNOR U833 ( .A(n725), .B(n785), .Z(n726) );
  AND U834 ( .A(n363), .B(n367), .Z(n785) );
  XOR U835 ( .A(n789), .B(n727), .Z(n784) );
  NAND U836 ( .A(n388), .B(n341), .Z(n727) );
  IV U837 ( .A(n729), .Z(n789) );
  XNOR U838 ( .A(n734), .B(n735), .Z(n731) );
  NAND U839 ( .A(n511), .B(n309), .Z(n735) );
  XNOR U840 ( .A(n733), .B(n793), .Z(n734) );
  AND U841 ( .A(n327), .B(n493), .Z(n793) );
  XNOR U842 ( .A(n747), .B(n736), .Z(n783) );
  XOR U843 ( .A(n797), .B(n798), .Z(n736) );
  XNOR U844 ( .A(n799), .B(n750), .Z(n747) );
  NAND U845 ( .A(n192), .B(n400), .Z(n745) );
  XNOR U846 ( .A(n743), .B(n800), .Z(n744) );
  AND U847 ( .A(n742), .B(n163), .Z(n800) );
  XNOR U848 ( .A(n749), .B(n746), .Z(n799) );
  XOR U849 ( .A(n804), .B(n805), .Z(n746) );
  AND U850 ( .A(n806), .B(n807), .Z(n805) );
  XOR U851 ( .A(n808), .B(n809), .Z(n807) );
  XOR U852 ( .A(n804), .B(n810), .Z(n809) );
  XOR U853 ( .A(n791), .B(n811), .Z(n806) );
  XOR U854 ( .A(n804), .B(n792), .Z(n811) );
  NAND U855 ( .A(n309), .B(n531), .Z(n796) );
  XNOR U856 ( .A(n794), .B(n812), .Z(n795) );
  AND U857 ( .A(n327), .B(n511), .Z(n812) );
  XNOR U858 ( .A(n786), .B(n817), .Z(n787) );
  AND U859 ( .A(n363), .B(n388), .Z(n817) );
  XOR U860 ( .A(n821), .B(n788), .Z(n816) );
  NAND U861 ( .A(n493), .B(n341), .Z(n788) );
  IV U862 ( .A(n790), .Z(n821) );
  XOR U863 ( .A(n825), .B(n826), .Z(n804) );
  AND U864 ( .A(n827), .B(n828), .Z(n826) );
  XOR U865 ( .A(n829), .B(n830), .Z(n828) );
  XOR U866 ( .A(n825), .B(n831), .Z(n830) );
  XOR U867 ( .A(n823), .B(n832), .Z(n827) );
  XOR U868 ( .A(n825), .B(n824), .Z(n832) );
  NAND U869 ( .A(n309), .B(n551), .Z(n815) );
  XNOR U870 ( .A(n813), .B(n833), .Z(n814) );
  AND U871 ( .A(n531), .B(n327), .Z(n833) );
  XOR U872 ( .A(n834), .B(n835), .Z(n813) );
  ANDN U873 ( .A(n836), .B(n837), .Z(n835) );
  XNOR U874 ( .A(n838), .B(n834), .Z(n836) );
  XNOR U875 ( .A(n818), .B(n840), .Z(n819) );
  AND U876 ( .A(n363), .B(n493), .Z(n840) );
  XOR U877 ( .A(n841), .B(n842), .Z(n818) );
  ANDN U878 ( .A(n843), .B(n844), .Z(n842) );
  XNOR U879 ( .A(n845), .B(n841), .Z(n843) );
  XOR U880 ( .A(n846), .B(n820), .Z(n839) );
  NAND U881 ( .A(n511), .B(n341), .Z(n820) );
  IV U882 ( .A(n822), .Z(n846) );
  XOR U883 ( .A(n850), .B(n851), .Z(n825) );
  AND U884 ( .A(n852), .B(n853), .Z(n851) );
  XOR U885 ( .A(n854), .B(n855), .Z(n853) );
  XOR U886 ( .A(n850), .B(n856), .Z(n855) );
  XOR U887 ( .A(n848), .B(n857), .Z(n852) );
  XOR U888 ( .A(n850), .B(n849), .Z(n857) );
  NAND U889 ( .A(n309), .B(n673), .Z(n838) );
  XNOR U890 ( .A(n834), .B(n858), .Z(n837) );
  AND U891 ( .A(n551), .B(n327), .Z(n858) );
  XOR U892 ( .A(n859), .B(n860), .Z(n834) );
  ANDN U893 ( .A(n861), .B(n862), .Z(n860) );
  XNOR U894 ( .A(n863), .B(n859), .Z(n861) );
  XNOR U895 ( .A(n864), .B(n865), .Z(n848) );
  IV U896 ( .A(n844), .Z(n865) );
  XNOR U897 ( .A(n841), .B(n866), .Z(n844) );
  AND U898 ( .A(n363), .B(n511), .Z(n866) );
  XOR U899 ( .A(n867), .B(n868), .Z(n841) );
  ANDN U900 ( .A(n869), .B(n870), .Z(n868) );
  XNOR U901 ( .A(n871), .B(n867), .Z(n869) );
  XOR U902 ( .A(n872), .B(n845), .Z(n864) );
  NAND U903 ( .A(n341), .B(n531), .Z(n845) );
  IV U904 ( .A(n847), .Z(n872) );
  XOR U905 ( .A(n876), .B(n877), .Z(n850) );
  AND U906 ( .A(n878), .B(n879), .Z(n877) );
  XOR U907 ( .A(n880), .B(n881), .Z(n879) );
  XOR U908 ( .A(n876), .B(n882), .Z(n881) );
  XOR U909 ( .A(n874), .B(n883), .Z(n878) );
  XOR U910 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U911 ( .A(n884), .B(n863), .Z(n875) );
  NAND U912 ( .A(n309), .B(n678), .Z(n863) );
  IV U913 ( .A(n862), .Z(n884) );
  XNOR U914 ( .A(n859), .B(n885), .Z(n862) );
  AND U915 ( .A(n673), .B(n327), .Z(n885) );
  XOR U916 ( .A(n886), .B(n887), .Z(n859) );
  ANDN U917 ( .A(n888), .B(n889), .Z(n887) );
  XNOR U918 ( .A(n890), .B(n886), .Z(n888) );
  XNOR U919 ( .A(n891), .B(n892), .Z(n874) );
  IV U920 ( .A(n870), .Z(n892) );
  XNOR U921 ( .A(n867), .B(n893), .Z(n870) );
  AND U922 ( .A(n531), .B(n363), .Z(n893) );
  XOR U923 ( .A(n894), .B(n895), .Z(n867) );
  ANDN U924 ( .A(n896), .B(n897), .Z(n895) );
  XNOR U925 ( .A(n898), .B(n894), .Z(n896) );
  XOR U926 ( .A(n899), .B(n871), .Z(n891) );
  NAND U927 ( .A(n341), .B(n551), .Z(n871) );
  IV U928 ( .A(n873), .Z(n899) );
  XOR U929 ( .A(n903), .B(n904), .Z(n876) );
  AND U930 ( .A(n905), .B(n906), .Z(n904) );
  XOR U931 ( .A(n907), .B(n908), .Z(n906) );
  XOR U932 ( .A(n903), .B(n909), .Z(n908) );
  XOR U933 ( .A(n901), .B(n910), .Z(n905) );
  XOR U934 ( .A(n903), .B(n902), .Z(n910) );
  XNOR U935 ( .A(n911), .B(n890), .Z(n902) );
  NANDN U936 ( .B(n708), .A(n309), .Z(n890) );
  IV U937 ( .A(n889), .Z(n911) );
  XNOR U938 ( .A(n886), .B(n912), .Z(n889) );
  AND U939 ( .A(n678), .B(n327), .Z(n912) );
  XOR U940 ( .A(n913), .B(n914), .Z(n886) );
  ANDN U941 ( .A(n915), .B(n916), .Z(n914) );
  XNOR U942 ( .A(n917), .B(n913), .Z(n915) );
  XNOR U943 ( .A(n918), .B(n919), .Z(n901) );
  IV U944 ( .A(n897), .Z(n919) );
  XNOR U945 ( .A(n894), .B(n920), .Z(n897) );
  AND U946 ( .A(n551), .B(n363), .Z(n920) );
  XOR U947 ( .A(n921), .B(n922), .Z(n894) );
  ANDN U948 ( .A(n923), .B(n924), .Z(n922) );
  XNOR U949 ( .A(n925), .B(n921), .Z(n923) );
  XOR U950 ( .A(n926), .B(n898), .Z(n918) );
  NAND U951 ( .A(n341), .B(n673), .Z(n898) );
  IV U952 ( .A(n900), .Z(n926) );
  XOR U953 ( .A(n930), .B(n931), .Z(n903) );
  AND U954 ( .A(n932), .B(n933), .Z(n931) );
  XOR U955 ( .A(n934), .B(n935), .Z(n933) );
  XOR U956 ( .A(n930), .B(n936), .Z(n935) );
  XOR U957 ( .A(n928), .B(n937), .Z(n932) );
  XOR U958 ( .A(n930), .B(n929), .Z(n937) );
  XNOR U959 ( .A(n938), .B(n917), .Z(n929) );
  NANDN U960 ( .B(n712), .A(n309), .Z(n917) );
  IV U961 ( .A(n916), .Z(n938) );
  XNOR U962 ( .A(n913), .B(n939), .Z(n916) );
  ANDN U963 ( .A(n327), .B(n708), .Z(n939) );
  XNOR U964 ( .A(n943), .B(n944), .Z(n928) );
  IV U965 ( .A(n924), .Z(n944) );
  XNOR U966 ( .A(n921), .B(n945), .Z(n924) );
  AND U967 ( .A(n673), .B(n363), .Z(n945) );
  XOR U968 ( .A(n946), .B(n947), .Z(n921) );
  ANDN U969 ( .A(n948), .B(n949), .Z(n947) );
  XNOR U970 ( .A(n950), .B(n946), .Z(n948) );
  XOR U971 ( .A(n951), .B(n925), .Z(n943) );
  NAND U972 ( .A(n341), .B(n678), .Z(n925) );
  IV U973 ( .A(n927), .Z(n951) );
  XOR U974 ( .A(n955), .B(n956), .Z(n930) );
  AND U975 ( .A(n957), .B(n958), .Z(n956) );
  XOR U976 ( .A(n959), .B(n960), .Z(n958) );
  XOR U977 ( .A(n955), .B(n961), .Z(n960) );
  XOR U978 ( .A(n953), .B(n962), .Z(n957) );
  XOR U979 ( .A(n955), .B(n954), .Z(n962) );
  XNOR U980 ( .A(n963), .B(n942), .Z(n954) );
  NAND U981 ( .A(n309), .B(n777), .Z(n942) );
  IV U982 ( .A(n941), .Z(n963) );
  XNOR U983 ( .A(n940), .B(n964), .Z(n941) );
  ANDN U984 ( .A(n327), .B(n712), .Z(n964) );
  XOR U985 ( .A(n965), .B(n966), .Z(n940) );
  ANDN U986 ( .A(n967), .B(n968), .Z(n966) );
  XNOR U987 ( .A(n969), .B(n965), .Z(n967) );
  XNOR U988 ( .A(n970), .B(n971), .Z(n953) );
  IV U989 ( .A(n949), .Z(n971) );
  XNOR U990 ( .A(n946), .B(n972), .Z(n949) );
  AND U991 ( .A(n678), .B(n363), .Z(n972) );
  XOR U992 ( .A(n973), .B(n974), .Z(n946) );
  ANDN U993 ( .A(n975), .B(n976), .Z(n974) );
  XNOR U994 ( .A(n977), .B(n973), .Z(n975) );
  XOR U995 ( .A(n978), .B(n950), .Z(n970) );
  NANDN U996 ( .B(n708), .A(n341), .Z(n950) );
  IV U997 ( .A(n952), .Z(n978) );
  XOR U998 ( .A(n983), .B(n984), .Z(n798) );
  XNOR U999 ( .A(n985), .B(n982), .Z(n983) );
  XNOR U1000 ( .A(n973), .B(n987), .Z(n976) );
  ANDN U1001 ( .A(n363), .B(n708), .Z(n987) );
  XOR U1002 ( .A(n990), .B(n988), .Z(n989) );
  ANDN U1003 ( .A(n363), .B(n712), .Z(n990) );
  AND U1004 ( .A(n777), .B(n341), .Z(n991) );
  XOR U1005 ( .A(n992), .B(n993), .Z(n988) );
  ANDN U1006 ( .A(n994), .B(n995), .Z(n993) );
  XNOR U1007 ( .A(n996), .B(n992), .Z(n994) );
  XOR U1008 ( .A(n997), .B(n977), .Z(n986) );
  NANDN U1009 ( .B(n712), .A(n341), .Z(n977) );
  IV U1010 ( .A(n979), .Z(n997) );
  NAND U1011 ( .A(n341), .B(n998), .Z(n996) );
  XNOR U1012 ( .A(n992), .B(n999), .Z(n995) );
  AND U1013 ( .A(n777), .B(n363), .Z(n999) );
  AND U1014 ( .A(n1000), .B(\_MAC/_MULT/A__[0] ), .Z(n992) );
  NANDN U1015 ( .B(n341), .A(n1001), .Z(n1000) );
  NAND U1016 ( .A(n998), .B(n363), .Z(n1001) );
  XNOR U1017 ( .A(n968), .B(n969), .Z(n981) );
  NAND U1018 ( .A(n309), .B(n998), .Z(n969) );
  XNOR U1019 ( .A(n965), .B(n1004), .Z(n968) );
  AND U1020 ( .A(n777), .B(n327), .Z(n1004) );
  AND U1021 ( .A(n1005), .B(\_MAC/_MULT/A__[0] ), .Z(n965) );
  NANDN U1022 ( .B(n309), .A(n1006), .Z(n1005) );
  NAND U1023 ( .A(n998), .B(n327), .Z(n1006) );
  XOR U1024 ( .A(n1009), .B(n1010), .Z(n982) );
  XOR U1025 ( .A(n1011), .B(n1012), .Z(n749) );
  AND U1026 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U1027 ( .B(n141), .A(n1015), .Z(n1014) );
  NANDN U1028 ( .B(n1016), .A(n1017), .Z(n141) );
  AND U1029 ( .A(n1018), .B(g_input[15]), .Z(n1017) );
  OR U1030 ( .A(n1019), .B(n1020), .Z(n1013) );
  AND U1031 ( .A(n810), .B(n1023), .Z(n1022) );
  XNOR U1032 ( .A(n1021), .B(n808), .Z(n1023) );
  NAND U1033 ( .A(n367), .B(n400), .Z(n803) );
  XNOR U1034 ( .A(n801), .B(n1024), .Z(n802) );
  AND U1035 ( .A(n742), .B(n192), .Z(n1024) );
  XOR U1036 ( .A(n1032), .B(n1019), .Z(n1028) );
  NAND U1037 ( .A(n163), .B(n1015), .Z(n1019) );
  IV U1038 ( .A(n1021), .Z(n1032) );
  NAND U1039 ( .A(n388), .B(n400), .Z(n1027) );
  XNOR U1040 ( .A(n1025), .B(n1034), .Z(n1026) );
  AND U1041 ( .A(n742), .B(n367), .Z(n1034) );
  XOR U1042 ( .A(n1035), .B(n1036), .Z(n1025) );
  ANDN U1043 ( .A(n1037), .B(n1038), .Z(n1036) );
  XNOR U1044 ( .A(n1039), .B(n1035), .Z(n1037) );
  XNOR U1045 ( .A(n1029), .B(n1041), .Z(n1030) );
  AND U1046 ( .A(n163), .B(\_MAC/_MULT/X__[0] ), .Z(n1041) );
  XNOR U1047 ( .A(n1018), .B(g_input[14]), .Z(n1016) );
  NOR U1048 ( .A(n1042), .B(n1043), .Z(n1018) );
  XOR U1049 ( .A(n1047), .B(n1031), .Z(n1040) );
  NAND U1050 ( .A(n192), .B(n1015), .Z(n1031) );
  IV U1051 ( .A(n1033), .Z(n1047) );
  NAND U1052 ( .A(n493), .B(n400), .Z(n1039) );
  XNOR U1053 ( .A(n1035), .B(n1049), .Z(n1038) );
  AND U1054 ( .A(n742), .B(n388), .Z(n1049) );
  XOR U1055 ( .A(n1050), .B(n1051), .Z(n1035) );
  ANDN U1056 ( .A(n1052), .B(n1053), .Z(n1051) );
  XNOR U1057 ( .A(n1054), .B(n1050), .Z(n1052) );
  XNOR U1058 ( .A(n1055), .B(n1056), .Z(n856) );
  IV U1059 ( .A(n1045), .Z(n1056) );
  XNOR U1060 ( .A(n1044), .B(n1057), .Z(n1045) );
  AND U1061 ( .A(n192), .B(\_MAC/_MULT/X__[0] ), .Z(n1057) );
  XOR U1062 ( .A(n1042), .B(g_input[13]), .Z(n1043) );
  NANDN U1063 ( .B(n1058), .A(n1059), .Z(n1042) );
  XOR U1064 ( .A(n1060), .B(n1061), .Z(n1044) );
  ANDN U1065 ( .A(n1062), .B(n1063), .Z(n1061) );
  XNOR U1066 ( .A(n1064), .B(n1060), .Z(n1062) );
  XOR U1067 ( .A(n1065), .B(n1046), .Z(n1055) );
  NAND U1068 ( .A(n367), .B(n1015), .Z(n1046) );
  IV U1069 ( .A(n1048), .Z(n1065) );
  XNOR U1070 ( .A(n1067), .B(n1054), .Z(n880) );
  NAND U1071 ( .A(n511), .B(n400), .Z(n1054) );
  IV U1072 ( .A(n1053), .Z(n1067) );
  XNOR U1073 ( .A(n1050), .B(n1068), .Z(n1053) );
  AND U1074 ( .A(n742), .B(n493), .Z(n1068) );
  XOR U1075 ( .A(n1069), .B(n1070), .Z(n1050) );
  ANDN U1076 ( .A(n1071), .B(n1072), .Z(n1070) );
  XNOR U1077 ( .A(n1073), .B(n1069), .Z(n1071) );
  XNOR U1078 ( .A(n1074), .B(n1075), .Z(n882) );
  IV U1079 ( .A(n1063), .Z(n1075) );
  XNOR U1080 ( .A(n1060), .B(n1076), .Z(n1063) );
  AND U1081 ( .A(n367), .B(\_MAC/_MULT/X__[0] ), .Z(n1076) );
  XNOR U1082 ( .A(n1059), .B(g_input[12]), .Z(n1058) );
  NOR U1083 ( .A(n1077), .B(n1078), .Z(n1059) );
  XOR U1084 ( .A(n1082), .B(n1064), .Z(n1074) );
  NAND U1085 ( .A(n388), .B(n1015), .Z(n1064) );
  IV U1086 ( .A(n1066), .Z(n1082) );
  NAND U1087 ( .A(n531), .B(n400), .Z(n1073) );
  XNOR U1088 ( .A(n1069), .B(n1084), .Z(n1072) );
  AND U1089 ( .A(n742), .B(n511), .Z(n1084) );
  XOR U1090 ( .A(n1085), .B(n1086), .Z(n1069) );
  ANDN U1091 ( .A(n1087), .B(n1088), .Z(n1086) );
  XNOR U1092 ( .A(n1089), .B(n1085), .Z(n1087) );
  XNOR U1093 ( .A(n1079), .B(n1091), .Z(n1080) );
  AND U1094 ( .A(n388), .B(\_MAC/_MULT/X__[0] ), .Z(n1091) );
  XOR U1095 ( .A(n1077), .B(g_input[11]), .Z(n1078) );
  NANDN U1096 ( .B(n1092), .A(n1093), .Z(n1077) );
  XOR U1097 ( .A(n1094), .B(n1095), .Z(n1079) );
  ANDN U1098 ( .A(n1096), .B(n1097), .Z(n1095) );
  XNOR U1099 ( .A(n1098), .B(n1094), .Z(n1096) );
  XOR U1100 ( .A(n1099), .B(n1081), .Z(n1090) );
  NAND U1101 ( .A(n493), .B(n1015), .Z(n1081) );
  IV U1102 ( .A(n1083), .Z(n1099) );
  XNOR U1103 ( .A(n1101), .B(n1089), .Z(n934) );
  NAND U1104 ( .A(n551), .B(n400), .Z(n1089) );
  IV U1105 ( .A(n1088), .Z(n1101) );
  XNOR U1106 ( .A(n1085), .B(n1102), .Z(n1088) );
  AND U1107 ( .A(n742), .B(n531), .Z(n1102) );
  XOR U1108 ( .A(n1103), .B(n1104), .Z(n1085) );
  ANDN U1109 ( .A(n1105), .B(n1106), .Z(n1104) );
  XNOR U1110 ( .A(n1107), .B(n1103), .Z(n1105) );
  XNOR U1111 ( .A(n1108), .B(n1109), .Z(n936) );
  IV U1112 ( .A(n1097), .Z(n1109) );
  XNOR U1113 ( .A(n1094), .B(n1110), .Z(n1097) );
  AND U1114 ( .A(n493), .B(\_MAC/_MULT/X__[0] ), .Z(n1110) );
  XNOR U1115 ( .A(n1093), .B(g_input[10]), .Z(n1092) );
  NOR U1116 ( .A(n1111), .B(n1112), .Z(n1093) );
  XOR U1117 ( .A(n1113), .B(n1114), .Z(n1094) );
  ANDN U1118 ( .A(n1115), .B(n1116), .Z(n1114) );
  XNOR U1119 ( .A(n1117), .B(n1113), .Z(n1115) );
  XOR U1120 ( .A(n1118), .B(n1098), .Z(n1108) );
  NAND U1121 ( .A(n511), .B(n1015), .Z(n1098) );
  IV U1122 ( .A(n1100), .Z(n1118) );
  XNOR U1123 ( .A(n1120), .B(n1107), .Z(n959) );
  NAND U1124 ( .A(n673), .B(n400), .Z(n1107) );
  IV U1125 ( .A(n1106), .Z(n1120) );
  XNOR U1126 ( .A(n1103), .B(n1121), .Z(n1106) );
  AND U1127 ( .A(n742), .B(n551), .Z(n1121) );
  XOR U1128 ( .A(n1122), .B(n1123), .Z(n1103) );
  ANDN U1129 ( .A(n1124), .B(n1125), .Z(n1123) );
  XNOR U1130 ( .A(n1126), .B(n1122), .Z(n1124) );
  XNOR U1131 ( .A(n1113), .B(n1128), .Z(n1116) );
  AND U1132 ( .A(n511), .B(\_MAC/_MULT/X__[0] ), .Z(n1128) );
  XOR U1133 ( .A(n1111), .B(g_input[9]), .Z(n1112) );
  NANDN U1134 ( .B(n1129), .A(n1130), .Z(n1111) );
  XOR U1135 ( .A(n1131), .B(n1132), .Z(n1113) );
  ANDN U1136 ( .A(n1133), .B(n1134), .Z(n1132) );
  XNOR U1137 ( .A(n1135), .B(n1131), .Z(n1133) );
  XOR U1138 ( .A(n1136), .B(n1117), .Z(n1127) );
  NAND U1139 ( .A(n531), .B(n1015), .Z(n1117) );
  IV U1140 ( .A(n1119), .Z(n1136) );
  NAND U1141 ( .A(n678), .B(n400), .Z(n1126) );
  XNOR U1142 ( .A(n1122), .B(n1138), .Z(n1125) );
  AND U1143 ( .A(n742), .B(n673), .Z(n1138) );
  XNOR U1144 ( .A(n1142), .B(n1139), .Z(n1141) );
  XNOR U1145 ( .A(n1131), .B(n1144), .Z(n1134) );
  AND U1146 ( .A(n531), .B(\_MAC/_MULT/X__[0] ), .Z(n1144) );
  XNOR U1147 ( .A(n1148), .B(n1145), .Z(n1147) );
  XOR U1148 ( .A(n1149), .B(n1135), .Z(n1143) );
  NAND U1149 ( .A(n551), .B(n1015), .Z(n1135) );
  IV U1150 ( .A(n1137), .Z(n1149) );
  XNOR U1151 ( .A(n1150), .B(n1151), .Z(n1137) );
  AND U1152 ( .A(n1152), .B(n1153), .Z(n1151) );
  XOR U1153 ( .A(n1146), .B(n1154), .Z(n1153) );
  XNOR U1154 ( .A(n1148), .B(n1150), .Z(n1154) );
  NAND U1155 ( .A(n673), .B(n1015), .Z(n1148) );
  XOR U1156 ( .A(n1145), .B(n1155), .Z(n1146) );
  AND U1157 ( .A(n551), .B(\_MAC/_MULT/X__[0] ), .Z(n1155) );
  XNOR U1158 ( .A(n1159), .B(n1156), .Z(n1158) );
  XOR U1159 ( .A(n1140), .B(n1160), .Z(n1152) );
  XNOR U1160 ( .A(n1142), .B(n1150), .Z(n1160) );
  NANDN U1161 ( .B(n708), .A(n400), .Z(n1142) );
  XOR U1162 ( .A(n1139), .B(n1161), .Z(n1140) );
  AND U1163 ( .A(n742), .B(n678), .Z(n1161) );
  XOR U1164 ( .A(n1162), .B(n1163), .Z(n1139) );
  AND U1165 ( .A(n1164), .B(n1165), .Z(n1163) );
  XNOR U1166 ( .A(n1166), .B(n1162), .Z(n1165) );
  XOR U1167 ( .A(n1167), .B(n1168), .Z(n1150) );
  AND U1168 ( .A(n1169), .B(n1170), .Z(n1168) );
  XOR U1169 ( .A(n1157), .B(n1171), .Z(n1170) );
  XNOR U1170 ( .A(n1159), .B(n1167), .Z(n1171) );
  NAND U1171 ( .A(n678), .B(n1015), .Z(n1159) );
  XOR U1172 ( .A(n1156), .B(n1172), .Z(n1157) );
  AND U1173 ( .A(n673), .B(\_MAC/_MULT/X__[0] ), .Z(n1172) );
  XNOR U1174 ( .A(n1176), .B(n1173), .Z(n1175) );
  XOR U1175 ( .A(n1164), .B(n1177), .Z(n1169) );
  XNOR U1176 ( .A(n1166), .B(n1167), .Z(n1177) );
  NANDN U1177 ( .B(n712), .A(n400), .Z(n1166) );
  XOR U1178 ( .A(n1162), .B(n1178), .Z(n1164) );
  ANDN U1179 ( .A(n742), .B(n708), .Z(n1178) );
  XNOR U1180 ( .A(n1182), .B(n1179), .Z(n1181) );
  XOR U1181 ( .A(n1183), .B(n1184), .Z(n1167) );
  AND U1182 ( .A(n1185), .B(n1186), .Z(n1184) );
  XOR U1183 ( .A(n1174), .B(n1187), .Z(n1186) );
  XNOR U1184 ( .A(n1176), .B(n1183), .Z(n1187) );
  NANDN U1185 ( .B(n708), .A(n1015), .Z(n1176) );
  XOR U1186 ( .A(n1173), .B(n1188), .Z(n1174) );
  AND U1187 ( .A(n678), .B(\_MAC/_MULT/X__[0] ), .Z(n1188) );
  XOR U1188 ( .A(n1189), .B(n1190), .Z(n1173) );
  ANDN U1189 ( .A(n1191), .B(n1192), .Z(n1190) );
  XNOR U1190 ( .A(n1193), .B(n1189), .Z(n1191) );
  XOR U1191 ( .A(n1180), .B(n1194), .Z(n1185) );
  XNOR U1192 ( .A(n1182), .B(n1183), .Z(n1194) );
  NAND U1193 ( .A(n400), .B(n777), .Z(n1182) );
  XOR U1194 ( .A(n1179), .B(n1195), .Z(n1180) );
  ANDN U1195 ( .A(n742), .B(n712), .Z(n1195) );
  XOR U1196 ( .A(n1196), .B(n1197), .Z(n1179) );
  ANDN U1197 ( .A(n1198), .B(n1199), .Z(n1197) );
  XNOR U1198 ( .A(n1200), .B(n1196), .Z(n1198) );
  NAND U1199 ( .A(n400), .B(n998), .Z(n1200) );
  XNOR U1200 ( .A(n1196), .B(n1202), .Z(n1199) );
  AND U1201 ( .A(n777), .B(n742), .Z(n1202) );
  AND U1202 ( .A(n1203), .B(\_MAC/_MULT/A__[0] ), .Z(n1196) );
  NANDN U1203 ( .B(n400), .A(n1204), .Z(n1203) );
  NAND U1204 ( .A(n998), .B(n742), .Z(n1204) );
  XNOR U1205 ( .A(n1189), .B(n1208), .Z(n1192) );
  ANDN U1206 ( .A(\_MAC/_MULT/X__[0] ), .B(n708), .Z(n1208) );
  XOR U1207 ( .A(n1211), .B(n1209), .Z(n1210) );
  ANDN U1208 ( .A(\_MAC/_MULT/X__[0] ), .B(n712), .Z(n1211) );
  AND U1209 ( .A(n1015), .B(n777), .Z(n1212) );
  XOR U1210 ( .A(n1216), .B(n1193), .Z(n1207) );
  NANDN U1211 ( .B(n712), .A(n1015), .Z(n1193) );
  IV U1212 ( .A(n1201), .Z(n1216) );
  NAND U1213 ( .A(n1015), .B(n998), .Z(n1215) );
  XNOR U1214 ( .A(n1213), .B(n1217), .Z(n1214) );
  AND U1215 ( .A(n777), .B(\_MAC/_MULT/X__[0] ), .Z(n1217) );
  AND U1216 ( .A(n1218), .B(\_MAC/_MULT/A__[0] ), .Z(n1213) );
  NANDN U1217 ( .B(n1015), .A(n1219), .Z(n1218) );
  NAND U1218 ( .A(n998), .B(\_MAC/_MULT/X__[0] ), .Z(n1219) );
  XNOR U1219 ( .A(n1221), .B(n767), .Z(n757) );
  XNOR U1220 ( .A(n754), .B(n755), .Z(n767) );
  NAND U1221 ( .A(n419), .B(n678), .Z(n755) );
  XNOR U1222 ( .A(n753), .B(n1222), .Z(n754) );
  AND U1223 ( .A(n673), .B(n428), .Z(n1222) );
  XNOR U1224 ( .A(n1226), .B(n1223), .Z(n1225) );
  XNOR U1225 ( .A(n766), .B(n756), .Z(n1221) );
  XOR U1226 ( .A(n1227), .B(n1228), .Z(n756) );
  XNOR U1227 ( .A(n761), .B(n1230), .Z(n762) );
  AND U1228 ( .A(n531), .B(n466), .Z(n1230) );
  XNOR U1229 ( .A(n1130), .B(g_input[8]), .Z(n1129) );
  NOR U1230 ( .A(n1231), .B(n1232), .Z(n1130) );
  XOR U1231 ( .A(n1233), .B(n1234), .Z(n761) );
  AND U1232 ( .A(n1235), .B(n1236), .Z(n1234) );
  XNOR U1233 ( .A(n1237), .B(n1233), .Z(n1236) );
  XOR U1234 ( .A(n1238), .B(n763), .Z(n1229) );
  NAND U1235 ( .A(n446), .B(n551), .Z(n763) );
  IV U1236 ( .A(n765), .Z(n1238) );
  XNOR U1237 ( .A(n1239), .B(n1240), .Z(n765) );
  AND U1238 ( .A(n1241), .B(n1242), .Z(n1240) );
  XOR U1239 ( .A(n1235), .B(n1243), .Z(n1242) );
  XNOR U1240 ( .A(n1237), .B(n1239), .Z(n1243) );
  NAND U1241 ( .A(n446), .B(n673), .Z(n1237) );
  XOR U1242 ( .A(n1233), .B(n1244), .Z(n1235) );
  AND U1243 ( .A(n551), .B(n466), .Z(n1244) );
  XOR U1244 ( .A(n1231), .B(g_input[7]), .Z(n1232) );
  NANDN U1245 ( .B(n1245), .A(n1246), .Z(n1231) );
  XOR U1246 ( .A(n1247), .B(n1248), .Z(n1233) );
  AND U1247 ( .A(n1249), .B(n1250), .Z(n1248) );
  XNOR U1248 ( .A(n1251), .B(n1247), .Z(n1250) );
  XOR U1249 ( .A(n1224), .B(n1252), .Z(n1241) );
  XNOR U1250 ( .A(n1226), .B(n1239), .Z(n1252) );
  NANDN U1251 ( .B(n708), .A(n419), .Z(n1226) );
  XOR U1252 ( .A(n1223), .B(n1253), .Z(n1224) );
  AND U1253 ( .A(n678), .B(n428), .Z(n1253) );
  XNOR U1254 ( .A(n1257), .B(n1254), .Z(n1256) );
  XOR U1255 ( .A(n1258), .B(n1259), .Z(n1239) );
  AND U1256 ( .A(n1260), .B(n1261), .Z(n1259) );
  XOR U1257 ( .A(n1249), .B(n1262), .Z(n1261) );
  XNOR U1258 ( .A(n1251), .B(n1258), .Z(n1262) );
  NAND U1259 ( .A(n446), .B(n678), .Z(n1251) );
  XOR U1260 ( .A(n1247), .B(n1263), .Z(n1249) );
  AND U1261 ( .A(n673), .B(n466), .Z(n1263) );
  XNOR U1262 ( .A(n1246), .B(g_input[6]), .Z(n1245) );
  NOR U1263 ( .A(n1264), .B(n1265), .Z(n1246) );
  XOR U1264 ( .A(n1266), .B(n1267), .Z(n1247) );
  AND U1265 ( .A(n1268), .B(n1269), .Z(n1267) );
  XNOR U1266 ( .A(n1270), .B(n1266), .Z(n1269) );
  XOR U1267 ( .A(n1255), .B(n1271), .Z(n1260) );
  XNOR U1268 ( .A(n1257), .B(n1258), .Z(n1271) );
  NANDN U1269 ( .B(n712), .A(n419), .Z(n1257) );
  XOR U1270 ( .A(n1254), .B(n1272), .Z(n1255) );
  ANDN U1271 ( .A(n428), .B(n708), .Z(n1272) );
  XNOR U1272 ( .A(n1276), .B(n1273), .Z(n1275) );
  XOR U1273 ( .A(n1277), .B(n1278), .Z(n1258) );
  AND U1274 ( .A(n1279), .B(n1280), .Z(n1278) );
  XOR U1275 ( .A(n1268), .B(n1281), .Z(n1280) );
  XNOR U1276 ( .A(n1270), .B(n1277), .Z(n1281) );
  NANDN U1277 ( .B(n708), .A(n446), .Z(n1270) );
  XOR U1278 ( .A(n1266), .B(n1282), .Z(n1268) );
  AND U1279 ( .A(n678), .B(n466), .Z(n1282) );
  XOR U1280 ( .A(n1264), .B(g_input[5]), .Z(n1265) );
  NANDN U1281 ( .B(n1283), .A(n1284), .Z(n1264) );
  XOR U1282 ( .A(n1285), .B(n1286), .Z(n1266) );
  ANDN U1283 ( .A(n1287), .B(n1288), .Z(n1286) );
  XNOR U1284 ( .A(n1289), .B(n1285), .Z(n1287) );
  XOR U1285 ( .A(n1274), .B(n1290), .Z(n1279) );
  XNOR U1286 ( .A(n1276), .B(n1277), .Z(n1290) );
  NAND U1287 ( .A(n419), .B(n777), .Z(n1276) );
  XOR U1288 ( .A(n1273), .B(n1291), .Z(n1274) );
  ANDN U1289 ( .A(n428), .B(n712), .Z(n1291) );
  XOR U1290 ( .A(n1292), .B(n1293), .Z(n1273) );
  ANDN U1291 ( .A(n1294), .B(n1295), .Z(n1293) );
  XNOR U1292 ( .A(n1296), .B(n1292), .Z(n1294) );
  NAND U1293 ( .A(n419), .B(n998), .Z(n1296) );
  XNOR U1294 ( .A(n1292), .B(n1298), .Z(n1295) );
  AND U1295 ( .A(n777), .B(n428), .Z(n1298) );
  AND U1296 ( .A(n1299), .B(\_MAC/_MULT/A__[0] ), .Z(n1292) );
  NANDN U1297 ( .B(n419), .A(n1300), .Z(n1299) );
  NAND U1298 ( .A(n998), .B(n428), .Z(n1300) );
  XNOR U1299 ( .A(n1285), .B(n1304), .Z(n1288) );
  ANDN U1300 ( .A(n466), .B(n708), .Z(n1304) );
  XOR U1301 ( .A(n1305), .B(n1306), .Z(n1285) );
  AND U1302 ( .A(n1307), .B(n1308), .Z(n1306) );
  XOR U1303 ( .A(n1309), .B(n1305), .Z(n1308) );
  ANDN U1304 ( .A(n466), .B(n712), .Z(n1309) );
  XOR U1305 ( .A(n1310), .B(n1305), .Z(n1307) );
  AND U1306 ( .A(n777), .B(n446), .Z(n1310) );
  XOR U1307 ( .A(n1311), .B(n1312), .Z(n1305) );
  ANDN U1308 ( .A(n1313), .B(n1314), .Z(n1312) );
  XNOR U1309 ( .A(n1315), .B(n1311), .Z(n1313) );
  XOR U1310 ( .A(n1316), .B(n1289), .Z(n1303) );
  NANDN U1311 ( .B(n712), .A(n446), .Z(n1289) );
  IV U1312 ( .A(n1297), .Z(n1316) );
  XOR U1313 ( .A(n1317), .B(n1315), .Z(n1297) );
  NAND U1314 ( .A(n446), .B(n998), .Z(n1315) );
  IV U1315 ( .A(n1314), .Z(n1317) );
  XNOR U1316 ( .A(n1311), .B(n1318), .Z(n1314) );
  AND U1317 ( .A(n777), .B(n466), .Z(n1318) );
  AND U1318 ( .A(n1319), .B(\_MAC/_MULT/A__[0] ), .Z(n1311) );
  NANDN U1319 ( .B(n446), .A(n1320), .Z(n1319) );
  NAND U1320 ( .A(n998), .B(n466), .Z(n1320) );
  XNOR U1321 ( .A(n770), .B(n1324), .Z(n771) );
  ANDN U1322 ( .A(n642), .B(n708), .Z(n1324) );
  XNOR U1323 ( .A(n1284), .B(g_input[4]), .Z(n1283) );
  NOR U1324 ( .A(n1325), .B(n1326), .Z(n1284) );
  XOR U1325 ( .A(n1327), .B(n1328), .Z(n770) );
  AND U1326 ( .A(n1329), .B(n1330), .Z(n1328) );
  XOR U1327 ( .A(n1331), .B(n1327), .Z(n1330) );
  ANDN U1328 ( .A(n642), .B(n712), .Z(n1331) );
  XOR U1329 ( .A(n1332), .B(n1327), .Z(n1329) );
  AND U1330 ( .A(n777), .B(n187), .Z(n1332) );
  XOR U1331 ( .A(n1333), .B(n1334), .Z(n1327) );
  ANDN U1332 ( .A(n1335), .B(n1336), .Z(n1334) );
  XNOR U1333 ( .A(n1337), .B(n1333), .Z(n1335) );
  XOR U1334 ( .A(n1338), .B(n772), .Z(n1323) );
  NANDN U1335 ( .B(n712), .A(n187), .Z(n772) );
  NANDN U1336 ( .B(n1339), .A(n1340), .Z(n1325) );
  IV U1337 ( .A(n774), .Z(n1338) );
  NAND U1338 ( .A(n187), .B(n998), .Z(n1337) );
  XNOR U1339 ( .A(n1333), .B(n1341), .Z(n1336) );
  AND U1340 ( .A(n777), .B(n642), .Z(n1341) );
  AND U1341 ( .A(n1342), .B(\_MAC/_MULT/A__[0] ), .Z(n1333) );
  NANDN U1342 ( .B(n187), .A(n1343), .Z(n1342) );
  NAND U1343 ( .A(n998), .B(n642), .Z(n1343) );
  XNOR U1344 ( .A(n1344), .B(e_input[12]), .Z(n642) );
  NAND U1345 ( .A(n1345), .B(e_input[15]), .Z(n1344) );
  XOR U1346 ( .A(n1346), .B(e_input[12]), .Z(n1345) );
  XNOR U1347 ( .A(n781), .B(n782), .Z(n776) );
  NANDN U1348 ( .B(n142), .A(n998), .Z(n782) );
  XNOR U1349 ( .A(n780), .B(n1348), .Z(n781) );
  AND U1350 ( .A(n777), .B(n162), .Z(n1348) );
  XNOR U1351 ( .A(n1340), .B(g_input[2]), .Z(n1339) );
  AND U1352 ( .A(n1350), .B(\_MAC/_MULT/A__[0] ), .Z(n780) );
  NAND U1353 ( .A(n1351), .B(n142), .Z(n1350) );
  NANDN U1354 ( .B(n1352), .A(n1353), .Z(n142) );
  ANDN U1355 ( .A(e_input[15]), .B(n1354), .Z(n1353) );
  NAND U1356 ( .A(n998), .B(n162), .Z(n1351) );
  XOR U1357 ( .A(n1354), .B(e_input[14]), .Z(n1352) );
  OR U1358 ( .A(n1347), .B(n1355), .Z(n1354) );
  XOR U1359 ( .A(n1355), .B(e_input[13]), .Z(n1347) );
  OR U1360 ( .A(n1346), .B(n1356), .Z(n1355) );
  XOR U1361 ( .A(n1356), .B(e_input[12]), .Z(n1346) );
  OR U1362 ( .A(n1302), .B(n1357), .Z(n1356) );
  XOR U1363 ( .A(n1357), .B(e_input[11]), .Z(n1302) );
  OR U1364 ( .A(n1301), .B(n1358), .Z(n1357) );
  XOR U1365 ( .A(n1358), .B(e_input[10]), .Z(n1301) );
  OR U1366 ( .A(n1322), .B(n1359), .Z(n1358) );
  XOR U1367 ( .A(n1359), .B(e_input[9]), .Z(n1322) );
  OR U1368 ( .A(n1321), .B(n1360), .Z(n1359) );
  XOR U1369 ( .A(n1360), .B(e_input[8]), .Z(n1321) );
  OR U1370 ( .A(n1008), .B(n1361), .Z(n1360) );
  XOR U1371 ( .A(n1361), .B(e_input[7]), .Z(n1008) );
  OR U1372 ( .A(n1007), .B(n1362), .Z(n1361) );
  XOR U1373 ( .A(n1362), .B(e_input[6]), .Z(n1007) );
  OR U1374 ( .A(n1003), .B(n1363), .Z(n1362) );
  XOR U1375 ( .A(n1363), .B(e_input[5]), .Z(n1003) );
  OR U1376 ( .A(n1002), .B(n1364), .Z(n1363) );
  XOR U1377 ( .A(n1364), .B(e_input[4]), .Z(n1002) );
  OR U1378 ( .A(n1206), .B(n1365), .Z(n1364) );
  XOR U1379 ( .A(n1365), .B(e_input[3]), .Z(n1206) );
  OR U1380 ( .A(n1205), .B(n1366), .Z(n1365) );
  XOR U1381 ( .A(n1366), .B(e_input[2]), .Z(n1205) );
  NANDN U1382 ( .B(\_MAC/_MULT/X__[0] ), .A(n1220), .Z(n1366) );
  XNOR U1383 ( .A(\_MAC/_MULT/X__[0] ), .B(e_input[1]), .Z(n1220) );
  XOR U1384 ( .A(\_MAC/_MULT/A__[0] ), .B(g_input[1]), .Z(n1349) );
endmodule

