
module MxM_TG_W32_N10000 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MxM/n184 , \_MxM/n181 , \_MxM/n178 , \_MxM/n175 , \_MxM/n172 ,
         \_MxM/n169 , \_MxM/n166 , \_MxM/n163 , \_MxM/n160 , \_MxM/n157 ,
         \_MxM/n154 , \_MxM/n151 , \_MxM/n148 , \_MxM/n145 , \_MxM/n142 ,
         \_MxM/n139 , \_MxM/n136 , \_MxM/n133 , \_MxM/n130 , \_MxM/n127 ,
         \_MxM/n124 , \_MxM/n121 , \_MxM/n118 , \_MxM/n115 , \_MxM/n112 ,
         \_MxM/n109 , \_MxM/n106 , \_MxM/n103 , \_MxM/n100 , \_MxM/n97 ,
         \_MxM/n94 , \_MxM/n91 , \_MxM/N31 , \_MxM/N30 , \_MxM/N29 ,
         \_MxM/N28 , \_MxM/N27 , \_MxM/N26 , \_MxM/N25 , \_MxM/N24 ,
         \_MxM/N23 , \_MxM/N22 , \_MxM/N21 , \_MxM/N20 , \_MxM/N19 ,
         \_MxM/N18 , \_MxM/N16 , \_MxM/N15 , \_MxM/N14 , \_MxM/N13 ,
         \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/N7 ,
         \_MxM/N6 , \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] ,
         \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/n[7] ,
         \_MxM/n[8] , \_MxM/n[9] , \_MxM/n[10] , \_MxM/n[11] , \_MxM/n[12] ,
         \_MxM/n[13] , \_MxM/Y1[0] , \_MxM/Y1[1] , \_MxM/Y1[2] , \_MxM/Y1[3] ,
         \_MxM/Y1[4] , \_MxM/Y1[5] , \_MxM/Y1[6] , \_MxM/Y1[7] , \_MxM/Y1[8] ,
         \_MxM/Y1[9] , \_MxM/Y1[10] , \_MxM/Y1[11] , \_MxM/Y1[12] ,
         \_MxM/Y1[13] , \_MxM/Y1[14] , \_MxM/Y1[15] , \_MxM/Y1[16] ,
         \_MxM/Y1[17] , \_MxM/Y1[18] , \_MxM/Y1[19] , \_MxM/Y1[20] ,
         \_MxM/Y1[21] , \_MxM/Y1[22] , \_MxM/Y1[23] , \_MxM/Y1[24] ,
         \_MxM/Y1[25] , \_MxM/Y1[26] , \_MxM/Y1[27] , \_MxM/Y1[28] ,
         \_MxM/Y1[29] , \_MxM/Y1[30] , \_MxM/Y1[31] , \_MxM/Y0[31] ,
         \_MxM/Y0[30] , \_MxM/Y0[29] , \_MxM/Y0[28] , \_MxM/Y0[27] ,
         \_MxM/Y0[26] , \_MxM/Y0[25] , \_MxM/Y0[24] , \_MxM/Y0[23] ,
         \_MxM/Y0[22] , \_MxM/Y0[21] , \_MxM/Y0[20] , \_MxM/Y0[19] ,
         \_MxM/Y0[18] , \_MxM/Y0[17] , \_MxM/Y0[16] , \_MxM/Y0[15] ,
         \_MxM/Y0[14] , \_MxM/Y0[13] , \_MxM/Y0[12] , \_MxM/Y0[11] ,
         \_MxM/Y0[10] , \_MxM/Y0[9] , \_MxM/Y0[8] , \_MxM/Y0[7] , \_MxM/Y0[6] ,
         \_MxM/Y0[5] , \_MxM/Y0[4] , \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] ,
         \_MxM/Y0[0] , \_MxM/add_43/carry[13] , \_MxM/add_43/carry[12] ,
         \_MxM/add_43/carry[11] , \_MxM/add_43/carry[10] ,
         \_MxM/add_43/carry[9] , \_MxM/add_43/carry[8] ,
         \_MxM/add_43/carry[7] , \_MxM/add_43/carry[6] ,
         \_MxM/add_43/carry[5] , \_MxM/add_43/carry[4] ,
         \_MxM/add_43/carry[3] , \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226;

  DFF \_MxM/Y_reg[31]  ( .D(\_MxM/n91 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[31]) );
  DFF \_MxM/Y0_reg[31]  ( .D(\_MxM/Y1[31] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[31] ) );
  DFF \_MxM/Y_reg[30]  ( .D(\_MxM/n94 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[30]) );
  DFF \_MxM/Y0_reg[30]  ( .D(\_MxM/Y1[30] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[30] ) );
  DFF \_MxM/Y_reg[29]  ( .D(\_MxM/n97 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[29]) );
  DFF \_MxM/Y0_reg[29]  ( .D(\_MxM/Y1[29] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[29] ) );
  DFF \_MxM/Y_reg[28]  ( .D(\_MxM/n100 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[28]) );
  DFF \_MxM/Y0_reg[28]  ( .D(\_MxM/Y1[28] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[28] ) );
  DFF \_MxM/Y_reg[27]  ( .D(\_MxM/n103 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[27]) );
  DFF \_MxM/Y0_reg[27]  ( .D(\_MxM/Y1[27] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[27] ) );
  DFF \_MxM/Y_reg[26]  ( .D(\_MxM/n106 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[26]) );
  DFF \_MxM/Y0_reg[26]  ( .D(\_MxM/Y1[26] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[26] ) );
  DFF \_MxM/Y_reg[25]  ( .D(\_MxM/n109 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[25]) );
  DFF \_MxM/Y0_reg[25]  ( .D(\_MxM/Y1[25] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[25] ) );
  DFF \_MxM/Y_reg[24]  ( .D(\_MxM/n112 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[24]) );
  DFF \_MxM/Y0_reg[24]  ( .D(\_MxM/Y1[24] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[24] ) );
  DFF \_MxM/Y_reg[23]  ( .D(\_MxM/n115 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[23]) );
  DFF \_MxM/Y0_reg[23]  ( .D(\_MxM/Y1[23] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[23] ) );
  DFF \_MxM/Y_reg[22]  ( .D(\_MxM/n118 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[22]) );
  DFF \_MxM/Y0_reg[22]  ( .D(\_MxM/Y1[22] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[22] ) );
  DFF \_MxM/Y_reg[21]  ( .D(\_MxM/n121 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[21]) );
  DFF \_MxM/Y0_reg[21]  ( .D(\_MxM/Y1[21] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[21] ) );
  DFF \_MxM/Y_reg[20]  ( .D(\_MxM/n124 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[20]) );
  DFF \_MxM/Y0_reg[20]  ( .D(\_MxM/Y1[20] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[20] ) );
  DFF \_MxM/Y_reg[19]  ( .D(\_MxM/n127 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[19]) );
  DFF \_MxM/Y0_reg[19]  ( .D(\_MxM/Y1[19] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[19] ) );
  DFF \_MxM/Y_reg[18]  ( .D(\_MxM/n130 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[18]) );
  DFF \_MxM/Y0_reg[18]  ( .D(\_MxM/Y1[18] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[18] ) );
  DFF \_MxM/Y_reg[17]  ( .D(\_MxM/n133 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[17]) );
  DFF \_MxM/Y0_reg[17]  ( .D(\_MxM/Y1[17] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[17] ) );
  DFF \_MxM/Y_reg[16]  ( .D(\_MxM/n136 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[16]) );
  DFF \_MxM/Y0_reg[16]  ( .D(\_MxM/Y1[16] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[16] ) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n139 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/Y1[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n142 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/Y1[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n145 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/Y1[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n148 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/Y1[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n151 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/Y1[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n154 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/Y1[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n157 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/Y1[9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n160 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/Y1[8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n163 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n166 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n169 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n172 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n175 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n178 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n181 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n184 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[13]  ( .D(\_MxM/N31 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[13] ) );
  DFF \_MxM/n_reg[12]  ( .D(\_MxM/N30 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[12] ) );
  DFF \_MxM/n_reg[11]  ( .D(\_MxM/N29 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[11] ) );
  DFF \_MxM/n_reg[10]  ( .D(\_MxM/N28 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[10] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N27 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N26 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N25 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N24 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_43/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_43/carry[6] ), .COUT(\_MxM/add_43/carry[7] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_43/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_43/carry[7] ), .COUT(\_MxM/add_43/carry[8] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_43/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_43/carry[8] ), .COUT(\_MxM/add_43/carry[9] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_43/U1_1_9  ( .IN0(\_MxM/n[9] ), .IN1(\_MxM/add_43/carry[9] ), .COUT(\_MxM/add_43/carry[10] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_43/U1_1_10  ( .IN0(\_MxM/n[10] ), .IN1(
        \_MxM/add_43/carry[10] ), .COUT(\_MxM/add_43/carry[11] ), .SUM(
        \_MxM/N14 ) );
  HADDER \_MxM/add_43/U1_1_11  ( .IN0(\_MxM/n[11] ), .IN1(
        \_MxM/add_43/carry[11] ), .COUT(\_MxM/add_43/carry[12] ), .SUM(
        \_MxM/N15 ) );
  HADDER \_MxM/add_43/U1_1_12  ( .IN0(\_MxM/n[12] ), .IN1(
        \_MxM/add_43/carry[12] ), .COUT(\_MxM/add_43/carry[13] ), .SUM(
        \_MxM/N16 ) );
  MUX U1 ( .IN0(n1), .IN1(n4127), .SEL(n4128), .F(n4110) );
  IV U2 ( .A(n4129), .Z(n1) );
  XOR U3 ( .A(n4522), .B(n4514), .Z(n4124) );
  XOR U4 ( .A(n4455), .B(n4456), .Z(n4055) );
  XOR U5 ( .A(n4984), .B(n4976), .Z(n4852) );
  MUX U6 ( .IN0(n4426), .IN1(n2), .SEL(n4005), .F(n4413) );
  IV U7 ( .A(n4004), .Z(n2) );
  MUX U8 ( .IN0(n4587), .IN1(n3), .SEL(n4245), .F(n4576) );
  IV U9 ( .A(n4243), .Z(n3) );
  MUX U10 ( .IN0(n4361), .IN1(n4), .SEL(n3920), .F(n4348) );
  IV U11 ( .A(n3919), .Z(n4) );
  MUX U12 ( .IN0(n3194), .IN1(n3192), .SEL(n3193), .F(n3063) );
  MUX U13 ( .IN0(n2783), .IN1(n2781), .SEL(n2782), .F(n2654) );
  MUX U14 ( .IN0(n2562), .IN1(n2560), .SEL(n2561), .F(n2438) );
  MUX U15 ( .IN0(n2369), .IN1(n2367), .SEL(n2368), .F(n2251) );
  MUX U16 ( .IN0(n1930), .IN1(n1928), .SEL(n1929), .F(n1828) );
  MUX U17 ( .IN0(n1466), .IN1(n1464), .SEL(n1465), .F(n1387) );
  MUX U18 ( .IN0(n5), .IN1(n102), .SEL(n1439), .F(n1359) );
  IV U19 ( .A(n1440), .Z(n5) );
  MUX U20 ( .IN0(n1115), .IN1(n1113), .SEL(n1114), .F(n1052) );
  MUX U21 ( .IN0(n1141), .IN1(n1139), .SEL(n1140), .F(n1073) );
  MUX U22 ( .IN0(n852), .IN1(n850), .SEL(n851), .F(n811) );
  MUX U23 ( .IN0(n6), .IN1(n3125), .SEL(n3126), .F(n2989) );
  IV U24 ( .A(n3127), .Z(n6) );
  MUX U25 ( .IN0(n7), .IN1(n1356), .SEL(n1357), .F(n1287) );
  IV U26 ( .A(n1358), .Z(n7) );
  MUX U27 ( .IN0(n8), .IN1(n1210), .SEL(n1211), .F(n1146) );
  IV U28 ( .A(n1212), .Z(n8) );
  MUX U29 ( .IN0(n1866), .IN1(n9), .SEL(n1867), .F(n1766) );
  IV U30 ( .A(n1868), .Z(n9) );
  MUX U31 ( .IN0(n914), .IN1(n10), .SEL(n913), .F(n868) );
  IV U32 ( .A(n912), .Z(n10) );
  OR U33 ( .A(n760), .B(n761), .Z(n731) );
  XNOR U34 ( .A(n712), .B(n711), .Z(n710) );
  MUX U35 ( .IN0(n4133), .IN1(n4131), .SEL(n4132), .F(n4114) );
  MUX U36 ( .IN0(n3766), .IN1(n3768), .SEL(n3767), .F(n3728) );
  XOR U37 ( .A(n4509), .B(n4501), .Z(n4107) );
  MUX U38 ( .IN0(n3595), .IN1(n3593), .SEL(n3594), .F(n3555) );
  XNOR U39 ( .A(n4074), .B(n4060), .Z(n4064) );
  XOR U40 ( .A(n4470), .B(n4462), .Z(n4056) );
  XOR U41 ( .A(n4442), .B(n4443), .Z(n4038) );
  MUX U42 ( .IN0(n4014), .IN1(n4012), .SEL(n4013), .F(n3995) );
  MUX U43 ( .IN0(n4620), .IN1(n11), .SEL(n4305), .F(n4609) );
  IV U44 ( .A(n4304), .Z(n11) );
  MUX U45 ( .IN0(n4278), .IN1(n12), .SEL(n4279), .F(n4257) );
  IV U46 ( .A(n4280), .Z(n12) );
  MUX U47 ( .IN0(n4979), .IN1(n13), .SEL(n4852), .F(n4966) );
  IV U48 ( .A(n4850), .Z(n13) );
  MUX U49 ( .IN0(n14), .IN1(n4572), .SEL(n4573), .F(n4561) );
  IV U50 ( .A(n4574), .Z(n14) );
  MUX U51 ( .IN0(n15), .IN1(n4211), .SEL(n4212), .F(n4190) );
  IV U52 ( .A(n4213), .Z(n15) );
  MUX U53 ( .IN0(n4400), .IN1(n16), .SEL(n3971), .F(n4387) );
  IV U54 ( .A(n3970), .Z(n16) );
  MUX U55 ( .IN0(n4801), .IN1(n17), .SEL(n4802), .F(n4780) );
  IV U56 ( .A(n4803), .Z(n17) );
  MUX U57 ( .IN0(n3946), .IN1(n3944), .SEL(n3945), .F(n3927) );
  MUX U58 ( .IN0(n4927), .IN1(n18), .SEL(n4768), .F(n4914) );
  IV U59 ( .A(n4766), .Z(n18) );
  MUX U60 ( .IN0(n3253), .IN1(n3251), .SEL(n3252), .F(n3213) );
  XOR U61 ( .A(n4353), .B(n4342), .Z(n3903) );
  MUX U62 ( .IN0(n19), .IN1(n3172), .SEL(n3173), .F(n3042) );
  IV U63 ( .A(n3174), .Z(n19) );
  MUX U64 ( .IN0(n20), .IN1(n2597), .SEL(n2598), .F(n2475) );
  IV U65 ( .A(n2599), .Z(n20) );
  MUX U66 ( .IN0(n21), .IN1(n2125), .SEL(n2126), .F(n2020) );
  IV U67 ( .A(n2127), .Z(n21) );
  MUX U68 ( .IN0(n22), .IN1(n1410), .SEL(n1411), .F(n1335) );
  IV U69 ( .A(n1412), .Z(n22) );
  MUX U70 ( .IN0(n23), .IN1(n1451), .SEL(n1452), .F(n1372) );
  IV U71 ( .A(n1453), .Z(n23) );
  MUX U72 ( .IN0(n24), .IN1(n1162), .SEL(n1163), .F(n1100) );
  IV U73 ( .A(n1164), .Z(n24) );
  MUX U74 ( .IN0(n3145), .IN1(n3143), .SEL(n3144), .F(n3007) );
  MUX U75 ( .IN0(n2959), .IN1(n2957), .SEL(n2958), .F(n2819) );
  MUX U76 ( .IN0(n2929), .IN1(n2927), .SEL(n2928), .F(n2793) );
  MUX U77 ( .IN0(n2656), .IN1(n2654), .SEL(n2655), .F(n2528) );
  MUX U78 ( .IN0(n2519), .IN1(n2521), .SEL(n2520), .F(n2398) );
  MUX U79 ( .IN0(n2253), .IN1(n2251), .SEL(n2252), .F(n2138) );
  MUX U80 ( .IN0(n2201), .IN1(n2199), .SEL(n2200), .F(n2088) );
  MUX U81 ( .IN0(n2112), .IN1(n2114), .SEL(n2113), .F(n2007) );
  MUX U82 ( .IN0(n1736), .IN1(n1734), .SEL(n1735), .F(n1643) );
  MUX U83 ( .IN0(n1686), .IN1(n1684), .SEL(n1685), .F(n1593) );
  MUX U84 ( .IN0(n1634), .IN1(n1636), .SEL(n1635), .F(n1540) );
  MUX U85 ( .IN0(n1389), .IN1(n1387), .SEL(n1388), .F(n1313) );
  MUX U86 ( .IN0(n1355), .IN1(n25), .SEL(n1354), .F(n1286) );
  IV U87 ( .A(n1353), .Z(n25) );
  MUX U88 ( .IN0(n1054), .IN1(n1052), .SEL(n1053), .F(n998) );
  MUX U89 ( .IN0(n881), .IN1(n883), .SEL(n882), .F(n841) );
  MUX U90 ( .IN0(n26), .IN1(n2722), .SEL(n2723), .F(n2592) );
  IV U91 ( .A(n2724), .Z(n26) );
  MUX U92 ( .IN0(n2160), .IN1(n27), .SEL(n2161), .F(n2057) );
  IV U93 ( .A(n2162), .Z(n27) );
  MUX U94 ( .IN0(n28), .IN1(n1910), .SEL(n1911), .F(n1810) );
  IV U95 ( .A(n1912), .Z(n28) );
  MUX U96 ( .IN0(n29), .IN1(n1095), .SEL(n1096), .F(n1034) );
  IV U97 ( .A(n1097), .Z(n29) );
  MUX U98 ( .IN0(n813), .IN1(n811), .SEL(n812), .F(n772) );
  MUX U99 ( .IN0(n2430), .IN1(n2428), .SEL(n2429), .F(n2303) );
  MUX U100 ( .IN0(n30), .IN1(n2445), .SEL(n2446), .F(n2324) );
  IV U101 ( .A(n2447), .Z(n30) );
  MUX U102 ( .IN0(n31), .IN1(n1505), .SEL(n1506), .F(n1421) );
  IV U103 ( .A(n1507), .Z(n31) );
  XNOR U104 ( .A(n1271), .B(n1270), .Z(n1289) );
  OR U105 ( .A(n1088), .B(n1089), .Z(n1027) );
  MUX U106 ( .IN0(n1672), .IN1(n32), .SEL(n1673), .F(n1583) );
  IV U107 ( .A(n1674), .Z(n32) );
  OR U108 ( .A(n868), .B(n869), .Z(n829) );
  AND U109 ( .A(n780), .B(n781), .Z(n750) );
  OR U110 ( .A(n1130), .B(n1131), .Z(n1068) );
  OR U111 ( .A(n758), .B(n759), .Z(n729) );
  OR U112 ( .A(n709), .B(n710), .Z(n687) );
  MUX U113 ( .IN0(n3747), .IN1(n3745), .SEL(n3746), .F(n3707) );
  MUX U114 ( .IN0(n4116), .IN1(n4114), .SEL(n4115), .F(n4097) );
  MUX U115 ( .IN0(n33), .IN1(n4506), .SEL(n4507), .F(n4493) );
  IV U116 ( .A(n4508), .Z(n33) );
  XOR U117 ( .A(n3722), .B(n3687), .Z(n3691) );
  XOR U118 ( .A(n4496), .B(n4488), .Z(n4090) );
  XOR U119 ( .A(n4457), .B(n4449), .Z(n4039) );
  MUX U120 ( .IN0(n4031), .IN1(n4029), .SEL(n4030), .F(n4012) );
  MUX U121 ( .IN0(n34), .IN1(n3496), .SEL(n3497), .F(n3458) );
  IV U122 ( .A(n3498), .Z(n34) );
  XNOR U123 ( .A(n3511), .B(n3476), .Z(n3480) );
  MUX U124 ( .IN0(n35), .IN1(n3991), .SEL(n3992), .F(n3974) );
  IV U125 ( .A(n3993), .Z(n35) );
  MUX U126 ( .IN0(n36), .IN1(n4600), .SEL(n4601), .F(n4589) );
  IV U127 ( .A(n4602), .Z(n36) );
  MUX U128 ( .IN0(n4301), .IN1(n4299), .SEL(n4300), .F(n4278) );
  MUX U129 ( .IN0(n37), .IN1(n4975), .SEL(n4976), .F(n4962) );
  IV U130 ( .A(n4977), .Z(n37) );
  MUX U131 ( .IN0(n4866), .IN1(n4864), .SEL(n4865), .F(n4843) );
  MUX U132 ( .IN0(n38), .IN1(n3982), .SEL(n3983), .F(n3965) );
  IV U133 ( .A(n3984), .Z(n38) );
  XNOR U134 ( .A(n3397), .B(n3362), .Z(n3366) );
  XOR U135 ( .A(n4405), .B(n4397), .Z(n3971) );
  XOR U136 ( .A(n3418), .B(n3383), .Z(n3387) );
  XOR U137 ( .A(n4377), .B(n4378), .Z(n3953) );
  XOR U138 ( .A(n4945), .B(n4937), .Z(n4789) );
  MUX U139 ( .IN0(n39), .IN1(n3923), .SEL(n3924), .F(n3906) );
  IV U140 ( .A(n3925), .Z(n39) );
  MUX U141 ( .IN0(n4576), .IN1(n40), .SEL(n4224), .F(n4565) );
  IV U142 ( .A(n4222), .Z(n40) );
  MUX U143 ( .IN0(n4215), .IN1(n41), .SEL(n4216), .F(n4194) );
  IV U144 ( .A(n4217), .Z(n41) );
  MUX U145 ( .IN0(n4759), .IN1(n42), .SEL(n4760), .F(n4738) );
  IV U146 ( .A(n4761), .Z(n42) );
  XOR U147 ( .A(n4346), .B(n4347), .Z(n3902) );
  XOR U148 ( .A(n4906), .B(n4898), .Z(n4726) );
  MUX U149 ( .IN0(n43), .IN1(n4710), .SEL(n4711), .F(n3097) );
  IV U150 ( .A(n4712), .Z(n43) );
  MUX U151 ( .IN0(n44), .IN1(n3180), .SEL(n3181), .F(n3050) );
  IV U152 ( .A(n3182), .Z(n44) );
  XNOR U153 ( .A(n3207), .B(n3173), .Z(n3177) );
  MUX U154 ( .IN0(n45), .IN1(n2994), .SEL(n2995), .F(n2856) );
  IV U155 ( .A(n2996), .Z(n45) );
  MUX U156 ( .IN0(n46), .IN1(n2768), .SEL(n2769), .F(n2641) );
  IV U157 ( .A(n2770), .Z(n46) );
  MUX U158 ( .IN0(n47), .IN1(n2524), .SEL(n2525), .F(n2403) );
  IV U159 ( .A(n2526), .Z(n47) );
  MUX U160 ( .IN0(n48), .IN1(n2580), .SEL(n2581), .F(n2458) );
  IV U161 ( .A(n2582), .Z(n48) );
  MUX U162 ( .IN0(n49), .IN1(n2065), .SEL(n2066), .F(n1960) );
  IV U163 ( .A(n2067), .Z(n49) );
  MUX U164 ( .IN0(n50), .IN1(n1798), .SEL(n1799), .F(n1704) );
  IV U165 ( .A(n1800), .Z(n50) );
  MUX U166 ( .IN0(n51), .IN1(n1335), .SEL(n1336), .F(n1265) );
  IV U167 ( .A(n1337), .Z(n51) );
  MUX U168 ( .IN0(n52), .IN1(n1300), .SEL(n1301), .F(n1230) );
  IV U169 ( .A(n1302), .Z(n52) );
  MUX U170 ( .IN0(n53), .IN1(n1239), .SEL(n1240), .F(n1171) );
  IV U171 ( .A(n1241), .Z(n53) );
  MUX U172 ( .IN0(n54), .IN1(n994), .SEL(n995), .F(n934) );
  IV U173 ( .A(n996), .Z(n54) );
  MUX U174 ( .IN0(n3037), .IN1(n3039), .SEL(n3038), .F(n2901) );
  MUX U175 ( .IN0(n3065), .IN1(n3063), .SEL(n3064), .F(n2927) );
  MUX U176 ( .IN0(n2843), .IN1(n2845), .SEL(n2844), .F(n2714) );
  MUX U177 ( .IN0(n2821), .IN1(n2819), .SEL(n2820), .F(n2690) );
  MUX U178 ( .IN0(n2871), .IN1(n2869), .SEL(n2870), .F(n2740) );
  MUX U179 ( .IN0(n2801), .IN1(n55), .SEL(n2800), .F(n2670) );
  IV U180 ( .A(n2799), .Z(n55) );
  MUX U181 ( .IN0(n2731), .IN1(n2733), .SEL(n2732), .F(n2601) );
  MUX U182 ( .IN0(n2398), .IN1(n2400), .SEL(n2399), .F(n2277) );
  MUX U183 ( .IN0(n2294), .IN1(n2292), .SEL(n2293), .F(n2178) );
  MUX U184 ( .IN0(n2319), .IN1(n2317), .SEL(n2318), .F(n2199) );
  MUX U185 ( .IN0(n2240), .IN1(n2242), .SEL(n2241), .F(n2129) );
  MUX U186 ( .IN0(n2140), .IN1(n2138), .SEL(n2139), .F(n2033) );
  MUX U187 ( .IN0(n2007), .IN1(n2009), .SEL(n2008), .F(n1902) );
  MUX U188 ( .IN0(n1880), .IN1(n1878), .SEL(n1879), .F(n1778) );
  MUX U189 ( .IN0(n1819), .IN1(n1821), .SEL(n1820), .F(n1725) );
  MUX U190 ( .IN0(n1500), .IN1(n1498), .SEL(n1499), .F(n1414) );
  MUX U191 ( .IN0(n1455), .IN1(n1457), .SEL(n1456), .F(n1376) );
  MUX U192 ( .IN0(n1104), .IN1(n1106), .SEL(n1105), .F(n1043) );
  MUX U193 ( .IN0(n56), .IN1(n2636), .SEL(n2637), .F(n2510) );
  IV U194 ( .A(n2638), .Z(n56) );
  MUX U195 ( .IN0(n57), .IN1(n2470), .SEL(n2471), .F(n2349) );
  IV U196 ( .A(n2472), .Z(n57) );
  MUX U197 ( .IN0(n58), .IN1(n1716), .SEL(n1717), .F(n1625) );
  IV U198 ( .A(n1718), .Z(n58) );
  XNOR U199 ( .A(n1728), .B(n1640), .Z(n1644) );
  MUX U200 ( .IN0(n59), .IN1(n1359), .SEL(n1360), .F(n1280) );
  IV U201 ( .A(n1361), .Z(n59) );
  MUX U202 ( .IN0(n60), .IN1(n1367), .SEL(n1368), .F(n1295) );
  IV U203 ( .A(n1369), .Z(n60) );
  MUX U204 ( .IN0(n61), .IN1(n1034), .SEL(n1035), .F(n979) );
  IV U205 ( .A(n1036), .Z(n61) );
  MUX U206 ( .IN0(n1075), .IN1(n1073), .SEL(n1074), .F(n1017) );
  MUX U207 ( .IN0(n803), .IN1(n62), .SEL(n802), .F(n763) );
  IV U208 ( .A(n801), .Z(n62) );
  MUX U209 ( .IN0(n63), .IN1(n3100), .SEL(n3101), .F(n2964) );
  IV U210 ( .A(n3102), .Z(n63) );
  MUX U211 ( .IN0(n2305), .IN1(n2303), .SEL(n2304), .F(n2188) );
  MUX U212 ( .IN0(n64), .IN1(n2206), .SEL(n2207), .F(n2095) );
  IV U213 ( .A(n2208), .Z(n64) );
  MUX U214 ( .IN0(n1149), .IN1(n1151), .SEL(n1150), .F(n1088) );
  MUX U215 ( .IN0(n774), .IN1(n772), .SEL(n773), .F(n739) );
  XNOR U216 ( .A(n715), .B(n714), .Z(n712) );
  MUX U217 ( .IN0(n2414), .IN1(n65), .SEL(n2415), .F(n2299) );
  IV U218 ( .A(n2416), .Z(n65) );
  MUX U219 ( .IN0(n1971), .IN1(n66), .SEL(n1972), .F(n1866) );
  IV U220 ( .A(n1973), .Z(n66) );
  NANDN U221 ( .B(n1769), .A(n1770), .Z(n1675) );
  MUX U222 ( .IN0(n1488), .IN1(n1490), .SEL(n1489), .F(n1404) );
  ANDN U223 ( .A(n1322), .B(n1323), .Z(n1252) );
  AND U224 ( .A(n1060), .B(n1061), .Z(n1006) );
  XNOR U225 ( .A(n878), .B(n877), .Z(n869) );
  OR U226 ( .A(n1014), .B(n1015), .Z(n954) );
  OR U227 ( .A(n788), .B(n789), .Z(n758) );
  XNOR U228 ( .A(n732), .B(n731), .Z(n730) );
  XNOR U229 ( .A(n688), .B(n687), .Z(n679) );
  MUX U230 ( .IN0(n67), .IN1(n3711), .SEL(n3712), .F(n3673) );
  IV U231 ( .A(n3713), .Z(n67) );
  MUX U232 ( .IN0(n68), .IN1(n3724), .SEL(n3725), .F(n3686) );
  IV U233 ( .A(n3726), .Z(n68) );
  MUX U234 ( .IN0(n69), .IN1(n4526), .SEL(n4527), .F(n4513) );
  IV U235 ( .A(n4528), .Z(n69) );
  XNOR U236 ( .A(n4125), .B(n4111), .Z(n4115) );
  MUX U237 ( .IN0(n70), .IN1(n3757), .SEL(n3758), .F(n3719) );
  IV U238 ( .A(n3759), .Z(n70) );
  XNOR U239 ( .A(n3701), .B(n3666), .Z(n3670) );
  MUX U240 ( .IN0(n4517), .IN1(n71), .SEL(n4124), .F(n4504) );
  IV U241 ( .A(n4123), .Z(n71) );
  MUX U242 ( .IN0(n72), .IN1(n4104), .SEL(n3699), .F(n4087) );
  IV U243 ( .A(n3697), .Z(n72) );
  XOR U244 ( .A(n4468), .B(n4469), .Z(n4072) );
  XOR U245 ( .A(n3646), .B(n3611), .Z(n3615) );
  MUX U246 ( .IN0(n4065), .IN1(n4063), .SEL(n4064), .F(n4046) );
  XNOR U247 ( .A(n3587), .B(n3552), .Z(n3556) );
  XOR U248 ( .A(n4444), .B(n4436), .Z(n4022) );
  XOR U249 ( .A(n3532), .B(n3497), .Z(n3501) );
  XOR U250 ( .A(n4270), .B(n4271), .Z(n4280) );
  MUX U251 ( .IN0(n3443), .IN1(n3441), .SEL(n3442), .F(n3403) );
  MUX U252 ( .IN0(n3997), .IN1(n3995), .SEL(n3996), .F(n3978) );
  MUX U253 ( .IN0(n73), .IN1(n3974), .SEL(n3975), .F(n3957) );
  IV U254 ( .A(n3976), .Z(n73) );
  MUX U255 ( .IN0(n4609), .IN1(n74), .SEL(n4287), .F(n4598) );
  IV U256 ( .A(n4285), .Z(n74) );
  MUX U257 ( .IN0(n75), .IN1(n4253), .SEL(n4254), .F(n4232) );
  IV U258 ( .A(n4255), .Z(n75) );
  XOR U259 ( .A(n4971), .B(n4963), .Z(n4831) );
  XOR U260 ( .A(n4837), .B(n4819), .Z(n4823) );
  MUX U261 ( .IN0(n76), .IN1(n4792), .SEL(n4793), .F(n4771) );
  IV U262 ( .A(n4794), .Z(n76) );
  XOR U263 ( .A(n4392), .B(n4384), .Z(n3954) );
  MUX U264 ( .IN0(n77), .IN1(n4776), .SEL(n4777), .F(n4755) );
  IV U265 ( .A(n4778), .Z(n77) );
  XNOR U266 ( .A(n3321), .B(n3286), .Z(n3290) );
  XOR U267 ( .A(n4930), .B(n4931), .Z(n4787) );
  MUX U268 ( .IN0(n3929), .IN1(n3927), .SEL(n3928), .F(n3910) );
  MUX U269 ( .IN0(n3310), .IN1(n3312), .SEL(n3311), .F(n3272) );
  MUX U270 ( .IN0(n4565), .IN1(n78), .SEL(n4203), .F(n4554) );
  IV U271 ( .A(n4201), .Z(n78) );
  MUX U272 ( .IN0(n4194), .IN1(n79), .SEL(n4195), .F(n4173) );
  IV U273 ( .A(n4196), .Z(n79) );
  MUX U274 ( .IN0(n80), .IN1(n3230), .SEL(n3231), .F(n3163) );
  IV U275 ( .A(n3232), .Z(n80) );
  MUX U276 ( .IN0(n81), .IN1(n4345), .SEL(n4346), .F(n3880) );
  IV U277 ( .A(n4347), .Z(n81) );
  MUX U278 ( .IN0(n4706), .IN1(n82), .SEL(n4707), .F(n3093) );
  IV U279 ( .A(n4708), .Z(n82) );
  MUX U280 ( .IN0(n83), .IN1(n3003), .SEL(n3004), .F(n2865) );
  IV U281 ( .A(n3005), .Z(n83) );
  MUX U282 ( .IN0(n84), .IN1(n2839), .SEL(n2840), .F(n2710) );
  IV U283 ( .A(n2841), .Z(n84) );
  MUX U284 ( .IN0(n85), .IN1(n2815), .SEL(n2816), .F(n2686) );
  IV U285 ( .A(n2817), .Z(n85) );
  MUX U286 ( .IN0(n86), .IN1(n2641), .SEL(n2642), .F(n2515) );
  IV U287 ( .A(n2643), .Z(n86) );
  MUX U288 ( .IN0(n87), .IN1(n2923), .SEL(n2924), .F(n2799) );
  IV U289 ( .A(n2925), .Z(n87) );
  MUX U290 ( .IN0(n88), .IN1(n2475), .SEL(n2476), .F(n2354) );
  IV U291 ( .A(n2477), .Z(n88) );
  MUX U292 ( .IN0(n89), .IN1(n2288), .SEL(n2289), .F(n2174) );
  IV U293 ( .A(n2290), .Z(n89) );
  MUX U294 ( .IN0(n90), .IN1(n2337), .SEL(n2338), .F(n2219) );
  IV U295 ( .A(n2339), .Z(n90) );
  MUX U296 ( .IN0(n91), .IN1(n1987), .SEL(n1988), .F(n1882) );
  IV U297 ( .A(n1989), .Z(n91) );
  MUX U298 ( .IN0(n92), .IN1(n1824), .SEL(n1825), .F(n1730) );
  IV U299 ( .A(n1826), .Z(n92) );
  MUX U300 ( .IN0(n93), .IN1(n1774), .SEL(n1775), .F(n1680) );
  IV U301 ( .A(n1776), .Z(n93) );
  MUX U302 ( .IN0(n94), .IN1(n1696), .SEL(n1697), .F(n1605) );
  IV U303 ( .A(n1698), .Z(n94) );
  MUX U304 ( .IN0(n95), .IN1(n1704), .SEL(n1705), .F(n1613) );
  IV U305 ( .A(n1706), .Z(n95) );
  MUX U306 ( .IN0(n96), .IN1(n1343), .SEL(n1344), .F(n1273) );
  IV U307 ( .A(n1345), .Z(n96) );
  MUX U308 ( .IN0(n97), .IN1(n1197), .SEL(n1198), .F(n1134) );
  IV U309 ( .A(n1199), .Z(n97) );
  MUX U310 ( .IN0(n98), .IN1(n888), .SEL(n889), .F(n846) );
  IV U311 ( .A(n890), .Z(n98) );
  MUX U312 ( .IN0(n3134), .IN1(n3136), .SEL(n3135), .F(n2998) );
  MUX U313 ( .IN0(n3117), .IN1(n3119), .SEL(n3118), .F(n2981) );
  MUX U314 ( .IN0(n3048), .IN1(n3046), .SEL(n3047), .F(n2910) );
  MUX U315 ( .IN0(n3883), .IN1(n99), .SEL(n3205), .F(n3080) );
  IV U316 ( .A(n3204), .Z(n99) );
  MUX U317 ( .IN0(n2901), .IN1(n2903), .SEL(n2902), .F(n2772) );
  MUX U318 ( .IN0(n2673), .IN1(n100), .SEL(n2672), .F(n2539) );
  IV U319 ( .A(n2671), .Z(n100) );
  MUX U320 ( .IN0(n2530), .IN1(n2528), .SEL(n2529), .F(n2407) );
  MUX U321 ( .IN0(n2584), .IN1(n2586), .SEL(n2585), .F(n2462) );
  MUX U322 ( .IN0(n2601), .IN1(n2603), .SEL(n2602), .F(n2479) );
  MUX U323 ( .IN0(n2440), .IN1(n2438), .SEL(n2439), .F(n2317) );
  MUX U324 ( .IN0(n2277), .IN1(n2279), .SEL(n2278), .F(n101) );
  IV U325 ( .A(n101), .Z(n2169) );
  MUX U326 ( .IN0(n2071), .IN1(n2069), .SEL(n2070), .F(n1964) );
  XOR U327 ( .A(n2039), .B(n2142), .Z(n2040) );
  MUX U328 ( .IN0(n2024), .IN1(n2026), .SEL(n2025), .F(n1919) );
  MUX U329 ( .IN0(n1902), .IN1(n1904), .SEL(n1903), .F(n1802) );
  MUX U330 ( .IN0(n1595), .IN1(n1593), .SEL(n1594), .F(n1498) );
  MUX U331 ( .IN0(n1517), .IN1(n1519), .SEL(n1518), .F(n102) );
  IV U332 ( .A(n102), .Z(n1438) );
  MUX U333 ( .IN0(n1540), .IN1(n1542), .SEL(n1541), .F(n1455) );
  MUX U334 ( .IN0(n1315), .IN1(n1313), .SEL(n1314), .F(n1243) );
  MUX U335 ( .IN0(n1234), .IN1(n1236), .SEL(n1235), .F(n1166) );
  MUX U336 ( .IN0(n989), .IN1(n991), .SEL(n990), .F(n929) );
  MUX U337 ( .IN0(n1000), .IN1(n998), .SEL(n999), .F(n938) );
  MUX U338 ( .IN0(n2972), .IN1(n103), .SEL(n2973), .F(n2834) );
  IV U339 ( .A(n2974), .Z(n103) );
  MUX U340 ( .IN0(n104), .IN1(n2989), .SEL(n2990), .F(n2851) );
  IV U341 ( .A(n2991), .Z(n104) );
  MUX U342 ( .IN0(n105), .IN1(n2763), .SEL(n2764), .F(n2636) );
  IV U343 ( .A(n2765), .Z(n105) );
  XNOR U344 ( .A(n2734), .B(n2607), .Z(n2613) );
  MUX U345 ( .IN0(n106), .IN1(n2349), .SEL(n2350), .F(n2231) );
  IV U346 ( .A(n2351), .Z(n106) );
  XNOR U347 ( .A(n2082), .B(n1980), .Z(n1984) );
  XNOR U348 ( .A(n2132), .B(n2030), .Z(n2034) );
  MUX U349 ( .IN0(n107), .IN1(n1810), .SEL(n1811), .F(n1716) );
  IV U350 ( .A(n1812), .Z(n107) );
  MUX U351 ( .IN0(n1793), .IN1(n108), .SEL(n1794), .F(n1699) );
  IV U352 ( .A(n1795), .Z(n108) );
  MUX U353 ( .IN0(n109), .IN1(n1429), .SEL(n1430), .F(n1356) );
  IV U354 ( .A(n1431), .Z(n109) );
  MUX U355 ( .IN0(n110), .IN1(n1157), .SEL(n1158), .F(n1095) );
  IV U356 ( .A(n1159), .Z(n110) );
  MUX U357 ( .IN0(n111), .IN1(n876), .SEL(n877), .F(n838) );
  IV U358 ( .A(n878), .Z(n111) );
  XNOR U359 ( .A(n804), .B(n768), .Z(n773) );
  MUX U360 ( .IN0(n112), .IN1(n2697), .SEL(n2698), .F(n2567) );
  IV U361 ( .A(n2699), .Z(n112) );
  MUX U362 ( .IN0(n2552), .IN1(n2550), .SEL(n2551), .F(n2428) );
  MUX U363 ( .IN0(n113), .IN1(n2095), .SEL(n2096), .F(n1990) );
  IV U364 ( .A(n2097), .Z(n113) );
  MUX U365 ( .IN0(n114), .IN1(n1600), .SEL(n1601), .F(n1505) );
  IV U366 ( .A(n1602), .Z(n114) );
  MUX U367 ( .IN0(n1665), .IN1(n1663), .SEL(n1664), .F(n1580) );
  NANDN U368 ( .B(n1218), .A(n1219), .Z(n1213) );
  MUX U369 ( .IN0(n115), .IN1(n1024), .SEL(n1025), .F(n969) );
  IV U370 ( .A(n1026), .Z(n115) );
  MUX U371 ( .IN0(n1019), .IN1(n1017), .SEL(n1018), .F(n964) );
  XNOR U372 ( .A(n741), .B(n740), .Z(n736) );
  ANDN U373 ( .A(n2622), .B(n2621), .Z(n2497) );
  MUX U374 ( .IN0(n2185), .IN1(n116), .SEL(n2186), .F(n2076) );
  IV U375 ( .A(n2187), .Z(n116) );
  NANDN U376 ( .B(n2079), .A(n2080), .Z(n1974) );
  MUX U377 ( .IN0(n1766), .IN1(n117), .SEL(n1767), .F(n1672) );
  IV U378 ( .A(n1768), .Z(n117) );
  NANDN U379 ( .B(n1675), .A(n1676), .Z(n1569) );
  ANDN U380 ( .A(n1652), .B(n1653), .Z(n1560) );
  AND U381 ( .A(n1121), .B(n1122), .Z(n1060) );
  AND U382 ( .A(n902), .B(n903), .Z(n858) );
  XNOR U383 ( .A(n694), .B(n693), .Z(n690) );
  MUX U384 ( .IN0(n1406), .IN1(n1404), .SEL(n1405), .F(n1330) );
  OR U385 ( .A(n1068), .B(n1069), .Z(n1014) );
  OR U386 ( .A(n866), .B(n867), .Z(n827) );
  XNOR U387 ( .A(n791), .B(n790), .Z(n789) );
  MUX U388 ( .IN0(n118), .IN1(n2749), .SEL(n702), .F(n2623) );
  IV U389 ( .A(\_MxM/Y0[3] ), .Z(n118) );
  MUX U390 ( .IN0(n2262), .IN1(n119), .SEL(n661), .F(n2149) );
  IV U391 ( .A(\_MxM/Y0[7] ), .Z(n119) );
  MUX U392 ( .IN0(n1839), .IN1(n120), .SEL(n1840), .F(n1745) );
  IV U393 ( .A(\_MxM/Y0[11] ), .Z(n120) );
  MUX U394 ( .IN0(n1475), .IN1(n121), .SEL(n1476), .F(n1398) );
  IV U395 ( .A(\_MxM/Y0[15] ), .Z(n121) );
  MUX U396 ( .IN0(n122), .IN1(n1185), .SEL(n1186), .F(n1123) );
  IV U397 ( .A(\_MxM/Y0[19] ), .Z(n122) );
  MUX U398 ( .IN0(n123), .IN1(n948), .SEL(n949), .F(n904) );
  IV U399 ( .A(\_MxM/Y0[23] ), .Z(n123) );
  MUX U400 ( .IN0(n124), .IN1(n782), .SEL(n783), .F(n752) );
  IV U401 ( .A(\_MxM/Y0[27] ), .Z(n124) );
  XNOR U402 ( .A(n708), .B(n707), .Z(n726) );
  MUX U403 ( .IN0(n125), .IN1(n3762), .SEL(n3763), .F(n3724) );
  IV U404 ( .A(n3764), .Z(n125) );
  MUX U405 ( .IN0(n126), .IN1(n4118), .SEL(n4119), .F(n4101) );
  IV U406 ( .A(n4120), .Z(n126) );
  MUX U407 ( .IN0(n127), .IN1(n3716), .SEL(n3717), .F(n3678) );
  IV U408 ( .A(n3718), .Z(n127) );
  MUX U409 ( .IN0(n128), .IN1(n3673), .SEL(n3674), .F(n3635) );
  IV U410 ( .A(n3675), .Z(n128) );
  MUX U411 ( .IN0(n129), .IN1(n4513), .SEL(n4514), .F(n4500) );
  IV U412 ( .A(n4515), .Z(n129) );
  MUX U413 ( .IN0(n130), .IN1(n4121), .SEL(n3737), .F(n4104) );
  IV U414 ( .A(n3735), .Z(n130) );
  MUX U415 ( .IN0(n3719), .IN1(n131), .SEL(n3720), .F(n3681) );
  IV U416 ( .A(n3721), .Z(n131) );
  XNOR U417 ( .A(n3663), .B(n3628), .Z(n3632) );
  MUX U418 ( .IN0(n132), .IN1(n4493), .SEL(n4494), .F(n4480) );
  IV U419 ( .A(n4495), .Z(n132) );
  XNOR U420 ( .A(n4091), .B(n4077), .Z(n4081) );
  XOR U421 ( .A(n3684), .B(n3649), .Z(n3653) );
  XOR U422 ( .A(n4483), .B(n4475), .Z(n4073) );
  MUX U423 ( .IN0(n133), .IN1(n4050), .SEL(n4051), .F(n4033) );
  IV U424 ( .A(n4052), .Z(n133) );
  MUX U425 ( .IN0(n134), .IN1(n3521), .SEL(n3522), .F(n3483) );
  IV U426 ( .A(n3523), .Z(n134) );
  XNOR U427 ( .A(n3549), .B(n3514), .Z(n3518) );
  XNOR U428 ( .A(n4040), .B(n4026), .Z(n4030) );
  XOR U429 ( .A(n3570), .B(n3535), .Z(n3539) );
  MUX U430 ( .IN0(n135), .IN1(n4295), .SEL(n4296), .F(n4274) );
  IV U431 ( .A(n4297), .Z(n135) );
  MUX U432 ( .IN0(n4439), .IN1(n136), .SEL(n4022), .F(n4426) );
  IV U433 ( .A(n4021), .Z(n136) );
  MUX U434 ( .IN0(n137), .IN1(n4968), .SEL(n4969), .F(n4955) );
  IV U435 ( .A(n4970), .Z(n137) );
  MUX U436 ( .IN0(n138), .IN1(n4834), .SEL(n4835), .F(n4813) );
  IV U437 ( .A(n4836), .Z(n138) );
  XNOR U438 ( .A(n3435), .B(n3400), .Z(n3404) );
  XOR U439 ( .A(n4603), .B(n4595), .Z(n4266) );
  MUX U440 ( .IN0(n139), .IN1(n4589), .SEL(n4590), .F(n4578) );
  IV U441 ( .A(n4591), .Z(n139) );
  XOR U442 ( .A(n4858), .B(n4840), .Z(n4844) );
  MUX U443 ( .IN0(n140), .IN1(n3369), .SEL(n3370), .F(n3331) );
  IV U444 ( .A(n3371), .Z(n140) );
  XOR U445 ( .A(n3456), .B(n3421), .Z(n3425) );
  MUX U446 ( .IN0(n3980), .IN1(n3978), .SEL(n3979), .F(n3961) );
  MUX U447 ( .IN0(n141), .IN1(n4676), .SEL(n4677), .F(n4661) );
  IV U448 ( .A(n4678), .Z(n141) );
  MUX U449 ( .IN0(n142), .IN1(n4671), .SEL(n4672), .F(n4655) );
  IV U450 ( .A(n4673), .Z(n142) );
  MUX U451 ( .IN0(n4257), .IN1(n143), .SEL(n4258), .F(n4236) );
  IV U452 ( .A(n4259), .Z(n143) );
  MUX U453 ( .IN0(n144), .IN1(n4402), .SEL(n4403), .F(n4389) );
  IV U454 ( .A(n4404), .Z(n144) );
  MUX U455 ( .IN0(n145), .IN1(n5048), .SEL(n5049), .F(n5033) );
  IV U456 ( .A(n5050), .Z(n145) );
  MUX U457 ( .IN0(n146), .IN1(n5043), .SEL(n5044), .F(n5027) );
  IV U458 ( .A(n5045), .Z(n146) );
  XOR U459 ( .A(n4958), .B(n4950), .Z(n4810) );
  MUX U460 ( .IN0(n147), .IN1(n3344), .SEL(n3345), .F(n3306) );
  IV U461 ( .A(n3346), .Z(n147) );
  MUX U462 ( .IN0(n148), .IN1(n3826), .SEL(n3827), .F(n3810) );
  IV U463 ( .A(n3828), .Z(n148) );
  XOR U464 ( .A(n4207), .B(n4208), .Z(n4217) );
  XOR U465 ( .A(n4186), .B(n4187), .Z(n4196) );
  XOR U466 ( .A(n4379), .B(n4371), .Z(n3937) );
  MUX U467 ( .IN0(n149), .IN1(n5153), .SEL(n5154), .F(n5149) );
  IV U468 ( .A(n5155), .Z(n149) );
  MUX U469 ( .IN0(n4780), .IN1(n150), .SEL(n4781), .F(n4759) );
  IV U470 ( .A(n4782), .Z(n150) );
  MUX U471 ( .IN0(n151), .IN1(n4755), .SEL(n4756), .F(n4734) );
  IV U472 ( .A(n4757), .Z(n151) );
  MUX U473 ( .IN0(n3291), .IN1(n3289), .SEL(n3290), .F(n3251) );
  MUX U474 ( .IN0(n152), .IN1(n3914), .SEL(n3915), .F(n3894) );
  IV U475 ( .A(n3916), .Z(n152) );
  XOR U476 ( .A(n4559), .B(n4551), .Z(n4182) );
  MUX U477 ( .IN0(n153), .IN1(n4545), .SEL(n4546), .F(n4534) );
  IV U478 ( .A(n4547), .Z(n153) );
  XOR U479 ( .A(n4165), .B(n4166), .Z(n4175) );
  MUX U480 ( .IN0(n154), .IN1(n4169), .SEL(n4170), .F(n4144) );
  IV U481 ( .A(n4171), .Z(n154) );
  MUX U482 ( .IN0(n155), .IN1(n4903), .SEL(n4904), .F(n4717) );
  IV U483 ( .A(n4905), .Z(n155) );
  XOR U484 ( .A(n4919), .B(n4911), .Z(n4747) );
  MUX U485 ( .IN0(n156), .IN1(n3209), .SEL(n3210), .F(n3172) );
  IV U486 ( .A(n3211), .Z(n156) );
  XNOR U487 ( .A(n3921), .B(n3907), .Z(n3911) );
  MUX U488 ( .IN0(n3272), .IN1(n3274), .SEL(n3273), .F(n3234) );
  MUX U489 ( .IN0(n157), .IN1(n3163), .SEL(n3164), .F(n3033) );
  IV U490 ( .A(n3165), .Z(n157) );
  MUX U491 ( .IN0(n158), .IN1(n2914), .SEL(n2915), .F(n2785) );
  IV U492 ( .A(n2916), .Z(n158) );
  MUX U493 ( .IN0(n159), .IN1(n2931), .SEL(n2932), .F(n2803) );
  IV U494 ( .A(n2933), .Z(n159) );
  MUX U495 ( .IN0(n160), .IN1(n2823), .SEL(n2824), .F(n2694) );
  IV U496 ( .A(n2825), .Z(n160) );
  MUX U497 ( .IN0(n161), .IN1(n2856), .SEL(n2857), .F(n2727) );
  IV U498 ( .A(n2858), .Z(n161) );
  MUX U499 ( .IN0(n162), .IN1(n2650), .SEL(n2651), .F(n2524) );
  IV U500 ( .A(n2652), .Z(n162) );
  MUX U501 ( .IN0(n163), .IN1(n2736), .SEL(n2737), .F(n2606) );
  IV U502 ( .A(n2738), .Z(n163) );
  MUX U503 ( .IN0(n164), .IN1(n2313), .SEL(n2314), .F(n2195) );
  IV U504 ( .A(n2315), .Z(n164) );
  MUX U505 ( .IN0(n165), .IN1(n2174), .SEL(n2175), .F(n2065) );
  IV U506 ( .A(n2176), .Z(n165) );
  MUX U507 ( .IN0(n166), .IN1(n2228), .SEL(n2229), .F(n2117) );
  IV U508 ( .A(n2230), .Z(n166) );
  MUX U509 ( .IN0(n167), .IN1(n2108), .SEL(n2109), .F(n2003) );
  IV U510 ( .A(n2110), .Z(n167) );
  MUX U511 ( .IN0(n168), .IN1(n2020), .SEL(n2021), .F(n1915) );
  IV U512 ( .A(n2022), .Z(n168) );
  MUX U513 ( .IN0(n169), .IN1(n1613), .SEL(n1614), .F(n1523) );
  IV U514 ( .A(n1615), .Z(n169) );
  MUX U515 ( .IN0(n170), .IN1(n1460), .SEL(n1461), .F(n1381) );
  IV U516 ( .A(n1462), .Z(n170) );
  MUX U517 ( .IN0(n171), .IN1(n1265), .SEL(n1266), .F(n1197) );
  IV U518 ( .A(n1267), .Z(n171) );
  MUX U519 ( .IN0(n172), .IN1(n1171), .SEL(n1172), .F(n1109) );
  IV U520 ( .A(n1173), .Z(n172) );
  MUX U521 ( .IN0(n173), .IN1(n1180), .SEL(n1181), .F(n1118) );
  IV U522 ( .A(n1182), .Z(n173) );
  MUX U523 ( .IN0(n174), .IN1(n1039), .SEL(n1040), .F(n985) );
  IV U524 ( .A(n1041), .Z(n174) );
  MUX U525 ( .IN0(n3898), .IN1(n4334), .SEL(n3899), .F(n175) );
  IV U526 ( .A(n175), .Z(n3083) );
  XNOR U527 ( .A(n4700), .B(n3090), .Z(n3094) );
  XNOR U528 ( .A(n3186), .B(n3060), .Z(n3064) );
  MUX U529 ( .IN0(n2981), .IN1(n2983), .SEL(n2982), .F(n2843) );
  MUX U530 ( .IN0(n2998), .IN1(n3000), .SEL(n2999), .F(n2860) );
  MUX U531 ( .IN0(n2772), .IN1(n2774), .SEL(n2773), .F(n2645) );
  MUX U532 ( .IN0(n2409), .IN1(n2407), .SEL(n2408), .F(n2292) );
  MUX U533 ( .IN0(n2479), .IN1(n2481), .SEL(n2480), .F(n2358) );
  MUX U534 ( .IN0(n2462), .IN1(n2464), .SEL(n2463), .F(n2341) );
  MUX U535 ( .IN0(n2285), .IN1(n176), .SEL(n2284), .F(n2168) );
  IV U536 ( .A(n2283), .Z(n176) );
  MUX U537 ( .IN0(n2090), .IN1(n2088), .SEL(n2089), .F(n1983) );
  MUX U538 ( .IN0(n1966), .IN1(n1964), .SEL(n1965), .F(n1851) );
  MUX U539 ( .IN0(n1802), .IN1(n1804), .SEL(n1803), .F(n1708) );
  MUX U540 ( .IN0(n1725), .IN1(n1727), .SEL(n1726), .F(n1634) );
  MUX U541 ( .IN0(n1416), .IN1(n1414), .SEL(n1415), .F(n1339) );
  MUX U542 ( .IN0(n1376), .IN1(n1378), .SEL(n1377), .F(n1304) );
  MUX U543 ( .IN0(n1245), .IN1(n1243), .SEL(n1244), .F(n1175) );
  MUX U544 ( .IN0(n940), .IN1(n938), .SEL(n939), .F(n892) );
  MUX U545 ( .IN0(n929), .IN1(n931), .SEL(n930), .F(n881) );
  MUX U546 ( .IN0(n177), .IN1(n846), .SEL(n847), .F(n807) );
  IV U547 ( .A(n848), .Z(n177) );
  XNOR U548 ( .A(n3137), .B(n3004), .Z(n3008) );
  XNOR U549 ( .A(n3040), .B(n2907), .Z(n2911) );
  MUX U550 ( .IN0(n178), .IN1(n3028), .SEL(n3029), .F(n2892) );
  IV U551 ( .A(n3030), .Z(n178) );
  MUX U552 ( .IN0(n2949), .IN1(n179), .SEL(n2948), .F(n2809) );
  IV U553 ( .A(n2947), .Z(n179) );
  MUX U554 ( .IN0(n2834), .IN1(n180), .SEL(n2835), .F(n2705) );
  IV U555 ( .A(n2836), .Z(n180) );
  XNOR U556 ( .A(n2813), .B(n2687), .Z(n2691) );
  MUX U557 ( .IN0(n181), .IN1(n2851), .SEL(n2852), .F(n2722) );
  IV U558 ( .A(n2853), .Z(n181) );
  MUX U559 ( .IN0(n2541), .IN1(n2539), .SEL(n2540), .F(n2427) );
  XNOR U560 ( .A(n2482), .B(n2364), .Z(n2368) );
  MUX U561 ( .IN0(n2332), .IN1(n182), .SEL(n2333), .F(n2214) );
  IV U562 ( .A(n2334), .Z(n182) );
  MUX U563 ( .IN0(n183), .IN1(n2231), .SEL(n2232), .F(n2120) );
  IV U564 ( .A(n2233), .Z(n183) );
  MUX U565 ( .IN0(n2057), .IN1(n184), .SEL(n2058), .F(n1955) );
  IV U566 ( .A(n2059), .Z(n184) );
  XNOR U567 ( .A(n2027), .B(n1925), .Z(n1929) );
  MUX U568 ( .IN0(n1893), .IN1(n185), .SEL(n1894), .F(n1793) );
  IV U569 ( .A(n1895), .Z(n185) );
  XNOR U570 ( .A(n1772), .B(n1681), .Z(n1685) );
  MUX U571 ( .IN0(n186), .IN1(n1625), .SEL(n1626), .F(n1531) );
  IV U572 ( .A(n1627), .Z(n186) );
  XOR U573 ( .A(n1427), .B(n1428), .Z(n1440) );
  MUX U574 ( .IN0(n1289), .IN1(n187), .SEL(n1288), .F(n1215) );
  IV U575 ( .A(n1287), .Z(n187) );
  MUX U576 ( .IN0(n188), .IN1(n1295), .SEL(n1296), .F(n1225) );
  IV U577 ( .A(n1297), .Z(n188) );
  XNOR U578 ( .A(n1133), .B(n1076), .Z(n1074) );
  MUX U579 ( .IN0(n189), .IN1(n838), .SEL(n839), .F(n801) );
  IV U580 ( .A(n840), .Z(n189) );
  AND U581 ( .A(n798), .B(n794), .Z(n797) );
  MUX U582 ( .IN0(n190), .IN1(n816), .SEL(n817), .F(n777) );
  IV U583 ( .A(n818), .Z(n190) );
  MUX U584 ( .IN0(n191), .IN1(n2806), .SEL(n2807), .F(n2680) );
  IV U585 ( .A(n2808), .Z(n191) );
  MUX U586 ( .IN0(n192), .IN1(n2567), .SEL(n2568), .F(n2445) );
  IV U587 ( .A(n2569), .Z(n192) );
  MUX U588 ( .IN0(n193), .IN1(n1990), .SEL(n1991), .F(n1885) );
  IV U589 ( .A(n1992), .Z(n193) );
  MUX U590 ( .IN0(n194), .IN1(n1421), .SEL(n1422), .F(n1346) );
  IV U591 ( .A(n1423), .Z(n194) );
  MUX U592 ( .IN0(n195), .IN1(n1146), .SEL(n1147), .F(n1083) );
  IV U593 ( .A(n1148), .Z(n195) );
  MUX U594 ( .IN0(n196), .IN1(n1021), .SEL(n1022), .F(n966) );
  IV U595 ( .A(n1023), .Z(n196) );
  XNOR U596 ( .A(n766), .B(n742), .Z(n740) );
  MUX U597 ( .IN0(n2917), .IN1(n197), .SEL(n2918), .F(n2788) );
  IV U598 ( .A(n2919), .Z(n197) );
  XNOR U599 ( .A(n2512), .B(n2511), .Z(n2552) );
  ANDN U600 ( .A(n2497), .B(n2498), .Z(n2376) );
  MUX U601 ( .IN0(n2299), .IN1(n198), .SEL(n2300), .F(n2185) );
  IV U602 ( .A(n2301), .Z(n198) );
  ANDN U603 ( .A(n2042), .B(n2043), .Z(n1937) );
  MUX U604 ( .IN0(n199), .IN1(n1585), .SEL(n1584), .F(n1488) );
  IV U605 ( .A(n1583), .Z(n199) );
  NOR U606 ( .A(n1486), .B(n1487), .Z(n1485) );
  ANDN U607 ( .A(n1473), .B(n1474), .Z(n1396) );
  AND U608 ( .A(n1183), .B(n1184), .Z(n1121) );
  AND U609 ( .A(n858), .B(n859), .Z(n819) );
  XOR U610 ( .A(n1869), .B(n1866), .Z(n1944) );
  OR U611 ( .A(n1260), .B(n1261), .Z(n1191) );
  XNOR U612 ( .A(n1026), .B(n1025), .Z(n1015) );
  XNOR U613 ( .A(n973), .B(n972), .Z(n955) );
  OR U614 ( .A(n827), .B(n828), .Z(n788) );
  XNOR U615 ( .A(n761), .B(n760), .Z(n759) );
  MUX U616 ( .IN0(n200), .IN1(n2623), .SEL(n664), .F(n2499) );
  IV U617 ( .A(\_MxM/Y0[4] ), .Z(n200) );
  MUX U618 ( .IN0(n2149), .IN1(n201), .SEL(n660), .F(n2044) );
  IV U619 ( .A(\_MxM/Y0[8] ), .Z(n201) );
  MUX U620 ( .IN0(n1745), .IN1(n202), .SEL(n1746), .F(n1654) );
  IV U621 ( .A(\_MxM/Y0[12] ), .Z(n202) );
  MUX U622 ( .IN0(n1398), .IN1(n203), .SEL(n1399), .F(n1324) );
  IV U623 ( .A(\_MxM/Y0[16] ), .Z(n203) );
  MUX U624 ( .IN0(n204), .IN1(n1123), .SEL(n1124), .F(n1062) );
  IV U625 ( .A(\_MxM/Y0[20] ), .Z(n204) );
  MUX U626 ( .IN0(n205), .IN1(n904), .SEL(n905), .F(n860) );
  IV U627 ( .A(\_MxM/Y0[24] ), .Z(n205) );
  MUX U628 ( .IN0(n206), .IN1(n752), .SEL(n753), .F(n723) );
  IV U629 ( .A(\_MxM/Y0[28] ), .Z(n206) );
  AND U630 ( .A(n695), .B(n696), .Z(n691) );
  MUX U631 ( .IN0(n207), .IN1(n3741), .SEL(n3742), .F(n3703) );
  IV U632 ( .A(n3743), .Z(n207) );
  MUX U633 ( .IN0(n208), .IN1(n3754), .SEL(n3755), .F(n3716) );
  IV U634 ( .A(n3756), .Z(n208) );
  MUX U635 ( .IN0(n209), .IN1(n4519), .SEL(n4520), .F(n4506) );
  IV U636 ( .A(n4521), .Z(n209) );
  MUX U637 ( .IN0(n3671), .IN1(n3669), .SEL(n3670), .F(n3631) );
  MUX U638 ( .IN0(n210), .IN1(n3769), .SEL(n3184), .F(n3731) );
  IV U639 ( .A(n3183), .Z(n210) );
  MUX U640 ( .IN0(n211), .IN1(n4084), .SEL(n4085), .F(n4067) );
  IV U641 ( .A(n4086), .Z(n211) );
  MUX U642 ( .IN0(n212), .IN1(n4076), .SEL(n4077), .F(n4059) );
  IV U643 ( .A(n4078), .Z(n212) );
  MUX U644 ( .IN0(n3690), .IN1(n3692), .SEL(n3691), .F(n3652) );
  MUX U645 ( .IN0(n4504), .IN1(n213), .SEL(n4107), .F(n4491) );
  IV U646 ( .A(n4106), .Z(n213) );
  MUX U647 ( .IN0(n214), .IN1(n3589), .SEL(n3590), .F(n3551) );
  IV U648 ( .A(n3591), .Z(n214) );
  MUX U649 ( .IN0(n215), .IN1(n3602), .SEL(n3603), .F(n3564) );
  IV U650 ( .A(n3604), .Z(n215) );
  MUX U651 ( .IN0(n216), .IN1(n3610), .SEL(n3611), .F(n3572) );
  IV U652 ( .A(n3612), .Z(n216) );
  MUX U653 ( .IN0(n217), .IN1(n4087), .SEL(n3661), .F(n4070) );
  IV U654 ( .A(n3659), .Z(n217) );
  MUX U655 ( .IN0(n4048), .IN1(n4046), .SEL(n4047), .F(n4029) );
  MUX U656 ( .IN0(n3605), .IN1(n218), .SEL(n3606), .F(n3567) );
  IV U657 ( .A(n3607), .Z(n218) );
  MUX U658 ( .IN0(n219), .IN1(n4454), .SEL(n4455), .F(n4441) );
  IV U659 ( .A(n4456), .Z(n219) );
  MUX U660 ( .IN0(n3519), .IN1(n3517), .SEL(n3518), .F(n3479) );
  MUX U661 ( .IN0(n220), .IN1(n4008), .SEL(n4009), .F(n3991) );
  IV U662 ( .A(n4010), .Z(n220) );
  MUX U663 ( .IN0(n3538), .IN1(n3540), .SEL(n3539), .F(n3500) );
  MUX U664 ( .IN0(n221), .IN1(n4611), .SEL(n4612), .F(n4600) );
  IV U665 ( .A(n4613), .Z(n221) );
  MUX U666 ( .IN0(n222), .IN1(n4981), .SEL(n4982), .F(n4968) );
  IV U667 ( .A(n4983), .Z(n222) );
  MUX U668 ( .IN0(n223), .IN1(n3437), .SEL(n3438), .F(n3399) );
  IV U669 ( .A(n3439), .Z(n223) );
  MUX U670 ( .IN0(n224), .IN1(n4448), .SEL(n4449), .F(n4435) );
  IV U671 ( .A(n4450), .Z(n224) );
  MUX U672 ( .IN0(n225), .IN1(n3450), .SEL(n3451), .F(n3412) );
  IV U673 ( .A(n3452), .Z(n225) );
  MUX U674 ( .IN0(n226), .IN1(n3458), .SEL(n3459), .F(n3420) );
  IV U675 ( .A(n3460), .Z(n226) );
  MUX U676 ( .IN0(n227), .IN1(n4605), .SEL(n4606), .F(n4594) );
  IV U677 ( .A(n4607), .Z(n227) );
  MUX U678 ( .IN0(n228), .IN1(n4839), .SEL(n4840), .F(n4818) );
  IV U679 ( .A(n4841), .Z(n228) );
  MUX U680 ( .IN0(n229), .IN1(n4019), .SEL(n3509), .F(n4002) );
  IV U681 ( .A(n3507), .Z(n229) );
  XOR U682 ( .A(n4293), .B(n4275), .Z(n4279) );
  XOR U683 ( .A(n4249), .B(n4250), .Z(n4259) );
  XOR U684 ( .A(n4418), .B(n4410), .Z(n3988) );
  MUX U685 ( .IN0(n3453), .IN1(n230), .SEL(n3454), .F(n3415) );
  IV U686 ( .A(n3455), .Z(n230) );
  MUX U687 ( .IN0(n4598), .IN1(n231), .SEL(n4266), .F(n4587) );
  IV U688 ( .A(n4264), .Z(n231) );
  XOR U689 ( .A(n4228), .B(n4229), .Z(n4238) );
  MUX U690 ( .IN0(n232), .IN1(n4232), .SEL(n4233), .F(n4211) );
  IV U691 ( .A(n4234), .Z(n232) );
  MUX U692 ( .IN0(n4966), .IN1(n233), .SEL(n4831), .F(n4953) );
  IV U693 ( .A(n4829), .Z(n233) );
  MUX U694 ( .IN0(n234), .IN1(n4949), .SEL(n4950), .F(n4936) );
  IV U695 ( .A(n4951), .Z(n234) );
  MUX U696 ( .IN0(n4822), .IN1(n235), .SEL(n4823), .F(n4801) );
  IV U697 ( .A(n4824), .Z(n235) );
  MUX U698 ( .IN0(n3367), .IN1(n3365), .SEL(n3366), .F(n3327) );
  XNOR U699 ( .A(n3972), .B(n3958), .Z(n3962) );
  MUX U700 ( .IN0(n236), .IN1(n3948), .SEL(n3949), .F(n3931) );
  IV U701 ( .A(n3950), .Z(n236) );
  MUX U702 ( .IN0(n3386), .IN1(n3388), .SEL(n3387), .F(n3348) );
  MUX U703 ( .IN0(n237), .IN1(n4326), .SEL(n4327), .F(n4665) );
  IV U704 ( .A(n4679), .Z(n237) );
  MUX U705 ( .IN0(n4655), .IN1(n4670), .SEL(n4657), .F(n4639) );
  MUX U706 ( .IN0(n238), .IN1(n5138), .SEL(n5139), .F(n5121) );
  IV U707 ( .A(n5140), .Z(n238) );
  MUX U708 ( .IN0(n239), .IN1(n4891), .SEL(n4892), .F(n5037) );
  IV U709 ( .A(n5051), .Z(n239) );
  MUX U710 ( .IN0(n5027), .IN1(n5042), .SEL(n5029), .F(n5011) );
  MUX U711 ( .IN0(n240), .IN1(n4929), .SEL(n4930), .F(n4916) );
  IV U712 ( .A(n4931), .Z(n240) );
  XOR U713 ( .A(n4772), .B(n4773), .Z(n4782) );
  MUX U714 ( .IN0(n241), .IN1(n3285), .SEL(n3286), .F(n3247) );
  IV U715 ( .A(n3287), .Z(n241) );
  MUX U716 ( .IN0(n242), .IN1(n3306), .SEL(n3307), .F(n3268) );
  IV U717 ( .A(n3308), .Z(n242) );
  MUX U718 ( .IN0(n243), .IN1(n3779), .SEL(n3780), .F(n3820) );
  IV U719 ( .A(n3834), .Z(n243) );
  MUX U720 ( .IN0(n3810), .IN1(n3825), .SEL(n3812), .F(n3794) );
  MUX U721 ( .IN0(n244), .IN1(n4376), .SEL(n4377), .F(n4363) );
  IV U722 ( .A(n4378), .Z(n244) );
  MUX U723 ( .IN0(n5115), .IN1(n5130), .SEL(n5117), .F(n5097) );
  XOR U724 ( .A(n4751), .B(n4752), .Z(n4761) );
  MUX U725 ( .IN0(n245), .IN1(n4383), .SEL(n4384), .F(n4370) );
  IV U726 ( .A(n4385), .Z(n245) );
  MUX U727 ( .IN0(n246), .IN1(n3951), .SEL(n3357), .F(n3934) );
  IV U728 ( .A(n3355), .Z(n246) );
  MUX U729 ( .IN0(n247), .IN1(n3906), .SEL(n3907), .F(n3886) );
  IV U730 ( .A(n3908), .Z(n247) );
  MUX U731 ( .IN0(n248), .IN1(n4550), .SEL(n4551), .F(n4539) );
  IV U732 ( .A(n4552), .Z(n248) );
  XOR U733 ( .A(n4730), .B(n4731), .Z(n4740) );
  MUX U734 ( .IN0(n249), .IN1(n4734), .SEL(n4735), .F(n4702) );
  IV U735 ( .A(n4736), .Z(n249) );
  MUX U736 ( .IN0(n3912), .IN1(n3910), .SEL(n3911), .F(n3890) );
  MUX U737 ( .IN0(n3301), .IN1(n250), .SEL(n3302), .F(n3263) );
  IV U738 ( .A(n3303), .Z(n250) );
  MUX U739 ( .IN0(n4554), .IN1(n251), .SEL(n4182), .F(n4543) );
  IV U740 ( .A(n4180), .Z(n251) );
  XOR U741 ( .A(n4188), .B(n4170), .Z(n4174) );
  XOR U742 ( .A(n4153), .B(n4154), .Z(n4150) );
  MUX U743 ( .IN0(n5166), .IN1(n5169), .SEL(n5167), .F(n3139) );
  MUX U744 ( .IN0(n4914), .IN1(n252), .SEL(n4747), .F(n4901) );
  IV U745 ( .A(n4745), .Z(n252) );
  XOR U746 ( .A(n4711), .B(n4712), .Z(n4708) );
  MUX U747 ( .IN0(n3215), .IN1(n3213), .SEL(n3214), .F(n3176) );
  MUX U748 ( .IN0(n3234), .IN1(n3236), .SEL(n3235), .F(n3167) );
  MUX U749 ( .IN0(n253), .IN1(n3113), .SEL(n3114), .F(n2977) );
  IV U750 ( .A(n3115), .Z(n253) );
  MUX U751 ( .IN0(n254), .IN1(n3042), .SEL(n3043), .F(n2906) );
  IV U752 ( .A(n3044), .Z(n254) );
  MUX U753 ( .IN0(n255), .IN1(n3025), .SEL(n3026), .F(n2889) );
  IV U754 ( .A(n3027), .Z(n255) );
  MUX U755 ( .IN0(n256), .IN1(n3033), .SEL(n3034), .F(n2897) );
  IV U756 ( .A(n3035), .Z(n256) );
  MUX U757 ( .IN0(n257), .IN1(n3902), .SEL(n3903), .F(n4334) );
  IV U758 ( .A(n4348), .Z(n257) );
  MUX U759 ( .IN0(n258), .IN1(n2719), .SEL(n2720), .F(n2589) );
  IV U760 ( .A(n2721), .Z(n258) );
  MUX U761 ( .IN0(n259), .IN1(n2694), .SEL(n2695), .F(n2564) );
  IV U762 ( .A(n2696), .Z(n259) );
  MUX U763 ( .IN0(n260), .IN1(n2532), .SEL(n2533), .F(n2411) );
  IV U764 ( .A(n2534), .Z(n260) );
  MUX U765 ( .IN0(n261), .IN1(n2515), .SEL(n2516), .F(n2394) );
  IV U766 ( .A(n2517), .Z(n261) );
  MUX U767 ( .IN0(n262), .IN1(n2450), .SEL(n2451), .F(n2329) );
  IV U768 ( .A(n2452), .Z(n262) );
  MUX U769 ( .IN0(n263), .IN1(n2458), .SEL(n2459), .F(n2337) );
  IV U770 ( .A(n2460), .Z(n263) );
  MUX U771 ( .IN0(n264), .IN1(n2354), .SEL(n2355), .F(n2236) );
  IV U772 ( .A(n2356), .Z(n264) );
  MUX U773 ( .IN0(n265), .IN1(n2203), .SEL(n2204), .F(n2092) );
  IV U774 ( .A(n2205), .Z(n265) );
  MUX U775 ( .IN0(n266), .IN1(n2195), .SEL(n2196), .F(n2084) );
  IV U776 ( .A(n2197), .Z(n266) );
  MUX U777 ( .IN0(n267), .IN1(n2003), .SEL(n2004), .F(n1898) );
  IV U778 ( .A(n2005), .Z(n267) );
  MUX U779 ( .IN0(n268), .IN1(n1915), .SEL(n1916), .F(n1815) );
  IV U780 ( .A(n1917), .Z(n268) );
  MUX U781 ( .IN0(n269), .IN1(n1807), .SEL(n1808), .F(n1713) );
  IV U782 ( .A(n1809), .Z(n269) );
  MUX U783 ( .IN0(n270), .IN1(n1782), .SEL(n1783), .F(n1688) );
  IV U784 ( .A(n1784), .Z(n270) );
  MUX U785 ( .IN0(n271), .IN1(n1968), .SEL(n1969), .F(n1863) );
  IV U786 ( .A(n1970), .Z(n271) );
  MUX U787 ( .IN0(n272), .IN1(n1960), .SEL(n1961), .F(n1859) );
  IV U788 ( .A(n1962), .Z(n272) );
  MUX U789 ( .IN0(n273), .IN1(n1418), .SEL(n1419), .F(n1343) );
  IV U790 ( .A(n1420), .Z(n273) );
  MUX U791 ( .IN0(n274), .IN1(n1230), .SEL(n1231), .F(n1162) );
  IV U792 ( .A(n1232), .Z(n274) );
  MUX U793 ( .IN0(n275), .IN1(n1154), .SEL(n1155), .F(n1092) );
  IV U794 ( .A(n1156), .Z(n275) );
  MUX U795 ( .IN0(n276), .IN1(n1109), .SEL(n1110), .F(n1048) );
  IV U796 ( .A(n1111), .Z(n276) );
  MUX U797 ( .IN0(n277), .IN1(n1057), .SEL(n1058), .F(n1003) );
  IV U798 ( .A(n1059), .Z(n277) );
  MUX U799 ( .IN0(n278), .IN1(n985), .SEL(n986), .F(n924) );
  IV U800 ( .A(n987), .Z(n278) );
  MUX U801 ( .IN0(n279), .IN1(n917), .SEL(n918), .F(n873) );
  IV U802 ( .A(n919), .Z(n279) );
  XOR U803 ( .A(n3078), .B(n3079), .Z(n3085) );
  MUX U804 ( .IN0(n2795), .IN1(n2793), .SEL(n2794), .F(n2671) );
  XOR U805 ( .A(n2746), .B(n2873), .Z(n2747) );
  MUX U806 ( .IN0(n2645), .IN1(n2647), .SEL(n2646), .F(n2519) );
  MUX U807 ( .IN0(n2714), .IN1(n2716), .SEL(n2715), .F(n2584) );
  MUX U808 ( .IN0(n2180), .IN1(n2178), .SEL(n2179), .F(n2069) );
  MUX U809 ( .IN0(n2223), .IN1(n2225), .SEL(n2224), .F(n2112) );
  MUX U810 ( .IN0(n2171), .IN1(n280), .SEL(n2170), .F(n2060) );
  IV U811 ( .A(n2169), .Z(n280) );
  MUX U812 ( .IN0(n2129), .IN1(n2131), .SEL(n2130), .F(n2024) );
  XOR U813 ( .A(n1649), .B(n1738), .Z(n1650) );
  MUX U814 ( .IN0(n1708), .IN1(n1710), .SEL(n1709), .F(n1617) );
  XNOR U815 ( .A(n1851), .B(n1852), .Z(n1850) );
  MUX U816 ( .IN0(n1271), .IN1(n1269), .SEL(n1270), .F(n1201) );
  MUX U817 ( .IN0(n1304), .IN1(n1306), .SEL(n1305), .F(n1234) );
  MUX U818 ( .IN0(n1043), .IN1(n1045), .SEL(n1044), .F(n989) );
  MUX U819 ( .IN0(n1136), .IN1(n281), .SEL(n1135), .F(n1076) );
  IV U820 ( .A(n1134), .Z(n281) );
  MUX U821 ( .IN0(n282), .IN1(n1143), .SEL(n1144), .F(n1080) );
  IV U822 ( .A(n1145), .Z(n282) );
  XOR U823 ( .A(n3128), .B(n2995), .Z(n2999) );
  XNOR U824 ( .A(n2951), .B(n2816), .Z(n2820) );
  XNOR U825 ( .A(n3001), .B(n2866), .Z(n2870) );
  MUX U826 ( .IN0(n283), .IN1(n2892), .SEL(n2893), .F(n2763) );
  IV U827 ( .A(n2894), .Z(n283) );
  XNOR U828 ( .A(n2775), .B(n2651), .Z(n2655) );
  MUX U829 ( .IN0(n2575), .IN1(n284), .SEL(n2576), .F(n2453) );
  IV U830 ( .A(n2577), .Z(n284) );
  XNOR U831 ( .A(n2554), .B(n2435), .Z(n2439) );
  XNOR U832 ( .A(n2604), .B(n2485), .Z(n2489) );
  MUX U833 ( .IN0(n285), .IN1(n2592), .SEL(n2593), .F(n2470) );
  IV U834 ( .A(n2594), .Z(n285) );
  MUX U835 ( .IN0(n286), .IN1(n2389), .SEL(n2390), .F(n2273) );
  IV U836 ( .A(n2391), .Z(n286) );
  XNOR U837 ( .A(n2243), .B(n2135), .Z(n2139) );
  MUX U838 ( .IN0(n2103), .IN1(n287), .SEL(n2104), .F(n1998) );
  IV U839 ( .A(n2105), .Z(n287) );
  MUX U840 ( .IN0(n288), .IN1(n2015), .SEL(n2016), .F(n1910) );
  IV U841 ( .A(n2017), .Z(n288) );
  XNOR U842 ( .A(n1977), .B(n1875), .Z(n1879) );
  MUX U843 ( .IN0(n1955), .IN1(n289), .SEL(n1956), .F(n1846) );
  IV U844 ( .A(n1957), .Z(n289) );
  XNOR U845 ( .A(n1822), .B(n1731), .Z(n1735) );
  XOR U846 ( .A(n1719), .B(n1631), .Z(n1635) );
  MUX U847 ( .IN0(n1608), .IN1(n290), .SEL(n1609), .F(n1513) );
  IV U848 ( .A(n1610), .Z(n290) );
  XNOR U849 ( .A(n1587), .B(n1495), .Z(n1499) );
  MUX U850 ( .IN0(n291), .IN1(n1531), .SEL(n1532), .F(n1446) );
  IV U851 ( .A(n1533), .Z(n291) );
  XNOR U852 ( .A(n1543), .B(n1461), .Z(n1465) );
  XNOR U853 ( .A(n1359), .B(n1432), .Z(n1360) );
  NAND U854 ( .A(n1286), .B(n1351), .Z(n1350) );
  MUX U855 ( .IN0(n292), .IN1(n1225), .SEL(n1226), .F(n1157) );
  IV U856 ( .A(n1227), .Z(n292) );
  MUX U857 ( .IN0(n293), .IN1(n979), .SEL(n980), .F(n920) );
  IV U858 ( .A(n981), .Z(n293) );
  XNOR U859 ( .A(n992), .B(n935), .Z(n939) );
  MUX U860 ( .IN0(n841), .IN1(n843), .SEL(n842), .F(n294) );
  IV U861 ( .A(n294), .Z(n794) );
  MUX U862 ( .IN0(n295), .IN1(n3070), .SEL(n3071), .F(n2934) );
  IV U863 ( .A(n3072), .Z(n295) );
  XNOR U864 ( .A(n3127), .B(n3126), .Z(n3102) );
  MUX U865 ( .IN0(n296), .IN1(n2324), .SEL(n2325), .F(n2206) );
  IV U866 ( .A(n2326), .Z(n296) );
  MUX U867 ( .IN0(n297), .IN1(n1785), .SEL(n1786), .F(n1691) );
  IV U868 ( .A(n1787), .Z(n297) );
  MUX U869 ( .IN0(n298), .IN1(n1346), .SEL(n1347), .F(n1276) );
  IV U870 ( .A(n1348), .Z(n298) );
  ANDN U871 ( .A(n960), .B(n961), .Z(n959) );
  XNOR U872 ( .A(n852), .B(n851), .Z(n840) );
  XNOR U873 ( .A(n813), .B(n812), .Z(n803) );
  MUX U874 ( .IN0(n2788), .IN1(n299), .SEL(n2789), .F(n2661) );
  IV U875 ( .A(n2790), .Z(n299) );
  XNOR U876 ( .A(n2550), .B(n2549), .Z(n2664) );
  XOR U877 ( .A(n2302), .B(n2188), .Z(n2189) );
  ANDN U878 ( .A(n2376), .B(n2377), .Z(n2260) );
  MUX U879 ( .IN0(n2076), .IN1(n300), .SEL(n2077), .F(n1971) );
  IV U880 ( .A(n2078), .Z(n300) );
  ANDN U881 ( .A(n1560), .B(n1561), .Z(n1473) );
  ANDN U882 ( .A(n1252), .B(n1253), .Z(n1183) );
  XOR U883 ( .A(n1088), .B(n1083), .Z(n1132) );
  AND U884 ( .A(n1006), .B(n1007), .Z(n946) );
  AND U885 ( .A(n819), .B(n820), .Z(n780) );
  OR U886 ( .A(n742), .B(n743), .Z(n737) );
  XOR U887 ( .A(n1675), .B(n1672), .Z(n1751) );
  XNOR U888 ( .A(n1404), .B(n1486), .Z(n1481) );
  OR U889 ( .A(n1191), .B(n1192), .Z(n1130) );
  OR U890 ( .A(n954), .B(n955), .Z(n910) );
  XNOR U891 ( .A(n869), .B(n868), .Z(n867) );
  ANDN U892 ( .A(n688), .B(n687), .Z(n686) );
  OR U893 ( .A(n729), .B(n730), .Z(n707) );
  MUX U894 ( .IN0(n2499), .IN1(n301), .SEL(n663), .F(n2378) );
  IV U895 ( .A(\_MxM/Y0[5] ), .Z(n301) );
  MUX U896 ( .IN0(n2044), .IN1(n302), .SEL(n659), .F(n1939) );
  IV U897 ( .A(\_MxM/Y0[9] ), .Z(n302) );
  MUX U898 ( .IN0(n1654), .IN1(n303), .SEL(n1655), .F(n1562) );
  IV U899 ( .A(\_MxM/Y0[13] ), .Z(n303) );
  MUX U900 ( .IN0(n1324), .IN1(n304), .SEL(n1325), .F(n1254) );
  IV U901 ( .A(\_MxM/Y0[17] ), .Z(n304) );
  MUX U902 ( .IN0(n305), .IN1(n1062), .SEL(n1063), .F(n1008) );
  IV U903 ( .A(\_MxM/Y0[21] ), .Z(n305) );
  MUX U904 ( .IN0(n306), .IN1(n860), .SEL(n861), .F(n821) );
  IV U905 ( .A(\_MxM/Y0[25] ), .Z(n306) );
  MUX U906 ( .IN0(\_MxM/Y0[29] ), .IN1(n307), .SEL(n724), .F(n701) );
  IV U907 ( .A(n723), .Z(n307) );
  NAND U908 ( .A(n676), .B(n677), .Z(n675) );
  MUX U909 ( .IN0(n308), .IN1(n4135), .SEL(n4136), .F(n4118) );
  IV U910 ( .A(n4137), .Z(n308) );
  MUX U911 ( .IN0(n3709), .IN1(n3707), .SEL(n3708), .F(n3669) );
  MUX U912 ( .IN0(n309), .IN1(n4138), .SEL(n3772), .F(n4121) );
  IV U913 ( .A(n3771), .Z(n309) );
  MUX U914 ( .IN0(n3728), .IN1(n3730), .SEL(n3729), .F(n3690) );
  XOR U915 ( .A(n4494), .B(n4495), .Z(n4106) );
  MUX U916 ( .IN0(n310), .IN1(n3635), .SEL(n3636), .F(n3597) );
  IV U917 ( .A(n3637), .Z(n310) );
  MUX U918 ( .IN0(n311), .IN1(n3627), .SEL(n3628), .F(n3589) );
  IV U919 ( .A(n3629), .Z(n311) );
  MUX U920 ( .IN0(n4099), .IN1(n4097), .SEL(n4098), .F(n4080) );
  MUX U921 ( .IN0(n312), .IN1(n3648), .SEL(n3649), .F(n3610) );
  IV U922 ( .A(n3650), .Z(n312) );
  XOR U923 ( .A(n4481), .B(n4482), .Z(n4089) );
  MUX U924 ( .IN0(n313), .IN1(n4500), .SEL(n4501), .F(n4487) );
  IV U925 ( .A(n4502), .Z(n313) );
  MUX U926 ( .IN0(n314), .IN1(n4059), .SEL(n4060), .F(n4042) );
  IV U927 ( .A(n4061), .Z(n314) );
  MUX U928 ( .IN0(n3643), .IN1(n315), .SEL(n3644), .F(n3605) );
  IV U929 ( .A(n3645), .Z(n315) );
  MUX U930 ( .IN0(n3557), .IN1(n3555), .SEL(n3556), .F(n3517) );
  MUX U931 ( .IN0(n316), .IN1(n4070), .SEL(n3623), .F(n4053) );
  IV U932 ( .A(n3621), .Z(n316) );
  MUX U933 ( .IN0(n3576), .IN1(n3578), .SEL(n3577), .F(n3538) );
  MUX U934 ( .IN0(n317), .IN1(n3483), .SEL(n3484), .F(n3445) );
  IV U935 ( .A(n3485), .Z(n317) );
  MUX U936 ( .IN0(n318), .IN1(n3475), .SEL(n3476), .F(n3437) );
  IV U937 ( .A(n3477), .Z(n318) );
  MUX U938 ( .IN0(n319), .IN1(n4016), .SEL(n4017), .F(n3999) );
  IV U939 ( .A(n4018), .Z(n319) );
  MUX U940 ( .IN0(n320), .IN1(n4290), .SEL(n4291), .F(n4269) );
  IV U941 ( .A(n4292), .Z(n320) );
  MUX U942 ( .IN0(n321), .IN1(n4616), .SEL(n4617), .F(n4605) );
  IV U943 ( .A(n4618), .Z(n321) );
  MUX U944 ( .IN0(n4452), .IN1(n322), .SEL(n4039), .F(n4439) );
  IV U945 ( .A(n4038), .Z(n322) );
  MUX U946 ( .IN0(n323), .IN1(n4988), .SEL(n4989), .F(n4975) );
  IV U947 ( .A(n4990), .Z(n323) );
  XNOR U948 ( .A(n4023), .B(n4009), .Z(n4013) );
  MUX U949 ( .IN0(n324), .IN1(n4435), .SEL(n4436), .F(n4422) );
  IV U950 ( .A(n4437), .Z(n324) );
  MUX U951 ( .IN0(n3491), .IN1(n325), .SEL(n3492), .F(n3453) );
  IV U952 ( .A(n3493), .Z(n325) );
  MUX U953 ( .IN0(n326), .IN1(n4302), .SEL(n3877), .F(n4281) );
  IV U954 ( .A(n3876), .Z(n326) );
  MUX U955 ( .IN0(n327), .IN1(n4415), .SEL(n4416), .F(n4402) );
  IV U956 ( .A(n4417), .Z(n327) );
  MUX U957 ( .IN0(n328), .IN1(n4867), .SEL(n4714), .F(n4846) );
  IV U958 ( .A(n4713), .Z(n328) );
  MUX U959 ( .IN0(n4843), .IN1(n329), .SEL(n4844), .F(n4822) );
  IV U960 ( .A(n4845), .Z(n329) );
  MUX U961 ( .IN0(n3405), .IN1(n3403), .SEL(n3404), .F(n3365) );
  MUX U962 ( .IN0(n330), .IN1(n4002), .SEL(n3471), .F(n3985) );
  IV U963 ( .A(n3469), .Z(n330) );
  MUX U964 ( .IN0(n3424), .IN1(n3426), .SEL(n3425), .F(n3386) );
  MUX U965 ( .IN0(n331), .IN1(n3382), .SEL(n3383), .F(n3344) );
  IV U966 ( .A(n3384), .Z(n331) );
  XOR U967 ( .A(n4592), .B(n4584), .Z(n4245) );
  XOR U968 ( .A(n4956), .B(n4957), .Z(n4829) );
  XOR U969 ( .A(n4793), .B(n4794), .Z(n4803) );
  MUX U970 ( .IN0(n332), .IN1(n4797), .SEL(n4798), .F(n4776) );
  IV U971 ( .A(n4799), .Z(n332) );
  MUX U972 ( .IN0(n333), .IN1(n3331), .SEL(n3332), .F(n3293) );
  IV U973 ( .A(n3333), .Z(n333) );
  MUX U974 ( .IN0(n334), .IN1(n3323), .SEL(n3324), .F(n3285) );
  IV U975 ( .A(n3325), .Z(n334) );
  MUX U976 ( .IN0(n3963), .IN1(n3961), .SEL(n3962), .F(n3944) );
  MUX U977 ( .IN0(n335), .IN1(n3940), .SEL(n3941), .F(n3923) );
  IV U978 ( .A(n3942), .Z(n335) );
  MUX U979 ( .IN0(n336), .IN1(n3831), .SEL(n3832), .F(n3816) );
  IV U980 ( .A(n3833), .Z(n336) );
  MUX U981 ( .IN0(n337), .IN1(n4206), .SEL(n4207), .F(n4185) );
  IV U982 ( .A(n4208), .Z(n337) );
  MUX U983 ( .IN0(n4661), .IN1(n4675), .SEL(n4663), .F(n4645) );
  MUX U984 ( .IN0(n338), .IN1(n4691), .SEL(n4692), .F(n4687) );
  IV U985 ( .A(n4693), .Z(n338) );
  XOR U986 ( .A(n4251), .B(n4233), .Z(n4237) );
  MUX U987 ( .IN0(n339), .IN1(n4567), .SEL(n4568), .F(n4556) );
  IV U988 ( .A(n4569), .Z(n339) );
  MUX U989 ( .IN0(n5033), .IN1(n5047), .SEL(n5035), .F(n5017) );
  MUX U990 ( .IN0(n340), .IN1(n5063), .SEL(n5064), .F(n5059) );
  IV U991 ( .A(n5065), .Z(n340) );
  XOR U992 ( .A(n4943), .B(n4944), .Z(n4808) );
  MUX U993 ( .IN0(n341), .IN1(n4936), .SEL(n4937), .F(n4923) );
  IV U994 ( .A(n4938), .Z(n341) );
  MUX U995 ( .IN0(n342), .IN1(n3298), .SEL(n3299), .F(n3260) );
  IV U996 ( .A(n3300), .Z(n342) );
  MUX U997 ( .IN0(n343), .IN1(n3847), .SEL(n3848), .F(n3843) );
  IV U998 ( .A(n3849), .Z(n343) );
  MUX U999 ( .IN0(n344), .IN1(n4312), .SEL(n4313), .F(n4308) );
  IV U1000 ( .A(n4314), .Z(n344) );
  MUX U1001 ( .IN0(n345), .IN1(n4561), .SEL(n4562), .F(n4550) );
  IV U1002 ( .A(n4563), .Z(n345) );
  MUX U1003 ( .IN0(n4387), .IN1(n346), .SEL(n3954), .F(n4374) );
  IV U1004 ( .A(n3953), .Z(n346) );
  MUX U1005 ( .IN0(n347), .IN1(n5078), .SEL(n5079), .F(n5125) );
  IV U1006 ( .A(n5141), .Z(n347) );
  MUX U1007 ( .IN0(n348), .IN1(n4877), .SEL(n4878), .F(n4873) );
  IV U1008 ( .A(n4879), .Z(n348) );
  MUX U1009 ( .IN0(n349), .IN1(n4916), .SEL(n4917), .F(n4903) );
  IV U1010 ( .A(n4918), .Z(n349) );
  MUX U1011 ( .IN0(n3339), .IN1(n350), .SEL(n3340), .F(n3301) );
  IV U1012 ( .A(n3341), .Z(n350) );
  MUX U1013 ( .IN0(n351), .IN1(n4363), .SEL(n4364), .F(n4350) );
  IV U1014 ( .A(n4365), .Z(n351) );
  MUX U1015 ( .IN0(n5097), .IN1(n5112), .SEL(n5099), .F(n5084) );
  MUX U1016 ( .IN0(n352), .IN1(n4370), .SEL(n4371), .F(n4357) );
  IV U1017 ( .A(n4372), .Z(n352) );
  MUX U1018 ( .IN0(n353), .IN1(n3934), .SEL(n3319), .F(n3917) );
  IV U1019 ( .A(n3317), .Z(n353) );
  XOR U1020 ( .A(n3304), .B(n3269), .Z(n3273) );
  XNOR U1021 ( .A(n3253), .B(n3252), .Z(n3265) );
  MUX U1022 ( .IN0(n3858), .IN1(n3861), .SEL(n3859), .F(n3741) );
  MUX U1023 ( .IN0(n354), .IN1(n4144), .SEL(n4145), .F(n4127) );
  IV U1024 ( .A(n4146), .Z(n354) );
  MUX U1025 ( .IN0(n4173), .IN1(n355), .SEL(n4174), .F(n4148) );
  IV U1026 ( .A(n4175), .Z(n355) );
  MUX U1027 ( .IN0(n5074), .IN1(n5102), .SEL(n5076), .F(n3122) );
  MUX U1028 ( .IN0(n4738), .IN1(n356), .SEL(n4739), .F(n4706) );
  IV U1029 ( .A(n4740), .Z(n356) );
  MUX U1030 ( .IN0(n357), .IN1(n4702), .SEL(n4703), .F(n3089) );
  IV U1031 ( .A(n4704), .Z(n357) );
  MUX U1032 ( .IN0(n358), .IN1(n3196), .SEL(n3197), .F(n3067) );
  IV U1033 ( .A(n3198), .Z(n358) );
  XNOR U1034 ( .A(n3904), .B(n3887), .Z(n3891) );
  XNOR U1035 ( .A(n3215), .B(n3214), .Z(n3227) );
  MUX U1036 ( .IN0(n4543), .IN1(n359), .SEL(n4161), .F(n4530) );
  IV U1037 ( .A(n4159), .Z(n359) );
  MUX U1038 ( .IN0(n360), .IN1(n3139), .SEL(n3140), .F(n3003) );
  IV U1039 ( .A(n3141), .Z(n360) );
  MUX U1040 ( .IN0(n361), .IN1(n3097), .SEL(n3098), .F(n2961) );
  IV U1041 ( .A(n3099), .Z(n361) );
  MUX U1042 ( .IN0(n362), .IN1(n3059), .SEL(n3060), .F(n2923) );
  IV U1043 ( .A(n3061), .Z(n362) );
  NAND U1044 ( .A(n4333), .B(n4337), .Z(n4336) );
  XNOR U1045 ( .A(n5171), .B(n5172), .Z(n3143) );
  MUX U1046 ( .IN0(n4901), .IN1(n363), .SEL(n4726), .F(n3117) );
  IV U1047 ( .A(n4724), .Z(n363) );
  MUX U1048 ( .IN0(n364), .IN1(n2969), .SEL(n2970), .F(n2831) );
  IV U1049 ( .A(n2971), .Z(n364) );
  MUX U1050 ( .IN0(n365), .IN1(n2977), .SEL(n2978), .F(n2839) );
  IV U1051 ( .A(n2979), .Z(n365) );
  MUX U1052 ( .IN0(n366), .IN1(n2889), .SEL(n2890), .F(n2760) );
  IV U1053 ( .A(n2891), .Z(n366) );
  MUX U1054 ( .IN0(n367), .IN1(n2777), .SEL(n2778), .F(n2650) );
  IV U1055 ( .A(n2779), .Z(n367) );
  MUX U1056 ( .IN0(n368), .IN1(n2727), .SEL(n2728), .F(n2597) );
  IV U1057 ( .A(n2729), .Z(n368) );
  MUX U1058 ( .IN0(n369), .IN1(n2564), .SEL(n2565), .F(n2442) );
  IV U1059 ( .A(n2566), .Z(n369) );
  MUX U1060 ( .IN0(n370), .IN1(n2386), .SEL(n2387), .F(n2270) );
  IV U1061 ( .A(n2388), .Z(n370) );
  MUX U1062 ( .IN0(n371), .IN1(n2411), .SEL(n2412), .F(n2296) );
  IV U1063 ( .A(n2413), .Z(n371) );
  MUX U1064 ( .IN0(n372), .IN1(n2675), .SEL(n2676), .F(n2545) );
  IV U1065 ( .A(n2677), .Z(n372) );
  MUX U1066 ( .IN0(n373), .IN1(n2394), .SEL(n2395), .F(n2283) );
  IV U1067 ( .A(n2396), .Z(n373) );
  MUX U1068 ( .IN0(n374), .IN1(n2236), .SEL(n2237), .F(n2125) );
  IV U1069 ( .A(n2238), .Z(n374) );
  MUX U1070 ( .IN0(n375), .IN1(n2100), .SEL(n2101), .F(n1995) );
  IV U1071 ( .A(n2102), .Z(n375) );
  MUX U1072 ( .IN0(n376), .IN1(n2092), .SEL(n2093), .F(n1987) );
  IV U1073 ( .A(n2094), .Z(n376) );
  MUX U1074 ( .IN0(n377), .IN1(n1898), .SEL(n1899), .F(n1798) );
  IV U1075 ( .A(n1900), .Z(n377) );
  MUX U1076 ( .IN0(n378), .IN1(n1874), .SEL(n1875), .F(n1774) );
  IV U1077 ( .A(n1876), .Z(n378) );
  MUX U1078 ( .IN0(n379), .IN1(n1815), .SEL(n1816), .F(n1721) );
  IV U1079 ( .A(n1817), .Z(n379) );
  MUX U1080 ( .IN0(n380), .IN1(n1688), .SEL(n1689), .F(n1597) );
  IV U1081 ( .A(n1690), .Z(n380) );
  MUX U1082 ( .IN0(n381), .IN1(n1605), .SEL(n1606), .F(n1510) );
  IV U1083 ( .A(n1607), .Z(n381) );
  MUX U1084 ( .IN0(n382), .IN1(n1443), .SEL(n1444), .F(n1364) );
  IV U1085 ( .A(n1445), .Z(n382) );
  MUX U1086 ( .IN0(n383), .IN1(n1372), .SEL(n1373), .F(n1300) );
  IV U1087 ( .A(n1374), .Z(n383) );
  MUX U1088 ( .IN0(n384), .IN1(n1309), .SEL(n1310), .F(n1239) );
  IV U1089 ( .A(n1311), .Z(n384) );
  MUX U1090 ( .IN0(n385), .IN1(n1100), .SEL(n1101), .F(n1039) );
  IV U1091 ( .A(n1102), .Z(n385) );
  MUX U1092 ( .IN0(n386), .IN1(n1048), .SEL(n1049), .F(n994) );
  IV U1093 ( .A(n1050), .Z(n386) );
  MUX U1094 ( .IN0(n387), .IN1(n1003), .SEL(n1004), .F(n943) );
  IV U1095 ( .A(n1005), .Z(n387) );
  XOR U1096 ( .A(n3013), .B(n3147), .Z(n3014) );
  XOR U1097 ( .A(n3161), .B(n3034), .Z(n3038) );
  MUX U1098 ( .IN0(n2912), .IN1(n2910), .SEL(n2911), .F(n2781) );
  MUX U1099 ( .IN0(n3079), .IN1(n388), .SEL(n3078), .F(n2941) );
  IV U1100 ( .A(n3077), .Z(n388) );
  MUX U1101 ( .IN0(n2860), .IN1(n2862), .SEL(n2861), .F(n2731) );
  XOR U1102 ( .A(n2494), .B(n2616), .Z(n2495) );
  MUX U1103 ( .IN0(n2358), .IN1(n2360), .SEL(n2359), .F(n2240) );
  XOR U1104 ( .A(n1834), .B(n1932), .Z(n1835) );
  MUX U1105 ( .IN0(n1919), .IN1(n1921), .SEL(n1920), .F(n1819) );
  MUX U1106 ( .IN0(n389), .IN1(n1863), .SEL(n1864), .F(n1763) );
  IV U1107 ( .A(n1865), .Z(n389) );
  MUX U1108 ( .IN0(n1341), .IN1(n1339), .SEL(n1340), .F(n1269) );
  MUX U1109 ( .IN0(n1177), .IN1(n1175), .SEL(n1176), .F(n1113) );
  MUX U1110 ( .IN0(n1166), .IN1(n1168), .SEL(n1167), .F(n1104) );
  MUX U1111 ( .IN0(n3108), .IN1(n390), .SEL(n3109), .F(n2972) );
  IV U1112 ( .A(n3110), .Z(n390) );
  MUX U1113 ( .IN0(n391), .IN1(n3080), .SEL(n3081), .F(n2947) );
  IV U1114 ( .A(n3082), .Z(n391) );
  XOR U1115 ( .A(n2766), .B(n2642), .Z(n2646) );
  NAND U1116 ( .A(n2670), .B(n2797), .Z(n2796) );
  XNOR U1117 ( .A(n2863), .B(n2737), .Z(n2741) );
  XNOR U1118 ( .A(n2684), .B(n2557), .Z(n2561) );
  XOR U1119 ( .A(n2708), .B(n2581), .Z(n2585) );
  XNOR U1120 ( .A(n2522), .B(n2404), .Z(n2408) );
  MUX U1121 ( .IN0(n2453), .IN1(n392), .SEL(n2454), .F(n2332) );
  IV U1122 ( .A(n2455), .Z(n392) );
  MUX U1123 ( .IN0(n393), .IN1(n2273), .SEL(n2274), .F(n2160) );
  IV U1124 ( .A(n2275), .Z(n393) );
  XOR U1125 ( .A(n2335), .B(n2220), .Z(n2224) );
  XNOR U1126 ( .A(n2311), .B(n2196), .Z(n2200) );
  XNOR U1127 ( .A(n2361), .B(n2248), .Z(n2252) );
  MUX U1128 ( .IN0(n2062), .IN1(n2060), .SEL(n2061), .F(n394) );
  IV U1129 ( .A(n394), .Z(n1954) );
  XNOR U1130 ( .A(n2063), .B(n1961), .Z(n1965) );
  MUX U1131 ( .IN0(n395), .IN1(n2120), .SEL(n2121), .F(n2015) );
  IV U1132 ( .A(n2122), .Z(n395) );
  MUX U1133 ( .IN0(n1998), .IN1(n396), .SEL(n1999), .F(n1893) );
  IV U1134 ( .A(n2000), .Z(n396) );
  NAND U1135 ( .A(n1759), .B(n1857), .Z(n1856) );
  XNOR U1136 ( .A(n1922), .B(n1825), .Z(n1829) );
  XNOR U1137 ( .A(n1678), .B(n1590), .Z(n1594) );
  XOR U1138 ( .A(n1702), .B(n1614), .Z(n1618) );
  XOR U1139 ( .A(n1628), .B(n1537), .Z(n1541) );
  XNOR U1140 ( .A(n1637), .B(n1546), .Z(n1552) );
  MUX U1141 ( .IN0(n1513), .IN1(n397), .SEL(n1514), .F(n1429) );
  IV U1142 ( .A(n1515), .Z(n397) );
  XOR U1143 ( .A(n1354), .B(n1355), .Z(n1361) );
  MUX U1144 ( .IN0(n398), .IN1(n1446), .SEL(n1447), .F(n1367) );
  IV U1145 ( .A(n1448), .Z(n398) );
  MUX U1146 ( .IN0(n1217), .IN1(n1215), .SEL(n1216), .F(n1149) );
  OR U1147 ( .A(n1076), .B(n1077), .Z(n1071) );
  MUX U1148 ( .IN0(n399), .IN1(n1080), .SEL(n1081), .F(n1021) );
  IV U1149 ( .A(n1082), .Z(n399) );
  XOR U1150 ( .A(n982), .B(n925), .Z(n930) );
  XNOR U1151 ( .A(n932), .B(n889), .Z(n895) );
  MUX U1152 ( .IN0(n400), .IN1(n2964), .SEL(n2965), .F(n2826) );
  IV U1153 ( .A(n2966), .Z(n400) );
  XNOR U1154 ( .A(n2871), .B(n2870), .Z(n2853) );
  MUX U1155 ( .IN0(n401), .IN1(n2934), .SEL(n2935), .F(n2806) );
  IV U1156 ( .A(n2936), .Z(n401) );
  MUX U1157 ( .IN0(n402), .IN1(n1885), .SEL(n1886), .F(n1785) );
  IV U1158 ( .A(n1887), .Z(n402) );
  MUX U1159 ( .IN0(n403), .IN1(n1276), .SEL(n1277), .F(n1210) );
  IV U1160 ( .A(n1278), .Z(n403) );
  XOR U1161 ( .A(n763), .B(n799), .Z(n792) );
  MUX U1162 ( .IN0(n769), .IN1(n404), .SEL(n768), .F(n742) );
  IV U1163 ( .A(n767), .Z(n404) );
  MUX U1164 ( .IN0(n2661), .IN1(n405), .SEL(n2662), .F(n2535) );
  IV U1165 ( .A(n2663), .Z(n405) );
  XNOR U1166 ( .A(n2594), .B(n2593), .Z(n2569) );
  XNOR U1167 ( .A(n2428), .B(n2422), .Z(n2538) );
  ANDN U1168 ( .A(n2260), .B(n2261), .Z(n2147) );
  NANDN U1169 ( .B(n1869), .A(n1870), .Z(n1769) );
  ANDN U1170 ( .A(n1837), .B(n1838), .Z(n1743) );
  ANDN U1171 ( .A(n1396), .B(n1397), .Z(n1322) );
  XNOR U1172 ( .A(n1036), .B(n1035), .Z(n1026) );
  AND U1173 ( .A(n946), .B(n947), .Z(n902) );
  MUX U1174 ( .IN0(n406), .IN1(n747), .SEL(n748), .F(n718) );
  IV U1175 ( .A(n749), .Z(n406) );
  AND U1176 ( .A(n750), .B(n751), .Z(n721) );
  XOR U1177 ( .A(n2079), .B(n2076), .Z(n2154) );
  XNOR U1178 ( .A(n1693), .B(n1692), .Z(n1674) );
  OR U1179 ( .A(n1330), .B(n1331), .Z(n1260) );
  XNOR U1180 ( .A(n1148), .B(n1147), .Z(n1131) );
  XNOR U1181 ( .A(n1087), .B(n1086), .Z(n1069) );
  OR U1182 ( .A(n910), .B(n911), .Z(n866) );
  XNOR U1183 ( .A(n832), .B(n829), .Z(n828) );
  ANDN U1184 ( .A(n690), .B(n689), .Z(n685) );
  MUX U1185 ( .IN0(n407), .IN1(n2878), .SEL(n1125), .F(n2749) );
  IV U1186 ( .A(\_MxM/Y0[2] ), .Z(n407) );
  MUX U1187 ( .IN0(n2378), .IN1(n408), .SEL(n662), .F(n2262) );
  IV U1188 ( .A(\_MxM/Y0[6] ), .Z(n408) );
  MUX U1189 ( .IN0(n1939), .IN1(n409), .SEL(n658), .F(n1839) );
  IV U1190 ( .A(\_MxM/Y0[10] ), .Z(n409) );
  MUX U1191 ( .IN0(n1562), .IN1(n410), .SEL(n1563), .F(n1475) );
  IV U1192 ( .A(\_MxM/Y0[14] ), .Z(n410) );
  MUX U1193 ( .IN0(n1254), .IN1(n411), .SEL(n1255), .F(n1185) );
  IV U1194 ( .A(\_MxM/Y0[18] ), .Z(n411) );
  MUX U1195 ( .IN0(n412), .IN1(n1008), .SEL(n1009), .F(n948) );
  IV U1196 ( .A(\_MxM/Y0[22] ), .Z(n412) );
  MUX U1197 ( .IN0(n413), .IN1(n821), .SEL(n822), .F(n782) );
  IV U1198 ( .A(\_MxM/Y0[26] ), .Z(n413) );
  OR U1199 ( .A(n707), .B(n708), .Z(n678) );
  MUX U1200 ( .IN0(n414), .IN1(n4110), .SEL(n4111), .F(n4093) );
  IV U1201 ( .A(n4112), .Z(n414) );
  XNOR U1202 ( .A(n3739), .B(n3704), .Z(n3708) );
  XOR U1203 ( .A(n3760), .B(n3725), .Z(n3729) );
  MUX U1204 ( .IN0(n415), .IN1(n3678), .SEL(n3679), .F(n3640) );
  IV U1205 ( .A(n3680), .Z(n415) );
  MUX U1206 ( .IN0(n416), .IN1(n4067), .SEL(n4068), .F(n4050) );
  IV U1207 ( .A(n4069), .Z(n416) );
  MUX U1208 ( .IN0(n4082), .IN1(n4080), .SEL(n4081), .F(n4063) );
  XNOR U1209 ( .A(n3625), .B(n3590), .Z(n3594) );
  MUX U1210 ( .IN0(n4491), .IN1(n417), .SEL(n4090), .F(n4478) );
  IV U1211 ( .A(n4089), .Z(n417) );
  MUX U1212 ( .IN0(n418), .IN1(n3559), .SEL(n3560), .F(n3521) );
  IV U1213 ( .A(n3561), .Z(n418) );
  MUX U1214 ( .IN0(n419), .IN1(n4487), .SEL(n4488), .F(n4474) );
  IV U1215 ( .A(n4489), .Z(n419) );
  MUX U1216 ( .IN0(n420), .IN1(n4042), .SEL(n4043), .F(n4025) );
  IV U1217 ( .A(n4044), .Z(n420) );
  MUX U1218 ( .IN0(n3614), .IN1(n3616), .SEL(n3615), .F(n3576) );
  MUX U1219 ( .IN0(n421), .IN1(n4467), .SEL(n4468), .F(n4454) );
  IV U1220 ( .A(n4469), .Z(n421) );
  MUX U1221 ( .IN0(n422), .IN1(n3526), .SEL(n3527), .F(n3488) );
  IV U1222 ( .A(n3528), .Z(n422) );
  MUX U1223 ( .IN0(n423), .IN1(n3534), .SEL(n3535), .F(n3496) );
  IV U1224 ( .A(n3536), .Z(n423) );
  MUX U1225 ( .IN0(n424), .IN1(n4053), .SEL(n3585), .F(n4036) );
  IV U1226 ( .A(n3583), .Z(n424) );
  MUX U1227 ( .IN0(n3567), .IN1(n425), .SEL(n3568), .F(n3529) );
  IV U1228 ( .A(n3569), .Z(n425) );
  XOR U1229 ( .A(n4429), .B(n4430), .Z(n4021) );
  MUX U1230 ( .IN0(n426), .IN1(n4855), .SEL(n4856), .F(n4834) );
  IV U1231 ( .A(n4857), .Z(n426) );
  MUX U1232 ( .IN0(n427), .IN1(n4860), .SEL(n4861), .F(n4839) );
  IV U1233 ( .A(n4862), .Z(n427) );
  MUX U1234 ( .IN0(n428), .IN1(n3999), .SEL(n4000), .F(n3982) );
  IV U1235 ( .A(n4001), .Z(n428) );
  XNOR U1236 ( .A(n3473), .B(n3438), .Z(n3442) );
  MUX U1237 ( .IN0(n429), .IN1(n4269), .SEL(n4270), .F(n4248) );
  IV U1238 ( .A(n4271), .Z(n429) );
  XOR U1239 ( .A(n4614), .B(n4606), .Z(n4287) );
  MUX U1240 ( .IN0(n430), .IN1(n4274), .SEL(n4275), .F(n4253) );
  IV U1241 ( .A(n4276), .Z(n430) );
  XOR U1242 ( .A(n4416), .B(n4417), .Z(n4004) );
  MUX U1243 ( .IN0(n4992), .IN1(n431), .SEL(n4870), .F(n4979) );
  IV U1244 ( .A(n4869), .Z(n431) );
  MUX U1245 ( .IN0(n432), .IN1(n3407), .SEL(n3408), .F(n3369) );
  IV U1246 ( .A(n3409), .Z(n432) );
  XNOR U1247 ( .A(n4006), .B(n3992), .Z(n3996) );
  MUX U1248 ( .IN0(n3462), .IN1(n3464), .SEL(n3463), .F(n3424) );
  MUX U1249 ( .IN0(n433), .IN1(n4955), .SEL(n4956), .F(n4942) );
  IV U1250 ( .A(n4957), .Z(n433) );
  MUX U1251 ( .IN0(n434), .IN1(n4962), .SEL(n4963), .F(n4949) );
  IV U1252 ( .A(n4964), .Z(n434) );
  MUX U1253 ( .IN0(n435), .IN1(n4422), .SEL(n4423), .F(n4409) );
  IV U1254 ( .A(n4424), .Z(n435) );
  MUX U1255 ( .IN0(n436), .IN1(n3374), .SEL(n3375), .F(n3336) );
  IV U1256 ( .A(n3376), .Z(n436) );
  MUX U1257 ( .IN0(n437), .IN1(n4583), .SEL(n4584), .F(n4572) );
  IV U1258 ( .A(n4585), .Z(n437) );
  XOR U1259 ( .A(n4590), .B(n4591), .Z(n4264) );
  MUX U1260 ( .IN0(n438), .IN1(n3985), .SEL(n3433), .F(n3968) );
  IV U1261 ( .A(n3431), .Z(n438) );
  MUX U1262 ( .IN0(n3415), .IN1(n439), .SEL(n3416), .F(n3377) );
  IV U1263 ( .A(n3417), .Z(n439) );
  XNOR U1264 ( .A(n3359), .B(n3324), .Z(n3328) );
  XOR U1265 ( .A(n4579), .B(n4580), .Z(n4243) );
  MUX U1266 ( .IN0(n4236), .IN1(n440), .SEL(n4237), .F(n4215) );
  IV U1267 ( .A(n4238), .Z(n440) );
  MUX U1268 ( .IN0(n441), .IN1(n4389), .SEL(n4390), .F(n4376) );
  IV U1269 ( .A(n4391), .Z(n441) );
  MUX U1270 ( .IN0(n442), .IN1(n5133), .SEL(n5134), .F(n5115) );
  IV U1271 ( .A(n5135), .Z(n442) );
  XOR U1272 ( .A(n4816), .B(n4798), .Z(n4802) );
  MUX U1273 ( .IN0(n443), .IN1(n4771), .SEL(n4772), .F(n4750) );
  IV U1274 ( .A(n4773), .Z(n443) );
  XNOR U1275 ( .A(n3955), .B(n3941), .Z(n3945) );
  MUX U1276 ( .IN0(n444), .IN1(n3931), .SEL(n3932), .F(n3914) );
  IV U1277 ( .A(n3933), .Z(n444) );
  MUX U1278 ( .IN0(n3816), .IN1(n3830), .SEL(n3818), .F(n3800) );
  MUX U1279 ( .IN0(n445), .IN1(n4185), .SEL(n4186), .F(n4164) );
  IV U1280 ( .A(n4187), .Z(n445) );
  MUX U1281 ( .IN0(n4645), .IN1(n4660), .SEL(n4647), .F(n4622) );
  MUX U1282 ( .IN0(n4639), .IN1(n4654), .SEL(n4641), .F(n4628) );
  XOR U1283 ( .A(n4568), .B(n4569), .Z(n4222) );
  MUX U1284 ( .IN0(n446), .IN1(n4190), .SEL(n4191), .F(n4169) );
  IV U1285 ( .A(n4192), .Z(n446) );
  MUX U1286 ( .IN0(n5017), .IN1(n5032), .SEL(n5019), .F(n4994) );
  MUX U1287 ( .IN0(n5011), .IN1(n5026), .SEL(n5013), .F(n5000) );
  MUX U1288 ( .IN0(n4940), .IN1(n447), .SEL(n4789), .F(n4927) );
  IV U1289 ( .A(n4787), .Z(n447) );
  MUX U1290 ( .IN0(n448), .IN1(n3255), .SEL(n3256), .F(n3217) );
  IV U1291 ( .A(n3257), .Z(n448) );
  XOR U1292 ( .A(n3342), .B(n3307), .Z(n3311) );
  MUX U1293 ( .IN0(n3794), .IN1(n3809), .SEL(n3796), .F(n3783) );
  MUX U1294 ( .IN0(n449), .IN1(n3862), .SEL(n3863), .F(n3858) );
  IV U1295 ( .A(n3864), .Z(n449) );
  XNOR U1296 ( .A(n4692), .B(n4693), .Z(n4679) );
  XOR U1297 ( .A(n4557), .B(n4558), .Z(n4201) );
  NOR U1298 ( .A(g_input[0]), .B(n5182), .Z(n5175) );
  MUX U1299 ( .IN0(n4374), .IN1(n450), .SEL(n3937), .F(n4361) );
  IV U1300 ( .A(n3936), .Z(n450) );
  MUX U1301 ( .IN0(n5103), .IN1(n5120), .SEL(n5105), .F(n5074) );
  XNOR U1302 ( .A(n5064), .B(n5065), .Z(n5051) );
  MUX U1303 ( .IN0(n451), .IN1(n4910), .SEL(n4911), .F(n4897) );
  IV U1304 ( .A(n4912), .Z(n451) );
  MUX U1305 ( .IN0(n452), .IN1(n3222), .SEL(n3223), .F(n3155) );
  IV U1306 ( .A(n3224), .Z(n452) );
  XNOR U1307 ( .A(n3245), .B(n3210), .Z(n3214) );
  XNOR U1308 ( .A(n3848), .B(n3849), .Z(n3834) );
  XNOR U1309 ( .A(n4313), .B(n4314), .Z(n4299) );
  MUX U1310 ( .IN0(n453), .IN1(n4539), .SEL(n4540), .F(n4526) );
  IV U1311 ( .A(n4541), .Z(n453) );
  XOR U1312 ( .A(n4546), .B(n4547), .Z(n4180) );
  XNOR U1313 ( .A(n5154), .B(n5155), .Z(n5141) );
  XNOR U1314 ( .A(n4878), .B(n4879), .Z(n4864) );
  XOR U1315 ( .A(n4753), .B(n4735), .Z(n4739) );
  MUX U1316 ( .IN0(n454), .IN1(n3188), .SEL(n3189), .F(n3059) );
  IV U1317 ( .A(n3190), .Z(n454) );
  MUX U1318 ( .IN0(n455), .IN1(n3917), .SEL(n3281), .F(n3900) );
  IV U1319 ( .A(n3279), .Z(n455) );
  MUX U1320 ( .IN0(n3892), .IN1(n3890), .SEL(n3891), .F(n3192) );
  MUX U1321 ( .IN0(n3263), .IN1(n456), .SEL(n3264), .F(n3225) );
  IV U1322 ( .A(n3265), .Z(n456) );
  MUX U1323 ( .IN0(n4148), .IN1(n457), .SEL(n4149), .F(n4131) );
  IV U1324 ( .A(n4150), .Z(n457) );
  XOR U1325 ( .A(n4535), .B(n4536), .Z(n4159) );
  MUX U1326 ( .IN0(n458), .IN1(n3130), .SEL(n3131), .F(n2994) );
  IV U1327 ( .A(n3132), .Z(n458) );
  MUX U1328 ( .IN0(n459), .IN1(n3105), .SEL(n3106), .F(n2969) );
  IV U1329 ( .A(n3107), .Z(n459) );
  XOR U1330 ( .A(n3881), .B(n3882), .Z(n3898) );
  MUX U1331 ( .IN0(n4343), .IN1(n460), .SEL(n4342), .F(n4333) );
  IV U1332 ( .A(n4341), .Z(n460) );
  XNOR U1333 ( .A(n3178), .B(n3177), .Z(n3160) );
  XOR U1334 ( .A(n3228), .B(n3164), .Z(n3168) );
  MUX U1335 ( .IN0(n461), .IN1(n2961), .SEL(n2962), .F(n2823) );
  IV U1336 ( .A(n2963), .Z(n461) );
  MUX U1337 ( .IN0(n462), .IN1(n2760), .SEL(n2761), .F(n2633) );
  IV U1338 ( .A(n2762), .Z(n462) );
  MUX U1339 ( .IN0(n463), .IN1(n2848), .SEL(n2849), .F(n2719) );
  IV U1340 ( .A(n2850), .Z(n463) );
  MUX U1341 ( .IN0(n464), .IN1(n2658), .SEL(n2659), .F(n2532) );
  IV U1342 ( .A(n2660), .Z(n464) );
  MUX U1343 ( .IN0(n465), .IN1(n2686), .SEL(n2687), .F(n2556) );
  IV U1344 ( .A(n2688), .Z(n465) );
  MUX U1345 ( .IN0(n466), .IN1(n2710), .SEL(n2711), .F(n2580) );
  IV U1346 ( .A(n2712), .Z(n466) );
  MUX U1347 ( .IN0(n467), .IN1(n2572), .SEL(n2573), .F(n2450) );
  IV U1348 ( .A(n2574), .Z(n467) );
  MUX U1349 ( .IN0(n468), .IN1(n2606), .SEL(n2607), .F(n2484) );
  IV U1350 ( .A(n2608), .Z(n468) );
  MUX U1351 ( .IN0(n469), .IN1(n2442), .SEL(n2443), .F(n2321) );
  IV U1352 ( .A(n2444), .Z(n469) );
  MUX U1353 ( .IN0(n470), .IN1(n2803), .SEL(n2804), .F(n2675) );
  IV U1354 ( .A(n2805), .Z(n470) );
  MUX U1355 ( .IN0(n471), .IN1(n2346), .SEL(n2347), .F(n2228) );
  IV U1356 ( .A(n2348), .Z(n471) );
  MUX U1357 ( .IN0(n472), .IN1(n2182), .SEL(n2183), .F(n2073) );
  IV U1358 ( .A(n2184), .Z(n472) );
  MUX U1359 ( .IN0(n473), .IN1(n2219), .SEL(n2220), .F(n2108) );
  IV U1360 ( .A(n2221), .Z(n473) );
  MUX U1361 ( .IN0(n474), .IN1(n2084), .SEL(n2085), .F(n1979) );
  IV U1362 ( .A(n2086), .Z(n474) );
  MUX U1363 ( .IN0(n475), .IN1(n2134), .SEL(n2135), .F(n2029) );
  IV U1364 ( .A(n2136), .Z(n475) );
  MUX U1365 ( .IN0(n476), .IN1(n2270), .SEL(n2271), .F(n2157) );
  IV U1366 ( .A(n2272), .Z(n476) );
  MUX U1367 ( .IN0(n477), .IN1(n1995), .SEL(n1996), .F(n1890) );
  IV U1368 ( .A(n1997), .Z(n477) );
  MUX U1369 ( .IN0(n478), .IN1(n1882), .SEL(n1883), .F(n1782) );
  IV U1370 ( .A(n1884), .Z(n478) );
  MUX U1371 ( .IN0(n479), .IN1(n1907), .SEL(n1908), .F(n1807) );
  IV U1372 ( .A(n1909), .Z(n479) );
  MUX U1373 ( .IN0(n480), .IN1(n1730), .SEL(n1731), .F(n1639) );
  IV U1374 ( .A(n1732), .Z(n480) );
  MUX U1375 ( .IN0(n481), .IN1(n1502), .SEL(n1503), .F(n1418) );
  IV U1376 ( .A(n1504), .Z(n481) );
  MUX U1377 ( .IN0(n482), .IN1(n1494), .SEL(n1495), .F(n1410) );
  IV U1378 ( .A(n1496), .Z(n482) );
  MUX U1379 ( .IN0(n483), .IN1(n1528), .SEL(n1529), .F(n1443) );
  IV U1380 ( .A(n1530), .Z(n483) );
  MUX U1381 ( .IN0(n484), .IN1(n1536), .SEL(n1537), .F(n1451) );
  IV U1382 ( .A(n1538), .Z(n484) );
  MUX U1383 ( .IN0(n485), .IN1(n1222), .SEL(n1223), .F(n1154) );
  IV U1384 ( .A(n1224), .Z(n485) );
  MUX U1385 ( .IN0(n486), .IN1(n1118), .SEL(n1119), .F(n1057) );
  IV U1386 ( .A(n1120), .Z(n486) );
  MUX U1387 ( .IN0(n487), .IN1(n976), .SEL(n977), .F(n917) );
  IV U1388 ( .A(n978), .Z(n487) );
  MUX U1389 ( .IN0(n488), .IN1(n934), .SEL(n935), .F(n888) );
  IV U1390 ( .A(n936), .Z(n488) );
  MUX U1391 ( .IN0(n489), .IN1(n899), .SEL(n900), .F(n855) );
  IV U1392 ( .A(n901), .Z(n489) );
  XNOR U1393 ( .A(n3747), .B(n3746), .Z(n3759) );
  MUX U1394 ( .IN0(n2341), .IN1(n2343), .SEL(n2342), .F(n2223) );
  MUX U1395 ( .IN0(n1617), .IN1(n1619), .SEL(n1618), .F(n1517) );
  MUX U1396 ( .IN0(n1645), .IN1(n1643), .SEL(n1644), .F(n1549) );
  XOR U1397 ( .A(n1470), .B(n1555), .Z(n1471) );
  MUX U1398 ( .IN0(n1525), .IN1(n490), .SEL(n1524), .F(n1437) );
  IV U1399 ( .A(n1523), .Z(n490) );
  MUX U1400 ( .IN0(n926), .IN1(n491), .SEL(n925), .F(n884) );
  IV U1401 ( .A(n924), .Z(n491) );
  XNOR U1402 ( .A(n3087), .B(n2954), .Z(n2958) );
  XOR U1403 ( .A(n3111), .B(n2978), .Z(n2982) );
  XNOR U1404 ( .A(n3145), .B(n3144), .Z(n3127) );
  XNOR U1405 ( .A(n3048), .B(n3047), .Z(n3030) );
  XNOR U1406 ( .A(n2904), .B(n2778), .Z(n2782) );
  XOR U1407 ( .A(n2895), .B(n2769), .Z(n2773) );
  XNOR U1408 ( .A(n2921), .B(n2800), .Z(n2794) );
  XOR U1409 ( .A(n2854), .B(n2728), .Z(n2732) );
  MUX U1410 ( .IN0(n2705), .IN1(n492), .SEL(n2706), .F(n2575) );
  IV U1411 ( .A(n2707), .Z(n492) );
  MUX U1412 ( .IN0(n493), .IN1(n2510), .SEL(n2511), .F(n2389) );
  IV U1413 ( .A(n2512), .Z(n493) );
  XOR U1414 ( .A(n2392), .B(n2284), .Z(n2278) );
  XNOR U1415 ( .A(n2401), .B(n2289), .Z(n2293) );
  XOR U1416 ( .A(n2473), .B(n2355), .Z(n2359) );
  XNOR U1417 ( .A(n2432), .B(n2314), .Z(n2318) );
  NAND U1418 ( .A(n2424), .B(n2543), .Z(n2542) );
  MUX U1419 ( .IN0(n2214), .IN1(n494), .SEL(n2215), .F(n2103) );
  IV U1420 ( .A(n2216), .Z(n494) );
  NAND U1421 ( .A(n1949), .B(n2052), .Z(n2051) );
  XOR U1422 ( .A(n2123), .B(n2021), .Z(n2025) );
  XNOR U1423 ( .A(n1958), .B(n1860), .Z(n1854) );
  XOR U1424 ( .A(n2001), .B(n1899), .Z(n1903) );
  XNOR U1425 ( .A(n1872), .B(n1775), .Z(n1779) );
  XOR U1426 ( .A(n1813), .B(n1722), .Z(n1726) );
  MUX U1427 ( .IN0(n1699), .IN1(n495), .SEL(n1700), .F(n1608) );
  IV U1428 ( .A(n1701), .Z(n495) );
  MUX U1429 ( .IN0(n496), .IN1(n1763), .SEL(n1764), .F(n1669) );
  IV U1430 ( .A(n1765), .Z(n496) );
  XNOR U1431 ( .A(n1333), .B(n1266), .Z(n1270) );
  XOR U1432 ( .A(n1370), .B(n1301), .Z(n1305) );
  XNOR U1433 ( .A(n1379), .B(n1310), .Z(n1314) );
  OR U1434 ( .A(n1280), .B(n1281), .Z(n1218) );
  XNOR U1435 ( .A(n1169), .B(n1110), .Z(n1114) );
  XOR U1436 ( .A(n1160), .B(n1101), .Z(n1105) );
  MUX U1437 ( .IN0(n497), .IN1(n920), .SEL(n921), .F(n876) );
  IV U1438 ( .A(n922), .Z(n497) );
  XNOR U1439 ( .A(n844), .B(n808), .Z(n812) );
  AND U1440 ( .A(n800), .B(n799), .Z(n796) );
  XNOR U1441 ( .A(n3009), .B(n3008), .Z(n2991) );
  XNOR U1442 ( .A(n2809), .B(n2937), .Z(n2810) );
  MUX U1443 ( .IN0(n498), .IN1(n2826), .SEL(n2827), .F(n2697) );
  IV U1444 ( .A(n2828), .Z(n498) );
  XNOR U1445 ( .A(n2742), .B(n2741), .Z(n2724) );
  MUX U1446 ( .IN0(n2682), .IN1(n499), .SEL(n2681), .F(n2550) );
  IV U1447 ( .A(n2680), .Z(n499) );
  XNOR U1448 ( .A(n2369), .B(n2368), .Z(n2351) );
  XNOR U1449 ( .A(n1966), .B(n1965), .Z(n1957) );
  XNOR U1450 ( .A(n2035), .B(n2034), .Z(n2017) );
  XNOR U1451 ( .A(n1736), .B(n1735), .Z(n1718) );
  XNOR U1452 ( .A(n1341), .B(n1340), .Z(n1358) );
  XNOR U1453 ( .A(n1205), .B(n1204), .Z(n1217) );
  XNOR U1454 ( .A(n1245), .B(n1244), .Z(n1227) );
  XNOR U1455 ( .A(n1141), .B(n1140), .Z(n1151) );
  XNOR U1456 ( .A(n1075), .B(n1074), .Z(n1089) );
  XNOR U1457 ( .A(n1019), .B(n1018), .Z(n1028) );
  XNOR U1458 ( .A(n965), .B(n964), .Z(n961) );
  XNOR U1459 ( .A(n774), .B(n773), .Z(n765) );
  MUX U1460 ( .IN0(n2535), .IN1(n500), .SEL(n2536), .F(n2414) );
  IV U1461 ( .A(n2537), .Z(n500) );
  XNOR U1462 ( .A(n2472), .B(n2471), .Z(n2447) );
  XNOR U1463 ( .A(n2233), .B(n2232), .Z(n2208) );
  MUX U1464 ( .IN0(n2188), .IN1(n2302), .SEL(n2190), .F(n2079) );
  XNOR U1465 ( .A(n1912), .B(n1911), .Z(n1887) );
  XNOR U1466 ( .A(n1812), .B(n1811), .Z(n1787) );
  ANDN U1467 ( .A(n1937), .B(n1938), .Z(n1837) );
  NANDN U1468 ( .B(n1569), .A(n1570), .Z(n1486) );
  XNOR U1469 ( .A(n1369), .B(n1368), .Z(n1348) );
  XNOR U1470 ( .A(n1159), .B(n1158), .Z(n1148) );
  XNOR U1471 ( .A(n981), .B(n980), .Z(n973) );
  XNOR U1472 ( .A(n840), .B(n839), .Z(n832) );
  OR U1473 ( .A(n731), .B(n732), .Z(n709) );
  XNOR U1474 ( .A(n2097), .B(n2096), .Z(n2078) );
  XOR U1475 ( .A(n1769), .B(n1766), .Z(n1845) );
  XNOR U1476 ( .A(n1602), .B(n1601), .Z(n1585) );
  XNOR U1477 ( .A(n1507), .B(n1506), .Z(n1490) );
  ANDN U1478 ( .A(n694), .B(n693), .Z(n692) );
  AND U1479 ( .A(n721), .B(n722), .Z(n676) );
  XOR U1480 ( .A(n1261), .B(n1260), .Z(n1327) );
  XNOR U1481 ( .A(n1069), .B(n1068), .Z(n1127) );
  XNOR U1482 ( .A(n911), .B(n910), .Z(n951) );
  XNOR U1483 ( .A(n789), .B(n788), .Z(n824) );
  ANDN U1484 ( .A(n679), .B(n678), .Z(n672) );
  MUX U1485 ( .IN0(\_MxM/Y0[30] ), .IN1(n701), .SEL(n700), .F(n668) );
  XOR U1486 ( .A(n2749), .B(n2752), .Z(n2750) );
  XOR U1487 ( .A(n2378), .B(n2381), .Z(n2379) );
  XOR U1488 ( .A(n2044), .B(n2047), .Z(n2045) );
  XOR U1489 ( .A(n1745), .B(n1749), .Z(n1747) );
  XOR U1490 ( .A(n1475), .B(n1479), .Z(n1477) );
  XOR U1491 ( .A(n1254), .B(n1258), .Z(n1256) );
  XOR U1492 ( .A(n1062), .B(n1066), .Z(n1064) );
  XOR U1493 ( .A(n904), .B(n908), .Z(n906) );
  XOR U1494 ( .A(n782), .B(n786), .Z(n784) );
  MUX U1495 ( .IN0(n501), .IN1(n3749), .SEL(n3750), .F(n3711) );
  IV U1496 ( .A(n3751), .Z(n501) );
  MUX U1497 ( .IN0(n502), .IN1(n3703), .SEL(n3704), .F(n3665) );
  IV U1498 ( .A(n3705), .Z(n502) );
  XOR U1499 ( .A(n4507), .B(n4508), .Z(n4123) );
  MUX U1500 ( .IN0(n503), .IN1(n4101), .SEL(n4102), .F(n4084) );
  IV U1501 ( .A(n4103), .Z(n503) );
  XNOR U1502 ( .A(n4108), .B(n4094), .Z(n4098) );
  MUX U1503 ( .IN0(n504), .IN1(n3597), .SEL(n3598), .F(n3559) );
  IV U1504 ( .A(n3599), .Z(n504) );
  MUX U1505 ( .IN0(n3633), .IN1(n3631), .SEL(n3632), .F(n3593) );
  MUX U1506 ( .IN0(n3652), .IN1(n3654), .SEL(n3653), .F(n3614) );
  MUX U1507 ( .IN0(n3681), .IN1(n505), .SEL(n3682), .F(n3643) );
  IV U1508 ( .A(n3683), .Z(n505) );
  MUX U1509 ( .IN0(n506), .IN1(n4480), .SEL(n4481), .F(n4467) );
  IV U1510 ( .A(n4482), .Z(n506) );
  MUX U1511 ( .IN0(n507), .IN1(n3551), .SEL(n3552), .F(n3513) );
  IV U1512 ( .A(n3553), .Z(n507) );
  MUX U1513 ( .IN0(n508), .IN1(n3564), .SEL(n3565), .F(n3526) );
  IV U1514 ( .A(n3566), .Z(n508) );
  MUX U1515 ( .IN0(n509), .IN1(n3572), .SEL(n3573), .F(n3534) );
  IV U1516 ( .A(n3574), .Z(n509) );
  MUX U1517 ( .IN0(n510), .IN1(n4474), .SEL(n4475), .F(n4461) );
  IV U1518 ( .A(n4476), .Z(n510) );
  XNOR U1519 ( .A(n4057), .B(n4043), .Z(n4047) );
  MUX U1520 ( .IN0(n511), .IN1(n4033), .SEL(n4034), .F(n4016) );
  IV U1521 ( .A(n4035), .Z(n511) );
  MUX U1522 ( .IN0(n4465), .IN1(n512), .SEL(n4056), .F(n4452) );
  IV U1523 ( .A(n4055), .Z(n512) );
  MUX U1524 ( .IN0(n513), .IN1(n3445), .SEL(n3446), .F(n3407) );
  IV U1525 ( .A(n3447), .Z(n513) );
  MUX U1526 ( .IN0(n3481), .IN1(n3479), .SEL(n3480), .F(n3441) );
  MUX U1527 ( .IN0(n514), .IN1(n4036), .SEL(n3547), .F(n4019) );
  IV U1528 ( .A(n3545), .Z(n514) );
  MUX U1529 ( .IN0(n3500), .IN1(n3502), .SEL(n3501), .F(n3462) );
  MUX U1530 ( .IN0(n3529), .IN1(n515), .SEL(n3530), .F(n3491) );
  IV U1531 ( .A(n3531), .Z(n515) );
  MUX U1532 ( .IN0(n516), .IN1(n4428), .SEL(n4429), .F(n4415) );
  IV U1533 ( .A(n4430), .Z(n516) );
  XOR U1534 ( .A(n4835), .B(n4836), .Z(n4845) );
  MUX U1535 ( .IN0(n517), .IN1(n3399), .SEL(n3400), .F(n3361) );
  IV U1536 ( .A(n3401), .Z(n517) );
  MUX U1537 ( .IN0(n518), .IN1(n3412), .SEL(n3413), .F(n3374) );
  IV U1538 ( .A(n3414), .Z(n518) );
  MUX U1539 ( .IN0(n519), .IN1(n3420), .SEL(n3421), .F(n3382) );
  IV U1540 ( .A(n3422), .Z(n519) );
  MUX U1541 ( .IN0(n520), .IN1(n4248), .SEL(n4249), .F(n4227) );
  IV U1542 ( .A(n4250), .Z(n520) );
  XOR U1543 ( .A(n4601), .B(n4602), .Z(n4285) );
  XOR U1544 ( .A(n4969), .B(n4970), .Z(n4850) );
  XOR U1545 ( .A(n4814), .B(n4815), .Z(n4824) );
  MUX U1546 ( .IN0(n521), .IN1(n4818), .SEL(n4819), .F(n4797) );
  IV U1547 ( .A(n4820), .Z(n521) );
  XNOR U1548 ( .A(n3989), .B(n3975), .Z(n3979) );
  MUX U1549 ( .IN0(n522), .IN1(n3965), .SEL(n3966), .F(n3948) );
  IV U1550 ( .A(n3967), .Z(n522) );
  MUX U1551 ( .IN0(n4413), .IN1(n523), .SEL(n3988), .F(n4400) );
  IV U1552 ( .A(n3987), .Z(n523) );
  MUX U1553 ( .IN0(n524), .IN1(n4942), .SEL(n4943), .F(n4929) );
  IV U1554 ( .A(n4944), .Z(n524) );
  MUX U1555 ( .IN0(n525), .IN1(n4409), .SEL(n4410), .F(n4396) );
  IV U1556 ( .A(n4411), .Z(n525) );
  XOR U1557 ( .A(n4581), .B(n4573), .Z(n4224) );
  MUX U1558 ( .IN0(n526), .IN1(n3293), .SEL(n3294), .F(n3255) );
  IV U1559 ( .A(n3295), .Z(n526) );
  MUX U1560 ( .IN0(n3329), .IN1(n3327), .SEL(n3328), .F(n3289) );
  MUX U1561 ( .IN0(n527), .IN1(n3968), .SEL(n3395), .F(n3951) );
  IV U1562 ( .A(n3393), .Z(n527) );
  MUX U1563 ( .IN0(n3348), .IN1(n3350), .SEL(n3349), .F(n3310) );
  MUX U1564 ( .IN0(n3377), .IN1(n528), .SEL(n3378), .F(n3339) );
  IV U1565 ( .A(n3379), .Z(n528) );
  MUX U1566 ( .IN0(n4687), .IN1(n4690), .SEL(n4688), .F(n4671) );
  XOR U1567 ( .A(n4230), .B(n4212), .Z(n4216) );
  MUX U1568 ( .IN0(n529), .IN1(n4556), .SEL(n4557), .F(n4545) );
  IV U1569 ( .A(n4558), .Z(n529) );
  XOR U1570 ( .A(n4364), .B(n4365), .Z(n3936) );
  MUX U1571 ( .IN0(n5059), .IN1(n5062), .SEL(n5060), .F(n5043) );
  XOR U1572 ( .A(n4932), .B(n4924), .Z(n4768) );
  MUX U1573 ( .IN0(n530), .IN1(n4750), .SEL(n4751), .F(n4729) );
  IV U1574 ( .A(n4752), .Z(n530) );
  MUX U1575 ( .IN0(n531), .IN1(n3247), .SEL(n3248), .F(n3209) );
  IV U1576 ( .A(n3249), .Z(n531) );
  XNOR U1577 ( .A(n3938), .B(n3924), .Z(n3928) );
  MUX U1578 ( .IN0(n532), .IN1(n3260), .SEL(n3261), .F(n3222) );
  IV U1579 ( .A(n3262), .Z(n532) );
  MUX U1580 ( .IN0(n533), .IN1(n3268), .SEL(n3269), .F(n3230) );
  IV U1581 ( .A(n3270), .Z(n533) );
  MUX U1582 ( .IN0(n3800), .IN1(n3815), .SEL(n3802), .F(n3775) );
  MUX U1583 ( .IN0(n3843), .IN1(n3846), .SEL(n3844), .F(n3826) );
  MUX U1584 ( .IN0(n534), .IN1(n4164), .SEL(n4165), .F(n4152) );
  IV U1585 ( .A(n4166), .Z(n534) );
  MUX U1586 ( .IN0(n4628), .IN1(n4638), .SEL(n4630), .F(n4616) );
  XOR U1587 ( .A(n4351), .B(n4352), .Z(n3919) );
  MUX U1588 ( .IN0(n535), .IN1(n5170), .SEL(n5171), .F(n5166) );
  IV U1589 ( .A(n5172), .Z(n535) );
  MUX U1590 ( .IN0(n5149), .IN1(n5152), .SEL(n5150), .F(n5133) );
  MUX U1591 ( .IN0(n5000), .IN1(n5010), .SEL(n5002), .F(n4988) );
  XOR U1592 ( .A(n4774), .B(n4756), .Z(n4760) );
  MUX U1593 ( .IN0(n536), .IN1(n3894), .SEL(n3895), .F(n3196) );
  IV U1594 ( .A(n3896), .Z(n536) );
  MUX U1595 ( .IN0(n3783), .IN1(n3793), .SEL(n3785), .F(n3762) );
  XOR U1596 ( .A(n4677), .B(n4678), .Z(n4326) );
  XOR U1597 ( .A(n4548), .B(n4540), .Z(n4161) );
  XOR U1598 ( .A(n5049), .B(n5050), .Z(n4891) );
  XOR U1599 ( .A(n4904), .B(n4905), .Z(n4745) );
  MUX U1600 ( .IN0(n537), .IN1(n4897), .SEL(n4898), .F(n3113) );
  IV U1601 ( .A(n4899), .Z(n537) );
  MUX U1602 ( .IN0(n538), .IN1(n4357), .SEL(n4358), .F(n4341) );
  IV U1603 ( .A(n4359), .Z(n538) );
  XOR U1604 ( .A(n3832), .B(n3833), .Z(n3779) );
  XNOR U1605 ( .A(n3863), .B(n3864), .Z(n3745) );
  XNOR U1606 ( .A(n4306), .B(n4296), .Z(n4300) );
  XOR U1607 ( .A(n4612), .B(n4613), .Z(n4304) );
  XOR U1608 ( .A(n4167), .B(n4145), .Z(n4149) );
  XOR U1609 ( .A(n5164), .B(g_input[3]), .Z(n5165) );
  MUX U1610 ( .IN0(n539), .IN1(n3122), .SEL(n3123), .F(n2986) );
  IV U1611 ( .A(n3124), .Z(n539) );
  MUX U1612 ( .IN0(n540), .IN1(n3089), .SEL(n3090), .F(n2953) );
  IV U1613 ( .A(n3091), .Z(n540) );
  MUX U1614 ( .IN0(n541), .IN1(n3050), .SEL(n3051), .F(n2914) );
  IV U1615 ( .A(n3052), .Z(n541) );
  XOR U1616 ( .A(n5139), .B(n5140), .Z(n5078) );
  XNOR U1617 ( .A(n4871), .B(n4861), .Z(n4865) );
  XOR U1618 ( .A(n4982), .B(n4983), .Z(n4869) );
  XOR U1619 ( .A(n4718), .B(n4719), .Z(n4724) );
  MUX U1620 ( .IN0(n3178), .IN1(n3176), .SEL(n3177), .F(n3046) );
  MUX U1621 ( .IN0(n3167), .IN1(n3169), .SEL(n3168), .F(n3037) );
  MUX U1622 ( .IN0(n542), .IN1(n3900), .SEL(n3243), .F(n3883) );
  IV U1623 ( .A(n3241), .Z(n542) );
  XNOR U1624 ( .A(n3884), .B(n3189), .Z(n3193) );
  MUX U1625 ( .IN0(n3225), .IN1(n543), .SEL(n3226), .F(n3158) );
  IV U1626 ( .A(n3227), .Z(n543) );
  XOR U1627 ( .A(n4520), .B(n4521), .Z(n4140) );
  MUX U1628 ( .IN0(n544), .IN1(n2906), .SEL(n2907), .F(n2777) );
  IV U1629 ( .A(n2908), .Z(n544) );
  MUX U1630 ( .IN0(n545), .IN1(n2897), .SEL(n2898), .F(n2768) );
  IV U1631 ( .A(n2899), .Z(n545) );
  MUX U1632 ( .IN0(n546), .IN1(n3880), .SEL(n3881), .F(n3077) );
  IV U1633 ( .A(n3882), .Z(n546) );
  MUX U1634 ( .IN0(n547), .IN1(n2831), .SEL(n2832), .F(n2702) );
  IV U1635 ( .A(n2833), .Z(n547) );
  MUX U1636 ( .IN0(n548), .IN1(n2865), .SEL(n2866), .F(n2736) );
  IV U1637 ( .A(n2867), .Z(n548) );
  MUX U1638 ( .IN0(n549), .IN1(n2507), .SEL(n2508), .F(n2386) );
  IV U1639 ( .A(n2509), .Z(n549) );
  MUX U1640 ( .IN0(n550), .IN1(n2556), .SEL(n2557), .F(n2434) );
  IV U1641 ( .A(n2558), .Z(n550) );
  MUX U1642 ( .IN0(n551), .IN1(n2589), .SEL(n2590), .F(n2467) );
  IV U1643 ( .A(n2591), .Z(n551) );
  MUX U1644 ( .IN0(n552), .IN1(n2296), .SEL(n2297), .F(n2182) );
  IV U1645 ( .A(n2298), .Z(n552) );
  MUX U1646 ( .IN0(n553), .IN1(n2329), .SEL(n2330), .F(n2211) );
  IV U1647 ( .A(n2331), .Z(n553) );
  MUX U1648 ( .IN0(n554), .IN1(n2363), .SEL(n2364), .F(n2245) );
  IV U1649 ( .A(n2365), .Z(n554) );
  MUX U1650 ( .IN0(n555), .IN1(n2117), .SEL(n2118), .F(n2012) );
  IV U1651 ( .A(n2119), .Z(n555) );
  MUX U1652 ( .IN0(n556), .IN1(n1890), .SEL(n1891), .F(n1790) );
  IV U1653 ( .A(n1892), .Z(n556) );
  MUX U1654 ( .IN0(n557), .IN1(n1924), .SEL(n1925), .F(n1824) );
  IV U1655 ( .A(n1926), .Z(n557) );
  MUX U1656 ( .IN0(n558), .IN1(n1721), .SEL(n1722), .F(n1630) );
  IV U1657 ( .A(n1723), .Z(n558) );
  MUX U1658 ( .IN0(n559), .IN1(n1713), .SEL(n1714), .F(n1622) );
  IV U1659 ( .A(n1715), .Z(n559) );
  MUX U1660 ( .IN0(n560), .IN1(n1680), .SEL(n1681), .F(n1589) );
  IV U1661 ( .A(n1682), .Z(n560) );
  MUX U1662 ( .IN0(n561), .IN1(n1597), .SEL(n1598), .F(n1502) );
  IV U1663 ( .A(n1599), .Z(n561) );
  MUX U1664 ( .IN0(n562), .IN1(n1510), .SEL(n1511), .F(n1426) );
  IV U1665 ( .A(n1512), .Z(n562) );
  MUX U1666 ( .IN0(n563), .IN1(n1545), .SEL(n1546), .F(n1460) );
  IV U1667 ( .A(n1547), .Z(n563) );
  MUX U1668 ( .IN0(n564), .IN1(n1364), .SEL(n1365), .F(n1292) );
  IV U1669 ( .A(n1366), .Z(n564) );
  MUX U1670 ( .IN0(n565), .IN1(n1273), .SEL(n1274), .F(n1207) );
  IV U1671 ( .A(n1275), .Z(n565) );
  MUX U1672 ( .IN0(n566), .IN1(n1092), .SEL(n1093), .F(n1031) );
  IV U1673 ( .A(n1094), .Z(n566) );
  MUX U1674 ( .IN0(n567), .IN1(n943), .SEL(n944), .F(n899) );
  IV U1675 ( .A(n945), .Z(n567) );
  MUX U1676 ( .IN0(n3095), .IN1(n3093), .SEL(n3094), .F(n2957) );
  XOR U1677 ( .A(n5080), .B(n3131), .Z(n3135) );
  XNOR U1678 ( .A(n4133), .B(n4132), .Z(n3771) );
  MUX U1679 ( .IN0(n3009), .IN1(n3007), .SEL(n3008), .F(n2869) );
  MUX U1680 ( .IN0(n2490), .IN1(n2488), .SEL(n2489), .F(n2367) );
  MUX U1681 ( .IN0(n1830), .IN1(n1828), .SEL(n1829), .F(n1734) );
  MUX U1682 ( .IN0(n1780), .IN1(n1778), .SEL(n1779), .F(n1684) );
  MUX U1683 ( .IN0(n1861), .IN1(n568), .SEL(n1860), .F(n1759) );
  IV U1684 ( .A(n1859), .Z(n568) );
  MUX U1685 ( .IN0(n569), .IN1(n873), .SEL(n874), .F(n835) );
  IV U1686 ( .A(n875), .Z(n569) );
  MUX U1687 ( .IN0(n3085), .IN1(n570), .SEL(n3084), .F(n2946) );
  IV U1688 ( .A(n3083), .Z(n570) );
  XNOR U1689 ( .A(n3065), .B(n3064), .Z(n3082) );
  XNOR U1690 ( .A(n3759), .B(n3758), .Z(n3183) );
  XOR U1691 ( .A(n2975), .B(n2840), .Z(n2844) );
  XOR U1692 ( .A(n2792), .B(n2671), .Z(n2672) );
  XOR U1693 ( .A(n2639), .B(n2516), .Z(n2520) );
  XNOR U1694 ( .A(n2648), .B(n2525), .Z(n2529) );
  XOR U1695 ( .A(n2725), .B(n2598), .Z(n2602) );
  XOR U1696 ( .A(n2578), .B(n2459), .Z(n2463) );
  MUX U1697 ( .IN0(n2547), .IN1(n571), .SEL(n2546), .F(n2424) );
  IV U1698 ( .A(n2545), .Z(n571) );
  NAND U1699 ( .A(n2168), .B(n2281), .Z(n2280) );
  XNOR U1700 ( .A(n2286), .B(n2175), .Z(n2179) );
  XOR U1701 ( .A(n2352), .B(n2237), .Z(n2241) );
  XNOR U1702 ( .A(n2193), .B(n2085), .Z(n2089) );
  XOR U1703 ( .A(n2217), .B(n2109), .Z(n2113) );
  MUX U1704 ( .IN0(n2056), .IN1(n572), .SEL(n2055), .F(n1949) );
  IV U1705 ( .A(n2054), .Z(n572) );
  XOR U1706 ( .A(n2018), .B(n1916), .Z(n1920) );
  XOR U1707 ( .A(n1764), .B(n1765), .Z(n1761) );
  XOR U1708 ( .A(n1896), .B(n1799), .Z(n1803) );
  XOR U1709 ( .A(n1611), .B(n1524), .Z(n1518) );
  XOR U1710 ( .A(n1670), .B(n1671), .Z(n1665) );
  XNOR U1711 ( .A(n1492), .B(n1411), .Z(n1415) );
  XOR U1712 ( .A(n1534), .B(n1452), .Z(n1456) );
  XNOR U1713 ( .A(n1263), .B(n1198), .Z(n1204) );
  XNOR U1714 ( .A(n1307), .B(n1240), .Z(n1244) );
  XOR U1715 ( .A(n1298), .B(n1231), .Z(n1235) );
  XOR U1716 ( .A(n1098), .B(n1040), .Z(n1044) );
  XNOR U1717 ( .A(n1107), .B(n1049), .Z(n1053) );
  XOR U1718 ( .A(n923), .B(n884), .Z(n882) );
  XNOR U1719 ( .A(n886), .B(n847), .Z(n851) );
  XNOR U1720 ( .A(n2929), .B(n2928), .Z(n2949) );
  XNOR U1721 ( .A(n3030), .B(n3029), .Z(n3072) );
  XNOR U1722 ( .A(n2821), .B(n2820), .Z(n2836) );
  XNOR U1723 ( .A(n2783), .B(n2782), .Z(n2765) );
  XNOR U1724 ( .A(n2795), .B(n2794), .Z(n2811) );
  XNOR U1725 ( .A(n2656), .B(n2655), .Z(n2638) );
  XNOR U1726 ( .A(n2692), .B(n2691), .Z(n2707) );
  XNOR U1727 ( .A(n2614), .B(n2613), .Z(n2594) );
  XNOR U1728 ( .A(n2562), .B(n2561), .Z(n2577) );
  XNOR U1729 ( .A(n2319), .B(n2318), .Z(n2334) );
  XNOR U1730 ( .A(n2201), .B(n2200), .Z(n2216) );
  XNOR U1731 ( .A(n2253), .B(n2252), .Z(n2233) );
  XNOR U1732 ( .A(n2071), .B(n2070), .Z(n2059) );
  XNOR U1733 ( .A(n1985), .B(n1984), .Z(n2000) );
  XNOR U1734 ( .A(n1855), .B(n1854), .Z(n1848) );
  XNOR U1735 ( .A(n1930), .B(n1929), .Z(n1912) );
  XNOR U1736 ( .A(n1880), .B(n1879), .Z(n1895) );
  XNOR U1737 ( .A(n1645), .B(n1644), .Z(n1627) );
  MUX U1738 ( .IN0(n573), .IN1(n1691), .SEL(n1692), .F(n1600) );
  IV U1739 ( .A(n1693), .Z(n573) );
  XNOR U1740 ( .A(n1466), .B(n1465), .Z(n1448) );
  XNOR U1741 ( .A(n1389), .B(n1388), .Z(n1369) );
  XOR U1742 ( .A(n1280), .B(n1287), .Z(n1349) );
  XNOR U1743 ( .A(n1177), .B(n1176), .Z(n1159) );
  NOR U1744 ( .A(n1027), .B(n1028), .Z(n960) );
  XNOR U1745 ( .A(n1000), .B(n999), .Z(n981) );
  ANDN U1746 ( .A(n965), .B(n964), .Z(n963) );
  MUX U1747 ( .IN0(n765), .IN1(n763), .SEL(n764), .F(n733) );
  MUX U1748 ( .IN0(n574), .IN1(n777), .SEL(n778), .F(n747) );
  IV U1749 ( .A(n779), .Z(n574) );
  XNOR U1750 ( .A(n2894), .B(n2893), .Z(n2936) );
  XNOR U1751 ( .A(n3102), .B(n3101), .Z(n3055) );
  XNOR U1752 ( .A(n2853), .B(n2852), .Z(n2828) );
  XNOR U1753 ( .A(n2724), .B(n2723), .Z(n2699) );
  XNOR U1754 ( .A(n2391), .B(n2390), .Z(n2430) );
  XNOR U1755 ( .A(n2275), .B(n2274), .Z(n2305) );
  XNOR U1756 ( .A(n2351), .B(n2350), .Z(n2326) );
  XNOR U1757 ( .A(n2122), .B(n2121), .Z(n2097) );
  XNOR U1758 ( .A(n2017), .B(n2016), .Z(n1992) );
  ANDN U1759 ( .A(n2147), .B(n2148), .Z(n2042) );
  XNOR U1760 ( .A(n1533), .B(n1532), .Z(n1507) );
  XNOR U1761 ( .A(n1297), .B(n1296), .Z(n1278) );
  XNOR U1762 ( .A(n1097), .B(n1096), .Z(n1087) );
  XNOR U1763 ( .A(n922), .B(n921), .Z(n914) );
  XNOR U1764 ( .A(n803), .B(n802), .Z(n791) );
  XNOR U1765 ( .A(n2966), .B(n2965), .Z(n2919) );
  XNOR U1766 ( .A(n2447), .B(n2446), .Z(n2416) );
  XOR U1767 ( .A(n1974), .B(n1971), .Z(n2049) );
  XNOR U1768 ( .A(n1787), .B(n1786), .Z(n1768) );
  XNOR U1769 ( .A(n1488), .B(n1487), .Z(n1568) );
  MUX U1770 ( .IN0(n715), .IN1(n713), .SEL(n714), .F(n693) );
  XNOR U1771 ( .A(n710), .B(n709), .Z(n708) );
  XOR U1772 ( .A(n1192), .B(n1191), .Z(n1257) );
  XNOR U1773 ( .A(n1015), .B(n1014), .Z(n1065) );
  XNOR U1774 ( .A(n867), .B(n866), .Z(n907) );
  XNOR U1775 ( .A(n759), .B(n758), .Z(n785) );
  XOR U1776 ( .A(n2623), .B(n2626), .Z(n2624) );
  XOR U1777 ( .A(n2262), .B(n2265), .Z(n2263) );
  XOR U1778 ( .A(n1939), .B(n1942), .Z(n1940) );
  XOR U1779 ( .A(n1654), .B(n1658), .Z(n1656) );
  XOR U1780 ( .A(n1398), .B(n1402), .Z(n1400) );
  XOR U1781 ( .A(n1185), .B(n1189), .Z(n1187) );
  XOR U1782 ( .A(n1008), .B(n1012), .Z(n1010) );
  XOR U1783 ( .A(n860), .B(n864), .Z(n862) );
  XOR U1784 ( .A(n752), .B(n756), .Z(n754) );
  MUX U1785 ( .IN0(\_MxM/Y0[31] ), .IN1(n668), .SEL(n669), .F(n665) );
  MUX U1786 ( .IN0(n575), .IN1(n3665), .SEL(n3666), .F(n3627) );
  IV U1787 ( .A(n3667), .Z(n575) );
  MUX U1788 ( .IN0(n576), .IN1(n4093), .SEL(n4094), .F(n4076) );
  IV U1789 ( .A(n4095), .Z(n576) );
  MUX U1790 ( .IN0(n577), .IN1(n3686), .SEL(n3687), .F(n3648) );
  IV U1791 ( .A(n3688), .Z(n577) );
  XNOR U1792 ( .A(n3709), .B(n3708), .Z(n3721) );
  XNOR U1793 ( .A(n4116), .B(n4115), .Z(n3735) );
  MUX U1794 ( .IN0(n578), .IN1(n3640), .SEL(n3641), .F(n3602) );
  IV U1795 ( .A(n3642), .Z(n578) );
  XNOR U1796 ( .A(n3671), .B(n3670), .Z(n3683) );
  XNOR U1797 ( .A(n4099), .B(n4098), .Z(n3697) );
  XNOR U1798 ( .A(n3633), .B(n3632), .Z(n3645) );
  XNOR U1799 ( .A(n4082), .B(n4081), .Z(n3659) );
  XNOR U1800 ( .A(n3595), .B(n3594), .Z(n3607) );
  MUX U1801 ( .IN0(n4478), .IN1(n579), .SEL(n4073), .F(n4465) );
  IV U1802 ( .A(n4072), .Z(n579) );
  MUX U1803 ( .IN0(n580), .IN1(n3513), .SEL(n3514), .F(n3475) );
  IV U1804 ( .A(n3515), .Z(n580) );
  XNOR U1805 ( .A(n4065), .B(n4064), .Z(n3621) );
  XOR U1806 ( .A(n3608), .B(n3573), .Z(n3577) );
  MUX U1807 ( .IN0(n581), .IN1(n4025), .SEL(n4026), .F(n4008) );
  IV U1808 ( .A(n4027), .Z(n581) );
  XNOR U1809 ( .A(n3557), .B(n3556), .Z(n3569) );
  MUX U1810 ( .IN0(n582), .IN1(n4461), .SEL(n4462), .F(n4448) );
  IV U1811 ( .A(n4463), .Z(n582) );
  XNOR U1812 ( .A(n4048), .B(n4047), .Z(n3583) );
  MUX U1813 ( .IN0(n583), .IN1(n3488), .SEL(n3489), .F(n3450) );
  IV U1814 ( .A(n3490), .Z(n583) );
  XNOR U1815 ( .A(n3519), .B(n3518), .Z(n3531) );
  MUX U1816 ( .IN0(n584), .IN1(n4441), .SEL(n4442), .F(n4428) );
  IV U1817 ( .A(n4443), .Z(n584) );
  XNOR U1818 ( .A(n4031), .B(n4030), .Z(n3545) );
  XNOR U1819 ( .A(n3481), .B(n3480), .Z(n3493) );
  XOR U1820 ( .A(n4431), .B(n4423), .Z(n4005) );
  XNOR U1821 ( .A(n4014), .B(n4013), .Z(n3507) );
  XOR U1822 ( .A(n3494), .B(n3459), .Z(n3463) );
  XNOR U1823 ( .A(n3443), .B(n3442), .Z(n3455) );
  MUX U1824 ( .IN0(n585), .IN1(n4594), .SEL(n4595), .F(n4583) );
  IV U1825 ( .A(n4596), .Z(n585) );
  XOR U1826 ( .A(n4403), .B(n4404), .Z(n3987) );
  MUX U1827 ( .IN0(n586), .IN1(n4813), .SEL(n4814), .F(n4792) );
  IV U1828 ( .A(n4815), .Z(n586) );
  MUX U1829 ( .IN0(n587), .IN1(n3361), .SEL(n3362), .F(n3323) );
  IV U1830 ( .A(n3363), .Z(n587) );
  XNOR U1831 ( .A(n3997), .B(n3996), .Z(n3469) );
  MUX U1832 ( .IN0(n588), .IN1(n3957), .SEL(n3958), .F(n3940) );
  IV U1833 ( .A(n3959), .Z(n588) );
  XNOR U1834 ( .A(n3405), .B(n3404), .Z(n3417) );
  MUX U1835 ( .IN0(n589), .IN1(n4227), .SEL(n4228), .F(n4206) );
  IV U1836 ( .A(n4229), .Z(n589) );
  XOR U1837 ( .A(n4272), .B(n4254), .Z(n4258) );
  MUX U1838 ( .IN0(n590), .IN1(n4578), .SEL(n4579), .F(n4567) );
  IV U1839 ( .A(n4580), .Z(n590) );
  XOR U1840 ( .A(n4390), .B(n4391), .Z(n3970) );
  XNOR U1841 ( .A(n3980), .B(n3979), .Z(n3431) );
  MUX U1842 ( .IN0(n591), .IN1(n3336), .SEL(n3337), .F(n3298) );
  IV U1843 ( .A(n3338), .Z(n591) );
  XNOR U1844 ( .A(n3367), .B(n3366), .Z(n3379) );
  MUX U1845 ( .IN0(n4953), .IN1(n592), .SEL(n4810), .F(n4940) );
  IV U1846 ( .A(n4808), .Z(n592) );
  MUX U1847 ( .IN0(n593), .IN1(n4396), .SEL(n4397), .F(n4383) );
  IV U1848 ( .A(n4398), .Z(n593) );
  XNOR U1849 ( .A(n3963), .B(n3962), .Z(n3393) );
  XOR U1850 ( .A(n3380), .B(n3345), .Z(n3349) );
  XNOR U1851 ( .A(n3329), .B(n3328), .Z(n3341) );
  XOR U1852 ( .A(n4570), .B(n4562), .Z(n4203) );
  MUX U1853 ( .IN0(n5121), .IN1(n5137), .SEL(n5123), .F(n5103) );
  XOR U1854 ( .A(n4795), .B(n4777), .Z(n4781) );
  MUX U1855 ( .IN0(n594), .IN1(n4923), .SEL(n4924), .F(n4910) );
  IV U1856 ( .A(n4925), .Z(n594) );
  XNOR U1857 ( .A(n3946), .B(n3945), .Z(n3355) );
  XNOR U1858 ( .A(n3291), .B(n3290), .Z(n3303) );
  XNOR U1859 ( .A(n3283), .B(n3248), .Z(n3252) );
  MUX U1860 ( .IN0(n4308), .IN1(n4311), .SEL(n4309), .F(n4295) );
  MUX U1861 ( .IN0(n4622), .IN1(n4644), .SEL(n4624), .F(n4611) );
  XOR U1862 ( .A(n4209), .B(n4191), .Z(n4195) );
  XOR U1863 ( .A(n4366), .B(n4358), .Z(n3920) );
  MUX U1864 ( .IN0(n4873), .IN1(n4876), .SEL(n4874), .F(n4860) );
  MUX U1865 ( .IN0(n4994), .IN1(n5016), .SEL(n4996), .F(n4981) );
  XOR U1866 ( .A(n4917), .B(n4918), .Z(n4766) );
  MUX U1867 ( .IN0(n595), .IN1(n4729), .SEL(n4730), .F(n4710) );
  IV U1868 ( .A(n4731), .Z(n595) );
  MUX U1869 ( .IN0(n596), .IN1(n3217), .SEL(n3218), .F(n3180) );
  IV U1870 ( .A(n3219), .Z(n596) );
  XNOR U1871 ( .A(n3929), .B(n3928), .Z(n3317) );
  MUX U1872 ( .IN0(n597), .IN1(n3886), .SEL(n3887), .F(n3188) );
  IV U1873 ( .A(n3888), .Z(n597) );
  MUX U1874 ( .IN0(n3775), .IN1(n3799), .SEL(n3777), .F(n3754) );
  MUX U1875 ( .IN0(n598), .IN1(n4152), .SEL(n4153), .F(n4135) );
  IV U1876 ( .A(n4154), .Z(n598) );
  XOR U1877 ( .A(n4685), .B(n4672), .Z(n4327) );
  MUX U1878 ( .IN0(n599), .IN1(n4534), .SEL(n4535), .F(n4519) );
  IV U1879 ( .A(n4536), .Z(n599) );
  MUX U1880 ( .IN0(n600), .IN1(n4350), .SEL(n4351), .F(n4345) );
  IV U1881 ( .A(n4352), .Z(n600) );
  MUX U1882 ( .IN0(g_input[1]), .IN1(n5182), .SEL(g_input[31]), .F(n3835) );
  MUX U1883 ( .IN0(n5084), .IN1(n5094), .SEL(n5086), .F(n3130) );
  XOR U1884 ( .A(n5057), .B(n5044), .Z(n4892) );
  MUX U1885 ( .IN0(n601), .IN1(n4717), .SEL(n4718), .F(n3105) );
  IV U1886 ( .A(n4719), .Z(n601) );
  MUX U1887 ( .IN0(n602), .IN1(n3155), .SEL(n3156), .F(n3025) );
  IV U1888 ( .A(n3157), .Z(n602) );
  MUX U1889 ( .IN0(e_input[1]), .IN1(n603), .SEL(e_input[31]), .F(n4331) );
  IV U1890 ( .A(n4698), .Z(n603) );
  XNOR U1891 ( .A(n3912), .B(n3911), .Z(n3279) );
  XOR U1892 ( .A(n3266), .B(n3231), .Z(n3235) );
  XOR U1893 ( .A(n3841), .B(n3827), .Z(n3780) );
  XOR U1894 ( .A(n4626), .B(n4617), .Z(n4305) );
  MUX U1895 ( .IN0(g_input[2]), .IN1(n5174), .SEL(g_input[31]), .F(n3146) );
  MUX U1896 ( .IN0(n604), .IN1(n3067), .SEL(n3068), .F(n2931) );
  IV U1897 ( .A(n3069), .Z(n604) );
  XOR U1898 ( .A(n5147), .B(n5134), .Z(n5079) );
  XOR U1899 ( .A(n4998), .B(n4989), .Z(n4870) );
  XOR U1900 ( .A(n4732), .B(n4703), .Z(n4707) );
  XNOR U1901 ( .A(n3892), .B(n3891), .Z(n3241) );
  XOR U1902 ( .A(n3781), .B(n3763), .Z(n3767) );
  XNOR U1903 ( .A(n3856), .B(n3742), .Z(n3746) );
  XNOR U1904 ( .A(n4142), .B(n4128), .Z(n4132) );
  XNOR U1905 ( .A(n4301), .B(n4300), .Z(n3876) );
  XOR U1906 ( .A(n4537), .B(n4527), .Z(n4141) );
  MUX U1907 ( .IN0(n605), .IN1(n2953), .SEL(n2954), .F(n2815) );
  IV U1908 ( .A(n2955), .Z(n605) );
  MUX U1909 ( .IN0(n606), .IN1(n2986), .SEL(n2987), .F(n2848) );
  IV U1910 ( .A(n2988), .Z(n606) );
  MUX U1911 ( .IN0(g_input[3]), .IN1(n5165), .SEL(g_input[31]), .F(n607) );
  IV U1912 ( .A(n607), .Z(n3010) );
  MUX U1913 ( .IN0(n608), .IN1(n2785), .SEL(n2786), .F(n2658) );
  IV U1914 ( .A(n2787), .Z(n608) );
  MUX U1915 ( .IN0(e_input[4]), .IN1(n4319), .SEL(e_input[31]), .F(n2798) );
  MUX U1916 ( .IN0(g_input[4]), .IN1(n5131), .SEL(g_input[31]), .F(n609) );
  IV U1917 ( .A(n609), .Z(n2872) );
  MUX U1918 ( .IN0(n610), .IN1(n2633), .SEL(n2634), .F(n2507) );
  IV U1919 ( .A(n2635), .Z(n610) );
  MUX U1920 ( .IN0(g_input[5]), .IN1(n5114), .SEL(g_input[31]), .F(n2743) );
  MUX U1921 ( .IN0(n611), .IN1(n2702), .SEL(n2703), .F(n2572) );
  IV U1922 ( .A(n2704), .Z(n611) );
  MUX U1923 ( .IN0(g_input[6]), .IN1(n5095), .SEL(g_input[31]), .F(n2615) );
  MUX U1924 ( .IN0(n612), .IN1(n2403), .SEL(n2404), .F(n2288) );
  IV U1925 ( .A(n2405), .Z(n612) );
  MUX U1926 ( .IN0(n613), .IN1(n2467), .SEL(n2468), .F(n2346) );
  IV U1927 ( .A(n2469), .Z(n613) );
  MUX U1928 ( .IN0(g_input[7]), .IN1(n5083), .SEL(g_input[31]), .F(n2491) );
  MUX U1929 ( .IN0(n614), .IN1(n2484), .SEL(n2485), .F(n2363) );
  IV U1930 ( .A(n2486), .Z(n614) );
  MUX U1931 ( .IN0(n615), .IN1(n2434), .SEL(n2435), .F(n2313) );
  IV U1932 ( .A(n2436), .Z(n615) );
  MUX U1933 ( .IN0(e_input[8]), .IN1(n3854), .SEL(e_input[31]), .F(n2282) );
  MUX U1934 ( .IN0(n616), .IN1(n2321), .SEL(n2322), .F(n2203) );
  IV U1935 ( .A(n2323), .Z(n616) );
  MUX U1936 ( .IN0(g_input[8]), .IN1(n4986), .SEL(g_input[31]), .F(n2370) );
  MUX U1937 ( .IN0(e_input[9]), .IN1(n3855), .SEL(e_input[31]), .F(n2166) );
  MUX U1938 ( .IN0(g_input[9]), .IN1(n4974), .SEL(g_input[31]), .F(n2254) );
  MUX U1939 ( .IN0(n617), .IN1(n2211), .SEL(n2212), .F(n2100) );
  IV U1940 ( .A(n2213), .Z(n617) );
  MUX U1941 ( .IN0(n618), .IN1(n2073), .SEL(n2074), .F(n1968) );
  IV U1942 ( .A(n2075), .Z(n618) );
  MUX U1943 ( .IN0(g_input[10]), .IN1(n4960), .SEL(g_input[31]), .F(n2141) );
  MUX U1944 ( .IN0(n619), .IN1(n2012), .SEL(n2013), .F(n1907) );
  IV U1945 ( .A(n2014), .Z(n619) );
  MUX U1946 ( .IN0(g_input[11]), .IN1(n4948), .SEL(g_input[31]), .F(n2036) );
  MUX U1947 ( .IN0(n620), .IN1(n2029), .SEL(n2030), .F(n1924) );
  IV U1948 ( .A(n2031), .Z(n620) );
  MUX U1949 ( .IN0(n621), .IN1(n1979), .SEL(n1980), .F(n1874) );
  IV U1950 ( .A(n1981), .Z(n621) );
  MUX U1951 ( .IN0(e_input[12]), .IN1(n3869), .SEL(e_input[31]), .F(n1858) );
  MUX U1952 ( .IN0(g_input[12]), .IN1(n4934), .SEL(g_input[31]), .F(n1931) );
  MUX U1953 ( .IN0(g_input[13]), .IN1(n4922), .SEL(g_input[31]), .F(n1831) );
  MUX U1954 ( .IN0(n622), .IN1(n1790), .SEL(n1791), .F(n1696) );
  IV U1955 ( .A(n1792), .Z(n622) );
  MUX U1956 ( .IN0(g_input[14]), .IN1(n4908), .SEL(g_input[31]), .F(n1737) );
  MUX U1957 ( .IN0(n623), .IN1(n1589), .SEL(n1590), .F(n1494) );
  IV U1958 ( .A(n1591), .Z(n623) );
  MUX U1959 ( .IN0(n624), .IN1(n1622), .SEL(n1623), .F(n1528) );
  IV U1960 ( .A(n1624), .Z(n624) );
  MUX U1961 ( .IN0(n625), .IN1(n1630), .SEL(n1631), .F(n1536) );
  IV U1962 ( .A(n1632), .Z(n625) );
  MUX U1963 ( .IN0(g_input[15]), .IN1(n4896), .SEL(g_input[31]), .F(n1646) );
  MUX U1964 ( .IN0(n626), .IN1(n1639), .SEL(n1640), .F(n1545) );
  IV U1965 ( .A(n1641), .Z(n626) );
  MUX U1966 ( .IN0(e_input[16]), .IN1(n5070), .SEL(e_input[31]), .F(n1522) );
  MUX U1967 ( .IN0(g_input[16]), .IN1(n4524), .SEL(g_input[31]), .F(n1554) );
  MUX U1968 ( .IN0(e_input[17]), .IN1(n5071), .SEL(e_input[31]), .F(n1435) );
  MUX U1969 ( .IN0(g_input[17]), .IN1(n4512), .SEL(g_input[31]), .F(n1467) );
  MUX U1970 ( .IN0(g_input[18]), .IN1(n4498), .SEL(g_input[31]), .F(n1390) );
  MUX U1971 ( .IN0(n627), .IN1(n1426), .SEL(n1427), .F(n1353) );
  IV U1972 ( .A(n1428), .Z(n627) );
  MUX U1973 ( .IN0(g_input[19]), .IN1(n4486), .SEL(g_input[31]), .F(n1316) );
  MUX U1974 ( .IN0(n628), .IN1(n1292), .SEL(n1293), .F(n1222) );
  IV U1975 ( .A(n1294), .Z(n628) );
  MUX U1976 ( .IN0(g_input[20]), .IN1(n4472), .SEL(g_input[31]), .F(n1246) );
  MUX U1977 ( .IN0(e_input[20]), .IN1(n4884), .SEL(e_input[31]), .F(n1196) );
  MUX U1978 ( .IN0(e_input[21]), .IN1(n4885), .SEL(e_input[31]), .F(n1138) );
  MUX U1979 ( .IN0(g_input[21]), .IN1(n4460), .SEL(g_input[31]), .F(n1178) );
  MUX U1980 ( .IN0(g_input[22]), .IN1(n4446), .SEL(g_input[31]), .F(n1116) );
  MUX U1981 ( .IN0(g_input[23]), .IN1(n4434), .SEL(g_input[31]), .F(n1055) );
  MUX U1982 ( .IN0(n629), .IN1(n1031), .SEL(n1032), .F(n976) );
  IV U1983 ( .A(n1033), .Z(n629) );
  MUX U1984 ( .IN0(n630), .IN1(n1207), .SEL(n1208), .F(n1143) );
  IV U1985 ( .A(n1209), .Z(n630) );
  MUX U1986 ( .IN0(e_input[24]), .IN1(n5160), .SEL(e_input[31]), .F(n984) );
  MUX U1987 ( .IN0(g_input[24]), .IN1(n4420), .SEL(g_input[31]), .F(n1001) );
  MUX U1988 ( .IN0(g_input[25]), .IN1(n4408), .SEL(g_input[31]), .F(n941) );
  MUX U1989 ( .IN0(e_input[25]), .IN1(n5161), .SEL(e_input[31]), .F(n928) );
  MUX U1990 ( .IN0(g_input[26]), .IN1(n4394), .SEL(g_input[31]), .F(n897) );
  MUX U1991 ( .IN0(e_input[27]), .IN1(n5145), .SEL(e_input[31]), .F(n631) );
  IV U1992 ( .A(n631), .Z(n834) );
  MUX U1993 ( .IN0(e_input[26]), .IN1(n5146), .SEL(e_input[31]), .F(n872) );
  MUX U1994 ( .IN0(g_input[27]), .IN1(n4382), .SEL(g_input[31]), .F(n853) );
  MUX U1995 ( .IN0(e_input[2]), .IN1(n4683), .SEL(e_input[31]), .F(n3076) );
  XNOR U1996 ( .A(n5162), .B(n3140), .Z(n3144) );
  XNOR U1997 ( .A(n4866), .B(n4865), .Z(n4713) );
  XOR U1998 ( .A(n4893), .B(n3114), .Z(n3118) );
  XNOR U1999 ( .A(n3170), .B(n3043), .Z(n3047) );
  MUX U2000 ( .IN0(n3158), .IN1(n632), .SEL(n3159), .F(n3028) );
  IV U2001 ( .A(n3160), .Z(n632) );
  XNOR U2002 ( .A(n3083), .B(n4328), .Z(n3084) );
  XNOR U2003 ( .A(n3194), .B(n3193), .Z(n3204) );
  MUX U2004 ( .IN0(e_input[3]), .IN1(n4684), .SEL(e_input[31]), .F(n2944) );
  MUX U2005 ( .IN0(e_input[5]), .IN1(n4320), .SEL(e_input[31]), .F(n2668) );
  MUX U2006 ( .IN0(n2742), .IN1(n2740), .SEL(n2741), .F(n2610) );
  MUX U2007 ( .IN0(n2692), .IN1(n2690), .SEL(n2691), .F(n2560) );
  MUX U2008 ( .IN0(e_input[6]), .IN1(n4324), .SEL(e_input[31]), .F(n2544) );
  XOR U2009 ( .A(n2257), .B(n2371), .Z(n2258) );
  MUX U2010 ( .IN0(e_input[10]), .IN1(n3839), .SEL(e_input[31]), .F(n2053) );
  MUX U2011 ( .IN0(n633), .IN1(n2157), .SEL(n2158), .F(n2054) );
  IV U2012 ( .A(n2159), .Z(n633) );
  MUX U2013 ( .IN0(e_input[11]), .IN1(n3840), .SEL(e_input[31]), .F(n1952) );
  MUX U2014 ( .IN0(n2035), .IN1(n2033), .SEL(n2034), .F(n1928) );
  MUX U2015 ( .IN0(n1985), .IN1(n1983), .SEL(n1984), .F(n1878) );
  MUX U2016 ( .IN0(e_input[13]), .IN1(n3870), .SEL(e_input[31]), .F(n1757) );
  MUX U2017 ( .IN0(e_input[18]), .IN1(n5055), .SEL(e_input[31]), .F(n1352) );
  MUX U2018 ( .IN0(e_input[19]), .IN1(n5056), .SEL(e_input[31]), .F(n1284) );
  MUX U2019 ( .IN0(e_input[22]), .IN1(n4890), .SEL(e_input[31]), .F(n1079) );
  MUX U2020 ( .IN0(e_input[23]), .IN1(n4889), .SEL(e_input[31]), .F(n634) );
  IV U2021 ( .A(n634), .Z(n1020) );
  MUX U2022 ( .IN0(e_input[28]), .IN1(n5179), .SEL(e_input[31]), .F(n806) );
  MUX U2023 ( .IN0(e_input[29]), .IN1(n5180), .SEL(e_input[31]), .F(n771) );
  MUX U2024 ( .IN0(n635), .IN1(n855), .SEL(n856), .F(n816) );
  IV U2025 ( .A(n857), .Z(n635) );
  MUX U2026 ( .IN0(g_input[28]), .IN1(n4368), .SEL(g_input[31]), .F(n814) );
  XOR U2027 ( .A(n3031), .B(n2898), .Z(n2902) );
  XNOR U2028 ( .A(n3057), .B(n2924), .Z(n2928) );
  NAND U2029 ( .A(n2941), .B(n3075), .Z(n3074) );
  XNOR U2030 ( .A(n3095), .B(n3094), .Z(n3110) );
  XOR U2031 ( .A(n2992), .B(n2857), .Z(n2861) );
  XOR U2032 ( .A(n2676), .B(n2677), .Z(n2673) );
  XOR U2033 ( .A(n2837), .B(n2711), .Z(n2715) );
  XOR U2034 ( .A(n2546), .B(n2547), .Z(n2541) );
  XOR U2035 ( .A(n2513), .B(n2395), .Z(n2399) );
  XOR U2036 ( .A(n2595), .B(n2476), .Z(n2480) );
  MUX U2037 ( .IN0(e_input[7]), .IN1(n4325), .SEL(e_input[31]), .F(n2421) );
  XOR U2038 ( .A(n2456), .B(n2338), .Z(n2342) );
  XNOR U2039 ( .A(n2060), .B(n2163), .Z(n2061) );
  XNOR U2040 ( .A(n2172), .B(n2066), .Z(n2070) );
  XOR U2041 ( .A(n2234), .B(n2126), .Z(n2130) );
  XOR U2042 ( .A(n2106), .B(n2004), .Z(n2008) );
  XOR U2043 ( .A(n1913), .B(n1816), .Z(n1820) );
  XOR U2044 ( .A(n1796), .B(n1705), .Z(n1709) );
  MUX U2045 ( .IN0(n1761), .IN1(n1850), .SEL(n1760), .F(n1663) );
  MUX U2046 ( .IN0(e_input[14]), .IN1(n3874), .SEL(e_input[31]), .F(n1668) );
  NAND U2047 ( .A(n1437), .B(n1521), .Z(n1520) );
  XNOR U2048 ( .A(n1408), .B(n1336), .Z(n1340) );
  XNOR U2049 ( .A(n1458), .B(n1384), .Z(n1388) );
  XOR U2050 ( .A(n1449), .B(n1373), .Z(n1377) );
  XOR U2051 ( .A(n1228), .B(n1163), .Z(n1167) );
  XNOR U2052 ( .A(n1237), .B(n1172), .Z(n1176) );
  XNOR U2053 ( .A(n1194), .B(n1135), .Z(n1140) );
  XNOR U2054 ( .A(n1046), .B(n995), .Z(n999) );
  XOR U2055 ( .A(n1037), .B(n986), .Z(n990) );
  OR U2056 ( .A(n884), .B(n885), .Z(n879) );
  MUX U2057 ( .IN0(n636), .IN1(n835), .SEL(n836), .F(n799) );
  IV U2058 ( .A(n837), .Z(n636) );
  MUX U2059 ( .IN0(n637), .IN1(n807), .SEL(n808), .F(n767) );
  IV U2060 ( .A(n809), .Z(n637) );
  MUX U2061 ( .IN0(g_input[29]), .IN1(n4356), .SEL(g_input[31]), .F(n775) );
  XNOR U2062 ( .A(n2959), .B(n2958), .Z(n2974) );
  XNOR U2063 ( .A(n2912), .B(n2911), .Z(n2894) );
  MUX U2064 ( .IN0(n2811), .IN1(n2809), .SEL(n2810), .F(n638) );
  IV U2065 ( .A(n638), .Z(n2679) );
  XNOR U2066 ( .A(n2530), .B(n2529), .Z(n2512) );
  XNOR U2067 ( .A(n2409), .B(n2408), .Z(n2391) );
  XNOR U2068 ( .A(n2440), .B(n2439), .Z(n2455) );
  XNOR U2069 ( .A(n2490), .B(n2489), .Z(n2472) );
  XNOR U2070 ( .A(n2294), .B(n2293), .Z(n2275) );
  XNOR U2071 ( .A(n2180), .B(n2179), .Z(n2162) );
  XNOR U2072 ( .A(n2140), .B(n2139), .Z(n2122) );
  XNOR U2073 ( .A(n2090), .B(n2089), .Z(n2105) );
  MUX U2074 ( .IN0(n1846), .IN1(n639), .SEL(n1847), .F(n1753) );
  IV U2075 ( .A(n1848), .Z(n639) );
  XNOR U2076 ( .A(n1780), .B(n1779), .Z(n1795) );
  XNOR U2077 ( .A(n1830), .B(n1829), .Z(n1812) );
  XNOR U2078 ( .A(n1686), .B(n1685), .Z(n1701) );
  XNOR U2079 ( .A(n1595), .B(n1594), .Z(n1610) );
  XNOR U2080 ( .A(n1500), .B(n1499), .Z(n1515) );
  XNOR U2081 ( .A(n1553), .B(n1552), .Z(n1533) );
  MUX U2082 ( .IN0(e_input[15]), .IN1(n3875), .SEL(e_input[31]), .F(n1574) );
  MUX U2083 ( .IN0(n640), .IN1(n1669), .SEL(n1670), .F(n1582) );
  IV U2084 ( .A(n1671), .Z(n640) );
  XNOR U2085 ( .A(n1416), .B(n1415), .Z(n1431) );
  XNOR U2086 ( .A(n1315), .B(n1314), .Z(n1297) );
  XNOR U2087 ( .A(n1215), .B(n1219), .Z(n1279) );
  XNOR U2088 ( .A(n1115), .B(n1114), .Z(n1097) );
  XNOR U2089 ( .A(n1054), .B(n1053), .Z(n1036) );
  AND U2090 ( .A(n966), .B(n967), .Z(n962) );
  XNOR U2091 ( .A(n940), .B(n939), .Z(n922) );
  XNOR U2092 ( .A(n896), .B(n895), .Z(n878) );
  MUX U2093 ( .IN0(g_input[30]), .IN1(n4338), .SEL(g_input[31]), .F(n744) );
  MUX U2094 ( .IN0(e_input[30]), .IN1(n5185), .SEL(e_input[31]), .F(n746) );
  XNOR U2095 ( .A(n2991), .B(n2990), .Z(n2966) );
  MUX U2096 ( .IN0(n3053), .IN1(n641), .SEL(n3054), .F(n2917) );
  IV U2097 ( .A(n3055), .Z(n641) );
  XNOR U2098 ( .A(n2765), .B(n2764), .Z(n2808) );
  XNOR U2099 ( .A(n2638), .B(n2637), .Z(n2682) );
  XNOR U2100 ( .A(n2303), .B(n2417), .Z(n2304) );
  NANDN U2101 ( .B(n1974), .A(n1975), .Z(n1869) );
  XNOR U2102 ( .A(n1718), .B(n1717), .Z(n1693) );
  XNOR U2103 ( .A(n1627), .B(n1626), .Z(n1602) );
  ANDN U2104 ( .A(n1743), .B(n1744), .Z(n1652) );
  XNOR U2105 ( .A(n1448), .B(n1447), .Z(n1423) );
  XNOR U2106 ( .A(n1227), .B(n1226), .Z(n1212) );
  XOR U2107 ( .A(n1027), .B(n1024), .Z(n1070) );
  OR U2108 ( .A(n790), .B(n791), .Z(n760) );
  MUX U2109 ( .IN0(n741), .IN1(n739), .SEL(n740), .F(n713) );
  OR U2110 ( .A(n711), .B(n712), .Z(n689) );
  XNOR U2111 ( .A(n2828), .B(n2827), .Z(n2790) );
  XNOR U2112 ( .A(n2699), .B(n2698), .Z(n2663) );
  XNOR U2113 ( .A(n2569), .B(n2568), .Z(n2537) );
  XNOR U2114 ( .A(n2326), .B(n2325), .Z(n2301) );
  XNOR U2115 ( .A(n2208), .B(n2207), .Z(n2187) );
  XNOR U2116 ( .A(n1992), .B(n1991), .Z(n1973) );
  XNOR U2117 ( .A(n1887), .B(n1886), .Z(n1868) );
  XOR U2118 ( .A(n1569), .B(n1583), .Z(n1660) );
  MUX U2119 ( .IN0(n642), .IN1(n718), .SEL(n719), .F(n695) );
  IV U2120 ( .A(n720), .Z(n642) );
  MUX U2121 ( .IN0(n3016), .IN1(n643), .SEL(n3017), .F(n2878) );
  IV U2122 ( .A(\_MxM/Y0[1] ), .Z(n643) );
  XOR U2123 ( .A(n1331), .B(n1330), .Z(n1401) );
  XNOR U2124 ( .A(n1131), .B(n1130), .Z(n1188) );
  XNOR U2125 ( .A(n955), .B(n954), .Z(n1011) );
  XNOR U2126 ( .A(n828), .B(n827), .Z(n863) );
  XNOR U2127 ( .A(n730), .B(n729), .Z(n755) );
  XNOR U2128 ( .A(n679), .B(n678), .Z(n704) );
  XOR U2129 ( .A(n2499), .B(n2502), .Z(n2500) );
  XOR U2130 ( .A(n2149), .B(n2152), .Z(n2150) );
  XOR U2131 ( .A(n1839), .B(n1843), .Z(n1841) );
  XOR U2132 ( .A(n1562), .B(n1566), .Z(n1564) );
  XOR U2133 ( .A(n1324), .B(n1328), .Z(n1326) );
  XOR U2134 ( .A(n1123), .B(n1128), .Z(n1126) );
  XOR U2135 ( .A(n948), .B(n952), .Z(n950) );
  XOR U2136 ( .A(n821), .B(n825), .Z(n823) );
  XOR U2137 ( .A(n723), .B(n727), .Z(n725) );
  MUX U2138 ( .IN0(n665), .IN1(\_MxM/Y1[30] ), .SEL(n666), .F(\_MxM/Y1[31] )
         );
  MUX U2139 ( .IN0(\_MxM/Y1[29] ), .IN1(o[29]), .SEL(n644), .F(\_MxM/n97 ) );
  MUX U2140 ( .IN0(\_MxM/Y1[30] ), .IN1(o[30]), .SEL(n644), .F(\_MxM/n94 ) );
  MUX U2141 ( .IN0(\_MxM/Y1[31] ), .IN1(o[31]), .SEL(n644), .F(\_MxM/n91 ) );
  MUX U2142 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n644), .F(\_MxM/n184 ) );
  MUX U2143 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n644), .F(\_MxM/n181 ) );
  MUX U2144 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n644), .F(\_MxM/n178 ) );
  MUX U2145 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n644), .F(\_MxM/n175 ) );
  MUX U2146 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n644), .F(\_MxM/n172 ) );
  MUX U2147 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n644), .F(\_MxM/n169 ) );
  MUX U2148 ( .IN0(\_MxM/Y1[6] ), .IN1(o[6]), .SEL(n644), .F(\_MxM/n166 ) );
  MUX U2149 ( .IN0(\_MxM/Y1[7] ), .IN1(o[7]), .SEL(n644), .F(\_MxM/n163 ) );
  MUX U2150 ( .IN0(\_MxM/Y1[8] ), .IN1(o[8]), .SEL(n644), .F(\_MxM/n160 ) );
  MUX U2151 ( .IN0(\_MxM/Y1[9] ), .IN1(o[9]), .SEL(n644), .F(\_MxM/n157 ) );
  MUX U2152 ( .IN0(\_MxM/Y1[10] ), .IN1(o[10]), .SEL(n644), .F(\_MxM/n154 ) );
  MUX U2153 ( .IN0(\_MxM/Y1[11] ), .IN1(o[11]), .SEL(n644), .F(\_MxM/n151 ) );
  MUX U2154 ( .IN0(\_MxM/Y1[12] ), .IN1(o[12]), .SEL(n644), .F(\_MxM/n148 ) );
  MUX U2155 ( .IN0(\_MxM/Y1[13] ), .IN1(o[13]), .SEL(n644), .F(\_MxM/n145 ) );
  MUX U2156 ( .IN0(\_MxM/Y1[14] ), .IN1(o[14]), .SEL(n644), .F(\_MxM/n142 ) );
  MUX U2157 ( .IN0(\_MxM/Y1[15] ), .IN1(o[15]), .SEL(n644), .F(\_MxM/n139 ) );
  MUX U2158 ( .IN0(\_MxM/Y1[16] ), .IN1(o[16]), .SEL(n644), .F(\_MxM/n136 ) );
  MUX U2159 ( .IN0(\_MxM/Y1[17] ), .IN1(o[17]), .SEL(n644), .F(\_MxM/n133 ) );
  MUX U2160 ( .IN0(\_MxM/Y1[18] ), .IN1(o[18]), .SEL(n644), .F(\_MxM/n130 ) );
  MUX U2161 ( .IN0(\_MxM/Y1[19] ), .IN1(o[19]), .SEL(n644), .F(\_MxM/n127 ) );
  MUX U2162 ( .IN0(\_MxM/Y1[20] ), .IN1(o[20]), .SEL(n644), .F(\_MxM/n124 ) );
  MUX U2163 ( .IN0(\_MxM/Y1[21] ), .IN1(o[21]), .SEL(n644), .F(\_MxM/n121 ) );
  MUX U2164 ( .IN0(\_MxM/Y1[22] ), .IN1(o[22]), .SEL(n644), .F(\_MxM/n118 ) );
  MUX U2165 ( .IN0(\_MxM/Y1[23] ), .IN1(o[23]), .SEL(n644), .F(\_MxM/n115 ) );
  MUX U2166 ( .IN0(\_MxM/Y1[24] ), .IN1(o[24]), .SEL(n644), .F(\_MxM/n112 ) );
  MUX U2167 ( .IN0(\_MxM/Y1[25] ), .IN1(o[25]), .SEL(n644), .F(\_MxM/n109 ) );
  MUX U2168 ( .IN0(\_MxM/Y1[26] ), .IN1(o[26]), .SEL(n644), .F(\_MxM/n106 ) );
  IV U2169 ( .A(n645), .Z(n644) );
  MUX U2170 ( .IN0(o[27]), .IN1(\_MxM/Y1[27] ), .SEL(n645), .F(\_MxM/n103 ) );
  MUX U2171 ( .IN0(o[28]), .IN1(\_MxM/Y1[28] ), .SEL(n645), .F(\_MxM/n100 ) );
  AND U2172 ( .A(n646), .B(n647), .Z(n645) );
  AND U2173 ( .A(n648), .B(n649), .Z(n647) );
  ANDN U2174 ( .A(n650), .B(\_MxM/n[3] ), .Z(n649) );
  NOR U2175 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n650) );
  ANDN U2176 ( .A(n651), .B(\_MxM/n[13] ), .Z(n648) );
  NOR U2177 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n651) );
  AND U2178 ( .A(n652), .B(n653), .Z(n646) );
  ANDN U2179 ( .A(n654), .B(\_MxM/n[10] ), .Z(n653) );
  ANDN U2180 ( .A(n655), .B(n656), .Z(n652) );
  NOR U2181 ( .A(\_MxM/n[0] ), .B(n657), .Z(n655) );
  XOR U2182 ( .A(n658), .B(\_MxM/Y0[10] ), .Z(\_MxM/Y1[9] ) );
  XOR U2183 ( .A(n659), .B(\_MxM/Y0[9] ), .Z(\_MxM/Y1[8] ) );
  XOR U2184 ( .A(n660), .B(\_MxM/Y0[8] ), .Z(\_MxM/Y1[7] ) );
  XOR U2185 ( .A(n661), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XOR U2186 ( .A(n662), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XOR U2187 ( .A(n663), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U2188 ( .A(n664), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U2189 ( .A(\_MxM/Y0[31] ), .B(n667), .Z(n666) );
  XNOR U2190 ( .A(n669), .B(\_MxM/Y0[31] ), .Z(\_MxM/Y1[30] ) );
  XOR U2191 ( .A(n668), .B(n667), .Z(n669) );
  XOR U2192 ( .A(n670), .B(n671), .Z(n667) );
  XOR U2193 ( .A(n672), .B(n673), .Z(n671) );
  AND U2194 ( .A(n674), .B(n675), .Z(n673) );
  XNOR U2195 ( .A(n680), .B(n678), .Z(n670) );
  XOR U2196 ( .A(n681), .B(n682), .Z(n680) );
  XOR U2197 ( .A(n683), .B(n684), .Z(n682) );
  XOR U2198 ( .A(n685), .B(n686), .Z(n684) );
  XOR U2199 ( .A(n691), .B(n692), .Z(n683) );
  XOR U2200 ( .A(n697), .B(n698), .Z(n681) );
  XNOR U2201 ( .A(n687), .B(n699), .Z(n698) );
  XOR U2202 ( .A(n695), .B(n693), .Z(n697) );
  XNOR U2203 ( .A(n702), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U2204 ( .A(n700), .B(\_MxM/Y0[30] ), .Z(\_MxM/Y1[29] ) );
  XNOR U2205 ( .A(n703), .B(n704), .Z(n700) );
  XNOR U2206 ( .A(n701), .B(n705), .Z(n703) );
  AND U2207 ( .A(n674), .B(n706), .Z(n705) );
  XOR U2208 ( .A(n677), .B(n704), .Z(n706) );
  XNOR U2209 ( .A(n676), .B(n704), .Z(n677) );
  XOR U2210 ( .A(n690), .B(n699), .Z(n688) );
  IV U2211 ( .A(n689), .Z(n699) );
  XOR U2212 ( .A(n695), .B(n696), .Z(n694) );
  OR U2213 ( .A(n716), .B(n717), .Z(n696) );
  XNOR U2214 ( .A(n724), .B(\_MxM/Y0[29] ), .Z(\_MxM/Y1[28] ) );
  XNOR U2215 ( .A(n725), .B(n726), .Z(n724) );
  AND U2216 ( .A(n674), .B(n728), .Z(n727) );
  XOR U2217 ( .A(n722), .B(n726), .Z(n728) );
  XNOR U2218 ( .A(n721), .B(n726), .Z(n722) );
  XOR U2219 ( .A(n733), .B(n734), .Z(n711) );
  ANDN U2220 ( .A(n735), .B(n733), .Z(n734) );
  XOR U2221 ( .A(n733), .B(n736), .Z(n735) );
  XOR U2222 ( .A(n737), .B(n738), .Z(n714) );
  IV U2223 ( .A(n713), .Z(n738) );
  XNOR U2224 ( .A(n719), .B(n720), .Z(n715) );
  NANDN U2225 ( .B(n716), .A(n744), .Z(n720) );
  XNOR U2226 ( .A(n718), .B(n745), .Z(n719) );
  ANDN U2227 ( .A(n746), .B(n717), .Z(n745) );
  XNOR U2228 ( .A(n753), .B(\_MxM/Y0[28] ), .Z(\_MxM/Y1[27] ) );
  XNOR U2229 ( .A(n754), .B(n755), .Z(n753) );
  AND U2230 ( .A(n674), .B(n757), .Z(n756) );
  XOR U2231 ( .A(n751), .B(n755), .Z(n757) );
  XNOR U2232 ( .A(n750), .B(n755), .Z(n751) );
  XOR U2233 ( .A(n736), .B(n762), .Z(n732) );
  IV U2234 ( .A(n733), .Z(n762) );
  XOR U2235 ( .A(n770), .B(n743), .Z(n766) );
  NANDN U2236 ( .B(n717), .A(n771), .Z(n743) );
  IV U2237 ( .A(n739), .Z(n770) );
  XNOR U2238 ( .A(n748), .B(n749), .Z(n741) );
  NANDN U2239 ( .B(n716), .A(n775), .Z(n749) );
  XNOR U2240 ( .A(n747), .B(n776), .Z(n748) );
  AND U2241 ( .A(n744), .B(n746), .Z(n776) );
  XNOR U2242 ( .A(n783), .B(\_MxM/Y0[27] ), .Z(\_MxM/Y1[26] ) );
  XNOR U2243 ( .A(n784), .B(n785), .Z(n783) );
  AND U2244 ( .A(n674), .B(n787), .Z(n786) );
  XOR U2245 ( .A(n781), .B(n785), .Z(n787) );
  XNOR U2246 ( .A(n780), .B(n785), .Z(n781) );
  XNOR U2247 ( .A(n765), .B(n764), .Z(n761) );
  XOR U2248 ( .A(n792), .B(n793), .Z(n764) );
  XOR U2249 ( .A(n794), .B(n795), .Z(n793) );
  XOR U2250 ( .A(n796), .B(n797), .Z(n795) );
  XNOR U2251 ( .A(n767), .B(n805), .Z(n768) );
  ANDN U2252 ( .A(n806), .B(n717), .Z(n805) );
  XOR U2253 ( .A(n810), .B(n769), .Z(n804) );
  NAND U2254 ( .A(n771), .B(n744), .Z(n769) );
  IV U2255 ( .A(n772), .Z(n810) );
  XNOR U2256 ( .A(n778), .B(n779), .Z(n774) );
  NANDN U2257 ( .B(n716), .A(n814), .Z(n779) );
  XNOR U2258 ( .A(n777), .B(n815), .Z(n778) );
  AND U2259 ( .A(n775), .B(n746), .Z(n815) );
  XNOR U2260 ( .A(n822), .B(\_MxM/Y0[26] ), .Z(\_MxM/Y1[25] ) );
  XNOR U2261 ( .A(n823), .B(n824), .Z(n822) );
  AND U2262 ( .A(n674), .B(n826), .Z(n825) );
  XOR U2263 ( .A(n820), .B(n824), .Z(n826) );
  XNOR U2264 ( .A(n819), .B(n824), .Z(n820) );
  XOR U2265 ( .A(n829), .B(n830), .Z(n790) );
  ANDN U2266 ( .A(n831), .B(n829), .Z(n830) );
  XOR U2267 ( .A(n829), .B(n832), .Z(n831) );
  XNOR U2268 ( .A(n833), .B(n798), .Z(n802) );
  XOR U2269 ( .A(n799), .B(n800), .Z(n798) );
  OR U2270 ( .A(n717), .B(n834), .Z(n800) );
  XNOR U2271 ( .A(n794), .B(n801), .Z(n833) );
  XNOR U2272 ( .A(n807), .B(n845), .Z(n808) );
  AND U2273 ( .A(n744), .B(n806), .Z(n845) );
  XOR U2274 ( .A(n849), .B(n809), .Z(n844) );
  NAND U2275 ( .A(n771), .B(n775), .Z(n809) );
  IV U2276 ( .A(n811), .Z(n849) );
  XNOR U2277 ( .A(n817), .B(n818), .Z(n813) );
  NANDN U2278 ( .B(n716), .A(n853), .Z(n818) );
  XNOR U2279 ( .A(n816), .B(n854), .Z(n817) );
  AND U2280 ( .A(n814), .B(n746), .Z(n854) );
  XNOR U2281 ( .A(n861), .B(\_MxM/Y0[25] ), .Z(\_MxM/Y1[24] ) );
  XNOR U2282 ( .A(n862), .B(n863), .Z(n861) );
  AND U2283 ( .A(n674), .B(n865), .Z(n864) );
  XOR U2284 ( .A(n859), .B(n863), .Z(n865) );
  XNOR U2285 ( .A(n858), .B(n863), .Z(n859) );
  XNOR U2286 ( .A(n870), .B(n843), .Z(n839) );
  XNOR U2287 ( .A(n836), .B(n837), .Z(n843) );
  NANDN U2288 ( .B(n834), .A(n744), .Z(n837) );
  XNOR U2289 ( .A(n835), .B(n871), .Z(n836) );
  ANDN U2290 ( .A(n872), .B(n717), .Z(n871) );
  XNOR U2291 ( .A(n842), .B(n838), .Z(n870) );
  XNOR U2292 ( .A(n879), .B(n880), .Z(n842) );
  IV U2293 ( .A(n841), .Z(n880) );
  XNOR U2294 ( .A(n846), .B(n887), .Z(n847) );
  AND U2295 ( .A(n775), .B(n806), .Z(n887) );
  XOR U2296 ( .A(n891), .B(n848), .Z(n886) );
  NAND U2297 ( .A(n771), .B(n814), .Z(n848) );
  IV U2298 ( .A(n850), .Z(n891) );
  XOR U2299 ( .A(n892), .B(n893), .Z(n850) );
  ANDN U2300 ( .A(n894), .B(n895), .Z(n893) );
  XOR U2301 ( .A(n892), .B(n896), .Z(n894) );
  XNOR U2302 ( .A(n856), .B(n857), .Z(n852) );
  NANDN U2303 ( .B(n716), .A(n897), .Z(n857) );
  XNOR U2304 ( .A(n855), .B(n898), .Z(n856) );
  AND U2305 ( .A(n853), .B(n746), .Z(n898) );
  XNOR U2306 ( .A(n905), .B(\_MxM/Y0[24] ), .Z(\_MxM/Y1[23] ) );
  XNOR U2307 ( .A(n906), .B(n907), .Z(n905) );
  AND U2308 ( .A(n674), .B(n909), .Z(n908) );
  XOR U2309 ( .A(n903), .B(n907), .Z(n909) );
  XNOR U2310 ( .A(n902), .B(n907), .Z(n903) );
  XNOR U2311 ( .A(n915), .B(n883), .Z(n877) );
  XNOR U2312 ( .A(n874), .B(n875), .Z(n883) );
  NANDN U2313 ( .B(n834), .A(n775), .Z(n875) );
  XNOR U2314 ( .A(n873), .B(n916), .Z(n874) );
  AND U2315 ( .A(n744), .B(n872), .Z(n916) );
  XNOR U2316 ( .A(n882), .B(n876), .Z(n915) );
  XOR U2317 ( .A(n927), .B(n885), .Z(n923) );
  NANDN U2318 ( .B(n717), .A(n928), .Z(n885) );
  IV U2319 ( .A(n881), .Z(n927) );
  XNOR U2320 ( .A(n888), .B(n933), .Z(n889) );
  AND U2321 ( .A(n814), .B(n806), .Z(n933) );
  XOR U2322 ( .A(n937), .B(n890), .Z(n932) );
  NAND U2323 ( .A(n771), .B(n853), .Z(n890) );
  IV U2324 ( .A(n892), .Z(n937) );
  XNOR U2325 ( .A(n900), .B(n901), .Z(n896) );
  NANDN U2326 ( .B(n716), .A(n941), .Z(n901) );
  XNOR U2327 ( .A(n899), .B(n942), .Z(n900) );
  AND U2328 ( .A(n897), .B(n746), .Z(n942) );
  XNOR U2329 ( .A(n949), .B(\_MxM/Y0[23] ), .Z(\_MxM/Y1[22] ) );
  XNOR U2330 ( .A(n950), .B(n951), .Z(n949) );
  AND U2331 ( .A(n674), .B(n953), .Z(n952) );
  XOR U2332 ( .A(n947), .B(n951), .Z(n953) );
  XNOR U2333 ( .A(n946), .B(n951), .Z(n947) );
  XNOR U2334 ( .A(n914), .B(n913), .Z(n911) );
  XOR U2335 ( .A(n956), .B(n957), .Z(n913) );
  XOR U2336 ( .A(n958), .B(n959), .Z(n957) );
  XOR U2337 ( .A(n962), .B(n963), .Z(n958) );
  XOR U2338 ( .A(n968), .B(n912), .Z(n956) );
  XOR U2339 ( .A(n969), .B(n970), .Z(n912) );
  ANDN U2340 ( .A(n971), .B(n972), .Z(n970) );
  XNOR U2341 ( .A(n969), .B(n973), .Z(n971) );
  XOR U2342 ( .A(n966), .B(n964), .Z(n968) );
  XNOR U2343 ( .A(n974), .B(n931), .Z(n921) );
  XNOR U2344 ( .A(n918), .B(n919), .Z(n931) );
  NANDN U2345 ( .B(n834), .A(n814), .Z(n919) );
  XNOR U2346 ( .A(n917), .B(n975), .Z(n918) );
  AND U2347 ( .A(n775), .B(n872), .Z(n975) );
  XNOR U2348 ( .A(n930), .B(n920), .Z(n974) );
  XNOR U2349 ( .A(n924), .B(n983), .Z(n925) );
  ANDN U2350 ( .A(n984), .B(n717), .Z(n983) );
  XOR U2351 ( .A(n988), .B(n926), .Z(n982) );
  NAND U2352 ( .A(n928), .B(n744), .Z(n926) );
  IV U2353 ( .A(n929), .Z(n988) );
  XNOR U2354 ( .A(n934), .B(n993), .Z(n935) );
  AND U2355 ( .A(n853), .B(n806), .Z(n993) );
  XOR U2356 ( .A(n997), .B(n936), .Z(n992) );
  NAND U2357 ( .A(n771), .B(n897), .Z(n936) );
  IV U2358 ( .A(n938), .Z(n997) );
  XNOR U2359 ( .A(n944), .B(n945), .Z(n940) );
  NANDN U2360 ( .B(n716), .A(n1001), .Z(n945) );
  XNOR U2361 ( .A(n943), .B(n1002), .Z(n944) );
  AND U2362 ( .A(n941), .B(n746), .Z(n1002) );
  XNOR U2363 ( .A(n1009), .B(\_MxM/Y0[22] ), .Z(\_MxM/Y1[21] ) );
  XNOR U2364 ( .A(n1010), .B(n1011), .Z(n1009) );
  AND U2365 ( .A(n674), .B(n1013), .Z(n1012) );
  XOR U2366 ( .A(n1007), .B(n1011), .Z(n1013) );
  XNOR U2367 ( .A(n1006), .B(n1011), .Z(n1007) );
  XNOR U2368 ( .A(n1016), .B(n961), .Z(n972) );
  XOR U2369 ( .A(n966), .B(n967), .Z(n965) );
  OR U2370 ( .A(n717), .B(n1020), .Z(n967) );
  XNOR U2371 ( .A(n960), .B(n969), .Z(n1016) );
  XNOR U2372 ( .A(n1029), .B(n991), .Z(n980) );
  XNOR U2373 ( .A(n977), .B(n978), .Z(n991) );
  NANDN U2374 ( .B(n834), .A(n853), .Z(n978) );
  XNOR U2375 ( .A(n976), .B(n1030), .Z(n977) );
  AND U2376 ( .A(n814), .B(n872), .Z(n1030) );
  XNOR U2377 ( .A(n990), .B(n979), .Z(n1029) );
  XNOR U2378 ( .A(n985), .B(n1038), .Z(n986) );
  AND U2379 ( .A(n744), .B(n984), .Z(n1038) );
  XOR U2380 ( .A(n1042), .B(n987), .Z(n1037) );
  NAND U2381 ( .A(n928), .B(n775), .Z(n987) );
  IV U2382 ( .A(n989), .Z(n1042) );
  XNOR U2383 ( .A(n994), .B(n1047), .Z(n995) );
  AND U2384 ( .A(n897), .B(n806), .Z(n1047) );
  XOR U2385 ( .A(n1051), .B(n996), .Z(n1046) );
  NAND U2386 ( .A(n771), .B(n941), .Z(n996) );
  IV U2387 ( .A(n998), .Z(n1051) );
  XNOR U2388 ( .A(n1004), .B(n1005), .Z(n1000) );
  NANDN U2389 ( .B(n716), .A(n1055), .Z(n1005) );
  XNOR U2390 ( .A(n1003), .B(n1056), .Z(n1004) );
  AND U2391 ( .A(n1001), .B(n746), .Z(n1056) );
  XNOR U2392 ( .A(n1063), .B(\_MxM/Y0[21] ), .Z(\_MxM/Y1[20] ) );
  XNOR U2393 ( .A(n1064), .B(n1065), .Z(n1063) );
  AND U2394 ( .A(n674), .B(n1067), .Z(n1066) );
  XOR U2395 ( .A(n1061), .B(n1065), .Z(n1067) );
  XNOR U2396 ( .A(n1060), .B(n1065), .Z(n1061) );
  XNOR U2397 ( .A(n1070), .B(n1028), .Z(n1025) );
  XOR U2398 ( .A(n1071), .B(n1072), .Z(n1018) );
  IV U2399 ( .A(n1017), .Z(n1072) );
  XNOR U2400 ( .A(n1022), .B(n1023), .Z(n1019) );
  NANDN U2401 ( .B(n1020), .A(n744), .Z(n1023) );
  XNOR U2402 ( .A(n1021), .B(n1078), .Z(n1022) );
  ANDN U2403 ( .A(n1079), .B(n717), .Z(n1078) );
  XOR U2404 ( .A(n1083), .B(n1084), .Z(n1024) );
  ANDN U2405 ( .A(n1085), .B(n1086), .Z(n1084) );
  XNOR U2406 ( .A(n1083), .B(n1087), .Z(n1085) );
  XNOR U2407 ( .A(n1090), .B(n1045), .Z(n1035) );
  XNOR U2408 ( .A(n1032), .B(n1033), .Z(n1045) );
  NANDN U2409 ( .B(n834), .A(n897), .Z(n1033) );
  XNOR U2410 ( .A(n1031), .B(n1091), .Z(n1032) );
  AND U2411 ( .A(n853), .B(n872), .Z(n1091) );
  XNOR U2412 ( .A(n1044), .B(n1034), .Z(n1090) );
  XNOR U2413 ( .A(n1039), .B(n1099), .Z(n1040) );
  AND U2414 ( .A(n775), .B(n984), .Z(n1099) );
  XOR U2415 ( .A(n1103), .B(n1041), .Z(n1098) );
  NAND U2416 ( .A(n928), .B(n814), .Z(n1041) );
  IV U2417 ( .A(n1043), .Z(n1103) );
  XNOR U2418 ( .A(n1048), .B(n1108), .Z(n1049) );
  AND U2419 ( .A(n941), .B(n806), .Z(n1108) );
  XOR U2420 ( .A(n1112), .B(n1050), .Z(n1107) );
  NAND U2421 ( .A(n771), .B(n1001), .Z(n1050) );
  IV U2422 ( .A(n1052), .Z(n1112) );
  XNOR U2423 ( .A(n1058), .B(n1059), .Z(n1054) );
  NANDN U2424 ( .B(n716), .A(n1116), .Z(n1059) );
  XNOR U2425 ( .A(n1057), .B(n1117), .Z(n1058) );
  AND U2426 ( .A(n1055), .B(n746), .Z(n1117) );
  XNOR U2427 ( .A(n1125), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U2428 ( .A(n1124), .B(\_MxM/Y0[20] ), .Z(\_MxM/Y1[19] ) );
  XNOR U2429 ( .A(n1126), .B(n1127), .Z(n1124) );
  AND U2430 ( .A(n674), .B(n1129), .Z(n1128) );
  XOR U2431 ( .A(n1122), .B(n1127), .Z(n1129) );
  XNOR U2432 ( .A(n1121), .B(n1127), .Z(n1122) );
  XNOR U2433 ( .A(n1132), .B(n1089), .Z(n1086) );
  XOR U2434 ( .A(n1137), .B(n1077), .Z(n1133) );
  NANDN U2435 ( .B(n717), .A(n1138), .Z(n1077) );
  IV U2436 ( .A(n1073), .Z(n1137) );
  XNOR U2437 ( .A(n1081), .B(n1082), .Z(n1075) );
  NANDN U2438 ( .B(n1020), .A(n775), .Z(n1082) );
  XNOR U2439 ( .A(n1080), .B(n1142), .Z(n1081) );
  AND U2440 ( .A(n744), .B(n1079), .Z(n1142) );
  XNOR U2441 ( .A(n1152), .B(n1106), .Z(n1096) );
  XNOR U2442 ( .A(n1093), .B(n1094), .Z(n1106) );
  NANDN U2443 ( .B(n834), .A(n941), .Z(n1094) );
  XNOR U2444 ( .A(n1092), .B(n1153), .Z(n1093) );
  AND U2445 ( .A(n897), .B(n872), .Z(n1153) );
  XNOR U2446 ( .A(n1105), .B(n1095), .Z(n1152) );
  XNOR U2447 ( .A(n1100), .B(n1161), .Z(n1101) );
  AND U2448 ( .A(n814), .B(n984), .Z(n1161) );
  XOR U2449 ( .A(n1165), .B(n1102), .Z(n1160) );
  NAND U2450 ( .A(n928), .B(n853), .Z(n1102) );
  IV U2451 ( .A(n1104), .Z(n1165) );
  XNOR U2452 ( .A(n1109), .B(n1170), .Z(n1110) );
  AND U2453 ( .A(n1001), .B(n806), .Z(n1170) );
  XOR U2454 ( .A(n1174), .B(n1111), .Z(n1169) );
  NAND U2455 ( .A(n771), .B(n1055), .Z(n1111) );
  IV U2456 ( .A(n1113), .Z(n1174) );
  XNOR U2457 ( .A(n1119), .B(n1120), .Z(n1115) );
  NANDN U2458 ( .B(n716), .A(n1178), .Z(n1120) );
  XNOR U2459 ( .A(n1118), .B(n1179), .Z(n1119) );
  AND U2460 ( .A(n1116), .B(n746), .Z(n1179) );
  XNOR U2461 ( .A(n1186), .B(\_MxM/Y0[19] ), .Z(\_MxM/Y1[18] ) );
  XNOR U2462 ( .A(n1187), .B(n1188), .Z(n1186) );
  AND U2463 ( .A(n674), .B(n1190), .Z(n1189) );
  XOR U2464 ( .A(n1184), .B(n1188), .Z(n1190) );
  XNOR U2465 ( .A(n1183), .B(n1188), .Z(n1184) );
  XNOR U2466 ( .A(n1193), .B(n1151), .Z(n1147) );
  XNOR U2467 ( .A(n1134), .B(n1195), .Z(n1135) );
  ANDN U2468 ( .A(n1196), .B(n717), .Z(n1195) );
  XOR U2469 ( .A(n1200), .B(n1136), .Z(n1194) );
  NAND U2470 ( .A(n1138), .B(n744), .Z(n1136) );
  IV U2471 ( .A(n1139), .Z(n1200) );
  XOR U2472 ( .A(n1201), .B(n1202), .Z(n1139) );
  ANDN U2473 ( .A(n1203), .B(n1204), .Z(n1202) );
  XOR U2474 ( .A(n1201), .B(n1205), .Z(n1203) );
  XNOR U2475 ( .A(n1144), .B(n1145), .Z(n1141) );
  NANDN U2476 ( .B(n1020), .A(n814), .Z(n1145) );
  XNOR U2477 ( .A(n1143), .B(n1206), .Z(n1144) );
  AND U2478 ( .A(n775), .B(n1079), .Z(n1206) );
  XNOR U2479 ( .A(n1150), .B(n1146), .Z(n1193) );
  XNOR U2480 ( .A(n1213), .B(n1214), .Z(n1150) );
  IV U2481 ( .A(n1149), .Z(n1214) );
  XNOR U2482 ( .A(n1220), .B(n1168), .Z(n1158) );
  XNOR U2483 ( .A(n1155), .B(n1156), .Z(n1168) );
  NANDN U2484 ( .B(n834), .A(n1001), .Z(n1156) );
  XNOR U2485 ( .A(n1154), .B(n1221), .Z(n1155) );
  AND U2486 ( .A(n941), .B(n872), .Z(n1221) );
  XNOR U2487 ( .A(n1167), .B(n1157), .Z(n1220) );
  XNOR U2488 ( .A(n1162), .B(n1229), .Z(n1163) );
  AND U2489 ( .A(n853), .B(n984), .Z(n1229) );
  XOR U2490 ( .A(n1233), .B(n1164), .Z(n1228) );
  NAND U2491 ( .A(n928), .B(n897), .Z(n1164) );
  IV U2492 ( .A(n1166), .Z(n1233) );
  XNOR U2493 ( .A(n1171), .B(n1238), .Z(n1172) );
  AND U2494 ( .A(n1055), .B(n806), .Z(n1238) );
  XOR U2495 ( .A(n1242), .B(n1173), .Z(n1237) );
  NAND U2496 ( .A(n771), .B(n1116), .Z(n1173) );
  IV U2497 ( .A(n1175), .Z(n1242) );
  XNOR U2498 ( .A(n1181), .B(n1182), .Z(n1177) );
  NANDN U2499 ( .B(n716), .A(n1246), .Z(n1182) );
  XNOR U2500 ( .A(n1180), .B(n1247), .Z(n1181) );
  AND U2501 ( .A(n1178), .B(n746), .Z(n1247) );
  ANDN U2502 ( .A(n1248), .B(n1249), .Z(n1180) );
  NANDN U2503 ( .B(n1250), .A(n1251), .Z(n1248) );
  XOR U2504 ( .A(n1255), .B(\_MxM/Y0[18] ), .Z(\_MxM/Y1[17] ) );
  XNOR U2505 ( .A(n1256), .B(n1257), .Z(n1255) );
  AND U2506 ( .A(n674), .B(n1259), .Z(n1258) );
  XOR U2507 ( .A(n1253), .B(n1257), .Z(n1259) );
  XNOR U2508 ( .A(n1252), .B(n1257), .Z(n1253) );
  XNOR U2509 ( .A(n1212), .B(n1211), .Z(n1192) );
  XOR U2510 ( .A(n1262), .B(n1217), .Z(n1211) );
  XNOR U2511 ( .A(n1197), .B(n1264), .Z(n1198) );
  AND U2512 ( .A(n744), .B(n1196), .Z(n1264) );
  XOR U2513 ( .A(n1268), .B(n1199), .Z(n1263) );
  NAND U2514 ( .A(n1138), .B(n775), .Z(n1199) );
  IV U2515 ( .A(n1201), .Z(n1268) );
  XNOR U2516 ( .A(n1208), .B(n1209), .Z(n1205) );
  NANDN U2517 ( .B(n1020), .A(n853), .Z(n1209) );
  XNOR U2518 ( .A(n1207), .B(n1272), .Z(n1208) );
  AND U2519 ( .A(n814), .B(n1079), .Z(n1272) );
  XNOR U2520 ( .A(n1216), .B(n1210), .Z(n1262) );
  XOR U2521 ( .A(n1279), .B(n1218), .Z(n1216) );
  NAND U2522 ( .A(n1282), .B(n1283), .Z(n1219) );
  NANDN U2523 ( .B(n717), .A(n1284), .Z(n1283) );
  OR U2524 ( .A(n1285), .B(n1286), .Z(n1282) );
  XNOR U2525 ( .A(n1290), .B(n1236), .Z(n1226) );
  XNOR U2526 ( .A(n1223), .B(n1224), .Z(n1236) );
  NANDN U2527 ( .B(n834), .A(n1055), .Z(n1224) );
  XNOR U2528 ( .A(n1222), .B(n1291), .Z(n1223) );
  AND U2529 ( .A(n1001), .B(n872), .Z(n1291) );
  XNOR U2530 ( .A(n1235), .B(n1225), .Z(n1290) );
  XNOR U2531 ( .A(n1230), .B(n1299), .Z(n1231) );
  AND U2532 ( .A(n897), .B(n984), .Z(n1299) );
  XOR U2533 ( .A(n1303), .B(n1232), .Z(n1298) );
  NAND U2534 ( .A(n928), .B(n941), .Z(n1232) );
  IV U2535 ( .A(n1234), .Z(n1303) );
  XNOR U2536 ( .A(n1239), .B(n1308), .Z(n1240) );
  AND U2537 ( .A(n1116), .B(n806), .Z(n1308) );
  XOR U2538 ( .A(n1312), .B(n1241), .Z(n1307) );
  NAND U2539 ( .A(n771), .B(n1178), .Z(n1241) );
  IV U2540 ( .A(n1243), .Z(n1312) );
  XNOR U2541 ( .A(n1250), .B(n1251), .Z(n1245) );
  NANDN U2542 ( .B(n716), .A(n1316), .Z(n1251) );
  XOR U2543 ( .A(n1249), .B(n1317), .Z(n1250) );
  AND U2544 ( .A(n1246), .B(n746), .Z(n1317) );
  NAND U2545 ( .A(n1318), .B(n1319), .Z(n1249) );
  NANDN U2546 ( .B(n1320), .A(n1321), .Z(n1318) );
  XOR U2547 ( .A(n1325), .B(\_MxM/Y0[17] ), .Z(\_MxM/Y1[16] ) );
  XNOR U2548 ( .A(n1326), .B(n1327), .Z(n1325) );
  AND U2549 ( .A(n674), .B(n1329), .Z(n1328) );
  XOR U2550 ( .A(n1323), .B(n1327), .Z(n1329) );
  XNOR U2551 ( .A(n1322), .B(n1327), .Z(n1323) );
  XNOR U2552 ( .A(n1278), .B(n1277), .Z(n1261) );
  XOR U2553 ( .A(n1332), .B(n1289), .Z(n1277) );
  XNOR U2554 ( .A(n1265), .B(n1334), .Z(n1266) );
  AND U2555 ( .A(n775), .B(n1196), .Z(n1334) );
  XOR U2556 ( .A(n1338), .B(n1267), .Z(n1333) );
  NAND U2557 ( .A(n1138), .B(n814), .Z(n1267) );
  IV U2558 ( .A(n1269), .Z(n1338) );
  XNOR U2559 ( .A(n1274), .B(n1275), .Z(n1271) );
  NANDN U2560 ( .B(n1020), .A(n897), .Z(n1275) );
  XNOR U2561 ( .A(n1273), .B(n1342), .Z(n1274) );
  AND U2562 ( .A(n853), .B(n1079), .Z(n1342) );
  XNOR U2563 ( .A(n1288), .B(n1276), .Z(n1332) );
  XNOR U2564 ( .A(n1349), .B(n1281), .Z(n1288) );
  XOR U2565 ( .A(n1350), .B(n1285), .Z(n1281) );
  NAND U2566 ( .A(n1284), .B(n744), .Z(n1285) );
  NANDN U2567 ( .B(n717), .A(n1352), .Z(n1351) );
  XNOR U2568 ( .A(n1362), .B(n1306), .Z(n1296) );
  XNOR U2569 ( .A(n1293), .B(n1294), .Z(n1306) );
  NANDN U2570 ( .B(n834), .A(n1116), .Z(n1294) );
  XNOR U2571 ( .A(n1292), .B(n1363), .Z(n1293) );
  AND U2572 ( .A(n1055), .B(n872), .Z(n1363) );
  XNOR U2573 ( .A(n1305), .B(n1295), .Z(n1362) );
  XNOR U2574 ( .A(n1300), .B(n1371), .Z(n1301) );
  AND U2575 ( .A(n941), .B(n984), .Z(n1371) );
  XOR U2576 ( .A(n1375), .B(n1302), .Z(n1370) );
  NAND U2577 ( .A(n928), .B(n1001), .Z(n1302) );
  IV U2578 ( .A(n1304), .Z(n1375) );
  XNOR U2579 ( .A(n1309), .B(n1380), .Z(n1310) );
  AND U2580 ( .A(n1178), .B(n806), .Z(n1380) );
  XOR U2581 ( .A(n1381), .B(n1382), .Z(n1309) );
  ANDN U2582 ( .A(n1383), .B(n1384), .Z(n1382) );
  XNOR U2583 ( .A(n1385), .B(n1381), .Z(n1383) );
  XOR U2584 ( .A(n1386), .B(n1311), .Z(n1379) );
  NAND U2585 ( .A(n771), .B(n1246), .Z(n1311) );
  IV U2586 ( .A(n1313), .Z(n1386) );
  XNOR U2587 ( .A(n1320), .B(n1321), .Z(n1315) );
  NANDN U2588 ( .B(n716), .A(n1390), .Z(n1321) );
  XNOR U2589 ( .A(n1319), .B(n1391), .Z(n1320) );
  AND U2590 ( .A(n1316), .B(n746), .Z(n1391) );
  AND U2591 ( .A(n1392), .B(n1393), .Z(n1319) );
  NANDN U2592 ( .B(n1394), .A(n1395), .Z(n1392) );
  XOR U2593 ( .A(n1399), .B(\_MxM/Y0[16] ), .Z(\_MxM/Y1[15] ) );
  XNOR U2594 ( .A(n1400), .B(n1401), .Z(n1399) );
  AND U2595 ( .A(n674), .B(n1403), .Z(n1402) );
  XOR U2596 ( .A(n1397), .B(n1401), .Z(n1403) );
  XNOR U2597 ( .A(n1396), .B(n1401), .Z(n1397) );
  XNOR U2598 ( .A(n1348), .B(n1347), .Z(n1331) );
  XOR U2599 ( .A(n1407), .B(n1358), .Z(n1347) );
  XNOR U2600 ( .A(n1335), .B(n1409), .Z(n1336) );
  AND U2601 ( .A(n814), .B(n1196), .Z(n1409) );
  XOR U2602 ( .A(n1413), .B(n1337), .Z(n1408) );
  NAND U2603 ( .A(n1138), .B(n853), .Z(n1337) );
  IV U2604 ( .A(n1339), .Z(n1413) );
  XNOR U2605 ( .A(n1344), .B(n1345), .Z(n1341) );
  NANDN U2606 ( .B(n1020), .A(n941), .Z(n1345) );
  XNOR U2607 ( .A(n1343), .B(n1417), .Z(n1344) );
  AND U2608 ( .A(n897), .B(n1079), .Z(n1417) );
  XNOR U2609 ( .A(n1357), .B(n1346), .Z(n1407) );
  XNOR U2610 ( .A(n1424), .B(n1361), .Z(n1357) );
  NAND U2611 ( .A(n1284), .B(n775), .Z(n1355) );
  XNOR U2612 ( .A(n1353), .B(n1425), .Z(n1354) );
  AND U2613 ( .A(n744), .B(n1352), .Z(n1425) );
  XNOR U2614 ( .A(n1360), .B(n1356), .Z(n1424) );
  AND U2615 ( .A(n1433), .B(n1434), .Z(n1432) );
  NANDN U2616 ( .B(n717), .A(n1435), .Z(n1434) );
  OR U2617 ( .A(n1436), .B(n1437), .Z(n1433) );
  XNOR U2618 ( .A(n1441), .B(n1378), .Z(n1368) );
  XNOR U2619 ( .A(n1365), .B(n1366), .Z(n1378) );
  NANDN U2620 ( .B(n834), .A(n1178), .Z(n1366) );
  XNOR U2621 ( .A(n1364), .B(n1442), .Z(n1365) );
  AND U2622 ( .A(n1116), .B(n872), .Z(n1442) );
  XNOR U2623 ( .A(n1377), .B(n1367), .Z(n1441) );
  XNOR U2624 ( .A(n1372), .B(n1450), .Z(n1373) );
  AND U2625 ( .A(n1001), .B(n984), .Z(n1450) );
  XOR U2626 ( .A(n1454), .B(n1374), .Z(n1449) );
  NAND U2627 ( .A(n928), .B(n1055), .Z(n1374) );
  IV U2628 ( .A(n1376), .Z(n1454) );
  XNOR U2629 ( .A(n1381), .B(n1459), .Z(n1384) );
  AND U2630 ( .A(n1246), .B(n806), .Z(n1459) );
  XOR U2631 ( .A(n1463), .B(n1385), .Z(n1458) );
  NAND U2632 ( .A(n771), .B(n1316), .Z(n1385) );
  IV U2633 ( .A(n1387), .Z(n1463) );
  XNOR U2634 ( .A(n1394), .B(n1395), .Z(n1389) );
  NANDN U2635 ( .B(n716), .A(n1467), .Z(n1395) );
  XNOR U2636 ( .A(n1393), .B(n1468), .Z(n1394) );
  AND U2637 ( .A(n1390), .B(n746), .Z(n1468) );
  ANDN U2638 ( .A(n1469), .B(n1470), .Z(n1393) );
  NANDN U2639 ( .B(n1471), .A(n1472), .Z(n1469) );
  XOR U2640 ( .A(n1476), .B(\_MxM/Y0[15] ), .Z(\_MxM/Y1[14] ) );
  XNOR U2641 ( .A(n1477), .B(n1478), .Z(n1476) );
  AND U2642 ( .A(n674), .B(n1480), .Z(n1479) );
  XOR U2643 ( .A(n1474), .B(n1478), .Z(n1480) );
  XNOR U2644 ( .A(n1473), .B(n1478), .Z(n1474) );
  XOR U2645 ( .A(n1406), .B(n1405), .Z(n1478) );
  XOR U2646 ( .A(n1481), .B(n1482), .Z(n1405) );
  XOR U2647 ( .A(n1483), .B(n1484), .Z(n1482) );
  XOR U2648 ( .A(n1485), .B(n1483), .Z(n1484) );
  XNOR U2649 ( .A(n1423), .B(n1422), .Z(n1406) );
  XOR U2650 ( .A(n1491), .B(n1431), .Z(n1422) );
  XNOR U2651 ( .A(n1410), .B(n1493), .Z(n1411) );
  AND U2652 ( .A(n853), .B(n1196), .Z(n1493) );
  XOR U2653 ( .A(n1497), .B(n1412), .Z(n1492) );
  NAND U2654 ( .A(n1138), .B(n897), .Z(n1412) );
  IV U2655 ( .A(n1414), .Z(n1497) );
  XNOR U2656 ( .A(n1419), .B(n1420), .Z(n1416) );
  NANDN U2657 ( .B(n1020), .A(n1001), .Z(n1420) );
  XNOR U2658 ( .A(n1418), .B(n1501), .Z(n1419) );
  AND U2659 ( .A(n941), .B(n1079), .Z(n1501) );
  XNOR U2660 ( .A(n1430), .B(n1421), .Z(n1491) );
  XNOR U2661 ( .A(n1508), .B(n1440), .Z(n1430) );
  NAND U2662 ( .A(n1284), .B(n814), .Z(n1428) );
  XNOR U2663 ( .A(n1426), .B(n1509), .Z(n1427) );
  AND U2664 ( .A(n775), .B(n1352), .Z(n1509) );
  XNOR U2665 ( .A(n1439), .B(n1429), .Z(n1508) );
  XNOR U2666 ( .A(n1516), .B(n1438), .Z(n1439) );
  XNOR U2667 ( .A(n1520), .B(n1436), .Z(n1516) );
  NAND U2668 ( .A(n1435), .B(n744), .Z(n1436) );
  NANDN U2669 ( .B(n717), .A(n1522), .Z(n1521) );
  XNOR U2670 ( .A(n1526), .B(n1457), .Z(n1447) );
  XNOR U2671 ( .A(n1444), .B(n1445), .Z(n1457) );
  NANDN U2672 ( .B(n834), .A(n1246), .Z(n1445) );
  XNOR U2673 ( .A(n1443), .B(n1527), .Z(n1444) );
  AND U2674 ( .A(n1178), .B(n872), .Z(n1527) );
  XNOR U2675 ( .A(n1456), .B(n1446), .Z(n1526) );
  XNOR U2676 ( .A(n1451), .B(n1535), .Z(n1452) );
  AND U2677 ( .A(n1055), .B(n984), .Z(n1535) );
  XOR U2678 ( .A(n1539), .B(n1453), .Z(n1534) );
  NAND U2679 ( .A(n928), .B(n1116), .Z(n1453) );
  IV U2680 ( .A(n1455), .Z(n1539) );
  XNOR U2681 ( .A(n1460), .B(n1544), .Z(n1461) );
  AND U2682 ( .A(n1316), .B(n806), .Z(n1544) );
  XOR U2683 ( .A(n1548), .B(n1462), .Z(n1543) );
  NAND U2684 ( .A(n771), .B(n1390), .Z(n1462) );
  IV U2685 ( .A(n1464), .Z(n1548) );
  XOR U2686 ( .A(n1549), .B(n1550), .Z(n1464) );
  ANDN U2687 ( .A(n1551), .B(n1552), .Z(n1550) );
  XOR U2688 ( .A(n1549), .B(n1553), .Z(n1551) );
  XNOR U2689 ( .A(n1471), .B(n1472), .Z(n1466) );
  NANDN U2690 ( .B(n716), .A(n1554), .Z(n1472) );
  AND U2691 ( .A(n1467), .B(n746), .Z(n1555) );
  NAND U2692 ( .A(n1556), .B(n1557), .Z(n1470) );
  NANDN U2693 ( .B(n1558), .A(n1559), .Z(n1556) );
  XOR U2694 ( .A(n1563), .B(\_MxM/Y0[14] ), .Z(\_MxM/Y1[13] ) );
  XNOR U2695 ( .A(n1564), .B(n1565), .Z(n1563) );
  AND U2696 ( .A(n674), .B(n1567), .Z(n1566) );
  XOR U2697 ( .A(n1561), .B(n1565), .Z(n1567) );
  XNOR U2698 ( .A(n1560), .B(n1565), .Z(n1561) );
  XNOR U2699 ( .A(n1490), .B(n1489), .Z(n1565) );
  XNOR U2700 ( .A(n1568), .B(n1486), .Z(n1489) );
  NAND U2701 ( .A(n1483), .B(n1571), .Z(n1487) );
  AND U2702 ( .A(n1572), .B(n1573), .Z(n1571) );
  NANDN U2703 ( .B(n717), .A(n1574), .Z(n1573) );
  NANDN U2704 ( .B(n1575), .A(n1576), .Z(n1572) );
  AND U2705 ( .A(n1577), .B(n1578), .Z(n1483) );
  NANDN U2706 ( .B(n1579), .A(n1580), .Z(n1578) );
  NANDN U2707 ( .B(n1581), .A(n1582), .Z(n1577) );
  XNOR U2708 ( .A(n1586), .B(n1515), .Z(n1506) );
  XNOR U2709 ( .A(n1494), .B(n1588), .Z(n1495) );
  AND U2710 ( .A(n897), .B(n1196), .Z(n1588) );
  XOR U2711 ( .A(n1592), .B(n1496), .Z(n1587) );
  NAND U2712 ( .A(n1138), .B(n941), .Z(n1496) );
  IV U2713 ( .A(n1498), .Z(n1592) );
  XNOR U2714 ( .A(n1503), .B(n1504), .Z(n1500) );
  NANDN U2715 ( .B(n1020), .A(n1055), .Z(n1504) );
  XNOR U2716 ( .A(n1502), .B(n1596), .Z(n1503) );
  AND U2717 ( .A(n1001), .B(n1079), .Z(n1596) );
  XNOR U2718 ( .A(n1514), .B(n1505), .Z(n1586) );
  XOR U2719 ( .A(n1603), .B(n1519), .Z(n1514) );
  XNOR U2720 ( .A(n1511), .B(n1512), .Z(n1519) );
  NAND U2721 ( .A(n1284), .B(n853), .Z(n1512) );
  XNOR U2722 ( .A(n1510), .B(n1604), .Z(n1511) );
  AND U2723 ( .A(n814), .B(n1352), .Z(n1604) );
  XNOR U2724 ( .A(n1518), .B(n1513), .Z(n1603) );
  XNOR U2725 ( .A(n1523), .B(n1612), .Z(n1524) );
  AND U2726 ( .A(n744), .B(n1522), .Z(n1612) );
  XOR U2727 ( .A(n1616), .B(n1525), .Z(n1611) );
  NAND U2728 ( .A(n1435), .B(n775), .Z(n1525) );
  IV U2729 ( .A(n1517), .Z(n1616) );
  XNOR U2730 ( .A(n1620), .B(n1542), .Z(n1532) );
  XNOR U2731 ( .A(n1529), .B(n1530), .Z(n1542) );
  NANDN U2732 ( .B(n834), .A(n1316), .Z(n1530) );
  XNOR U2733 ( .A(n1528), .B(n1621), .Z(n1529) );
  AND U2734 ( .A(n1246), .B(n872), .Z(n1621) );
  XNOR U2735 ( .A(n1541), .B(n1531), .Z(n1620) );
  XNOR U2736 ( .A(n1536), .B(n1629), .Z(n1537) );
  AND U2737 ( .A(n1116), .B(n984), .Z(n1629) );
  XOR U2738 ( .A(n1633), .B(n1538), .Z(n1628) );
  NAND U2739 ( .A(n928), .B(n1178), .Z(n1538) );
  IV U2740 ( .A(n1540), .Z(n1633) );
  XNOR U2741 ( .A(n1545), .B(n1638), .Z(n1546) );
  AND U2742 ( .A(n1390), .B(n806), .Z(n1638) );
  XOR U2743 ( .A(n1642), .B(n1547), .Z(n1637) );
  NAND U2744 ( .A(n771), .B(n1467), .Z(n1547) );
  IV U2745 ( .A(n1549), .Z(n1642) );
  XNOR U2746 ( .A(n1558), .B(n1559), .Z(n1553) );
  NANDN U2747 ( .B(n716), .A(n1646), .Z(n1559) );
  XNOR U2748 ( .A(n1557), .B(n1647), .Z(n1558) );
  AND U2749 ( .A(n1554), .B(n746), .Z(n1647) );
  ANDN U2750 ( .A(n1648), .B(n1649), .Z(n1557) );
  NANDN U2751 ( .B(n1650), .A(n1651), .Z(n1648) );
  XOR U2752 ( .A(n1655), .B(\_MxM/Y0[13] ), .Z(\_MxM/Y1[12] ) );
  XNOR U2753 ( .A(n1656), .B(n1657), .Z(n1655) );
  AND U2754 ( .A(n674), .B(n1659), .Z(n1658) );
  XOR U2755 ( .A(n1653), .B(n1657), .Z(n1659) );
  XNOR U2756 ( .A(n1652), .B(n1657), .Z(n1653) );
  XNOR U2757 ( .A(n1585), .B(n1584), .Z(n1657) );
  XNOR U2758 ( .A(n1660), .B(n1570), .Z(n1584) );
  XNOR U2759 ( .A(n1576), .B(n1575), .Z(n1570) );
  OR U2760 ( .A(n1661), .B(n1662), .Z(n1575) );
  XNOR U2761 ( .A(n1579), .B(n1580), .Z(n1576) );
  XOR U2762 ( .A(n1666), .B(n1581), .Z(n1579) );
  NAND U2763 ( .A(n744), .B(n1574), .Z(n1581) );
  NANDN U2764 ( .B(n1582), .A(n1667), .Z(n1666) );
  NANDN U2765 ( .B(n717), .A(n1668), .Z(n1667) );
  XNOR U2766 ( .A(n1677), .B(n1610), .Z(n1601) );
  XNOR U2767 ( .A(n1589), .B(n1679), .Z(n1590) );
  AND U2768 ( .A(n941), .B(n1196), .Z(n1679) );
  XOR U2769 ( .A(n1683), .B(n1591), .Z(n1678) );
  NAND U2770 ( .A(n1138), .B(n1001), .Z(n1591) );
  IV U2771 ( .A(n1593), .Z(n1683) );
  XNOR U2772 ( .A(n1598), .B(n1599), .Z(n1595) );
  NANDN U2773 ( .B(n1020), .A(n1116), .Z(n1599) );
  XNOR U2774 ( .A(n1597), .B(n1687), .Z(n1598) );
  AND U2775 ( .A(n1055), .B(n1079), .Z(n1687) );
  XNOR U2776 ( .A(n1609), .B(n1600), .Z(n1677) );
  XOR U2777 ( .A(n1694), .B(n1619), .Z(n1609) );
  XNOR U2778 ( .A(n1606), .B(n1607), .Z(n1619) );
  NAND U2779 ( .A(n1284), .B(n897), .Z(n1607) );
  XNOR U2780 ( .A(n1605), .B(n1695), .Z(n1606) );
  AND U2781 ( .A(n853), .B(n1352), .Z(n1695) );
  XNOR U2782 ( .A(n1618), .B(n1608), .Z(n1694) );
  XNOR U2783 ( .A(n1613), .B(n1703), .Z(n1614) );
  AND U2784 ( .A(n775), .B(n1522), .Z(n1703) );
  XOR U2785 ( .A(n1707), .B(n1615), .Z(n1702) );
  NAND U2786 ( .A(n1435), .B(n814), .Z(n1615) );
  IV U2787 ( .A(n1617), .Z(n1707) );
  XNOR U2788 ( .A(n1711), .B(n1636), .Z(n1626) );
  XNOR U2789 ( .A(n1623), .B(n1624), .Z(n1636) );
  NANDN U2790 ( .B(n834), .A(n1390), .Z(n1624) );
  XNOR U2791 ( .A(n1622), .B(n1712), .Z(n1623) );
  AND U2792 ( .A(n1316), .B(n872), .Z(n1712) );
  XNOR U2793 ( .A(n1635), .B(n1625), .Z(n1711) );
  XNOR U2794 ( .A(n1630), .B(n1720), .Z(n1631) );
  AND U2795 ( .A(n1178), .B(n984), .Z(n1720) );
  XOR U2796 ( .A(n1724), .B(n1632), .Z(n1719) );
  NAND U2797 ( .A(n928), .B(n1246), .Z(n1632) );
  IV U2798 ( .A(n1634), .Z(n1724) );
  XNOR U2799 ( .A(n1639), .B(n1729), .Z(n1640) );
  AND U2800 ( .A(n1467), .B(n806), .Z(n1729) );
  XOR U2801 ( .A(n1733), .B(n1641), .Z(n1728) );
  NAND U2802 ( .A(n771), .B(n1554), .Z(n1641) );
  IV U2803 ( .A(n1643), .Z(n1733) );
  XNOR U2804 ( .A(n1650), .B(n1651), .Z(n1645) );
  NANDN U2805 ( .B(n716), .A(n1737), .Z(n1651) );
  AND U2806 ( .A(n1646), .B(n746), .Z(n1738) );
  NAND U2807 ( .A(n1739), .B(n1740), .Z(n1649) );
  NANDN U2808 ( .B(n1741), .A(n1742), .Z(n1739) );
  XOR U2809 ( .A(n1746), .B(\_MxM/Y0[12] ), .Z(\_MxM/Y1[11] ) );
  XNOR U2810 ( .A(n1747), .B(n1748), .Z(n1746) );
  AND U2811 ( .A(n674), .B(n1750), .Z(n1749) );
  XOR U2812 ( .A(n1744), .B(n1748), .Z(n1750) );
  XNOR U2813 ( .A(n1743), .B(n1748), .Z(n1744) );
  XNOR U2814 ( .A(n1674), .B(n1673), .Z(n1748) );
  XNOR U2815 ( .A(n1751), .B(n1676), .Z(n1673) );
  XOR U2816 ( .A(n1662), .B(n1661), .Z(n1676) );
  NANDN U2817 ( .B(n1752), .A(n1753), .Z(n1661) );
  XOR U2818 ( .A(n1665), .B(n1664), .Z(n1662) );
  XOR U2819 ( .A(n1663), .B(n1754), .Z(n1664) );
  AND U2820 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U2821 ( .B(n717), .A(n1757), .Z(n1756) );
  OR U2822 ( .A(n1758), .B(n1759), .Z(n1755) );
  NAND U2823 ( .A(n775), .B(n1574), .Z(n1671) );
  XNOR U2824 ( .A(n1669), .B(n1762), .Z(n1670) );
  AND U2825 ( .A(n1668), .B(n744), .Z(n1762) );
  XNOR U2826 ( .A(n1771), .B(n1701), .Z(n1692) );
  XNOR U2827 ( .A(n1680), .B(n1773), .Z(n1681) );
  AND U2828 ( .A(n1001), .B(n1196), .Z(n1773) );
  XOR U2829 ( .A(n1777), .B(n1682), .Z(n1772) );
  NAND U2830 ( .A(n1138), .B(n1055), .Z(n1682) );
  IV U2831 ( .A(n1684), .Z(n1777) );
  XNOR U2832 ( .A(n1689), .B(n1690), .Z(n1686) );
  NANDN U2833 ( .B(n1020), .A(n1178), .Z(n1690) );
  XNOR U2834 ( .A(n1688), .B(n1781), .Z(n1689) );
  AND U2835 ( .A(n1116), .B(n1079), .Z(n1781) );
  XNOR U2836 ( .A(n1700), .B(n1691), .Z(n1771) );
  XOR U2837 ( .A(n1788), .B(n1710), .Z(n1700) );
  XNOR U2838 ( .A(n1697), .B(n1698), .Z(n1710) );
  NAND U2839 ( .A(n1284), .B(n941), .Z(n1698) );
  XNOR U2840 ( .A(n1696), .B(n1789), .Z(n1697) );
  AND U2841 ( .A(n897), .B(n1352), .Z(n1789) );
  XNOR U2842 ( .A(n1709), .B(n1699), .Z(n1788) );
  XNOR U2843 ( .A(n1704), .B(n1797), .Z(n1705) );
  AND U2844 ( .A(n814), .B(n1522), .Z(n1797) );
  XOR U2845 ( .A(n1801), .B(n1706), .Z(n1796) );
  NAND U2846 ( .A(n1435), .B(n853), .Z(n1706) );
  IV U2847 ( .A(n1708), .Z(n1801) );
  XNOR U2848 ( .A(n1805), .B(n1727), .Z(n1717) );
  XNOR U2849 ( .A(n1714), .B(n1715), .Z(n1727) );
  NANDN U2850 ( .B(n834), .A(n1467), .Z(n1715) );
  XNOR U2851 ( .A(n1713), .B(n1806), .Z(n1714) );
  AND U2852 ( .A(n1390), .B(n872), .Z(n1806) );
  XNOR U2853 ( .A(n1726), .B(n1716), .Z(n1805) );
  XNOR U2854 ( .A(n1721), .B(n1814), .Z(n1722) );
  AND U2855 ( .A(n1246), .B(n984), .Z(n1814) );
  XOR U2856 ( .A(n1818), .B(n1723), .Z(n1813) );
  NAND U2857 ( .A(n928), .B(n1316), .Z(n1723) );
  IV U2858 ( .A(n1725), .Z(n1818) );
  XNOR U2859 ( .A(n1730), .B(n1823), .Z(n1731) );
  AND U2860 ( .A(n1554), .B(n806), .Z(n1823) );
  XOR U2861 ( .A(n1827), .B(n1732), .Z(n1822) );
  NAND U2862 ( .A(n771), .B(n1646), .Z(n1732) );
  IV U2863 ( .A(n1734), .Z(n1827) );
  XNOR U2864 ( .A(n1741), .B(n1742), .Z(n1736) );
  NANDN U2865 ( .B(n716), .A(n1831), .Z(n1742) );
  XNOR U2866 ( .A(n1740), .B(n1832), .Z(n1741) );
  AND U2867 ( .A(n1737), .B(n746), .Z(n1832) );
  ANDN U2868 ( .A(n1833), .B(n1834), .Z(n1740) );
  NANDN U2869 ( .B(n1835), .A(n1836), .Z(n1833) );
  XOR U2870 ( .A(n1840), .B(\_MxM/Y0[11] ), .Z(\_MxM/Y1[10] ) );
  XNOR U2871 ( .A(n1841), .B(n1842), .Z(n1840) );
  AND U2872 ( .A(n674), .B(n1844), .Z(n1843) );
  XOR U2873 ( .A(n1838), .B(n1842), .Z(n1844) );
  XNOR U2874 ( .A(n1837), .B(n1842), .Z(n1838) );
  XNOR U2875 ( .A(n1768), .B(n1767), .Z(n1842) );
  XNOR U2876 ( .A(n1845), .B(n1770), .Z(n1767) );
  XNOR U2877 ( .A(n1752), .B(n1753), .Z(n1770) );
  XOR U2878 ( .A(n1761), .B(n1760), .Z(n1752) );
  XNOR U2879 ( .A(n1849), .B(n1850), .Z(n1760) );
  ANDN U2880 ( .A(n1853), .B(n1854), .Z(n1852) );
  XOR U2881 ( .A(n1851), .B(n1855), .Z(n1853) );
  XNOR U2882 ( .A(n1856), .B(n1758), .Z(n1849) );
  NAND U2883 ( .A(n744), .B(n1757), .Z(n1758) );
  NANDN U2884 ( .B(n717), .A(n1858), .Z(n1857) );
  NAND U2885 ( .A(n814), .B(n1574), .Z(n1765) );
  XNOR U2886 ( .A(n1763), .B(n1862), .Z(n1764) );
  AND U2887 ( .A(n1668), .B(n775), .Z(n1862) );
  XNOR U2888 ( .A(n1871), .B(n1795), .Z(n1786) );
  XNOR U2889 ( .A(n1774), .B(n1873), .Z(n1775) );
  AND U2890 ( .A(n1055), .B(n1196), .Z(n1873) );
  XOR U2891 ( .A(n1877), .B(n1776), .Z(n1872) );
  NAND U2892 ( .A(n1138), .B(n1116), .Z(n1776) );
  IV U2893 ( .A(n1778), .Z(n1877) );
  XNOR U2894 ( .A(n1783), .B(n1784), .Z(n1780) );
  NANDN U2895 ( .B(n1020), .A(n1246), .Z(n1784) );
  XNOR U2896 ( .A(n1782), .B(n1881), .Z(n1783) );
  AND U2897 ( .A(n1178), .B(n1079), .Z(n1881) );
  XNOR U2898 ( .A(n1794), .B(n1785), .Z(n1871) );
  XOR U2899 ( .A(n1888), .B(n1804), .Z(n1794) );
  XNOR U2900 ( .A(n1791), .B(n1792), .Z(n1804) );
  NAND U2901 ( .A(n1284), .B(n1001), .Z(n1792) );
  XNOR U2902 ( .A(n1790), .B(n1889), .Z(n1791) );
  AND U2903 ( .A(n941), .B(n1352), .Z(n1889) );
  XNOR U2904 ( .A(n1803), .B(n1793), .Z(n1888) );
  XNOR U2905 ( .A(n1798), .B(n1897), .Z(n1799) );
  AND U2906 ( .A(n853), .B(n1522), .Z(n1897) );
  XOR U2907 ( .A(n1901), .B(n1800), .Z(n1896) );
  NAND U2908 ( .A(n1435), .B(n897), .Z(n1800) );
  IV U2909 ( .A(n1802), .Z(n1901) );
  XNOR U2910 ( .A(n1905), .B(n1821), .Z(n1811) );
  XNOR U2911 ( .A(n1808), .B(n1809), .Z(n1821) );
  NANDN U2912 ( .B(n834), .A(n1554), .Z(n1809) );
  XNOR U2913 ( .A(n1807), .B(n1906), .Z(n1808) );
  AND U2914 ( .A(n1467), .B(n872), .Z(n1906) );
  XNOR U2915 ( .A(n1820), .B(n1810), .Z(n1905) );
  XNOR U2916 ( .A(n1815), .B(n1914), .Z(n1816) );
  AND U2917 ( .A(n1316), .B(n984), .Z(n1914) );
  XOR U2918 ( .A(n1918), .B(n1817), .Z(n1913) );
  NAND U2919 ( .A(n928), .B(n1390), .Z(n1817) );
  IV U2920 ( .A(n1819), .Z(n1918) );
  XNOR U2921 ( .A(n1824), .B(n1923), .Z(n1825) );
  AND U2922 ( .A(n1646), .B(n806), .Z(n1923) );
  XOR U2923 ( .A(n1927), .B(n1826), .Z(n1922) );
  NAND U2924 ( .A(n771), .B(n1737), .Z(n1826) );
  IV U2925 ( .A(n1828), .Z(n1927) );
  XNOR U2926 ( .A(n1835), .B(n1836), .Z(n1830) );
  NANDN U2927 ( .B(n716), .A(n1931), .Z(n1836) );
  AND U2928 ( .A(n1831), .B(n746), .Z(n1932) );
  NAND U2929 ( .A(n1933), .B(n1934), .Z(n1834) );
  NANDN U2930 ( .B(n1935), .A(n1936), .Z(n1933) );
  XNOR U2931 ( .A(n1940), .B(n1941), .Z(n658) );
  AND U2932 ( .A(n674), .B(n1943), .Z(n1942) );
  XOR U2933 ( .A(n1938), .B(n1941), .Z(n1943) );
  XNOR U2934 ( .A(n1937), .B(n1941), .Z(n1938) );
  XNOR U2935 ( .A(n1868), .B(n1867), .Z(n1941) );
  XNOR U2936 ( .A(n1944), .B(n1870), .Z(n1867) );
  XNOR U2937 ( .A(n1848), .B(n1847), .Z(n1870) );
  XNOR U2938 ( .A(n1846), .B(n1945), .Z(n1847) );
  AND U2939 ( .A(n1946), .B(n1947), .Z(n1945) );
  OR U2940 ( .A(n1948), .B(n1949), .Z(n1947) );
  AND U2941 ( .A(n1950), .B(n1951), .Z(n1946) );
  NANDN U2942 ( .B(n717), .A(n1952), .Z(n1951) );
  NAND U2943 ( .A(n1953), .B(n1954), .Z(n1950) );
  XNOR U2944 ( .A(n1859), .B(n1959), .Z(n1860) );
  AND U2945 ( .A(n1858), .B(n744), .Z(n1959) );
  XOR U2946 ( .A(n1963), .B(n1861), .Z(n1958) );
  NAND U2947 ( .A(n775), .B(n1757), .Z(n1861) );
  IV U2948 ( .A(n1851), .Z(n1963) );
  XNOR U2949 ( .A(n1864), .B(n1865), .Z(n1855) );
  NAND U2950 ( .A(n853), .B(n1574), .Z(n1865) );
  XNOR U2951 ( .A(n1863), .B(n1967), .Z(n1864) );
  AND U2952 ( .A(n1668), .B(n814), .Z(n1967) );
  XNOR U2953 ( .A(n1976), .B(n1895), .Z(n1886) );
  XNOR U2954 ( .A(n1874), .B(n1978), .Z(n1875) );
  AND U2955 ( .A(n1116), .B(n1196), .Z(n1978) );
  XOR U2956 ( .A(n1982), .B(n1876), .Z(n1977) );
  NAND U2957 ( .A(n1138), .B(n1178), .Z(n1876) );
  IV U2958 ( .A(n1878), .Z(n1982) );
  XNOR U2959 ( .A(n1883), .B(n1884), .Z(n1880) );
  NANDN U2960 ( .B(n1020), .A(n1316), .Z(n1884) );
  XNOR U2961 ( .A(n1882), .B(n1986), .Z(n1883) );
  AND U2962 ( .A(n1246), .B(n1079), .Z(n1986) );
  XNOR U2963 ( .A(n1894), .B(n1885), .Z(n1976) );
  XOR U2964 ( .A(n1993), .B(n1904), .Z(n1894) );
  XNOR U2965 ( .A(n1891), .B(n1892), .Z(n1904) );
  NAND U2966 ( .A(n1284), .B(n1055), .Z(n1892) );
  XNOR U2967 ( .A(n1890), .B(n1994), .Z(n1891) );
  AND U2968 ( .A(n1001), .B(n1352), .Z(n1994) );
  XNOR U2969 ( .A(n1903), .B(n1893), .Z(n1993) );
  XNOR U2970 ( .A(n1898), .B(n2002), .Z(n1899) );
  AND U2971 ( .A(n897), .B(n1522), .Z(n2002) );
  XOR U2972 ( .A(n2006), .B(n1900), .Z(n2001) );
  NAND U2973 ( .A(n1435), .B(n941), .Z(n1900) );
  IV U2974 ( .A(n1902), .Z(n2006) );
  XNOR U2975 ( .A(n2010), .B(n1921), .Z(n1911) );
  XNOR U2976 ( .A(n1908), .B(n1909), .Z(n1921) );
  NANDN U2977 ( .B(n834), .A(n1646), .Z(n1909) );
  XNOR U2978 ( .A(n1907), .B(n2011), .Z(n1908) );
  AND U2979 ( .A(n1554), .B(n872), .Z(n2011) );
  XNOR U2980 ( .A(n1920), .B(n1910), .Z(n2010) );
  XNOR U2981 ( .A(n1915), .B(n2019), .Z(n1916) );
  AND U2982 ( .A(n1390), .B(n984), .Z(n2019) );
  XOR U2983 ( .A(n2023), .B(n1917), .Z(n2018) );
  NAND U2984 ( .A(n928), .B(n1467), .Z(n1917) );
  IV U2985 ( .A(n1919), .Z(n2023) );
  XNOR U2986 ( .A(n1924), .B(n2028), .Z(n1925) );
  AND U2987 ( .A(n1737), .B(n806), .Z(n2028) );
  XOR U2988 ( .A(n2032), .B(n1926), .Z(n2027) );
  NAND U2989 ( .A(n771), .B(n1831), .Z(n1926) );
  IV U2990 ( .A(n1928), .Z(n2032) );
  XNOR U2991 ( .A(n1935), .B(n1936), .Z(n1930) );
  NANDN U2992 ( .B(n716), .A(n2036), .Z(n1936) );
  XNOR U2993 ( .A(n1934), .B(n2037), .Z(n1935) );
  AND U2994 ( .A(n1931), .B(n746), .Z(n2037) );
  ANDN U2995 ( .A(n2038), .B(n2039), .Z(n1934) );
  NANDN U2996 ( .B(n2040), .A(n2041), .Z(n2038) );
  XNOR U2997 ( .A(n2045), .B(n2046), .Z(n659) );
  AND U2998 ( .A(n674), .B(n2048), .Z(n2047) );
  XOR U2999 ( .A(n2043), .B(n2046), .Z(n2048) );
  XNOR U3000 ( .A(n2042), .B(n2046), .Z(n2043) );
  XNOR U3001 ( .A(n1973), .B(n1972), .Z(n2046) );
  XNOR U3002 ( .A(n2049), .B(n1975), .Z(n1972) );
  XNOR U3003 ( .A(n1957), .B(n1956), .Z(n1975) );
  XNOR U3004 ( .A(n2050), .B(n1953), .Z(n1956) );
  XNOR U3005 ( .A(n2051), .B(n1948), .Z(n1953) );
  NAND U3006 ( .A(n744), .B(n1952), .Z(n1948) );
  NANDN U3007 ( .B(n717), .A(n2053), .Z(n2052) );
  XNOR U3008 ( .A(n1954), .B(n1955), .Z(n2050) );
  XNOR U3009 ( .A(n1960), .B(n2064), .Z(n1961) );
  AND U3010 ( .A(n1858), .B(n775), .Z(n2064) );
  XOR U3011 ( .A(n2068), .B(n1962), .Z(n2063) );
  NAND U3012 ( .A(n814), .B(n1757), .Z(n1962) );
  IV U3013 ( .A(n1964), .Z(n2068) );
  XNOR U3014 ( .A(n1969), .B(n1970), .Z(n1966) );
  NAND U3015 ( .A(n897), .B(n1574), .Z(n1970) );
  XNOR U3016 ( .A(n1968), .B(n2072), .Z(n1969) );
  AND U3017 ( .A(n1668), .B(n853), .Z(n2072) );
  XNOR U3018 ( .A(n2081), .B(n2000), .Z(n1991) );
  XNOR U3019 ( .A(n1979), .B(n2083), .Z(n1980) );
  AND U3020 ( .A(n1178), .B(n1196), .Z(n2083) );
  XOR U3021 ( .A(n2087), .B(n1981), .Z(n2082) );
  NAND U3022 ( .A(n1138), .B(n1246), .Z(n1981) );
  IV U3023 ( .A(n1983), .Z(n2087) );
  XNOR U3024 ( .A(n1988), .B(n1989), .Z(n1985) );
  NANDN U3025 ( .B(n1020), .A(n1390), .Z(n1989) );
  XNOR U3026 ( .A(n1987), .B(n2091), .Z(n1988) );
  AND U3027 ( .A(n1316), .B(n1079), .Z(n2091) );
  XNOR U3028 ( .A(n1999), .B(n1990), .Z(n2081) );
  XOR U3029 ( .A(n2098), .B(n2009), .Z(n1999) );
  XNOR U3030 ( .A(n1996), .B(n1997), .Z(n2009) );
  NAND U3031 ( .A(n1284), .B(n1116), .Z(n1997) );
  XNOR U3032 ( .A(n1995), .B(n2099), .Z(n1996) );
  AND U3033 ( .A(n1055), .B(n1352), .Z(n2099) );
  XNOR U3034 ( .A(n2008), .B(n1998), .Z(n2098) );
  XNOR U3035 ( .A(n2003), .B(n2107), .Z(n2004) );
  AND U3036 ( .A(n941), .B(n1522), .Z(n2107) );
  XOR U3037 ( .A(n2111), .B(n2005), .Z(n2106) );
  NAND U3038 ( .A(n1435), .B(n1001), .Z(n2005) );
  IV U3039 ( .A(n2007), .Z(n2111) );
  XNOR U3040 ( .A(n2115), .B(n2026), .Z(n2016) );
  XNOR U3041 ( .A(n2013), .B(n2014), .Z(n2026) );
  NANDN U3042 ( .B(n834), .A(n1737), .Z(n2014) );
  XNOR U3043 ( .A(n2012), .B(n2116), .Z(n2013) );
  AND U3044 ( .A(n1646), .B(n872), .Z(n2116) );
  XNOR U3045 ( .A(n2025), .B(n2015), .Z(n2115) );
  XNOR U3046 ( .A(n2020), .B(n2124), .Z(n2021) );
  AND U3047 ( .A(n1467), .B(n984), .Z(n2124) );
  XOR U3048 ( .A(n2128), .B(n2022), .Z(n2123) );
  NAND U3049 ( .A(n928), .B(n1554), .Z(n2022) );
  IV U3050 ( .A(n2024), .Z(n2128) );
  XNOR U3051 ( .A(n2029), .B(n2133), .Z(n2030) );
  AND U3052 ( .A(n1831), .B(n806), .Z(n2133) );
  XOR U3053 ( .A(n2137), .B(n2031), .Z(n2132) );
  NAND U3054 ( .A(n771), .B(n1931), .Z(n2031) );
  IV U3055 ( .A(n2033), .Z(n2137) );
  XNOR U3056 ( .A(n2040), .B(n2041), .Z(n2035) );
  NANDN U3057 ( .B(n716), .A(n2141), .Z(n2041) );
  AND U3058 ( .A(n2036), .B(n746), .Z(n2142) );
  NAND U3059 ( .A(n2143), .B(n2144), .Z(n2039) );
  NANDN U3060 ( .B(n2145), .A(n2146), .Z(n2143) );
  XNOR U3061 ( .A(n2150), .B(n2151), .Z(n660) );
  AND U3062 ( .A(n674), .B(n2153), .Z(n2152) );
  XOR U3063 ( .A(n2148), .B(n2151), .Z(n2153) );
  XNOR U3064 ( .A(n2147), .B(n2151), .Z(n2148) );
  XNOR U3065 ( .A(n2078), .B(n2077), .Z(n2151) );
  XNOR U3066 ( .A(n2154), .B(n2080), .Z(n2077) );
  XNOR U3067 ( .A(n2059), .B(n2058), .Z(n2080) );
  XNOR U3068 ( .A(n2155), .B(n2062), .Z(n2058) );
  XNOR U3069 ( .A(n2055), .B(n2056), .Z(n2062) );
  NAND U3070 ( .A(n775), .B(n1952), .Z(n2056) );
  XNOR U3071 ( .A(n2054), .B(n2156), .Z(n2055) );
  AND U3072 ( .A(n2053), .B(n744), .Z(n2156) );
  XNOR U3073 ( .A(n2061), .B(n2057), .Z(n2155) );
  AND U3074 ( .A(n2164), .B(n2165), .Z(n2163) );
  NANDN U3075 ( .B(n717), .A(n2166), .Z(n2165) );
  OR U3076 ( .A(n2167), .B(n2168), .Z(n2164) );
  XNOR U3077 ( .A(n2065), .B(n2173), .Z(n2066) );
  AND U3078 ( .A(n1858), .B(n814), .Z(n2173) );
  XOR U3079 ( .A(n2177), .B(n2067), .Z(n2172) );
  NAND U3080 ( .A(n853), .B(n1757), .Z(n2067) );
  IV U3081 ( .A(n2069), .Z(n2177) );
  XNOR U3082 ( .A(n2074), .B(n2075), .Z(n2071) );
  NAND U3083 ( .A(n941), .B(n1574), .Z(n2075) );
  XNOR U3084 ( .A(n2073), .B(n2181), .Z(n2074) );
  AND U3085 ( .A(n1668), .B(n897), .Z(n2181) );
  XNOR U3086 ( .A(n2191), .B(n2188), .Z(n2190) );
  XNOR U3087 ( .A(n2192), .B(n2105), .Z(n2096) );
  XNOR U3088 ( .A(n2084), .B(n2194), .Z(n2085) );
  AND U3089 ( .A(n1246), .B(n1196), .Z(n2194) );
  XOR U3090 ( .A(n2198), .B(n2086), .Z(n2193) );
  NAND U3091 ( .A(n1138), .B(n1316), .Z(n2086) );
  IV U3092 ( .A(n2088), .Z(n2198) );
  XNOR U3093 ( .A(n2093), .B(n2094), .Z(n2090) );
  NANDN U3094 ( .B(n1020), .A(n1467), .Z(n2094) );
  XNOR U3095 ( .A(n2092), .B(n2202), .Z(n2093) );
  AND U3096 ( .A(n1390), .B(n1079), .Z(n2202) );
  XNOR U3097 ( .A(n2104), .B(n2095), .Z(n2192) );
  XOR U3098 ( .A(n2209), .B(n2114), .Z(n2104) );
  XNOR U3099 ( .A(n2101), .B(n2102), .Z(n2114) );
  NAND U3100 ( .A(n1284), .B(n1178), .Z(n2102) );
  XNOR U3101 ( .A(n2100), .B(n2210), .Z(n2101) );
  AND U3102 ( .A(n1116), .B(n1352), .Z(n2210) );
  XNOR U3103 ( .A(n2113), .B(n2103), .Z(n2209) );
  XNOR U3104 ( .A(n2108), .B(n2218), .Z(n2109) );
  AND U3105 ( .A(n1001), .B(n1522), .Z(n2218) );
  XOR U3106 ( .A(n2222), .B(n2110), .Z(n2217) );
  NAND U3107 ( .A(n1435), .B(n1055), .Z(n2110) );
  IV U3108 ( .A(n2112), .Z(n2222) );
  XNOR U3109 ( .A(n2226), .B(n2131), .Z(n2121) );
  XNOR U3110 ( .A(n2118), .B(n2119), .Z(n2131) );
  NANDN U3111 ( .B(n834), .A(n1831), .Z(n2119) );
  XNOR U3112 ( .A(n2117), .B(n2227), .Z(n2118) );
  AND U3113 ( .A(n1737), .B(n872), .Z(n2227) );
  XNOR U3114 ( .A(n2130), .B(n2120), .Z(n2226) );
  XNOR U3115 ( .A(n2125), .B(n2235), .Z(n2126) );
  AND U3116 ( .A(n1554), .B(n984), .Z(n2235) );
  XOR U3117 ( .A(n2239), .B(n2127), .Z(n2234) );
  NAND U3118 ( .A(n928), .B(n1646), .Z(n2127) );
  IV U3119 ( .A(n2129), .Z(n2239) );
  XNOR U3120 ( .A(n2134), .B(n2244), .Z(n2135) );
  AND U3121 ( .A(n1931), .B(n806), .Z(n2244) );
  XOR U3122 ( .A(n2245), .B(n2246), .Z(n2134) );
  ANDN U3123 ( .A(n2247), .B(n2248), .Z(n2246) );
  XNOR U3124 ( .A(n2249), .B(n2245), .Z(n2247) );
  XOR U3125 ( .A(n2250), .B(n2136), .Z(n2243) );
  NAND U3126 ( .A(n771), .B(n2036), .Z(n2136) );
  IV U3127 ( .A(n2138), .Z(n2250) );
  XNOR U3128 ( .A(n2145), .B(n2146), .Z(n2140) );
  NANDN U3129 ( .B(n716), .A(n2254), .Z(n2146) );
  XNOR U3130 ( .A(n2144), .B(n2255), .Z(n2145) );
  AND U3131 ( .A(n2141), .B(n746), .Z(n2255) );
  ANDN U3132 ( .A(n2256), .B(n2257), .Z(n2144) );
  NANDN U3133 ( .B(n2258), .A(n2259), .Z(n2256) );
  XNOR U3134 ( .A(n2263), .B(n2264), .Z(n661) );
  AND U3135 ( .A(n674), .B(n2266), .Z(n2265) );
  XOR U3136 ( .A(n2261), .B(n2264), .Z(n2266) );
  XNOR U3137 ( .A(n2260), .B(n2264), .Z(n2261) );
  XNOR U3138 ( .A(n2187), .B(n2186), .Z(n2264) );
  XNOR U3139 ( .A(n2267), .B(n2191), .Z(n2186) );
  XNOR U3140 ( .A(n2162), .B(n2161), .Z(n2191) );
  XNOR U3141 ( .A(n2268), .B(n2171), .Z(n2161) );
  XNOR U3142 ( .A(n2158), .B(n2159), .Z(n2171) );
  NAND U3143 ( .A(n814), .B(n1952), .Z(n2159) );
  XNOR U3144 ( .A(n2157), .B(n2269), .Z(n2158) );
  AND U3145 ( .A(n2053), .B(n775), .Z(n2269) );
  XNOR U3146 ( .A(n2170), .B(n2160), .Z(n2268) );
  XNOR U3147 ( .A(n2276), .B(n2169), .Z(n2170) );
  XNOR U3148 ( .A(n2280), .B(n2167), .Z(n2276) );
  NAND U3149 ( .A(n744), .B(n2166), .Z(n2167) );
  NANDN U3150 ( .B(n717), .A(n2282), .Z(n2281) );
  XNOR U3151 ( .A(n2174), .B(n2287), .Z(n2175) );
  AND U3152 ( .A(n1858), .B(n853), .Z(n2287) );
  XOR U3153 ( .A(n2291), .B(n2176), .Z(n2286) );
  NAND U3154 ( .A(n897), .B(n1757), .Z(n2176) );
  IV U3155 ( .A(n2178), .Z(n2291) );
  XNOR U3156 ( .A(n2183), .B(n2184), .Z(n2180) );
  NAND U3157 ( .A(n1001), .B(n1574), .Z(n2184) );
  XNOR U3158 ( .A(n2182), .B(n2295), .Z(n2183) );
  AND U3159 ( .A(n1668), .B(n941), .Z(n2295) );
  XNOR U3160 ( .A(n2189), .B(n2185), .Z(n2267) );
  XOR U3161 ( .A(n2306), .B(n2307), .Z(n2302) );
  NANDN U3162 ( .B(n2308), .A(n2309), .Z(n2306) );
  XNOR U3163 ( .A(n2310), .B(n2216), .Z(n2207) );
  XNOR U3164 ( .A(n2195), .B(n2312), .Z(n2196) );
  AND U3165 ( .A(n1316), .B(n1196), .Z(n2312) );
  XOR U3166 ( .A(n2316), .B(n2197), .Z(n2311) );
  NAND U3167 ( .A(n1138), .B(n1390), .Z(n2197) );
  IV U3168 ( .A(n2199), .Z(n2316) );
  XNOR U3169 ( .A(n2204), .B(n2205), .Z(n2201) );
  NANDN U3170 ( .B(n1020), .A(n1554), .Z(n2205) );
  XNOR U3171 ( .A(n2203), .B(n2320), .Z(n2204) );
  AND U3172 ( .A(n1467), .B(n1079), .Z(n2320) );
  XNOR U3173 ( .A(n2215), .B(n2206), .Z(n2310) );
  XOR U3174 ( .A(n2327), .B(n2225), .Z(n2215) );
  XNOR U3175 ( .A(n2212), .B(n2213), .Z(n2225) );
  NAND U3176 ( .A(n1284), .B(n1246), .Z(n2213) );
  XNOR U3177 ( .A(n2211), .B(n2328), .Z(n2212) );
  AND U3178 ( .A(n1178), .B(n1352), .Z(n2328) );
  XNOR U3179 ( .A(n2224), .B(n2214), .Z(n2327) );
  XNOR U3180 ( .A(n2219), .B(n2336), .Z(n2220) );
  AND U3181 ( .A(n1055), .B(n1522), .Z(n2336) );
  XOR U3182 ( .A(n2340), .B(n2221), .Z(n2335) );
  NAND U3183 ( .A(n1435), .B(n1116), .Z(n2221) );
  IV U3184 ( .A(n2223), .Z(n2340) );
  XNOR U3185 ( .A(n2344), .B(n2242), .Z(n2232) );
  XNOR U3186 ( .A(n2229), .B(n2230), .Z(n2242) );
  NANDN U3187 ( .B(n834), .A(n1931), .Z(n2230) );
  XNOR U3188 ( .A(n2228), .B(n2345), .Z(n2229) );
  AND U3189 ( .A(n1831), .B(n872), .Z(n2345) );
  XNOR U3190 ( .A(n2241), .B(n2231), .Z(n2344) );
  XNOR U3191 ( .A(n2236), .B(n2353), .Z(n2237) );
  AND U3192 ( .A(n1646), .B(n984), .Z(n2353) );
  XOR U3193 ( .A(n2357), .B(n2238), .Z(n2352) );
  NAND U3194 ( .A(n928), .B(n1737), .Z(n2238) );
  IV U3195 ( .A(n2240), .Z(n2357) );
  XNOR U3196 ( .A(n2245), .B(n2362), .Z(n2248) );
  AND U3197 ( .A(n2036), .B(n806), .Z(n2362) );
  XOR U3198 ( .A(n2366), .B(n2249), .Z(n2361) );
  NAND U3199 ( .A(n771), .B(n2141), .Z(n2249) );
  IV U3200 ( .A(n2251), .Z(n2366) );
  XNOR U3201 ( .A(n2258), .B(n2259), .Z(n2253) );
  NANDN U3202 ( .B(n716), .A(n2370), .Z(n2259) );
  AND U3203 ( .A(n2254), .B(n746), .Z(n2371) );
  NAND U3204 ( .A(n2372), .B(n2373), .Z(n2257) );
  NANDN U3205 ( .B(n2374), .A(n2375), .Z(n2372) );
  XNOR U3206 ( .A(n2379), .B(n2380), .Z(n662) );
  AND U3207 ( .A(n674), .B(n2382), .Z(n2381) );
  XOR U3208 ( .A(n2377), .B(n2380), .Z(n2382) );
  XNOR U3209 ( .A(n2376), .B(n2380), .Z(n2377) );
  XNOR U3210 ( .A(n2301), .B(n2300), .Z(n2380) );
  XNOR U3211 ( .A(n2383), .B(n2305), .Z(n2300) );
  XNOR U3212 ( .A(n2384), .B(n2279), .Z(n2274) );
  XNOR U3213 ( .A(n2271), .B(n2272), .Z(n2279) );
  NAND U3214 ( .A(n853), .B(n1952), .Z(n2272) );
  XNOR U3215 ( .A(n2270), .B(n2385), .Z(n2271) );
  AND U3216 ( .A(n2053), .B(n814), .Z(n2385) );
  XNOR U3217 ( .A(n2278), .B(n2273), .Z(n2384) );
  XNOR U3218 ( .A(n2283), .B(n2393), .Z(n2284) );
  AND U3219 ( .A(n2282), .B(n744), .Z(n2393) );
  XOR U3220 ( .A(n2397), .B(n2285), .Z(n2392) );
  NAND U3221 ( .A(n775), .B(n2166), .Z(n2285) );
  IV U3222 ( .A(n2277), .Z(n2397) );
  XNOR U3223 ( .A(n2288), .B(n2402), .Z(n2289) );
  AND U3224 ( .A(n1858), .B(n897), .Z(n2402) );
  XOR U3225 ( .A(n2406), .B(n2290), .Z(n2401) );
  NAND U3226 ( .A(n941), .B(n1757), .Z(n2290) );
  IV U3227 ( .A(n2292), .Z(n2406) );
  XNOR U3228 ( .A(n2297), .B(n2298), .Z(n2294) );
  NAND U3229 ( .A(n1055), .B(n1574), .Z(n2298) );
  XNOR U3230 ( .A(n2296), .B(n2410), .Z(n2297) );
  AND U3231 ( .A(n1668), .B(n1001), .Z(n2410) );
  XNOR U3232 ( .A(n2304), .B(n2299), .Z(n2383) );
  AND U3233 ( .A(n2307), .B(n2418), .Z(n2417) );
  AND U3234 ( .A(n2419), .B(n2420), .Z(n2418) );
  NANDN U3235 ( .B(n717), .A(n2421), .Z(n2420) );
  NANDN U3236 ( .B(n2422), .A(n2423), .Z(n2419) );
  ANDN U3237 ( .A(n2309), .B(n2308), .Z(n2307) );
  NOR U3238 ( .A(n2424), .B(n2425), .Z(n2308) );
  NANDN U3239 ( .B(n2426), .A(n2427), .Z(n2309) );
  XNOR U3240 ( .A(n2431), .B(n2334), .Z(n2325) );
  XNOR U3241 ( .A(n2313), .B(n2433), .Z(n2314) );
  AND U3242 ( .A(n1390), .B(n1196), .Z(n2433) );
  XOR U3243 ( .A(n2437), .B(n2315), .Z(n2432) );
  NAND U3244 ( .A(n1138), .B(n1467), .Z(n2315) );
  IV U3245 ( .A(n2317), .Z(n2437) );
  XNOR U3246 ( .A(n2322), .B(n2323), .Z(n2319) );
  NANDN U3247 ( .B(n1020), .A(n1646), .Z(n2323) );
  XNOR U3248 ( .A(n2321), .B(n2441), .Z(n2322) );
  AND U3249 ( .A(n1554), .B(n1079), .Z(n2441) );
  XNOR U3250 ( .A(n2333), .B(n2324), .Z(n2431) );
  XOR U3251 ( .A(n2448), .B(n2343), .Z(n2333) );
  XNOR U3252 ( .A(n2330), .B(n2331), .Z(n2343) );
  NAND U3253 ( .A(n1284), .B(n1316), .Z(n2331) );
  XNOR U3254 ( .A(n2329), .B(n2449), .Z(n2330) );
  AND U3255 ( .A(n1246), .B(n1352), .Z(n2449) );
  XNOR U3256 ( .A(n2342), .B(n2332), .Z(n2448) );
  XNOR U3257 ( .A(n2337), .B(n2457), .Z(n2338) );
  AND U3258 ( .A(n1116), .B(n1522), .Z(n2457) );
  XOR U3259 ( .A(n2461), .B(n2339), .Z(n2456) );
  NAND U3260 ( .A(n1435), .B(n1178), .Z(n2339) );
  IV U3261 ( .A(n2341), .Z(n2461) );
  XNOR U3262 ( .A(n2465), .B(n2360), .Z(n2350) );
  XNOR U3263 ( .A(n2347), .B(n2348), .Z(n2360) );
  NANDN U3264 ( .B(n834), .A(n2036), .Z(n2348) );
  XNOR U3265 ( .A(n2346), .B(n2466), .Z(n2347) );
  AND U3266 ( .A(n1931), .B(n872), .Z(n2466) );
  XNOR U3267 ( .A(n2359), .B(n2349), .Z(n2465) );
  XNOR U3268 ( .A(n2354), .B(n2474), .Z(n2355) );
  AND U3269 ( .A(n1737), .B(n984), .Z(n2474) );
  XOR U3270 ( .A(n2478), .B(n2356), .Z(n2473) );
  NAND U3271 ( .A(n928), .B(n1831), .Z(n2356) );
  IV U3272 ( .A(n2358), .Z(n2478) );
  XNOR U3273 ( .A(n2363), .B(n2483), .Z(n2364) );
  AND U3274 ( .A(n2141), .B(n806), .Z(n2483) );
  XOR U3275 ( .A(n2487), .B(n2365), .Z(n2482) );
  NAND U3276 ( .A(n771), .B(n2254), .Z(n2365) );
  IV U3277 ( .A(n2367), .Z(n2487) );
  XNOR U3278 ( .A(n2374), .B(n2375), .Z(n2369) );
  NANDN U3279 ( .B(n716), .A(n2491), .Z(n2375) );
  XNOR U3280 ( .A(n2373), .B(n2492), .Z(n2374) );
  AND U3281 ( .A(n2370), .B(n746), .Z(n2492) );
  ANDN U3282 ( .A(n2493), .B(n2494), .Z(n2373) );
  NANDN U3283 ( .B(n2495), .A(n2496), .Z(n2493) );
  XNOR U3284 ( .A(n2500), .B(n2501), .Z(n663) );
  AND U3285 ( .A(n674), .B(n2503), .Z(n2502) );
  XOR U3286 ( .A(n2498), .B(n2501), .Z(n2503) );
  XNOR U3287 ( .A(n2497), .B(n2501), .Z(n2498) );
  XNOR U3288 ( .A(n2416), .B(n2415), .Z(n2501) );
  XNOR U3289 ( .A(n2504), .B(n2430), .Z(n2415) );
  XNOR U3290 ( .A(n2505), .B(n2400), .Z(n2390) );
  XNOR U3291 ( .A(n2387), .B(n2388), .Z(n2400) );
  NAND U3292 ( .A(n897), .B(n1952), .Z(n2388) );
  XNOR U3293 ( .A(n2386), .B(n2506), .Z(n2387) );
  AND U3294 ( .A(n2053), .B(n853), .Z(n2506) );
  XNOR U3295 ( .A(n2399), .B(n2389), .Z(n2505) );
  XNOR U3296 ( .A(n2394), .B(n2514), .Z(n2395) );
  AND U3297 ( .A(n2282), .B(n775), .Z(n2514) );
  XOR U3298 ( .A(n2518), .B(n2396), .Z(n2513) );
  NAND U3299 ( .A(n814), .B(n2166), .Z(n2396) );
  IV U3300 ( .A(n2398), .Z(n2518) );
  XNOR U3301 ( .A(n2403), .B(n2523), .Z(n2404) );
  AND U3302 ( .A(n1858), .B(n941), .Z(n2523) );
  XOR U3303 ( .A(n2527), .B(n2405), .Z(n2522) );
  NAND U3304 ( .A(n1001), .B(n1757), .Z(n2405) );
  IV U3305 ( .A(n2407), .Z(n2527) );
  XNOR U3306 ( .A(n2412), .B(n2413), .Z(n2409) );
  NAND U3307 ( .A(n1116), .B(n1574), .Z(n2413) );
  XNOR U3308 ( .A(n2411), .B(n2531), .Z(n2412) );
  AND U3309 ( .A(n1668), .B(n1055), .Z(n2531) );
  XNOR U3310 ( .A(n2429), .B(n2414), .Z(n2504) );
  XOR U3311 ( .A(n2538), .B(n2423), .Z(n2429) );
  XNOR U3312 ( .A(n2426), .B(n2427), .Z(n2423) );
  XOR U3313 ( .A(n2542), .B(n2425), .Z(n2426) );
  NAND U3314 ( .A(n744), .B(n2421), .Z(n2425) );
  NANDN U3315 ( .B(n717), .A(n2544), .Z(n2543) );
  OR U3316 ( .A(n2548), .B(n2549), .Z(n2422) );
  XNOR U3317 ( .A(n2553), .B(n2455), .Z(n2446) );
  XNOR U3318 ( .A(n2434), .B(n2555), .Z(n2435) );
  AND U3319 ( .A(n1467), .B(n1196), .Z(n2555) );
  XOR U3320 ( .A(n2559), .B(n2436), .Z(n2554) );
  NAND U3321 ( .A(n1138), .B(n1554), .Z(n2436) );
  IV U3322 ( .A(n2438), .Z(n2559) );
  XNOR U3323 ( .A(n2443), .B(n2444), .Z(n2440) );
  NANDN U3324 ( .B(n1020), .A(n1737), .Z(n2444) );
  XNOR U3325 ( .A(n2442), .B(n2563), .Z(n2443) );
  AND U3326 ( .A(n1646), .B(n1079), .Z(n2563) );
  XNOR U3327 ( .A(n2454), .B(n2445), .Z(n2553) );
  XOR U3328 ( .A(n2570), .B(n2464), .Z(n2454) );
  XNOR U3329 ( .A(n2451), .B(n2452), .Z(n2464) );
  NAND U3330 ( .A(n1284), .B(n1390), .Z(n2452) );
  XNOR U3331 ( .A(n2450), .B(n2571), .Z(n2451) );
  AND U3332 ( .A(n1316), .B(n1352), .Z(n2571) );
  XNOR U3333 ( .A(n2463), .B(n2453), .Z(n2570) );
  XNOR U3334 ( .A(n2458), .B(n2579), .Z(n2459) );
  AND U3335 ( .A(n1178), .B(n1522), .Z(n2579) );
  XOR U3336 ( .A(n2583), .B(n2460), .Z(n2578) );
  NAND U3337 ( .A(n1435), .B(n1246), .Z(n2460) );
  IV U3338 ( .A(n2462), .Z(n2583) );
  XNOR U3339 ( .A(n2587), .B(n2481), .Z(n2471) );
  XNOR U3340 ( .A(n2468), .B(n2469), .Z(n2481) );
  NANDN U3341 ( .B(n834), .A(n2141), .Z(n2469) );
  XNOR U3342 ( .A(n2467), .B(n2588), .Z(n2468) );
  AND U3343 ( .A(n2036), .B(n872), .Z(n2588) );
  XNOR U3344 ( .A(n2480), .B(n2470), .Z(n2587) );
  XNOR U3345 ( .A(n2475), .B(n2596), .Z(n2476) );
  AND U3346 ( .A(n1831), .B(n984), .Z(n2596) );
  XOR U3347 ( .A(n2600), .B(n2477), .Z(n2595) );
  NAND U3348 ( .A(n928), .B(n1931), .Z(n2477) );
  IV U3349 ( .A(n2479), .Z(n2600) );
  XNOR U3350 ( .A(n2484), .B(n2605), .Z(n2485) );
  AND U3351 ( .A(n2254), .B(n806), .Z(n2605) );
  XOR U3352 ( .A(n2609), .B(n2486), .Z(n2604) );
  NAND U3353 ( .A(n771), .B(n2370), .Z(n2486) );
  IV U3354 ( .A(n2488), .Z(n2609) );
  XOR U3355 ( .A(n2610), .B(n2611), .Z(n2488) );
  ANDN U3356 ( .A(n2612), .B(n2613), .Z(n2611) );
  XOR U3357 ( .A(n2610), .B(n2614), .Z(n2612) );
  XNOR U3358 ( .A(n2495), .B(n2496), .Z(n2490) );
  NANDN U3359 ( .B(n716), .A(n2615), .Z(n2496) );
  AND U3360 ( .A(n2491), .B(n746), .Z(n2616) );
  NAND U3361 ( .A(n2617), .B(n2618), .Z(n2494) );
  NANDN U3362 ( .B(n2619), .A(n2620), .Z(n2617) );
  XOR U3363 ( .A(n2624), .B(n2625), .Z(n664) );
  AND U3364 ( .A(n674), .B(n2627), .Z(n2626) );
  XNOR U3365 ( .A(n2622), .B(n2625), .Z(n2627) );
  XNOR U3366 ( .A(n2625), .B(n2621), .Z(n2622) );
  OR U3367 ( .A(n2628), .B(n2629), .Z(n2621) );
  XNOR U3368 ( .A(n2537), .B(n2536), .Z(n2625) );
  XNOR U3369 ( .A(n2630), .B(n2552), .Z(n2536) );
  XNOR U3370 ( .A(n2631), .B(n2521), .Z(n2511) );
  XNOR U3371 ( .A(n2508), .B(n2509), .Z(n2521) );
  NAND U3372 ( .A(n941), .B(n1952), .Z(n2509) );
  XNOR U3373 ( .A(n2507), .B(n2632), .Z(n2508) );
  AND U3374 ( .A(n2053), .B(n897), .Z(n2632) );
  XNOR U3375 ( .A(n2520), .B(n2510), .Z(n2631) );
  XNOR U3376 ( .A(n2515), .B(n2640), .Z(n2516) );
  AND U3377 ( .A(n2282), .B(n814), .Z(n2640) );
  XOR U3378 ( .A(n2644), .B(n2517), .Z(n2639) );
  NAND U3379 ( .A(n853), .B(n2166), .Z(n2517) );
  IV U3380 ( .A(n2519), .Z(n2644) );
  XNOR U3381 ( .A(n2524), .B(n2649), .Z(n2525) );
  AND U3382 ( .A(n1858), .B(n1001), .Z(n2649) );
  XOR U3383 ( .A(n2653), .B(n2526), .Z(n2648) );
  NAND U3384 ( .A(n1055), .B(n1757), .Z(n2526) );
  IV U3385 ( .A(n2528), .Z(n2653) );
  XNOR U3386 ( .A(n2533), .B(n2534), .Z(n2530) );
  NAND U3387 ( .A(n1178), .B(n1574), .Z(n2534) );
  XNOR U3388 ( .A(n2532), .B(n2657), .Z(n2533) );
  AND U3389 ( .A(n1668), .B(n1116), .Z(n2657) );
  XNOR U3390 ( .A(n2551), .B(n2535), .Z(n2630) );
  XNOR U3391 ( .A(n2664), .B(n2548), .Z(n2551) );
  XOR U3392 ( .A(n2541), .B(n2540), .Z(n2548) );
  XOR U3393 ( .A(n2539), .B(n2665), .Z(n2540) );
  AND U3394 ( .A(n2666), .B(n2667), .Z(n2665) );
  NANDN U3395 ( .B(n717), .A(n2668), .Z(n2667) );
  OR U3396 ( .A(n2669), .B(n2670), .Z(n2666) );
  NAND U3397 ( .A(n775), .B(n2421), .Z(n2547) );
  XNOR U3398 ( .A(n2545), .B(n2674), .Z(n2546) );
  AND U3399 ( .A(n2544), .B(n744), .Z(n2674) );
  NANDN U3400 ( .B(n2678), .A(n2679), .Z(n2549) );
  XNOR U3401 ( .A(n2683), .B(n2577), .Z(n2568) );
  XNOR U3402 ( .A(n2556), .B(n2685), .Z(n2557) );
  AND U3403 ( .A(n1554), .B(n1196), .Z(n2685) );
  XOR U3404 ( .A(n2689), .B(n2558), .Z(n2684) );
  NAND U3405 ( .A(n1138), .B(n1646), .Z(n2558) );
  IV U3406 ( .A(n2560), .Z(n2689) );
  XNOR U3407 ( .A(n2565), .B(n2566), .Z(n2562) );
  NANDN U3408 ( .B(n1020), .A(n1831), .Z(n2566) );
  XNOR U3409 ( .A(n2564), .B(n2693), .Z(n2565) );
  AND U3410 ( .A(n1737), .B(n1079), .Z(n2693) );
  XNOR U3411 ( .A(n2576), .B(n2567), .Z(n2683) );
  XOR U3412 ( .A(n2700), .B(n2586), .Z(n2576) );
  XNOR U3413 ( .A(n2573), .B(n2574), .Z(n2586) );
  NAND U3414 ( .A(n1284), .B(n1467), .Z(n2574) );
  XNOR U3415 ( .A(n2572), .B(n2701), .Z(n2573) );
  AND U3416 ( .A(n1390), .B(n1352), .Z(n2701) );
  XNOR U3417 ( .A(n2585), .B(n2575), .Z(n2700) );
  XNOR U3418 ( .A(n2580), .B(n2709), .Z(n2581) );
  AND U3419 ( .A(n1246), .B(n1522), .Z(n2709) );
  XOR U3420 ( .A(n2713), .B(n2582), .Z(n2708) );
  NAND U3421 ( .A(n1435), .B(n1316), .Z(n2582) );
  IV U3422 ( .A(n2584), .Z(n2713) );
  XNOR U3423 ( .A(n2717), .B(n2603), .Z(n2593) );
  XNOR U3424 ( .A(n2590), .B(n2591), .Z(n2603) );
  NANDN U3425 ( .B(n834), .A(n2254), .Z(n2591) );
  XNOR U3426 ( .A(n2589), .B(n2718), .Z(n2590) );
  AND U3427 ( .A(n2141), .B(n872), .Z(n2718) );
  XNOR U3428 ( .A(n2602), .B(n2592), .Z(n2717) );
  XNOR U3429 ( .A(n2597), .B(n2726), .Z(n2598) );
  AND U3430 ( .A(n1931), .B(n984), .Z(n2726) );
  XOR U3431 ( .A(n2730), .B(n2599), .Z(n2725) );
  NAND U3432 ( .A(n928), .B(n2036), .Z(n2599) );
  IV U3433 ( .A(n2601), .Z(n2730) );
  XNOR U3434 ( .A(n2606), .B(n2735), .Z(n2607) );
  AND U3435 ( .A(n2370), .B(n806), .Z(n2735) );
  XOR U3436 ( .A(n2739), .B(n2608), .Z(n2734) );
  NAND U3437 ( .A(n771), .B(n2491), .Z(n2608) );
  IV U3438 ( .A(n2610), .Z(n2739) );
  XNOR U3439 ( .A(n2619), .B(n2620), .Z(n2614) );
  NANDN U3440 ( .B(n716), .A(n2743), .Z(n2620) );
  XNOR U3441 ( .A(n2618), .B(n2744), .Z(n2619) );
  AND U3442 ( .A(n2615), .B(n746), .Z(n2744) );
  ANDN U3443 ( .A(n2745), .B(n2746), .Z(n2618) );
  NANDN U3444 ( .B(n2747), .A(n2748), .Z(n2745) );
  XNOR U3445 ( .A(n2750), .B(n2751), .Z(n702) );
  AND U3446 ( .A(n674), .B(n2753), .Z(n2752) );
  XOR U3447 ( .A(n2628), .B(n2754), .Z(n2753) );
  XOR U3448 ( .A(n2754), .B(n2629), .Z(n2628) );
  OR U3449 ( .A(n2755), .B(n2756), .Z(n2629) );
  IV U3450 ( .A(n2751), .Z(n2754) );
  XOR U3451 ( .A(n2663), .B(n2662), .Z(n2751) );
  XNOR U3452 ( .A(n2757), .B(n2682), .Z(n2662) );
  XNOR U3453 ( .A(n2758), .B(n2647), .Z(n2637) );
  XNOR U3454 ( .A(n2634), .B(n2635), .Z(n2647) );
  NAND U3455 ( .A(n1001), .B(n1952), .Z(n2635) );
  XNOR U3456 ( .A(n2633), .B(n2759), .Z(n2634) );
  AND U3457 ( .A(n2053), .B(n941), .Z(n2759) );
  XNOR U3458 ( .A(n2646), .B(n2636), .Z(n2758) );
  XNOR U3459 ( .A(n2641), .B(n2767), .Z(n2642) );
  AND U3460 ( .A(n2282), .B(n853), .Z(n2767) );
  XOR U3461 ( .A(n2771), .B(n2643), .Z(n2766) );
  NAND U3462 ( .A(n897), .B(n2166), .Z(n2643) );
  IV U3463 ( .A(n2645), .Z(n2771) );
  XNOR U3464 ( .A(n2650), .B(n2776), .Z(n2651) );
  AND U3465 ( .A(n1858), .B(n1055), .Z(n2776) );
  XOR U3466 ( .A(n2780), .B(n2652), .Z(n2775) );
  NAND U3467 ( .A(n1116), .B(n1757), .Z(n2652) );
  IV U3468 ( .A(n2654), .Z(n2780) );
  XNOR U3469 ( .A(n2659), .B(n2660), .Z(n2656) );
  NAND U3470 ( .A(n1246), .B(n1574), .Z(n2660) );
  XNOR U3471 ( .A(n2658), .B(n2784), .Z(n2659) );
  AND U3472 ( .A(n1668), .B(n1178), .Z(n2784) );
  XNOR U3473 ( .A(n2681), .B(n2661), .Z(n2757) );
  XNOR U3474 ( .A(n2791), .B(n2678), .Z(n2681) );
  XOR U3475 ( .A(n2673), .B(n2672), .Z(n2678) );
  XNOR U3476 ( .A(n2796), .B(n2669), .Z(n2792) );
  NAND U3477 ( .A(n744), .B(n2668), .Z(n2669) );
  NANDN U3478 ( .B(n717), .A(n2798), .Z(n2797) );
  NAND U3479 ( .A(n814), .B(n2421), .Z(n2677) );
  XNOR U3480 ( .A(n2675), .B(n2802), .Z(n2676) );
  AND U3481 ( .A(n2544), .B(n775), .Z(n2802) );
  XNOR U3482 ( .A(n2679), .B(n2680), .Z(n2791) );
  XNOR U3483 ( .A(n2812), .B(n2707), .Z(n2698) );
  XNOR U3484 ( .A(n2686), .B(n2814), .Z(n2687) );
  AND U3485 ( .A(n1646), .B(n1196), .Z(n2814) );
  XOR U3486 ( .A(n2818), .B(n2688), .Z(n2813) );
  NAND U3487 ( .A(n1138), .B(n1737), .Z(n2688) );
  IV U3488 ( .A(n2690), .Z(n2818) );
  XNOR U3489 ( .A(n2695), .B(n2696), .Z(n2692) );
  NANDN U3490 ( .B(n1020), .A(n1931), .Z(n2696) );
  XNOR U3491 ( .A(n2694), .B(n2822), .Z(n2695) );
  AND U3492 ( .A(n1831), .B(n1079), .Z(n2822) );
  XNOR U3493 ( .A(n2706), .B(n2697), .Z(n2812) );
  XOR U3494 ( .A(n2829), .B(n2716), .Z(n2706) );
  XNOR U3495 ( .A(n2703), .B(n2704), .Z(n2716) );
  NAND U3496 ( .A(n1284), .B(n1554), .Z(n2704) );
  XNOR U3497 ( .A(n2702), .B(n2830), .Z(n2703) );
  AND U3498 ( .A(n1467), .B(n1352), .Z(n2830) );
  XNOR U3499 ( .A(n2715), .B(n2705), .Z(n2829) );
  XNOR U3500 ( .A(n2710), .B(n2838), .Z(n2711) );
  AND U3501 ( .A(n1316), .B(n1522), .Z(n2838) );
  XOR U3502 ( .A(n2842), .B(n2712), .Z(n2837) );
  NAND U3503 ( .A(n1435), .B(n1390), .Z(n2712) );
  IV U3504 ( .A(n2714), .Z(n2842) );
  XNOR U3505 ( .A(n2846), .B(n2733), .Z(n2723) );
  XNOR U3506 ( .A(n2720), .B(n2721), .Z(n2733) );
  NANDN U3507 ( .B(n834), .A(n2370), .Z(n2721) );
  XNOR U3508 ( .A(n2719), .B(n2847), .Z(n2720) );
  AND U3509 ( .A(n2254), .B(n872), .Z(n2847) );
  XNOR U3510 ( .A(n2732), .B(n2722), .Z(n2846) );
  XNOR U3511 ( .A(n2727), .B(n2855), .Z(n2728) );
  AND U3512 ( .A(n2036), .B(n984), .Z(n2855) );
  XOR U3513 ( .A(n2859), .B(n2729), .Z(n2854) );
  NAND U3514 ( .A(n928), .B(n2141), .Z(n2729) );
  IV U3515 ( .A(n2731), .Z(n2859) );
  XNOR U3516 ( .A(n2736), .B(n2864), .Z(n2737) );
  AND U3517 ( .A(n2491), .B(n806), .Z(n2864) );
  XOR U3518 ( .A(n2868), .B(n2738), .Z(n2863) );
  NAND U3519 ( .A(n771), .B(n2615), .Z(n2738) );
  IV U3520 ( .A(n2740), .Z(n2868) );
  XNOR U3521 ( .A(n2747), .B(n2748), .Z(n2742) );
  OR U3522 ( .A(n2872), .B(n716), .Z(n2748) );
  AND U3523 ( .A(n2743), .B(n746), .Z(n2873) );
  NAND U3524 ( .A(n2874), .B(n2875), .Z(n2746) );
  NANDN U3525 ( .B(n2876), .A(n2877), .Z(n2874) );
  XNOR U3526 ( .A(n2879), .B(n2880), .Z(n1125) );
  XOR U3527 ( .A(n2878), .B(n2881), .Z(n2879) );
  AND U3528 ( .A(n674), .B(n2882), .Z(n2881) );
  XOR U3529 ( .A(n2755), .B(n2883), .Z(n2882) );
  XOR U3530 ( .A(n2883), .B(n2756), .Z(n2755) );
  NANDN U3531 ( .B(n2884), .A(n2885), .Z(n2756) );
  IV U3532 ( .A(n2880), .Z(n2883) );
  XOR U3533 ( .A(n2790), .B(n2789), .Z(n2880) );
  XNOR U3534 ( .A(n2886), .B(n2808), .Z(n2789) );
  XNOR U3535 ( .A(n2887), .B(n2774), .Z(n2764) );
  XNOR U3536 ( .A(n2761), .B(n2762), .Z(n2774) );
  NAND U3537 ( .A(n1055), .B(n1952), .Z(n2762) );
  XNOR U3538 ( .A(n2760), .B(n2888), .Z(n2761) );
  AND U3539 ( .A(n2053), .B(n1001), .Z(n2888) );
  XNOR U3540 ( .A(n2773), .B(n2763), .Z(n2887) );
  XNOR U3541 ( .A(n2768), .B(n2896), .Z(n2769) );
  AND U3542 ( .A(n2282), .B(n897), .Z(n2896) );
  XOR U3543 ( .A(n2900), .B(n2770), .Z(n2895) );
  NAND U3544 ( .A(n941), .B(n2166), .Z(n2770) );
  IV U3545 ( .A(n2772), .Z(n2900) );
  XNOR U3546 ( .A(n2777), .B(n2905), .Z(n2778) );
  AND U3547 ( .A(n1858), .B(n1116), .Z(n2905) );
  XOR U3548 ( .A(n2909), .B(n2779), .Z(n2904) );
  NAND U3549 ( .A(n1178), .B(n1757), .Z(n2779) );
  IV U3550 ( .A(n2781), .Z(n2909) );
  XNOR U3551 ( .A(n2786), .B(n2787), .Z(n2783) );
  NAND U3552 ( .A(n1316), .B(n1574), .Z(n2787) );
  XNOR U3553 ( .A(n2785), .B(n2913), .Z(n2786) );
  AND U3554 ( .A(n1668), .B(n1246), .Z(n2913) );
  XNOR U3555 ( .A(n2807), .B(n2788), .Z(n2886) );
  XOR U3556 ( .A(n2920), .B(n2811), .Z(n2807) );
  XNOR U3557 ( .A(n2799), .B(n2922), .Z(n2800) );
  AND U3558 ( .A(n2798), .B(n744), .Z(n2922) );
  XOR U3559 ( .A(n2926), .B(n2801), .Z(n2921) );
  NAND U3560 ( .A(n775), .B(n2668), .Z(n2801) );
  IV U3561 ( .A(n2793), .Z(n2926) );
  XNOR U3562 ( .A(n2804), .B(n2805), .Z(n2795) );
  NAND U3563 ( .A(n853), .B(n2421), .Z(n2805) );
  XNOR U3564 ( .A(n2803), .B(n2930), .Z(n2804) );
  AND U3565 ( .A(n2544), .B(n814), .Z(n2930) );
  XNOR U3566 ( .A(n2810), .B(n2806), .Z(n2920) );
  AND U3567 ( .A(n2938), .B(n2939), .Z(n2937) );
  OR U3568 ( .A(n2940), .B(n2941), .Z(n2939) );
  AND U3569 ( .A(n2942), .B(n2943), .Z(n2938) );
  NANDN U3570 ( .B(n717), .A(n2944), .Z(n2943) );
  NANDN U3571 ( .B(n2945), .A(n2946), .Z(n2942) );
  XNOR U3572 ( .A(n2950), .B(n2836), .Z(n2827) );
  XNOR U3573 ( .A(n2815), .B(n2952), .Z(n2816) );
  AND U3574 ( .A(n1737), .B(n1196), .Z(n2952) );
  XOR U3575 ( .A(n2956), .B(n2817), .Z(n2951) );
  NAND U3576 ( .A(n1138), .B(n1831), .Z(n2817) );
  IV U3577 ( .A(n2819), .Z(n2956) );
  XNOR U3578 ( .A(n2824), .B(n2825), .Z(n2821) );
  NANDN U3579 ( .B(n1020), .A(n2036), .Z(n2825) );
  XNOR U3580 ( .A(n2823), .B(n2960), .Z(n2824) );
  AND U3581 ( .A(n1931), .B(n1079), .Z(n2960) );
  XNOR U3582 ( .A(n2835), .B(n2826), .Z(n2950) );
  XOR U3583 ( .A(n2967), .B(n2845), .Z(n2835) );
  XNOR U3584 ( .A(n2832), .B(n2833), .Z(n2845) );
  NAND U3585 ( .A(n1284), .B(n1646), .Z(n2833) );
  XNOR U3586 ( .A(n2831), .B(n2968), .Z(n2832) );
  AND U3587 ( .A(n1554), .B(n1352), .Z(n2968) );
  XNOR U3588 ( .A(n2844), .B(n2834), .Z(n2967) );
  XNOR U3589 ( .A(n2839), .B(n2976), .Z(n2840) );
  AND U3590 ( .A(n1390), .B(n1522), .Z(n2976) );
  XOR U3591 ( .A(n2980), .B(n2841), .Z(n2975) );
  NAND U3592 ( .A(n1435), .B(n1467), .Z(n2841) );
  IV U3593 ( .A(n2843), .Z(n2980) );
  XNOR U3594 ( .A(n2984), .B(n2862), .Z(n2852) );
  XNOR U3595 ( .A(n2849), .B(n2850), .Z(n2862) );
  NANDN U3596 ( .B(n834), .A(n2491), .Z(n2850) );
  XNOR U3597 ( .A(n2848), .B(n2985), .Z(n2849) );
  AND U3598 ( .A(n2370), .B(n872), .Z(n2985) );
  XNOR U3599 ( .A(n2861), .B(n2851), .Z(n2984) );
  XNOR U3600 ( .A(n2856), .B(n2993), .Z(n2857) );
  AND U3601 ( .A(n2141), .B(n984), .Z(n2993) );
  XOR U3602 ( .A(n2997), .B(n2858), .Z(n2992) );
  NAND U3603 ( .A(n928), .B(n2254), .Z(n2858) );
  IV U3604 ( .A(n2860), .Z(n2997) );
  XNOR U3605 ( .A(n2865), .B(n3002), .Z(n2866) );
  AND U3606 ( .A(n2615), .B(n806), .Z(n3002) );
  XOR U3607 ( .A(n3006), .B(n2867), .Z(n3001) );
  NAND U3608 ( .A(n771), .B(n2743), .Z(n2867) );
  IV U3609 ( .A(n2869), .Z(n3006) );
  XNOR U3610 ( .A(n2876), .B(n2877), .Z(n2871) );
  OR U3611 ( .A(n3010), .B(n716), .Z(n2877) );
  XNOR U3612 ( .A(n2875), .B(n3011), .Z(n2876) );
  ANDN U3613 ( .A(n746), .B(n2872), .Z(n3011) );
  ANDN U3614 ( .A(n3012), .B(n3013), .Z(n2875) );
  NANDN U3615 ( .B(n3014), .A(n3015), .Z(n3012) );
  XOR U3616 ( .A(n3017), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U3617 ( .A(n3018), .B(n3019), .Z(n3017) );
  XNOR U3618 ( .A(n3020), .B(n3016), .Z(n3018) );
  NANDN U3619 ( .B(n2885), .A(\_MxM/Y0[0] ), .Z(n3016) );
  NAND U3620 ( .A(n3021), .B(n674), .Z(n3020) );
  XOR U3621 ( .A(e_input[31]), .B(g_input[31]), .Z(n674) );
  XNOR U3622 ( .A(n2884), .B(n3019), .Z(n3021) );
  XOR U3623 ( .A(n2885), .B(n3019), .Z(n2884) );
  XOR U3624 ( .A(n2919), .B(n2918), .Z(n3019) );
  XNOR U3625 ( .A(n3022), .B(n2936), .Z(n2918) );
  XNOR U3626 ( .A(n3023), .B(n2903), .Z(n2893) );
  XNOR U3627 ( .A(n2890), .B(n2891), .Z(n2903) );
  NAND U3628 ( .A(n1116), .B(n1952), .Z(n2891) );
  XNOR U3629 ( .A(n2889), .B(n3024), .Z(n2890) );
  AND U3630 ( .A(n2053), .B(n1055), .Z(n3024) );
  XNOR U3631 ( .A(n2902), .B(n2892), .Z(n3023) );
  XNOR U3632 ( .A(n2897), .B(n3032), .Z(n2898) );
  AND U3633 ( .A(n2282), .B(n941), .Z(n3032) );
  XOR U3634 ( .A(n3036), .B(n2899), .Z(n3031) );
  NAND U3635 ( .A(n1001), .B(n2166), .Z(n2899) );
  IV U3636 ( .A(n2901), .Z(n3036) );
  XNOR U3637 ( .A(n2906), .B(n3041), .Z(n2907) );
  AND U3638 ( .A(n1858), .B(n1178), .Z(n3041) );
  XOR U3639 ( .A(n3045), .B(n2908), .Z(n3040) );
  NAND U3640 ( .A(n1246), .B(n1757), .Z(n2908) );
  IV U3641 ( .A(n2910), .Z(n3045) );
  XNOR U3642 ( .A(n2915), .B(n2916), .Z(n2912) );
  NAND U3643 ( .A(n1390), .B(n1574), .Z(n2916) );
  XNOR U3644 ( .A(n2914), .B(n3049), .Z(n2915) );
  AND U3645 ( .A(n1668), .B(n1316), .Z(n3049) );
  XNOR U3646 ( .A(n2935), .B(n2917), .Z(n3022) );
  XOR U3647 ( .A(n3056), .B(n2949), .Z(n2935) );
  XNOR U3648 ( .A(n2923), .B(n3058), .Z(n2924) );
  AND U3649 ( .A(n2798), .B(n775), .Z(n3058) );
  XOR U3650 ( .A(n3062), .B(n2925), .Z(n3057) );
  NAND U3651 ( .A(n814), .B(n2668), .Z(n2925) );
  IV U3652 ( .A(n2927), .Z(n3062) );
  XNOR U3653 ( .A(n2932), .B(n2933), .Z(n2929) );
  NAND U3654 ( .A(n897), .B(n2421), .Z(n2933) );
  XNOR U3655 ( .A(n2931), .B(n3066), .Z(n2932) );
  AND U3656 ( .A(n2544), .B(n853), .Z(n3066) );
  XNOR U3657 ( .A(n2948), .B(n2934), .Z(n3056) );
  XNOR U3658 ( .A(n3073), .B(n2945), .Z(n2948) );
  XOR U3659 ( .A(n3074), .B(n2940), .Z(n2945) );
  NAND U3660 ( .A(n744), .B(n2944), .Z(n2940) );
  NANDN U3661 ( .B(n717), .A(n3076), .Z(n3075) );
  XNOR U3662 ( .A(n2946), .B(n2947), .Z(n3073) );
  XNOR U3663 ( .A(n3086), .B(n2974), .Z(n2965) );
  XNOR U3664 ( .A(n2953), .B(n3088), .Z(n2954) );
  AND U3665 ( .A(n1831), .B(n1196), .Z(n3088) );
  XOR U3666 ( .A(n3092), .B(n2955), .Z(n3087) );
  NAND U3667 ( .A(n1138), .B(n1931), .Z(n2955) );
  IV U3668 ( .A(n2957), .Z(n3092) );
  XNOR U3669 ( .A(n2962), .B(n2963), .Z(n2959) );
  NANDN U3670 ( .B(n1020), .A(n2141), .Z(n2963) );
  XNOR U3671 ( .A(n2961), .B(n3096), .Z(n2962) );
  AND U3672 ( .A(n2036), .B(n1079), .Z(n3096) );
  XNOR U3673 ( .A(n2973), .B(n2964), .Z(n3086) );
  XOR U3674 ( .A(n3103), .B(n2983), .Z(n2973) );
  XNOR U3675 ( .A(n2970), .B(n2971), .Z(n2983) );
  NAND U3676 ( .A(n1284), .B(n1737), .Z(n2971) );
  XNOR U3677 ( .A(n2969), .B(n3104), .Z(n2970) );
  AND U3678 ( .A(n1646), .B(n1352), .Z(n3104) );
  XNOR U3679 ( .A(n2982), .B(n2972), .Z(n3103) );
  XNOR U3680 ( .A(n2977), .B(n3112), .Z(n2978) );
  AND U3681 ( .A(n1467), .B(n1522), .Z(n3112) );
  XOR U3682 ( .A(n3116), .B(n2979), .Z(n3111) );
  NAND U3683 ( .A(n1435), .B(n1554), .Z(n2979) );
  IV U3684 ( .A(n2981), .Z(n3116) );
  XNOR U3685 ( .A(n3120), .B(n3000), .Z(n2990) );
  XNOR U3686 ( .A(n2987), .B(n2988), .Z(n3000) );
  NANDN U3687 ( .B(n834), .A(n2615), .Z(n2988) );
  XNOR U3688 ( .A(n2986), .B(n3121), .Z(n2987) );
  AND U3689 ( .A(n2491), .B(n872), .Z(n3121) );
  XNOR U3690 ( .A(n2999), .B(n2989), .Z(n3120) );
  XNOR U3691 ( .A(n2994), .B(n3129), .Z(n2995) );
  AND U3692 ( .A(n2254), .B(n984), .Z(n3129) );
  XOR U3693 ( .A(n3133), .B(n2996), .Z(n3128) );
  NAND U3694 ( .A(n928), .B(n2370), .Z(n2996) );
  IV U3695 ( .A(n2998), .Z(n3133) );
  XNOR U3696 ( .A(n3003), .B(n3138), .Z(n3004) );
  AND U3697 ( .A(n2743), .B(n806), .Z(n3138) );
  XOR U3698 ( .A(n3142), .B(n3005), .Z(n3137) );
  NANDN U3699 ( .B(n2872), .A(n771), .Z(n3005) );
  IV U3700 ( .A(n3007), .Z(n3142) );
  XNOR U3701 ( .A(n3014), .B(n3015), .Z(n3009) );
  NANDN U3702 ( .B(n716), .A(n3146), .Z(n3015) );
  ANDN U3703 ( .A(n746), .B(n3010), .Z(n3147) );
  NAND U3704 ( .A(n3148), .B(n3149), .Z(n3013) );
  NANDN U3705 ( .B(n3150), .A(n3151), .Z(n3148) );
  XOR U3706 ( .A(n3055), .B(n3054), .Z(n2885) );
  XNOR U3707 ( .A(n3152), .B(n3072), .Z(n3054) );
  XNOR U3708 ( .A(n3153), .B(n3039), .Z(n3029) );
  XNOR U3709 ( .A(n3026), .B(n3027), .Z(n3039) );
  NAND U3710 ( .A(n1178), .B(n1952), .Z(n3027) );
  XNOR U3711 ( .A(n3025), .B(n3154), .Z(n3026) );
  AND U3712 ( .A(n2053), .B(n1116), .Z(n3154) );
  XNOR U3713 ( .A(n3038), .B(n3028), .Z(n3153) );
  XNOR U3714 ( .A(n3033), .B(n3162), .Z(n3034) );
  AND U3715 ( .A(n2282), .B(n1001), .Z(n3162) );
  XOR U3716 ( .A(n3166), .B(n3035), .Z(n3161) );
  NAND U3717 ( .A(n1055), .B(n2166), .Z(n3035) );
  IV U3718 ( .A(n3037), .Z(n3166) );
  XNOR U3719 ( .A(n3042), .B(n3171), .Z(n3043) );
  AND U3720 ( .A(n1858), .B(n1246), .Z(n3171) );
  XOR U3721 ( .A(n3175), .B(n3044), .Z(n3170) );
  NAND U3722 ( .A(n1316), .B(n1757), .Z(n3044) );
  IV U3723 ( .A(n3046), .Z(n3175) );
  XNOR U3724 ( .A(n3051), .B(n3052), .Z(n3048) );
  NAND U3725 ( .A(n1467), .B(n1574), .Z(n3052) );
  XNOR U3726 ( .A(n3050), .B(n3179), .Z(n3051) );
  AND U3727 ( .A(n1668), .B(n1390), .Z(n3179) );
  XNOR U3728 ( .A(n3071), .B(n3053), .Z(n3152) );
  XOR U3729 ( .A(n3183), .B(n3184), .Z(n3053) );
  XOR U3730 ( .A(n3185), .B(n3082), .Z(n3071) );
  XNOR U3731 ( .A(n3059), .B(n3187), .Z(n3060) );
  AND U3732 ( .A(n2798), .B(n814), .Z(n3187) );
  XOR U3733 ( .A(n3191), .B(n3061), .Z(n3186) );
  NAND U3734 ( .A(n853), .B(n2668), .Z(n3061) );
  IV U3735 ( .A(n3063), .Z(n3191) );
  XNOR U3736 ( .A(n3068), .B(n3069), .Z(n3065) );
  NAND U3737 ( .A(n941), .B(n2421), .Z(n3069) );
  XNOR U3738 ( .A(n3067), .B(n3195), .Z(n3068) );
  AND U3739 ( .A(n2544), .B(n897), .Z(n3195) );
  XNOR U3740 ( .A(n3081), .B(n3070), .Z(n3185) );
  XOR U3741 ( .A(n3199), .B(n3200), .Z(n3070) );
  AND U3742 ( .A(n3201), .B(n3202), .Z(n3200) );
  XNOR U3743 ( .A(n3203), .B(n3204), .Z(n3202) );
  XOR U3744 ( .A(n3205), .B(n3199), .Z(n3203) );
  XOR U3745 ( .A(n3159), .B(n3206), .Z(n3201) );
  XNOR U3746 ( .A(n3199), .B(n3160), .Z(n3206) );
  XNOR U3747 ( .A(n3172), .B(n3208), .Z(n3173) );
  AND U3748 ( .A(n1858), .B(n1316), .Z(n3208) );
  XOR U3749 ( .A(n3212), .B(n3174), .Z(n3207) );
  NAND U3750 ( .A(n1390), .B(n1757), .Z(n3174) );
  IV U3751 ( .A(n3176), .Z(n3212) );
  XNOR U3752 ( .A(n3181), .B(n3182), .Z(n3178) );
  NAND U3753 ( .A(n1574), .B(n1554), .Z(n3182) );
  XNOR U3754 ( .A(n3180), .B(n3216), .Z(n3181) );
  AND U3755 ( .A(n1668), .B(n1467), .Z(n3216) );
  XOR U3756 ( .A(n3220), .B(n3169), .Z(n3159) );
  XNOR U3757 ( .A(n3156), .B(n3157), .Z(n3169) );
  NAND U3758 ( .A(n1246), .B(n1952), .Z(n3157) );
  XNOR U3759 ( .A(n3155), .B(n3221), .Z(n3156) );
  AND U3760 ( .A(n2053), .B(n1178), .Z(n3221) );
  XNOR U3761 ( .A(n3168), .B(n3158), .Z(n3220) );
  XNOR U3762 ( .A(n3163), .B(n3229), .Z(n3164) );
  AND U3763 ( .A(n2282), .B(n1055), .Z(n3229) );
  XOR U3764 ( .A(n3233), .B(n3165), .Z(n3228) );
  NAND U3765 ( .A(n1116), .B(n2166), .Z(n3165) );
  IV U3766 ( .A(n3167), .Z(n3233) );
  XOR U3767 ( .A(n3237), .B(n3238), .Z(n3199) );
  AND U3768 ( .A(n3239), .B(n3240), .Z(n3238) );
  XNOR U3769 ( .A(n3241), .B(n3242), .Z(n3240) );
  XNOR U3770 ( .A(n3237), .B(n3243), .Z(n3242) );
  XOR U3771 ( .A(n3226), .B(n3244), .Z(n3239) );
  XNOR U3772 ( .A(n3237), .B(n3227), .Z(n3244) );
  XNOR U3773 ( .A(n3209), .B(n3246), .Z(n3210) );
  AND U3774 ( .A(n1858), .B(n1390), .Z(n3246) );
  XOR U3775 ( .A(n3250), .B(n3211), .Z(n3245) );
  NAND U3776 ( .A(n1467), .B(n1757), .Z(n3211) );
  IV U3777 ( .A(n3213), .Z(n3250) );
  XNOR U3778 ( .A(n3218), .B(n3219), .Z(n3215) );
  NAND U3779 ( .A(n1574), .B(n1646), .Z(n3219) );
  XNOR U3780 ( .A(n3217), .B(n3254), .Z(n3218) );
  AND U3781 ( .A(n1554), .B(n1668), .Z(n3254) );
  XOR U3782 ( .A(n3258), .B(n3236), .Z(n3226) );
  XNOR U3783 ( .A(n3223), .B(n3224), .Z(n3236) );
  NAND U3784 ( .A(n1316), .B(n1952), .Z(n3224) );
  XNOR U3785 ( .A(n3222), .B(n3259), .Z(n3223) );
  AND U3786 ( .A(n2053), .B(n1246), .Z(n3259) );
  XNOR U3787 ( .A(n3235), .B(n3225), .Z(n3258) );
  XNOR U3788 ( .A(n3230), .B(n3267), .Z(n3231) );
  AND U3789 ( .A(n2282), .B(n1116), .Z(n3267) );
  XOR U3790 ( .A(n3271), .B(n3232), .Z(n3266) );
  NAND U3791 ( .A(n1178), .B(n2166), .Z(n3232) );
  IV U3792 ( .A(n3234), .Z(n3271) );
  XOR U3793 ( .A(n3275), .B(n3276), .Z(n3237) );
  AND U3794 ( .A(n3277), .B(n3278), .Z(n3276) );
  XNOR U3795 ( .A(n3279), .B(n3280), .Z(n3278) );
  XNOR U3796 ( .A(n3275), .B(n3281), .Z(n3280) );
  XOR U3797 ( .A(n3264), .B(n3282), .Z(n3277) );
  XNOR U3798 ( .A(n3275), .B(n3265), .Z(n3282) );
  XNOR U3799 ( .A(n3247), .B(n3284), .Z(n3248) );
  AND U3800 ( .A(n1858), .B(n1467), .Z(n3284) );
  XOR U3801 ( .A(n3288), .B(n3249), .Z(n3283) );
  NAND U3802 ( .A(n1757), .B(n1554), .Z(n3249) );
  IV U3803 ( .A(n3251), .Z(n3288) );
  XNOR U3804 ( .A(n3256), .B(n3257), .Z(n3253) );
  NAND U3805 ( .A(n1574), .B(n1737), .Z(n3257) );
  XNOR U3806 ( .A(n3255), .B(n3292), .Z(n3256) );
  AND U3807 ( .A(n1646), .B(n1668), .Z(n3292) );
  XOR U3808 ( .A(n3296), .B(n3274), .Z(n3264) );
  XNOR U3809 ( .A(n3261), .B(n3262), .Z(n3274) );
  NAND U3810 ( .A(n1390), .B(n1952), .Z(n3262) );
  XNOR U3811 ( .A(n3260), .B(n3297), .Z(n3261) );
  AND U3812 ( .A(n2053), .B(n1316), .Z(n3297) );
  XNOR U3813 ( .A(n3273), .B(n3263), .Z(n3296) );
  XNOR U3814 ( .A(n3268), .B(n3305), .Z(n3269) );
  AND U3815 ( .A(n2282), .B(n1178), .Z(n3305) );
  XOR U3816 ( .A(n3309), .B(n3270), .Z(n3304) );
  NAND U3817 ( .A(n1246), .B(n2166), .Z(n3270) );
  IV U3818 ( .A(n3272), .Z(n3309) );
  XOR U3819 ( .A(n3313), .B(n3314), .Z(n3275) );
  AND U3820 ( .A(n3315), .B(n3316), .Z(n3314) );
  XNOR U3821 ( .A(n3317), .B(n3318), .Z(n3316) );
  XNOR U3822 ( .A(n3313), .B(n3319), .Z(n3318) );
  XOR U3823 ( .A(n3302), .B(n3320), .Z(n3315) );
  XNOR U3824 ( .A(n3313), .B(n3303), .Z(n3320) );
  XNOR U3825 ( .A(n3285), .B(n3322), .Z(n3286) );
  AND U3826 ( .A(n1554), .B(n1858), .Z(n3322) );
  XOR U3827 ( .A(n3326), .B(n3287), .Z(n3321) );
  NAND U3828 ( .A(n1757), .B(n1646), .Z(n3287) );
  IV U3829 ( .A(n3289), .Z(n3326) );
  XNOR U3830 ( .A(n3294), .B(n3295), .Z(n3291) );
  NAND U3831 ( .A(n1574), .B(n1831), .Z(n3295) );
  XNOR U3832 ( .A(n3293), .B(n3330), .Z(n3294) );
  AND U3833 ( .A(n1737), .B(n1668), .Z(n3330) );
  XOR U3834 ( .A(n3334), .B(n3312), .Z(n3302) );
  XNOR U3835 ( .A(n3299), .B(n3300), .Z(n3312) );
  NAND U3836 ( .A(n1467), .B(n1952), .Z(n3300) );
  XNOR U3837 ( .A(n3298), .B(n3335), .Z(n3299) );
  AND U3838 ( .A(n2053), .B(n1390), .Z(n3335) );
  XNOR U3839 ( .A(n3311), .B(n3301), .Z(n3334) );
  XNOR U3840 ( .A(n3306), .B(n3343), .Z(n3307) );
  AND U3841 ( .A(n2282), .B(n1246), .Z(n3343) );
  XOR U3842 ( .A(n3347), .B(n3308), .Z(n3342) );
  NAND U3843 ( .A(n1316), .B(n2166), .Z(n3308) );
  IV U3844 ( .A(n3310), .Z(n3347) );
  XOR U3845 ( .A(n3351), .B(n3352), .Z(n3313) );
  AND U3846 ( .A(n3353), .B(n3354), .Z(n3352) );
  XNOR U3847 ( .A(n3355), .B(n3356), .Z(n3354) );
  XNOR U3848 ( .A(n3351), .B(n3357), .Z(n3356) );
  XOR U3849 ( .A(n3340), .B(n3358), .Z(n3353) );
  XNOR U3850 ( .A(n3351), .B(n3341), .Z(n3358) );
  XNOR U3851 ( .A(n3323), .B(n3360), .Z(n3324) );
  AND U3852 ( .A(n1646), .B(n1858), .Z(n3360) );
  XOR U3853 ( .A(n3364), .B(n3325), .Z(n3359) );
  NAND U3854 ( .A(n1757), .B(n1737), .Z(n3325) );
  IV U3855 ( .A(n3327), .Z(n3364) );
  XNOR U3856 ( .A(n3332), .B(n3333), .Z(n3329) );
  NAND U3857 ( .A(n1574), .B(n1931), .Z(n3333) );
  XNOR U3858 ( .A(n3331), .B(n3368), .Z(n3332) );
  AND U3859 ( .A(n1831), .B(n1668), .Z(n3368) );
  XOR U3860 ( .A(n3372), .B(n3350), .Z(n3340) );
  XNOR U3861 ( .A(n3337), .B(n3338), .Z(n3350) );
  NAND U3862 ( .A(n1952), .B(n1554), .Z(n3338) );
  XNOR U3863 ( .A(n3336), .B(n3373), .Z(n3337) );
  AND U3864 ( .A(n2053), .B(n1467), .Z(n3373) );
  XNOR U3865 ( .A(n3349), .B(n3339), .Z(n3372) );
  XNOR U3866 ( .A(n3344), .B(n3381), .Z(n3345) );
  AND U3867 ( .A(n2282), .B(n1316), .Z(n3381) );
  XOR U3868 ( .A(n3385), .B(n3346), .Z(n3380) );
  NAND U3869 ( .A(n1390), .B(n2166), .Z(n3346) );
  IV U3870 ( .A(n3348), .Z(n3385) );
  XOR U3871 ( .A(n3389), .B(n3390), .Z(n3351) );
  AND U3872 ( .A(n3391), .B(n3392), .Z(n3390) );
  XNOR U3873 ( .A(n3393), .B(n3394), .Z(n3392) );
  XNOR U3874 ( .A(n3389), .B(n3395), .Z(n3394) );
  XOR U3875 ( .A(n3378), .B(n3396), .Z(n3391) );
  XNOR U3876 ( .A(n3389), .B(n3379), .Z(n3396) );
  XNOR U3877 ( .A(n3361), .B(n3398), .Z(n3362) );
  AND U3878 ( .A(n1737), .B(n1858), .Z(n3398) );
  XOR U3879 ( .A(n3402), .B(n3363), .Z(n3397) );
  NAND U3880 ( .A(n1757), .B(n1831), .Z(n3363) );
  IV U3881 ( .A(n3365), .Z(n3402) );
  XNOR U3882 ( .A(n3370), .B(n3371), .Z(n3367) );
  NAND U3883 ( .A(n1574), .B(n2036), .Z(n3371) );
  XNOR U3884 ( .A(n3369), .B(n3406), .Z(n3370) );
  AND U3885 ( .A(n1931), .B(n1668), .Z(n3406) );
  XOR U3886 ( .A(n3410), .B(n3388), .Z(n3378) );
  XNOR U3887 ( .A(n3375), .B(n3376), .Z(n3388) );
  NAND U3888 ( .A(n1952), .B(n1646), .Z(n3376) );
  XNOR U3889 ( .A(n3374), .B(n3411), .Z(n3375) );
  AND U3890 ( .A(n1554), .B(n2053), .Z(n3411) );
  XNOR U3891 ( .A(n3387), .B(n3377), .Z(n3410) );
  XNOR U3892 ( .A(n3382), .B(n3419), .Z(n3383) );
  AND U3893 ( .A(n2282), .B(n1390), .Z(n3419) );
  XOR U3894 ( .A(n3423), .B(n3384), .Z(n3418) );
  NAND U3895 ( .A(n1467), .B(n2166), .Z(n3384) );
  IV U3896 ( .A(n3386), .Z(n3423) );
  XOR U3897 ( .A(n3427), .B(n3428), .Z(n3389) );
  AND U3898 ( .A(n3429), .B(n3430), .Z(n3428) );
  XNOR U3899 ( .A(n3431), .B(n3432), .Z(n3430) );
  XNOR U3900 ( .A(n3427), .B(n3433), .Z(n3432) );
  XOR U3901 ( .A(n3416), .B(n3434), .Z(n3429) );
  XNOR U3902 ( .A(n3427), .B(n3417), .Z(n3434) );
  XNOR U3903 ( .A(n3399), .B(n3436), .Z(n3400) );
  AND U3904 ( .A(n1831), .B(n1858), .Z(n3436) );
  XOR U3905 ( .A(n3440), .B(n3401), .Z(n3435) );
  NAND U3906 ( .A(n1757), .B(n1931), .Z(n3401) );
  IV U3907 ( .A(n3403), .Z(n3440) );
  XNOR U3908 ( .A(n3408), .B(n3409), .Z(n3405) );
  NAND U3909 ( .A(n1574), .B(n2141), .Z(n3409) );
  XNOR U3910 ( .A(n3407), .B(n3444), .Z(n3408) );
  AND U3911 ( .A(n2036), .B(n1668), .Z(n3444) );
  XOR U3912 ( .A(n3448), .B(n3426), .Z(n3416) );
  XNOR U3913 ( .A(n3413), .B(n3414), .Z(n3426) );
  NAND U3914 ( .A(n1952), .B(n1737), .Z(n3414) );
  XNOR U3915 ( .A(n3412), .B(n3449), .Z(n3413) );
  AND U3916 ( .A(n1646), .B(n2053), .Z(n3449) );
  XNOR U3917 ( .A(n3425), .B(n3415), .Z(n3448) );
  XNOR U3918 ( .A(n3420), .B(n3457), .Z(n3421) );
  AND U3919 ( .A(n2282), .B(n1467), .Z(n3457) );
  XOR U3920 ( .A(n3461), .B(n3422), .Z(n3456) );
  NAND U3921 ( .A(n2166), .B(n1554), .Z(n3422) );
  IV U3922 ( .A(n3424), .Z(n3461) );
  XOR U3923 ( .A(n3465), .B(n3466), .Z(n3427) );
  AND U3924 ( .A(n3467), .B(n3468), .Z(n3466) );
  XNOR U3925 ( .A(n3469), .B(n3470), .Z(n3468) );
  XNOR U3926 ( .A(n3465), .B(n3471), .Z(n3470) );
  XOR U3927 ( .A(n3454), .B(n3472), .Z(n3467) );
  XNOR U3928 ( .A(n3465), .B(n3455), .Z(n3472) );
  XNOR U3929 ( .A(n3437), .B(n3474), .Z(n3438) );
  AND U3930 ( .A(n1931), .B(n1858), .Z(n3474) );
  XOR U3931 ( .A(n3478), .B(n3439), .Z(n3473) );
  NAND U3932 ( .A(n1757), .B(n2036), .Z(n3439) );
  IV U3933 ( .A(n3441), .Z(n3478) );
  XNOR U3934 ( .A(n3446), .B(n3447), .Z(n3443) );
  NAND U3935 ( .A(n1574), .B(n2254), .Z(n3447) );
  XNOR U3936 ( .A(n3445), .B(n3482), .Z(n3446) );
  AND U3937 ( .A(n2141), .B(n1668), .Z(n3482) );
  XOR U3938 ( .A(n3486), .B(n3464), .Z(n3454) );
  XNOR U3939 ( .A(n3451), .B(n3452), .Z(n3464) );
  NAND U3940 ( .A(n1952), .B(n1831), .Z(n3452) );
  XNOR U3941 ( .A(n3450), .B(n3487), .Z(n3451) );
  AND U3942 ( .A(n1737), .B(n2053), .Z(n3487) );
  XNOR U3943 ( .A(n3463), .B(n3453), .Z(n3486) );
  XNOR U3944 ( .A(n3458), .B(n3495), .Z(n3459) );
  AND U3945 ( .A(n1554), .B(n2282), .Z(n3495) );
  XOR U3946 ( .A(n3499), .B(n3460), .Z(n3494) );
  NAND U3947 ( .A(n2166), .B(n1646), .Z(n3460) );
  IV U3948 ( .A(n3462), .Z(n3499) );
  XOR U3949 ( .A(n3503), .B(n3504), .Z(n3465) );
  AND U3950 ( .A(n3505), .B(n3506), .Z(n3504) );
  XNOR U3951 ( .A(n3507), .B(n3508), .Z(n3506) );
  XNOR U3952 ( .A(n3503), .B(n3509), .Z(n3508) );
  XOR U3953 ( .A(n3492), .B(n3510), .Z(n3505) );
  XNOR U3954 ( .A(n3503), .B(n3493), .Z(n3510) );
  XNOR U3955 ( .A(n3475), .B(n3512), .Z(n3476) );
  AND U3956 ( .A(n2036), .B(n1858), .Z(n3512) );
  XOR U3957 ( .A(n3516), .B(n3477), .Z(n3511) );
  NAND U3958 ( .A(n1757), .B(n2141), .Z(n3477) );
  IV U3959 ( .A(n3479), .Z(n3516) );
  XNOR U3960 ( .A(n3484), .B(n3485), .Z(n3481) );
  NAND U3961 ( .A(n1574), .B(n2370), .Z(n3485) );
  XNOR U3962 ( .A(n3483), .B(n3520), .Z(n3484) );
  AND U3963 ( .A(n2254), .B(n1668), .Z(n3520) );
  XOR U3964 ( .A(n3524), .B(n3502), .Z(n3492) );
  XNOR U3965 ( .A(n3489), .B(n3490), .Z(n3502) );
  NAND U3966 ( .A(n1952), .B(n1931), .Z(n3490) );
  XNOR U3967 ( .A(n3488), .B(n3525), .Z(n3489) );
  AND U3968 ( .A(n1831), .B(n2053), .Z(n3525) );
  XNOR U3969 ( .A(n3501), .B(n3491), .Z(n3524) );
  XNOR U3970 ( .A(n3496), .B(n3533), .Z(n3497) );
  AND U3971 ( .A(n1646), .B(n2282), .Z(n3533) );
  XOR U3972 ( .A(n3537), .B(n3498), .Z(n3532) );
  NAND U3973 ( .A(n2166), .B(n1737), .Z(n3498) );
  IV U3974 ( .A(n3500), .Z(n3537) );
  XOR U3975 ( .A(n3541), .B(n3542), .Z(n3503) );
  AND U3976 ( .A(n3543), .B(n3544), .Z(n3542) );
  XNOR U3977 ( .A(n3545), .B(n3546), .Z(n3544) );
  XNOR U3978 ( .A(n3541), .B(n3547), .Z(n3546) );
  XOR U3979 ( .A(n3530), .B(n3548), .Z(n3543) );
  XNOR U3980 ( .A(n3541), .B(n3531), .Z(n3548) );
  XNOR U3981 ( .A(n3513), .B(n3550), .Z(n3514) );
  AND U3982 ( .A(n2141), .B(n1858), .Z(n3550) );
  XOR U3983 ( .A(n3554), .B(n3515), .Z(n3549) );
  NAND U3984 ( .A(n1757), .B(n2254), .Z(n3515) );
  IV U3985 ( .A(n3517), .Z(n3554) );
  XNOR U3986 ( .A(n3522), .B(n3523), .Z(n3519) );
  NAND U3987 ( .A(n1574), .B(n2491), .Z(n3523) );
  XNOR U3988 ( .A(n3521), .B(n3558), .Z(n3522) );
  AND U3989 ( .A(n2370), .B(n1668), .Z(n3558) );
  XOR U3990 ( .A(n3562), .B(n3540), .Z(n3530) );
  XNOR U3991 ( .A(n3527), .B(n3528), .Z(n3540) );
  NAND U3992 ( .A(n1952), .B(n2036), .Z(n3528) );
  XNOR U3993 ( .A(n3526), .B(n3563), .Z(n3527) );
  AND U3994 ( .A(n1931), .B(n2053), .Z(n3563) );
  XNOR U3995 ( .A(n3539), .B(n3529), .Z(n3562) );
  XNOR U3996 ( .A(n3534), .B(n3571), .Z(n3535) );
  AND U3997 ( .A(n1737), .B(n2282), .Z(n3571) );
  XOR U3998 ( .A(n3575), .B(n3536), .Z(n3570) );
  NAND U3999 ( .A(n2166), .B(n1831), .Z(n3536) );
  IV U4000 ( .A(n3538), .Z(n3575) );
  XOR U4001 ( .A(n3579), .B(n3580), .Z(n3541) );
  AND U4002 ( .A(n3581), .B(n3582), .Z(n3580) );
  XNOR U4003 ( .A(n3583), .B(n3584), .Z(n3582) );
  XNOR U4004 ( .A(n3579), .B(n3585), .Z(n3584) );
  XOR U4005 ( .A(n3568), .B(n3586), .Z(n3581) );
  XNOR U4006 ( .A(n3579), .B(n3569), .Z(n3586) );
  XNOR U4007 ( .A(n3551), .B(n3588), .Z(n3552) );
  AND U4008 ( .A(n2254), .B(n1858), .Z(n3588) );
  XOR U4009 ( .A(n3592), .B(n3553), .Z(n3587) );
  NAND U4010 ( .A(n1757), .B(n2370), .Z(n3553) );
  IV U4011 ( .A(n3555), .Z(n3592) );
  XNOR U4012 ( .A(n3560), .B(n3561), .Z(n3557) );
  NAND U4013 ( .A(n1574), .B(n2615), .Z(n3561) );
  XNOR U4014 ( .A(n3559), .B(n3596), .Z(n3560) );
  AND U4015 ( .A(n2491), .B(n1668), .Z(n3596) );
  XOR U4016 ( .A(n3600), .B(n3578), .Z(n3568) );
  XNOR U4017 ( .A(n3565), .B(n3566), .Z(n3578) );
  NAND U4018 ( .A(n1952), .B(n2141), .Z(n3566) );
  XNOR U4019 ( .A(n3564), .B(n3601), .Z(n3565) );
  AND U4020 ( .A(n2036), .B(n2053), .Z(n3601) );
  XNOR U4021 ( .A(n3577), .B(n3567), .Z(n3600) );
  XNOR U4022 ( .A(n3572), .B(n3609), .Z(n3573) );
  AND U4023 ( .A(n1831), .B(n2282), .Z(n3609) );
  XOR U4024 ( .A(n3613), .B(n3574), .Z(n3608) );
  NAND U4025 ( .A(n2166), .B(n1931), .Z(n3574) );
  IV U4026 ( .A(n3576), .Z(n3613) );
  XOR U4027 ( .A(n3617), .B(n3618), .Z(n3579) );
  AND U4028 ( .A(n3619), .B(n3620), .Z(n3618) );
  XNOR U4029 ( .A(n3621), .B(n3622), .Z(n3620) );
  XNOR U4030 ( .A(n3617), .B(n3623), .Z(n3622) );
  XOR U4031 ( .A(n3606), .B(n3624), .Z(n3619) );
  XNOR U4032 ( .A(n3617), .B(n3607), .Z(n3624) );
  XNOR U4033 ( .A(n3589), .B(n3626), .Z(n3590) );
  AND U4034 ( .A(n2370), .B(n1858), .Z(n3626) );
  XOR U4035 ( .A(n3630), .B(n3591), .Z(n3625) );
  NAND U4036 ( .A(n1757), .B(n2491), .Z(n3591) );
  IV U4037 ( .A(n3593), .Z(n3630) );
  XNOR U4038 ( .A(n3598), .B(n3599), .Z(n3595) );
  NAND U4039 ( .A(n1574), .B(n2743), .Z(n3599) );
  XNOR U4040 ( .A(n3597), .B(n3634), .Z(n3598) );
  AND U4041 ( .A(n2615), .B(n1668), .Z(n3634) );
  XOR U4042 ( .A(n3638), .B(n3616), .Z(n3606) );
  XNOR U4043 ( .A(n3603), .B(n3604), .Z(n3616) );
  NAND U4044 ( .A(n1952), .B(n2254), .Z(n3604) );
  XNOR U4045 ( .A(n3602), .B(n3639), .Z(n3603) );
  AND U4046 ( .A(n2141), .B(n2053), .Z(n3639) );
  XNOR U4047 ( .A(n3615), .B(n3605), .Z(n3638) );
  XNOR U4048 ( .A(n3610), .B(n3647), .Z(n3611) );
  AND U4049 ( .A(n1931), .B(n2282), .Z(n3647) );
  XOR U4050 ( .A(n3651), .B(n3612), .Z(n3646) );
  NAND U4051 ( .A(n2166), .B(n2036), .Z(n3612) );
  IV U4052 ( .A(n3614), .Z(n3651) );
  XOR U4053 ( .A(n3655), .B(n3656), .Z(n3617) );
  AND U4054 ( .A(n3657), .B(n3658), .Z(n3656) );
  XNOR U4055 ( .A(n3659), .B(n3660), .Z(n3658) );
  XNOR U4056 ( .A(n3655), .B(n3661), .Z(n3660) );
  XOR U4057 ( .A(n3644), .B(n3662), .Z(n3657) );
  XNOR U4058 ( .A(n3655), .B(n3645), .Z(n3662) );
  XNOR U4059 ( .A(n3627), .B(n3664), .Z(n3628) );
  AND U4060 ( .A(n2491), .B(n1858), .Z(n3664) );
  XOR U4061 ( .A(n3668), .B(n3629), .Z(n3663) );
  NAND U4062 ( .A(n1757), .B(n2615), .Z(n3629) );
  IV U4063 ( .A(n3631), .Z(n3668) );
  XNOR U4064 ( .A(n3636), .B(n3637), .Z(n3633) );
  NANDN U4065 ( .B(n2872), .A(n1574), .Z(n3637) );
  XNOR U4066 ( .A(n3635), .B(n3672), .Z(n3636) );
  AND U4067 ( .A(n2743), .B(n1668), .Z(n3672) );
  XOR U4068 ( .A(n3676), .B(n3654), .Z(n3644) );
  XNOR U4069 ( .A(n3641), .B(n3642), .Z(n3654) );
  NAND U4070 ( .A(n1952), .B(n2370), .Z(n3642) );
  XNOR U4071 ( .A(n3640), .B(n3677), .Z(n3641) );
  AND U4072 ( .A(n2254), .B(n2053), .Z(n3677) );
  XNOR U4073 ( .A(n3653), .B(n3643), .Z(n3676) );
  XNOR U4074 ( .A(n3648), .B(n3685), .Z(n3649) );
  AND U4075 ( .A(n2036), .B(n2282), .Z(n3685) );
  XOR U4076 ( .A(n3689), .B(n3650), .Z(n3684) );
  NAND U4077 ( .A(n2166), .B(n2141), .Z(n3650) );
  IV U4078 ( .A(n3652), .Z(n3689) );
  XOR U4079 ( .A(n3693), .B(n3694), .Z(n3655) );
  AND U4080 ( .A(n3695), .B(n3696), .Z(n3694) );
  XNOR U4081 ( .A(n3697), .B(n3698), .Z(n3696) );
  XNOR U4082 ( .A(n3693), .B(n3699), .Z(n3698) );
  XOR U4083 ( .A(n3682), .B(n3700), .Z(n3695) );
  XNOR U4084 ( .A(n3693), .B(n3683), .Z(n3700) );
  XNOR U4085 ( .A(n3665), .B(n3702), .Z(n3666) );
  AND U4086 ( .A(n2615), .B(n1858), .Z(n3702) );
  XOR U4087 ( .A(n3706), .B(n3667), .Z(n3701) );
  NAND U4088 ( .A(n1757), .B(n2743), .Z(n3667) );
  IV U4089 ( .A(n3669), .Z(n3706) );
  XNOR U4090 ( .A(n3674), .B(n3675), .Z(n3671) );
  NANDN U4091 ( .B(n3010), .A(n1574), .Z(n3675) );
  XNOR U4092 ( .A(n3673), .B(n3710), .Z(n3674) );
  ANDN U4093 ( .A(n1668), .B(n2872), .Z(n3710) );
  XOR U4094 ( .A(n3714), .B(n3692), .Z(n3682) );
  XNOR U4095 ( .A(n3679), .B(n3680), .Z(n3692) );
  NAND U4096 ( .A(n1952), .B(n2491), .Z(n3680) );
  XNOR U4097 ( .A(n3678), .B(n3715), .Z(n3679) );
  AND U4098 ( .A(n2370), .B(n2053), .Z(n3715) );
  XNOR U4099 ( .A(n3691), .B(n3681), .Z(n3714) );
  XNOR U4100 ( .A(n3686), .B(n3723), .Z(n3687) );
  AND U4101 ( .A(n2141), .B(n2282), .Z(n3723) );
  XOR U4102 ( .A(n3727), .B(n3688), .Z(n3722) );
  NAND U4103 ( .A(n2166), .B(n2254), .Z(n3688) );
  IV U4104 ( .A(n3690), .Z(n3727) );
  XOR U4105 ( .A(n3731), .B(n3732), .Z(n3693) );
  AND U4106 ( .A(n3733), .B(n3734), .Z(n3732) );
  XNOR U4107 ( .A(n3735), .B(n3736), .Z(n3734) );
  XNOR U4108 ( .A(n3731), .B(n3737), .Z(n3736) );
  XOR U4109 ( .A(n3720), .B(n3738), .Z(n3733) );
  XNOR U4110 ( .A(n3731), .B(n3721), .Z(n3738) );
  XNOR U4111 ( .A(n3703), .B(n3740), .Z(n3704) );
  AND U4112 ( .A(n2743), .B(n1858), .Z(n3740) );
  XOR U4113 ( .A(n3744), .B(n3705), .Z(n3739) );
  NANDN U4114 ( .B(n2872), .A(n1757), .Z(n3705) );
  IV U4115 ( .A(n3707), .Z(n3744) );
  XNOR U4116 ( .A(n3712), .B(n3713), .Z(n3709) );
  NAND U4117 ( .A(n1574), .B(n3146), .Z(n3713) );
  XNOR U4118 ( .A(n3711), .B(n3748), .Z(n3712) );
  ANDN U4119 ( .A(n1668), .B(n3010), .Z(n3748) );
  XOR U4120 ( .A(n3752), .B(n3730), .Z(n3720) );
  XNOR U4121 ( .A(n3717), .B(n3718), .Z(n3730) );
  NAND U4122 ( .A(n1952), .B(n2615), .Z(n3718) );
  XNOR U4123 ( .A(n3716), .B(n3753), .Z(n3717) );
  AND U4124 ( .A(n2491), .B(n2053), .Z(n3753) );
  XNOR U4125 ( .A(n3729), .B(n3719), .Z(n3752) );
  XNOR U4126 ( .A(n3724), .B(n3761), .Z(n3725) );
  AND U4127 ( .A(n2254), .B(n2282), .Z(n3761) );
  XOR U4128 ( .A(n3765), .B(n3726), .Z(n3760) );
  NAND U4129 ( .A(n2166), .B(n2370), .Z(n3726) );
  IV U4130 ( .A(n3728), .Z(n3765) );
  XNOR U4131 ( .A(n3770), .B(n3771), .Z(n3184) );
  XOR U4132 ( .A(n3772), .B(n3769), .Z(n3770) );
  XNOR U4133 ( .A(n3773), .B(n3768), .Z(n3758) );
  XNOR U4134 ( .A(n3755), .B(n3756), .Z(n3768) );
  NAND U4135 ( .A(n1952), .B(n2743), .Z(n3756) );
  XNOR U4136 ( .A(n3754), .B(n3774), .Z(n3755) );
  AND U4137 ( .A(n2615), .B(n2053), .Z(n3774) );
  XNOR U4138 ( .A(n3778), .B(n3775), .Z(n3777) );
  XNOR U4139 ( .A(n3767), .B(n3757), .Z(n3773) );
  XOR U4140 ( .A(n3779), .B(n3780), .Z(n3757) );
  XNOR U4141 ( .A(n3762), .B(n3782), .Z(n3763) );
  AND U4142 ( .A(n2370), .B(n2282), .Z(n3782) );
  XNOR U4143 ( .A(n3786), .B(n3783), .Z(n3785) );
  XOR U4144 ( .A(n3787), .B(n3764), .Z(n3781) );
  NAND U4145 ( .A(n2166), .B(n2491), .Z(n3764) );
  IV U4146 ( .A(n3766), .Z(n3787) );
  XNOR U4147 ( .A(n3788), .B(n3789), .Z(n3766) );
  AND U4148 ( .A(n3790), .B(n3791), .Z(n3789) );
  XOR U4149 ( .A(n3784), .B(n3792), .Z(n3791) );
  XNOR U4150 ( .A(n3786), .B(n3788), .Z(n3792) );
  NAND U4151 ( .A(n2166), .B(n2615), .Z(n3786) );
  XOR U4152 ( .A(n3783), .B(n3793), .Z(n3784) );
  AND U4153 ( .A(n2491), .B(n2282), .Z(n3793) );
  XNOR U4154 ( .A(n3797), .B(n3794), .Z(n3796) );
  XOR U4155 ( .A(n3776), .B(n3798), .Z(n3790) );
  XNOR U4156 ( .A(n3778), .B(n3788), .Z(n3798) );
  NANDN U4157 ( .B(n2872), .A(n1952), .Z(n3778) );
  XOR U4158 ( .A(n3775), .B(n3799), .Z(n3776) );
  AND U4159 ( .A(n2743), .B(n2053), .Z(n3799) );
  XNOR U4160 ( .A(n3803), .B(n3800), .Z(n3802) );
  XOR U4161 ( .A(n3804), .B(n3805), .Z(n3788) );
  AND U4162 ( .A(n3806), .B(n3807), .Z(n3805) );
  XOR U4163 ( .A(n3795), .B(n3808), .Z(n3807) );
  XNOR U4164 ( .A(n3797), .B(n3804), .Z(n3808) );
  NAND U4165 ( .A(n2166), .B(n2743), .Z(n3797) );
  XOR U4166 ( .A(n3794), .B(n3809), .Z(n3795) );
  AND U4167 ( .A(n2615), .B(n2282), .Z(n3809) );
  XNOR U4168 ( .A(n3813), .B(n3810), .Z(n3812) );
  XOR U4169 ( .A(n3801), .B(n3814), .Z(n3806) );
  XNOR U4170 ( .A(n3803), .B(n3804), .Z(n3814) );
  NANDN U4171 ( .B(n3010), .A(n1952), .Z(n3803) );
  XOR U4172 ( .A(n3800), .B(n3815), .Z(n3801) );
  ANDN U4173 ( .A(n2053), .B(n2872), .Z(n3815) );
  XNOR U4174 ( .A(n3819), .B(n3816), .Z(n3818) );
  XOR U4175 ( .A(n3820), .B(n3821), .Z(n3804) );
  AND U4176 ( .A(n3822), .B(n3823), .Z(n3821) );
  XOR U4177 ( .A(n3811), .B(n3824), .Z(n3823) );
  XNOR U4178 ( .A(n3813), .B(n3820), .Z(n3824) );
  NANDN U4179 ( .B(n2872), .A(n2166), .Z(n3813) );
  XOR U4180 ( .A(n3810), .B(n3825), .Z(n3811) );
  AND U4181 ( .A(n2743), .B(n2282), .Z(n3825) );
  XOR U4182 ( .A(n3817), .B(n3829), .Z(n3822) );
  XNOR U4183 ( .A(n3819), .B(n3820), .Z(n3829) );
  NAND U4184 ( .A(n1952), .B(n3146), .Z(n3819) );
  XOR U4185 ( .A(n3816), .B(n3830), .Z(n3817) );
  ANDN U4186 ( .A(n2053), .B(n3010), .Z(n3830) );
  NAND U4187 ( .A(n1952), .B(n3835), .Z(n3833) );
  XNOR U4188 ( .A(n3831), .B(n3836), .Z(n3832) );
  AND U4189 ( .A(n3146), .B(n2053), .Z(n3836) );
  AND U4190 ( .A(n3837), .B(g_input[0]), .Z(n3831) );
  NANDN U4191 ( .B(n1952), .A(n3838), .Z(n3837) );
  NAND U4192 ( .A(n3835), .B(n2053), .Z(n3838) );
  XNOR U4193 ( .A(n3826), .B(n3842), .Z(n3827) );
  ANDN U4194 ( .A(n2282), .B(n2872), .Z(n3842) );
  XOR U4195 ( .A(n3845), .B(n3843), .Z(n3844) );
  ANDN U4196 ( .A(n2282), .B(n3010), .Z(n3845) );
  AND U4197 ( .A(n3146), .B(n2166), .Z(n3846) );
  XOR U4198 ( .A(n3850), .B(n3828), .Z(n3841) );
  NANDN U4199 ( .B(n3010), .A(n2166), .Z(n3828) );
  IV U4200 ( .A(n3834), .Z(n3850) );
  NAND U4201 ( .A(n2166), .B(n3835), .Z(n3849) );
  XNOR U4202 ( .A(n3847), .B(n3851), .Z(n3848) );
  AND U4203 ( .A(n3146), .B(n2282), .Z(n3851) );
  AND U4204 ( .A(n3852), .B(g_input[0]), .Z(n3847) );
  NANDN U4205 ( .B(n2166), .A(n3853), .Z(n3852) );
  NAND U4206 ( .A(n3835), .B(n2282), .Z(n3853) );
  XNOR U4207 ( .A(n3741), .B(n3857), .Z(n3742) );
  ANDN U4208 ( .A(n1858), .B(n2872), .Z(n3857) );
  XOR U4209 ( .A(n3860), .B(n3858), .Z(n3859) );
  ANDN U4210 ( .A(n1858), .B(n3010), .Z(n3860) );
  AND U4211 ( .A(n3146), .B(n1757), .Z(n3861) );
  XOR U4212 ( .A(n3865), .B(n3743), .Z(n3856) );
  NANDN U4213 ( .B(n3010), .A(n1757), .Z(n3743) );
  IV U4214 ( .A(n3745), .Z(n3865) );
  NAND U4215 ( .A(n1757), .B(n3835), .Z(n3864) );
  XNOR U4216 ( .A(n3862), .B(n3866), .Z(n3863) );
  AND U4217 ( .A(n3146), .B(n1858), .Z(n3866) );
  AND U4218 ( .A(n3867), .B(g_input[0]), .Z(n3862) );
  NANDN U4219 ( .B(n1757), .A(n3868), .Z(n3867) );
  NAND U4220 ( .A(n3835), .B(n1858), .Z(n3868) );
  XNOR U4221 ( .A(n3750), .B(n3751), .Z(n3747) );
  NAND U4222 ( .A(n1574), .B(n3835), .Z(n3751) );
  XNOR U4223 ( .A(n3749), .B(n3871), .Z(n3750) );
  AND U4224 ( .A(n3146), .B(n1668), .Z(n3871) );
  AND U4225 ( .A(n3872), .B(g_input[0]), .Z(n3749) );
  NANDN U4226 ( .B(n1574), .A(n3873), .Z(n3872) );
  NAND U4227 ( .A(n3835), .B(n1668), .Z(n3873) );
  XOR U4228 ( .A(n3876), .B(n3877), .Z(n3769) );
  XNOR U4229 ( .A(n3878), .B(n3085), .Z(n3081) );
  NAND U4230 ( .A(n775), .B(n2944), .Z(n3079) );
  XNOR U4231 ( .A(n3077), .B(n3879), .Z(n3078) );
  AND U4232 ( .A(n3076), .B(n744), .Z(n3879) );
  XNOR U4233 ( .A(n3084), .B(n3080), .Z(n3878) );
  XNOR U4234 ( .A(n3188), .B(n3885), .Z(n3189) );
  AND U4235 ( .A(n2798), .B(n853), .Z(n3885) );
  XOR U4236 ( .A(n3889), .B(n3190), .Z(n3884) );
  NAND U4237 ( .A(n897), .B(n2668), .Z(n3190) );
  IV U4238 ( .A(n3192), .Z(n3889) );
  XNOR U4239 ( .A(n3197), .B(n3198), .Z(n3194) );
  NAND U4240 ( .A(n1001), .B(n2421), .Z(n3198) );
  XNOR U4241 ( .A(n3196), .B(n3893), .Z(n3197) );
  AND U4242 ( .A(n2544), .B(n941), .Z(n3893) );
  XOR U4243 ( .A(n3897), .B(n3898), .Z(n3205) );
  XNOR U4244 ( .A(n3899), .B(n3883), .Z(n3897) );
  XOR U4245 ( .A(n3901), .B(n3902), .Z(n3243) );
  XNOR U4246 ( .A(n3903), .B(n3900), .Z(n3901) );
  XNOR U4247 ( .A(n3886), .B(n3905), .Z(n3887) );
  AND U4248 ( .A(n2798), .B(n897), .Z(n3905) );
  XOR U4249 ( .A(n3909), .B(n3888), .Z(n3904) );
  NAND U4250 ( .A(n941), .B(n2668), .Z(n3888) );
  IV U4251 ( .A(n3890), .Z(n3909) );
  XNOR U4252 ( .A(n3895), .B(n3896), .Z(n3892) );
  NAND U4253 ( .A(n1055), .B(n2421), .Z(n3896) );
  XNOR U4254 ( .A(n3894), .B(n3913), .Z(n3895) );
  AND U4255 ( .A(n2544), .B(n1001), .Z(n3913) );
  XOR U4256 ( .A(n3918), .B(n3919), .Z(n3281) );
  XNOR U4257 ( .A(n3920), .B(n3917), .Z(n3918) );
  XNOR U4258 ( .A(n3906), .B(n3922), .Z(n3907) );
  AND U4259 ( .A(n2798), .B(n941), .Z(n3922) );
  XOR U4260 ( .A(n3926), .B(n3908), .Z(n3921) );
  NAND U4261 ( .A(n1001), .B(n2668), .Z(n3908) );
  IV U4262 ( .A(n3910), .Z(n3926) );
  XNOR U4263 ( .A(n3915), .B(n3916), .Z(n3912) );
  NAND U4264 ( .A(n1116), .B(n2421), .Z(n3916) );
  XNOR U4265 ( .A(n3914), .B(n3930), .Z(n3915) );
  AND U4266 ( .A(n2544), .B(n1055), .Z(n3930) );
  XOR U4267 ( .A(n3935), .B(n3936), .Z(n3319) );
  XNOR U4268 ( .A(n3937), .B(n3934), .Z(n3935) );
  XNOR U4269 ( .A(n3923), .B(n3939), .Z(n3924) );
  AND U4270 ( .A(n2798), .B(n1001), .Z(n3939) );
  XOR U4271 ( .A(n3943), .B(n3925), .Z(n3938) );
  NAND U4272 ( .A(n1055), .B(n2668), .Z(n3925) );
  IV U4273 ( .A(n3927), .Z(n3943) );
  XNOR U4274 ( .A(n3932), .B(n3933), .Z(n3929) );
  NAND U4275 ( .A(n1178), .B(n2421), .Z(n3933) );
  XNOR U4276 ( .A(n3931), .B(n3947), .Z(n3932) );
  AND U4277 ( .A(n2544), .B(n1116), .Z(n3947) );
  XOR U4278 ( .A(n3952), .B(n3953), .Z(n3357) );
  XNOR U4279 ( .A(n3954), .B(n3951), .Z(n3952) );
  XNOR U4280 ( .A(n3940), .B(n3956), .Z(n3941) );
  AND U4281 ( .A(n2798), .B(n1055), .Z(n3956) );
  XOR U4282 ( .A(n3960), .B(n3942), .Z(n3955) );
  NAND U4283 ( .A(n1116), .B(n2668), .Z(n3942) );
  IV U4284 ( .A(n3944), .Z(n3960) );
  XNOR U4285 ( .A(n3949), .B(n3950), .Z(n3946) );
  NAND U4286 ( .A(n1246), .B(n2421), .Z(n3950) );
  XNOR U4287 ( .A(n3948), .B(n3964), .Z(n3949) );
  AND U4288 ( .A(n2544), .B(n1178), .Z(n3964) );
  XOR U4289 ( .A(n3969), .B(n3970), .Z(n3395) );
  XNOR U4290 ( .A(n3971), .B(n3968), .Z(n3969) );
  XNOR U4291 ( .A(n3957), .B(n3973), .Z(n3958) );
  AND U4292 ( .A(n2798), .B(n1116), .Z(n3973) );
  XOR U4293 ( .A(n3977), .B(n3959), .Z(n3972) );
  NAND U4294 ( .A(n1178), .B(n2668), .Z(n3959) );
  IV U4295 ( .A(n3961), .Z(n3977) );
  XNOR U4296 ( .A(n3966), .B(n3967), .Z(n3963) );
  NAND U4297 ( .A(n1316), .B(n2421), .Z(n3967) );
  XNOR U4298 ( .A(n3965), .B(n3981), .Z(n3966) );
  AND U4299 ( .A(n2544), .B(n1246), .Z(n3981) );
  XOR U4300 ( .A(n3986), .B(n3987), .Z(n3433) );
  XNOR U4301 ( .A(n3988), .B(n3985), .Z(n3986) );
  XNOR U4302 ( .A(n3974), .B(n3990), .Z(n3975) );
  AND U4303 ( .A(n2798), .B(n1178), .Z(n3990) );
  XOR U4304 ( .A(n3994), .B(n3976), .Z(n3989) );
  NAND U4305 ( .A(n1246), .B(n2668), .Z(n3976) );
  IV U4306 ( .A(n3978), .Z(n3994) );
  XNOR U4307 ( .A(n3983), .B(n3984), .Z(n3980) );
  NAND U4308 ( .A(n1390), .B(n2421), .Z(n3984) );
  XNOR U4309 ( .A(n3982), .B(n3998), .Z(n3983) );
  AND U4310 ( .A(n2544), .B(n1316), .Z(n3998) );
  XOR U4311 ( .A(n4003), .B(n4004), .Z(n3471) );
  XNOR U4312 ( .A(n4005), .B(n4002), .Z(n4003) );
  XNOR U4313 ( .A(n3991), .B(n4007), .Z(n3992) );
  AND U4314 ( .A(n2798), .B(n1246), .Z(n4007) );
  XOR U4315 ( .A(n4011), .B(n3993), .Z(n4006) );
  NAND U4316 ( .A(n1316), .B(n2668), .Z(n3993) );
  IV U4317 ( .A(n3995), .Z(n4011) );
  XNOR U4318 ( .A(n4000), .B(n4001), .Z(n3997) );
  NAND U4319 ( .A(n1467), .B(n2421), .Z(n4001) );
  XNOR U4320 ( .A(n3999), .B(n4015), .Z(n4000) );
  AND U4321 ( .A(n2544), .B(n1390), .Z(n4015) );
  XOR U4322 ( .A(n4020), .B(n4021), .Z(n3509) );
  XNOR U4323 ( .A(n4022), .B(n4019), .Z(n4020) );
  XNOR U4324 ( .A(n4008), .B(n4024), .Z(n4009) );
  AND U4325 ( .A(n2798), .B(n1316), .Z(n4024) );
  XOR U4326 ( .A(n4028), .B(n4010), .Z(n4023) );
  NAND U4327 ( .A(n1390), .B(n2668), .Z(n4010) );
  IV U4328 ( .A(n4012), .Z(n4028) );
  XNOR U4329 ( .A(n4017), .B(n4018), .Z(n4014) );
  NAND U4330 ( .A(n1554), .B(n2421), .Z(n4018) );
  XNOR U4331 ( .A(n4016), .B(n4032), .Z(n4017) );
  AND U4332 ( .A(n2544), .B(n1467), .Z(n4032) );
  XOR U4333 ( .A(n4037), .B(n4038), .Z(n3547) );
  XNOR U4334 ( .A(n4039), .B(n4036), .Z(n4037) );
  XNOR U4335 ( .A(n4025), .B(n4041), .Z(n4026) );
  AND U4336 ( .A(n2798), .B(n1390), .Z(n4041) );
  XOR U4337 ( .A(n4045), .B(n4027), .Z(n4040) );
  NAND U4338 ( .A(n1467), .B(n2668), .Z(n4027) );
  IV U4339 ( .A(n4029), .Z(n4045) );
  XNOR U4340 ( .A(n4034), .B(n4035), .Z(n4031) );
  NAND U4341 ( .A(n1646), .B(n2421), .Z(n4035) );
  XNOR U4342 ( .A(n4033), .B(n4049), .Z(n4034) );
  AND U4343 ( .A(n2544), .B(n1554), .Z(n4049) );
  XOR U4344 ( .A(n4054), .B(n4055), .Z(n3585) );
  XNOR U4345 ( .A(n4056), .B(n4053), .Z(n4054) );
  XNOR U4346 ( .A(n4042), .B(n4058), .Z(n4043) );
  AND U4347 ( .A(n2798), .B(n1467), .Z(n4058) );
  XOR U4348 ( .A(n4062), .B(n4044), .Z(n4057) );
  NAND U4349 ( .A(n1554), .B(n2668), .Z(n4044) );
  IV U4350 ( .A(n4046), .Z(n4062) );
  XNOR U4351 ( .A(n4051), .B(n4052), .Z(n4048) );
  NAND U4352 ( .A(n1737), .B(n2421), .Z(n4052) );
  XNOR U4353 ( .A(n4050), .B(n4066), .Z(n4051) );
  AND U4354 ( .A(n2544), .B(n1646), .Z(n4066) );
  XOR U4355 ( .A(n4071), .B(n4072), .Z(n3623) );
  XNOR U4356 ( .A(n4073), .B(n4070), .Z(n4071) );
  XNOR U4357 ( .A(n4059), .B(n4075), .Z(n4060) );
  AND U4358 ( .A(n2798), .B(n1554), .Z(n4075) );
  XOR U4359 ( .A(n4079), .B(n4061), .Z(n4074) );
  NAND U4360 ( .A(n1646), .B(n2668), .Z(n4061) );
  IV U4361 ( .A(n4063), .Z(n4079) );
  XNOR U4362 ( .A(n4068), .B(n4069), .Z(n4065) );
  NAND U4363 ( .A(n1831), .B(n2421), .Z(n4069) );
  XNOR U4364 ( .A(n4067), .B(n4083), .Z(n4068) );
  AND U4365 ( .A(n2544), .B(n1737), .Z(n4083) );
  XOR U4366 ( .A(n4088), .B(n4089), .Z(n3661) );
  XNOR U4367 ( .A(n4090), .B(n4087), .Z(n4088) );
  XNOR U4368 ( .A(n4076), .B(n4092), .Z(n4077) );
  AND U4369 ( .A(n2798), .B(n1646), .Z(n4092) );
  XOR U4370 ( .A(n4096), .B(n4078), .Z(n4091) );
  NAND U4371 ( .A(n1737), .B(n2668), .Z(n4078) );
  IV U4372 ( .A(n4080), .Z(n4096) );
  XNOR U4373 ( .A(n4085), .B(n4086), .Z(n4082) );
  NAND U4374 ( .A(n1931), .B(n2421), .Z(n4086) );
  XNOR U4375 ( .A(n4084), .B(n4100), .Z(n4085) );
  AND U4376 ( .A(n2544), .B(n1831), .Z(n4100) );
  XOR U4377 ( .A(n4105), .B(n4106), .Z(n3699) );
  XNOR U4378 ( .A(n4107), .B(n4104), .Z(n4105) );
  XNOR U4379 ( .A(n4093), .B(n4109), .Z(n4094) );
  AND U4380 ( .A(n2798), .B(n1737), .Z(n4109) );
  XOR U4381 ( .A(n4113), .B(n4095), .Z(n4108) );
  NAND U4382 ( .A(n1831), .B(n2668), .Z(n4095) );
  IV U4383 ( .A(n4097), .Z(n4113) );
  XNOR U4384 ( .A(n4102), .B(n4103), .Z(n4099) );
  NAND U4385 ( .A(n2036), .B(n2421), .Z(n4103) );
  XNOR U4386 ( .A(n4101), .B(n4117), .Z(n4102) );
  AND U4387 ( .A(n2544), .B(n1931), .Z(n4117) );
  XOR U4388 ( .A(n4122), .B(n4123), .Z(n3737) );
  XNOR U4389 ( .A(n4124), .B(n4121), .Z(n4122) );
  XNOR U4390 ( .A(n4110), .B(n4126), .Z(n4111) );
  AND U4391 ( .A(n2798), .B(n1831), .Z(n4126) );
  XOR U4392 ( .A(n4130), .B(n4112), .Z(n4125) );
  NAND U4393 ( .A(n1931), .B(n2668), .Z(n4112) );
  IV U4394 ( .A(n4114), .Z(n4130) );
  XNOR U4395 ( .A(n4119), .B(n4120), .Z(n4116) );
  NAND U4396 ( .A(n2141), .B(n2421), .Z(n4120) );
  XNOR U4397 ( .A(n4118), .B(n4134), .Z(n4119) );
  AND U4398 ( .A(n2544), .B(n2036), .Z(n4134) );
  XOR U4399 ( .A(n4139), .B(n4140), .Z(n3772) );
  XNOR U4400 ( .A(n4141), .B(n4138), .Z(n4139) );
  XNOR U4401 ( .A(n4127), .B(n4143), .Z(n4128) );
  AND U4402 ( .A(n2798), .B(n1931), .Z(n4143) );
  XOR U4403 ( .A(n4147), .B(n4129), .Z(n4142) );
  NAND U4404 ( .A(n2036), .B(n2668), .Z(n4129) );
  IV U4405 ( .A(n4131), .Z(n4147) );
  XNOR U4406 ( .A(n4136), .B(n4137), .Z(n4133) );
  NAND U4407 ( .A(n2254), .B(n2421), .Z(n4137) );
  XNOR U4408 ( .A(n4135), .B(n4151), .Z(n4136) );
  AND U4409 ( .A(n2544), .B(n2141), .Z(n4151) );
  XOR U4410 ( .A(n4155), .B(n4156), .Z(n4138) );
  AND U4411 ( .A(n4157), .B(n4158), .Z(n4156) );
  XOR U4412 ( .A(n4159), .B(n4160), .Z(n4158) );
  XOR U4413 ( .A(n4155), .B(n4161), .Z(n4160) );
  XOR U4414 ( .A(n4149), .B(n4162), .Z(n4157) );
  XOR U4415 ( .A(n4155), .B(n4150), .Z(n4162) );
  NAND U4416 ( .A(n2421), .B(n2370), .Z(n4154) );
  XNOR U4417 ( .A(n4152), .B(n4163), .Z(n4153) );
  AND U4418 ( .A(n2544), .B(n2254), .Z(n4163) );
  XNOR U4419 ( .A(n4144), .B(n4168), .Z(n4145) );
  AND U4420 ( .A(n2798), .B(n2036), .Z(n4168) );
  XOR U4421 ( .A(n4172), .B(n4146), .Z(n4167) );
  NAND U4422 ( .A(n2141), .B(n2668), .Z(n4146) );
  IV U4423 ( .A(n4148), .Z(n4172) );
  XOR U4424 ( .A(n4176), .B(n4177), .Z(n4155) );
  AND U4425 ( .A(n4178), .B(n4179), .Z(n4177) );
  XOR U4426 ( .A(n4180), .B(n4181), .Z(n4179) );
  XOR U4427 ( .A(n4176), .B(n4182), .Z(n4181) );
  XOR U4428 ( .A(n4174), .B(n4183), .Z(n4178) );
  XOR U4429 ( .A(n4176), .B(n4175), .Z(n4183) );
  NAND U4430 ( .A(n2421), .B(n2491), .Z(n4166) );
  XNOR U4431 ( .A(n4164), .B(n4184), .Z(n4165) );
  AND U4432 ( .A(n2370), .B(n2544), .Z(n4184) );
  XNOR U4433 ( .A(n4169), .B(n4189), .Z(n4170) );
  AND U4434 ( .A(n2798), .B(n2141), .Z(n4189) );
  XOR U4435 ( .A(n4193), .B(n4171), .Z(n4188) );
  NAND U4436 ( .A(n2254), .B(n2668), .Z(n4171) );
  IV U4437 ( .A(n4173), .Z(n4193) );
  XOR U4438 ( .A(n4197), .B(n4198), .Z(n4176) );
  AND U4439 ( .A(n4199), .B(n4200), .Z(n4198) );
  XOR U4440 ( .A(n4201), .B(n4202), .Z(n4200) );
  XOR U4441 ( .A(n4197), .B(n4203), .Z(n4202) );
  XOR U4442 ( .A(n4195), .B(n4204), .Z(n4199) );
  XOR U4443 ( .A(n4197), .B(n4196), .Z(n4204) );
  NAND U4444 ( .A(n2421), .B(n2615), .Z(n4187) );
  XNOR U4445 ( .A(n4185), .B(n4205), .Z(n4186) );
  AND U4446 ( .A(n2491), .B(n2544), .Z(n4205) );
  XNOR U4447 ( .A(n4190), .B(n4210), .Z(n4191) );
  AND U4448 ( .A(n2798), .B(n2254), .Z(n4210) );
  XOR U4449 ( .A(n4214), .B(n4192), .Z(n4209) );
  NAND U4450 ( .A(n2668), .B(n2370), .Z(n4192) );
  IV U4451 ( .A(n4194), .Z(n4214) );
  XOR U4452 ( .A(n4218), .B(n4219), .Z(n4197) );
  AND U4453 ( .A(n4220), .B(n4221), .Z(n4219) );
  XOR U4454 ( .A(n4222), .B(n4223), .Z(n4221) );
  XOR U4455 ( .A(n4218), .B(n4224), .Z(n4223) );
  XOR U4456 ( .A(n4216), .B(n4225), .Z(n4220) );
  XOR U4457 ( .A(n4218), .B(n4217), .Z(n4225) );
  NAND U4458 ( .A(n2421), .B(n2743), .Z(n4208) );
  XNOR U4459 ( .A(n4206), .B(n4226), .Z(n4207) );
  AND U4460 ( .A(n2615), .B(n2544), .Z(n4226) );
  XNOR U4461 ( .A(n4211), .B(n4231), .Z(n4212) );
  AND U4462 ( .A(n2370), .B(n2798), .Z(n4231) );
  XOR U4463 ( .A(n4235), .B(n4213), .Z(n4230) );
  NAND U4464 ( .A(n2668), .B(n2491), .Z(n4213) );
  IV U4465 ( .A(n4215), .Z(n4235) );
  XOR U4466 ( .A(n4239), .B(n4240), .Z(n4218) );
  AND U4467 ( .A(n4241), .B(n4242), .Z(n4240) );
  XOR U4468 ( .A(n4243), .B(n4244), .Z(n4242) );
  XOR U4469 ( .A(n4239), .B(n4245), .Z(n4244) );
  XOR U4470 ( .A(n4237), .B(n4246), .Z(n4241) );
  XOR U4471 ( .A(n4239), .B(n4238), .Z(n4246) );
  NANDN U4472 ( .B(n2872), .A(n2421), .Z(n4229) );
  XNOR U4473 ( .A(n4227), .B(n4247), .Z(n4228) );
  AND U4474 ( .A(n2743), .B(n2544), .Z(n4247) );
  XNOR U4475 ( .A(n4232), .B(n4252), .Z(n4233) );
  AND U4476 ( .A(n2491), .B(n2798), .Z(n4252) );
  XOR U4477 ( .A(n4256), .B(n4234), .Z(n4251) );
  NAND U4478 ( .A(n2668), .B(n2615), .Z(n4234) );
  IV U4479 ( .A(n4236), .Z(n4256) );
  XOR U4480 ( .A(n4260), .B(n4261), .Z(n4239) );
  AND U4481 ( .A(n4262), .B(n4263), .Z(n4261) );
  XOR U4482 ( .A(n4264), .B(n4265), .Z(n4263) );
  XOR U4483 ( .A(n4260), .B(n4266), .Z(n4265) );
  XOR U4484 ( .A(n4258), .B(n4267), .Z(n4262) );
  XOR U4485 ( .A(n4260), .B(n4259), .Z(n4267) );
  NANDN U4486 ( .B(n3010), .A(n2421), .Z(n4250) );
  XNOR U4487 ( .A(n4248), .B(n4268), .Z(n4249) );
  ANDN U4488 ( .A(n2544), .B(n2872), .Z(n4268) );
  XNOR U4489 ( .A(n4253), .B(n4273), .Z(n4254) );
  AND U4490 ( .A(n2615), .B(n2798), .Z(n4273) );
  XOR U4491 ( .A(n4277), .B(n4255), .Z(n4272) );
  NAND U4492 ( .A(n2668), .B(n2743), .Z(n4255) );
  IV U4493 ( .A(n4257), .Z(n4277) );
  XOR U4494 ( .A(n4281), .B(n4282), .Z(n4260) );
  AND U4495 ( .A(n4283), .B(n4284), .Z(n4282) );
  XOR U4496 ( .A(n4285), .B(n4286), .Z(n4284) );
  XOR U4497 ( .A(n4281), .B(n4287), .Z(n4286) );
  XOR U4498 ( .A(n4279), .B(n4288), .Z(n4283) );
  XOR U4499 ( .A(n4281), .B(n4280), .Z(n4288) );
  NAND U4500 ( .A(n2421), .B(n3146), .Z(n4271) );
  XNOR U4501 ( .A(n4269), .B(n4289), .Z(n4270) );
  ANDN U4502 ( .A(n2544), .B(n3010), .Z(n4289) );
  XNOR U4503 ( .A(n4274), .B(n4294), .Z(n4275) );
  AND U4504 ( .A(n2743), .B(n2798), .Z(n4294) );
  XOR U4505 ( .A(n4298), .B(n4276), .Z(n4293) );
  NANDN U4506 ( .B(n2872), .A(n2668), .Z(n4276) );
  IV U4507 ( .A(n4278), .Z(n4298) );
  XOR U4508 ( .A(n4303), .B(n4304), .Z(n3877) );
  XNOR U4509 ( .A(n4305), .B(n4302), .Z(n4303) );
  XNOR U4510 ( .A(n4295), .B(n4307), .Z(n4296) );
  ANDN U4511 ( .A(n2798), .B(n2872), .Z(n4307) );
  XOR U4512 ( .A(n4310), .B(n4308), .Z(n4309) );
  ANDN U4513 ( .A(n2798), .B(n3010), .Z(n4310) );
  AND U4514 ( .A(n3146), .B(n2668), .Z(n4311) );
  XOR U4515 ( .A(n4315), .B(n4297), .Z(n4306) );
  NANDN U4516 ( .B(n3010), .A(n2668), .Z(n4297) );
  IV U4517 ( .A(n4299), .Z(n4315) );
  NAND U4518 ( .A(n2668), .B(n3835), .Z(n4314) );
  XNOR U4519 ( .A(n4312), .B(n4316), .Z(n4313) );
  AND U4520 ( .A(n3146), .B(n2798), .Z(n4316) );
  AND U4521 ( .A(n4317), .B(g_input[0]), .Z(n4312) );
  NANDN U4522 ( .B(n2668), .A(n4318), .Z(n4317) );
  NAND U4523 ( .A(n3835), .B(n2798), .Z(n4318) );
  XNOR U4524 ( .A(n4291), .B(n4292), .Z(n4301) );
  NAND U4525 ( .A(n2421), .B(n3835), .Z(n4292) );
  XNOR U4526 ( .A(n4290), .B(n4321), .Z(n4291) );
  AND U4527 ( .A(n3146), .B(n2544), .Z(n4321) );
  AND U4528 ( .A(n4322), .B(g_input[0]), .Z(n4290) );
  NANDN U4529 ( .B(n2421), .A(n4323), .Z(n4322) );
  NAND U4530 ( .A(n3835), .B(n2544), .Z(n4323) );
  XOR U4531 ( .A(n4326), .B(n4327), .Z(n4302) );
  AND U4532 ( .A(n4329), .B(n4330), .Z(n4328) );
  NANDN U4533 ( .B(n717), .A(n4331), .Z(n4330) );
  OR U4534 ( .A(n4332), .B(n4333), .Z(n4329) );
  XNOR U4535 ( .A(n4335), .B(n4334), .Z(n3899) );
  XNOR U4536 ( .A(n4336), .B(n4332), .Z(n4335) );
  NAND U4537 ( .A(n744), .B(n4331), .Z(n4332) );
  NANDN U4538 ( .B(n717), .A(e_input[0]), .Z(n4337) );
  NANDN U4539 ( .B(n4338), .A(n4339), .Z(n717) );
  AND U4540 ( .A(n4340), .B(g_input[31]), .Z(n4339) );
  NAND U4541 ( .A(n814), .B(n2944), .Z(n3882) );
  XNOR U4542 ( .A(n3880), .B(n4344), .Z(n3881) );
  AND U4543 ( .A(n3076), .B(n775), .Z(n4344) );
  NAND U4544 ( .A(n853), .B(n2944), .Z(n4347) );
  XNOR U4545 ( .A(n4345), .B(n4349), .Z(n4346) );
  AND U4546 ( .A(n3076), .B(n814), .Z(n4349) );
  XNOR U4547 ( .A(n4341), .B(n4354), .Z(n4342) );
  AND U4548 ( .A(n744), .B(e_input[0]), .Z(n4354) );
  XNOR U4549 ( .A(n4340), .B(g_input[30]), .Z(n4338) );
  NOR U4550 ( .A(n4355), .B(n4356), .Z(n4340) );
  XOR U4551 ( .A(n4360), .B(n4343), .Z(n4353) );
  NAND U4552 ( .A(n775), .B(n4331), .Z(n4343) );
  IV U4553 ( .A(n4348), .Z(n4360) );
  NAND U4554 ( .A(n897), .B(n2944), .Z(n4352) );
  XNOR U4555 ( .A(n4350), .B(n4362), .Z(n4351) );
  AND U4556 ( .A(n3076), .B(n853), .Z(n4362) );
  XNOR U4557 ( .A(n4357), .B(n4367), .Z(n4358) );
  AND U4558 ( .A(n775), .B(e_input[0]), .Z(n4367) );
  XOR U4559 ( .A(n4355), .B(g_input[29]), .Z(n4356) );
  NANDN U4560 ( .B(n4368), .A(n4369), .Z(n4355) );
  XOR U4561 ( .A(n4373), .B(n4359), .Z(n4366) );
  NAND U4562 ( .A(n814), .B(n4331), .Z(n4359) );
  IV U4563 ( .A(n4361), .Z(n4373) );
  NAND U4564 ( .A(n941), .B(n2944), .Z(n4365) );
  XNOR U4565 ( .A(n4363), .B(n4375), .Z(n4364) );
  AND U4566 ( .A(n3076), .B(n897), .Z(n4375) );
  XNOR U4567 ( .A(n4370), .B(n4380), .Z(n4371) );
  AND U4568 ( .A(n814), .B(e_input[0]), .Z(n4380) );
  XNOR U4569 ( .A(n4369), .B(g_input[28]), .Z(n4368) );
  NOR U4570 ( .A(n4381), .B(n4382), .Z(n4369) );
  XOR U4571 ( .A(n4386), .B(n4372), .Z(n4379) );
  NAND U4572 ( .A(n853), .B(n4331), .Z(n4372) );
  IV U4573 ( .A(n4374), .Z(n4386) );
  NAND U4574 ( .A(n1001), .B(n2944), .Z(n4378) );
  XNOR U4575 ( .A(n4376), .B(n4388), .Z(n4377) );
  AND U4576 ( .A(n3076), .B(n941), .Z(n4388) );
  XNOR U4577 ( .A(n4383), .B(n4393), .Z(n4384) );
  AND U4578 ( .A(n853), .B(e_input[0]), .Z(n4393) );
  XOR U4579 ( .A(n4381), .B(g_input[27]), .Z(n4382) );
  NANDN U4580 ( .B(n4394), .A(n4395), .Z(n4381) );
  XOR U4581 ( .A(n4399), .B(n4385), .Z(n4392) );
  NAND U4582 ( .A(n897), .B(n4331), .Z(n4385) );
  IV U4583 ( .A(n4387), .Z(n4399) );
  NAND U4584 ( .A(n1055), .B(n2944), .Z(n4391) );
  XNOR U4585 ( .A(n4389), .B(n4401), .Z(n4390) );
  AND U4586 ( .A(n3076), .B(n1001), .Z(n4401) );
  XNOR U4587 ( .A(n4396), .B(n4406), .Z(n4397) );
  AND U4588 ( .A(n897), .B(e_input[0]), .Z(n4406) );
  XNOR U4589 ( .A(n4395), .B(g_input[26]), .Z(n4394) );
  NOR U4590 ( .A(n4407), .B(n4408), .Z(n4395) );
  XOR U4591 ( .A(n4412), .B(n4398), .Z(n4405) );
  NAND U4592 ( .A(n941), .B(n4331), .Z(n4398) );
  IV U4593 ( .A(n4400), .Z(n4412) );
  NAND U4594 ( .A(n1116), .B(n2944), .Z(n4404) );
  XNOR U4595 ( .A(n4402), .B(n4414), .Z(n4403) );
  AND U4596 ( .A(n3076), .B(n1055), .Z(n4414) );
  XNOR U4597 ( .A(n4409), .B(n4419), .Z(n4410) );
  AND U4598 ( .A(n941), .B(e_input[0]), .Z(n4419) );
  XOR U4599 ( .A(n4407), .B(g_input[25]), .Z(n4408) );
  NANDN U4600 ( .B(n4420), .A(n4421), .Z(n4407) );
  XOR U4601 ( .A(n4425), .B(n4411), .Z(n4418) );
  NAND U4602 ( .A(n1001), .B(n4331), .Z(n4411) );
  IV U4603 ( .A(n4413), .Z(n4425) );
  NAND U4604 ( .A(n1178), .B(n2944), .Z(n4417) );
  XNOR U4605 ( .A(n4415), .B(n4427), .Z(n4416) );
  AND U4606 ( .A(n3076), .B(n1116), .Z(n4427) );
  XNOR U4607 ( .A(n4422), .B(n4432), .Z(n4423) );
  AND U4608 ( .A(n1001), .B(e_input[0]), .Z(n4432) );
  XNOR U4609 ( .A(n4421), .B(g_input[24]), .Z(n4420) );
  NOR U4610 ( .A(n4433), .B(n4434), .Z(n4421) );
  XOR U4611 ( .A(n4438), .B(n4424), .Z(n4431) );
  NAND U4612 ( .A(n1055), .B(n4331), .Z(n4424) );
  IV U4613 ( .A(n4426), .Z(n4438) );
  NAND U4614 ( .A(n1246), .B(n2944), .Z(n4430) );
  XNOR U4615 ( .A(n4428), .B(n4440), .Z(n4429) );
  AND U4616 ( .A(n3076), .B(n1178), .Z(n4440) );
  XNOR U4617 ( .A(n4435), .B(n4445), .Z(n4436) );
  AND U4618 ( .A(n1055), .B(e_input[0]), .Z(n4445) );
  XOR U4619 ( .A(n4433), .B(g_input[23]), .Z(n4434) );
  NANDN U4620 ( .B(n4446), .A(n4447), .Z(n4433) );
  XOR U4621 ( .A(n4451), .B(n4437), .Z(n4444) );
  NAND U4622 ( .A(n1116), .B(n4331), .Z(n4437) );
  IV U4623 ( .A(n4439), .Z(n4451) );
  NAND U4624 ( .A(n1316), .B(n2944), .Z(n4443) );
  XNOR U4625 ( .A(n4441), .B(n4453), .Z(n4442) );
  AND U4626 ( .A(n3076), .B(n1246), .Z(n4453) );
  XNOR U4627 ( .A(n4448), .B(n4458), .Z(n4449) );
  AND U4628 ( .A(n1116), .B(e_input[0]), .Z(n4458) );
  XNOR U4629 ( .A(n4447), .B(g_input[22]), .Z(n4446) );
  NOR U4630 ( .A(n4459), .B(n4460), .Z(n4447) );
  XOR U4631 ( .A(n4464), .B(n4450), .Z(n4457) );
  NAND U4632 ( .A(n1178), .B(n4331), .Z(n4450) );
  IV U4633 ( .A(n4452), .Z(n4464) );
  NAND U4634 ( .A(n1390), .B(n2944), .Z(n4456) );
  XNOR U4635 ( .A(n4454), .B(n4466), .Z(n4455) );
  AND U4636 ( .A(n3076), .B(n1316), .Z(n4466) );
  XNOR U4637 ( .A(n4461), .B(n4471), .Z(n4462) );
  AND U4638 ( .A(n1178), .B(e_input[0]), .Z(n4471) );
  XOR U4639 ( .A(n4459), .B(g_input[21]), .Z(n4460) );
  NANDN U4640 ( .B(n4472), .A(n4473), .Z(n4459) );
  XOR U4641 ( .A(n4477), .B(n4463), .Z(n4470) );
  NAND U4642 ( .A(n1246), .B(n4331), .Z(n4463) );
  IV U4643 ( .A(n4465), .Z(n4477) );
  NAND U4644 ( .A(n1467), .B(n2944), .Z(n4469) );
  XNOR U4645 ( .A(n4467), .B(n4479), .Z(n4468) );
  AND U4646 ( .A(n3076), .B(n1390), .Z(n4479) );
  XNOR U4647 ( .A(n4474), .B(n4484), .Z(n4475) );
  AND U4648 ( .A(n1246), .B(e_input[0]), .Z(n4484) );
  XNOR U4649 ( .A(n4473), .B(g_input[20]), .Z(n4472) );
  NOR U4650 ( .A(n4485), .B(n4486), .Z(n4473) );
  XOR U4651 ( .A(n4490), .B(n4476), .Z(n4483) );
  NAND U4652 ( .A(n1316), .B(n4331), .Z(n4476) );
  IV U4653 ( .A(n4478), .Z(n4490) );
  NAND U4654 ( .A(n1554), .B(n2944), .Z(n4482) );
  XNOR U4655 ( .A(n4480), .B(n4492), .Z(n4481) );
  AND U4656 ( .A(n3076), .B(n1467), .Z(n4492) );
  XNOR U4657 ( .A(n4487), .B(n4497), .Z(n4488) );
  AND U4658 ( .A(n1316), .B(e_input[0]), .Z(n4497) );
  XOR U4659 ( .A(n4485), .B(g_input[19]), .Z(n4486) );
  NANDN U4660 ( .B(n4498), .A(n4499), .Z(n4485) );
  XOR U4661 ( .A(n4503), .B(n4489), .Z(n4496) );
  NAND U4662 ( .A(n1390), .B(n4331), .Z(n4489) );
  IV U4663 ( .A(n4491), .Z(n4503) );
  NAND U4664 ( .A(n1646), .B(n2944), .Z(n4495) );
  XNOR U4665 ( .A(n4493), .B(n4505), .Z(n4494) );
  AND U4666 ( .A(n3076), .B(n1554), .Z(n4505) );
  XNOR U4667 ( .A(n4500), .B(n4510), .Z(n4501) );
  AND U4668 ( .A(n1390), .B(e_input[0]), .Z(n4510) );
  XNOR U4669 ( .A(n4499), .B(g_input[18]), .Z(n4498) );
  NOR U4670 ( .A(n4511), .B(n4512), .Z(n4499) );
  XOR U4671 ( .A(n4516), .B(n4502), .Z(n4509) );
  NAND U4672 ( .A(n1467), .B(n4331), .Z(n4502) );
  IV U4673 ( .A(n4504), .Z(n4516) );
  NAND U4674 ( .A(n1737), .B(n2944), .Z(n4508) );
  XNOR U4675 ( .A(n4506), .B(n4518), .Z(n4507) );
  AND U4676 ( .A(n3076), .B(n1646), .Z(n4518) );
  XNOR U4677 ( .A(n4513), .B(n4523), .Z(n4514) );
  AND U4678 ( .A(n1467), .B(e_input[0]), .Z(n4523) );
  XOR U4679 ( .A(n4511), .B(g_input[17]), .Z(n4512) );
  NANDN U4680 ( .B(n4524), .A(n4525), .Z(n4511) );
  XOR U4681 ( .A(n4529), .B(n4515), .Z(n4522) );
  NAND U4682 ( .A(n1554), .B(n4331), .Z(n4515) );
  IV U4683 ( .A(n4517), .Z(n4529) );
  XOR U4684 ( .A(n4530), .B(n4531), .Z(n4517) );
  AND U4685 ( .A(n4141), .B(n4532), .Z(n4531) );
  XNOR U4686 ( .A(n4530), .B(n4140), .Z(n4532) );
  NAND U4687 ( .A(n1831), .B(n2944), .Z(n4521) );
  XNOR U4688 ( .A(n4519), .B(n4533), .Z(n4520) );
  AND U4689 ( .A(n3076), .B(n1737), .Z(n4533) );
  XNOR U4690 ( .A(n4526), .B(n4538), .Z(n4527) );
  AND U4691 ( .A(n1554), .B(e_input[0]), .Z(n4538) );
  XOR U4692 ( .A(n4542), .B(n4528), .Z(n4537) );
  NAND U4693 ( .A(n1646), .B(n4331), .Z(n4528) );
  IV U4694 ( .A(n4530), .Z(n4542) );
  NAND U4695 ( .A(n1931), .B(n2944), .Z(n4536) );
  XNOR U4696 ( .A(n4534), .B(n4544), .Z(n4535) );
  AND U4697 ( .A(n3076), .B(n1831), .Z(n4544) );
  XNOR U4698 ( .A(n4539), .B(n4549), .Z(n4540) );
  AND U4699 ( .A(n1646), .B(e_input[0]), .Z(n4549) );
  XOR U4700 ( .A(n4553), .B(n4541), .Z(n4548) );
  NAND U4701 ( .A(n1737), .B(n4331), .Z(n4541) );
  IV U4702 ( .A(n4543), .Z(n4553) );
  NAND U4703 ( .A(n2036), .B(n2944), .Z(n4547) );
  XNOR U4704 ( .A(n4545), .B(n4555), .Z(n4546) );
  AND U4705 ( .A(n3076), .B(n1931), .Z(n4555) );
  XNOR U4706 ( .A(n4550), .B(n4560), .Z(n4551) );
  AND U4707 ( .A(n1737), .B(e_input[0]), .Z(n4560) );
  XOR U4708 ( .A(n4564), .B(n4552), .Z(n4559) );
  NAND U4709 ( .A(n1831), .B(n4331), .Z(n4552) );
  IV U4710 ( .A(n4554), .Z(n4564) );
  NAND U4711 ( .A(n2141), .B(n2944), .Z(n4558) );
  XNOR U4712 ( .A(n4556), .B(n4566), .Z(n4557) );
  AND U4713 ( .A(n3076), .B(n2036), .Z(n4566) );
  XNOR U4714 ( .A(n4561), .B(n4571), .Z(n4562) );
  AND U4715 ( .A(n1831), .B(e_input[0]), .Z(n4571) );
  XOR U4716 ( .A(n4575), .B(n4563), .Z(n4570) );
  NAND U4717 ( .A(n1931), .B(n4331), .Z(n4563) );
  IV U4718 ( .A(n4565), .Z(n4575) );
  NAND U4719 ( .A(n2254), .B(n2944), .Z(n4569) );
  XNOR U4720 ( .A(n4567), .B(n4577), .Z(n4568) );
  AND U4721 ( .A(n3076), .B(n2141), .Z(n4577) );
  XNOR U4722 ( .A(n4572), .B(n4582), .Z(n4573) );
  AND U4723 ( .A(n1931), .B(e_input[0]), .Z(n4582) );
  XOR U4724 ( .A(n4586), .B(n4574), .Z(n4581) );
  NAND U4725 ( .A(n2036), .B(n4331), .Z(n4574) );
  IV U4726 ( .A(n4576), .Z(n4586) );
  NAND U4727 ( .A(n2370), .B(n2944), .Z(n4580) );
  XNOR U4728 ( .A(n4578), .B(n4588), .Z(n4579) );
  AND U4729 ( .A(n3076), .B(n2254), .Z(n4588) );
  XNOR U4730 ( .A(n4583), .B(n4593), .Z(n4584) );
  AND U4731 ( .A(n2036), .B(e_input[0]), .Z(n4593) );
  XOR U4732 ( .A(n4597), .B(n4585), .Z(n4592) );
  NAND U4733 ( .A(n2141), .B(n4331), .Z(n4585) );
  IV U4734 ( .A(n4587), .Z(n4597) );
  NAND U4735 ( .A(n2491), .B(n2944), .Z(n4591) );
  XNOR U4736 ( .A(n4589), .B(n4599), .Z(n4590) );
  AND U4737 ( .A(n3076), .B(n2370), .Z(n4599) );
  XNOR U4738 ( .A(n4594), .B(n4604), .Z(n4595) );
  AND U4739 ( .A(n2141), .B(e_input[0]), .Z(n4604) );
  XOR U4740 ( .A(n4608), .B(n4596), .Z(n4603) );
  NAND U4741 ( .A(n2254), .B(n4331), .Z(n4596) );
  IV U4742 ( .A(n4598), .Z(n4608) );
  NAND U4743 ( .A(n2615), .B(n2944), .Z(n4602) );
  XNOR U4744 ( .A(n4600), .B(n4610), .Z(n4601) );
  AND U4745 ( .A(n3076), .B(n2491), .Z(n4610) );
  XNOR U4746 ( .A(n4605), .B(n4615), .Z(n4606) );
  AND U4747 ( .A(n2254), .B(e_input[0]), .Z(n4615) );
  XOR U4748 ( .A(n4619), .B(n4607), .Z(n4614) );
  NAND U4749 ( .A(n2370), .B(n4331), .Z(n4607) );
  IV U4750 ( .A(n4609), .Z(n4619) );
  NAND U4751 ( .A(n2743), .B(n2944), .Z(n4613) );
  XNOR U4752 ( .A(n4611), .B(n4621), .Z(n4612) );
  AND U4753 ( .A(n3076), .B(n2615), .Z(n4621) );
  XNOR U4754 ( .A(n4625), .B(n4622), .Z(n4624) );
  XNOR U4755 ( .A(n4616), .B(n4627), .Z(n4617) );
  AND U4756 ( .A(n2370), .B(e_input[0]), .Z(n4627) );
  XNOR U4757 ( .A(n4631), .B(n4628), .Z(n4630) );
  XOR U4758 ( .A(n4632), .B(n4618), .Z(n4626) );
  NAND U4759 ( .A(n2491), .B(n4331), .Z(n4618) );
  IV U4760 ( .A(n4620), .Z(n4632) );
  XNOR U4761 ( .A(n4633), .B(n4634), .Z(n4620) );
  AND U4762 ( .A(n4635), .B(n4636), .Z(n4634) );
  XOR U4763 ( .A(n4629), .B(n4637), .Z(n4636) );
  XNOR U4764 ( .A(n4631), .B(n4633), .Z(n4637) );
  NAND U4765 ( .A(n2615), .B(n4331), .Z(n4631) );
  XOR U4766 ( .A(n4628), .B(n4638), .Z(n4629) );
  AND U4767 ( .A(n2491), .B(e_input[0]), .Z(n4638) );
  XNOR U4768 ( .A(n4642), .B(n4639), .Z(n4641) );
  XOR U4769 ( .A(n4623), .B(n4643), .Z(n4635) );
  XNOR U4770 ( .A(n4625), .B(n4633), .Z(n4643) );
  NANDN U4771 ( .B(n2872), .A(n2944), .Z(n4625) );
  XOR U4772 ( .A(n4622), .B(n4644), .Z(n4623) );
  AND U4773 ( .A(n3076), .B(n2743), .Z(n4644) );
  XNOR U4774 ( .A(n4648), .B(n4645), .Z(n4647) );
  XOR U4775 ( .A(n4649), .B(n4650), .Z(n4633) );
  AND U4776 ( .A(n4651), .B(n4652), .Z(n4650) );
  XOR U4777 ( .A(n4640), .B(n4653), .Z(n4652) );
  XNOR U4778 ( .A(n4642), .B(n4649), .Z(n4653) );
  NAND U4779 ( .A(n2743), .B(n4331), .Z(n4642) );
  XOR U4780 ( .A(n4639), .B(n4654), .Z(n4640) );
  AND U4781 ( .A(n2615), .B(e_input[0]), .Z(n4654) );
  XNOR U4782 ( .A(n4658), .B(n4655), .Z(n4657) );
  XOR U4783 ( .A(n4646), .B(n4659), .Z(n4651) );
  XNOR U4784 ( .A(n4648), .B(n4649), .Z(n4659) );
  NANDN U4785 ( .B(n3010), .A(n2944), .Z(n4648) );
  XOR U4786 ( .A(n4645), .B(n4660), .Z(n4646) );
  ANDN U4787 ( .A(n3076), .B(n2872), .Z(n4660) );
  XNOR U4788 ( .A(n4664), .B(n4661), .Z(n4663) );
  XOR U4789 ( .A(n4665), .B(n4666), .Z(n4649) );
  AND U4790 ( .A(n4667), .B(n4668), .Z(n4666) );
  XOR U4791 ( .A(n4656), .B(n4669), .Z(n4668) );
  XNOR U4792 ( .A(n4658), .B(n4665), .Z(n4669) );
  NANDN U4793 ( .B(n2872), .A(n4331), .Z(n4658) );
  XOR U4794 ( .A(n4655), .B(n4670), .Z(n4656) );
  AND U4795 ( .A(n2743), .B(e_input[0]), .Z(n4670) );
  XOR U4796 ( .A(n4662), .B(n4674), .Z(n4667) );
  XNOR U4797 ( .A(n4664), .B(n4665), .Z(n4674) );
  NAND U4798 ( .A(n2944), .B(n3146), .Z(n4664) );
  XOR U4799 ( .A(n4661), .B(n4675), .Z(n4662) );
  ANDN U4800 ( .A(n3076), .B(n3010), .Z(n4675) );
  NAND U4801 ( .A(n2944), .B(n3835), .Z(n4678) );
  XNOR U4802 ( .A(n4676), .B(n4680), .Z(n4677) );
  AND U4803 ( .A(n3146), .B(n3076), .Z(n4680) );
  AND U4804 ( .A(n4681), .B(g_input[0]), .Z(n4676) );
  NANDN U4805 ( .B(n2944), .A(n4682), .Z(n4681) );
  NAND U4806 ( .A(n3835), .B(n3076), .Z(n4682) );
  XNOR U4807 ( .A(n4671), .B(n4686), .Z(n4672) );
  ANDN U4808 ( .A(e_input[0]), .B(n2872), .Z(n4686) );
  XOR U4809 ( .A(n4689), .B(n4687), .Z(n4688) );
  ANDN U4810 ( .A(e_input[0]), .B(n3010), .Z(n4689) );
  AND U4811 ( .A(n4331), .B(n3146), .Z(n4690) );
  XOR U4812 ( .A(n4694), .B(n4673), .Z(n4685) );
  NANDN U4813 ( .B(n3010), .A(n4331), .Z(n4673) );
  IV U4814 ( .A(n4679), .Z(n4694) );
  NAND U4815 ( .A(n4331), .B(n3835), .Z(n4693) );
  XNOR U4816 ( .A(n4691), .B(n4695), .Z(n4692) );
  AND U4817 ( .A(n3146), .B(e_input[0]), .Z(n4695) );
  AND U4818 ( .A(n4696), .B(g_input[0]), .Z(n4691) );
  NANDN U4819 ( .B(n4331), .A(n4697), .Z(n4696) );
  NAND U4820 ( .A(n3835), .B(e_input[0]), .Z(n4697) );
  XNOR U4821 ( .A(n4699), .B(n3110), .Z(n3101) );
  XNOR U4822 ( .A(n3089), .B(n4701), .Z(n3090) );
  AND U4823 ( .A(n1931), .B(n1196), .Z(n4701) );
  XOR U4824 ( .A(n4705), .B(n3091), .Z(n4700) );
  NAND U4825 ( .A(n1138), .B(n2036), .Z(n3091) );
  IV U4826 ( .A(n3093), .Z(n4705) );
  XNOR U4827 ( .A(n3098), .B(n3099), .Z(n3095) );
  NANDN U4828 ( .B(n1020), .A(n2254), .Z(n3099) );
  XNOR U4829 ( .A(n3097), .B(n4709), .Z(n3098) );
  AND U4830 ( .A(n2141), .B(n1079), .Z(n4709) );
  XNOR U4831 ( .A(n3109), .B(n3100), .Z(n4699) );
  XOR U4832 ( .A(n4713), .B(n4714), .Z(n3100) );
  XOR U4833 ( .A(n4715), .B(n3119), .Z(n3109) );
  XNOR U4834 ( .A(n3106), .B(n3107), .Z(n3119) );
  NAND U4835 ( .A(n1284), .B(n1831), .Z(n3107) );
  XNOR U4836 ( .A(n3105), .B(n4716), .Z(n3106) );
  AND U4837 ( .A(n1737), .B(n1352), .Z(n4716) );
  XNOR U4838 ( .A(n3118), .B(n3108), .Z(n4715) );
  XOR U4839 ( .A(n4720), .B(n4721), .Z(n3108) );
  AND U4840 ( .A(n4722), .B(n4723), .Z(n4721) );
  XOR U4841 ( .A(n4724), .B(n4725), .Z(n4723) );
  XOR U4842 ( .A(n4720), .B(n4726), .Z(n4725) );
  XOR U4843 ( .A(n4707), .B(n4727), .Z(n4722) );
  XOR U4844 ( .A(n4720), .B(n4708), .Z(n4727) );
  NANDN U4845 ( .B(n1020), .A(n2370), .Z(n4712) );
  XNOR U4846 ( .A(n4710), .B(n4728), .Z(n4711) );
  AND U4847 ( .A(n2254), .B(n1079), .Z(n4728) );
  XNOR U4848 ( .A(n4702), .B(n4733), .Z(n4703) );
  AND U4849 ( .A(n2036), .B(n1196), .Z(n4733) );
  XOR U4850 ( .A(n4737), .B(n4704), .Z(n4732) );
  NAND U4851 ( .A(n1138), .B(n2141), .Z(n4704) );
  IV U4852 ( .A(n4706), .Z(n4737) );
  XOR U4853 ( .A(n4741), .B(n4742), .Z(n4720) );
  AND U4854 ( .A(n4743), .B(n4744), .Z(n4742) );
  XOR U4855 ( .A(n4745), .B(n4746), .Z(n4744) );
  XOR U4856 ( .A(n4741), .B(n4747), .Z(n4746) );
  XOR U4857 ( .A(n4739), .B(n4748), .Z(n4743) );
  XOR U4858 ( .A(n4741), .B(n4740), .Z(n4748) );
  NANDN U4859 ( .B(n1020), .A(n2491), .Z(n4731) );
  XNOR U4860 ( .A(n4729), .B(n4749), .Z(n4730) );
  AND U4861 ( .A(n2370), .B(n1079), .Z(n4749) );
  XNOR U4862 ( .A(n4734), .B(n4754), .Z(n4735) );
  AND U4863 ( .A(n2141), .B(n1196), .Z(n4754) );
  XOR U4864 ( .A(n4758), .B(n4736), .Z(n4753) );
  NAND U4865 ( .A(n1138), .B(n2254), .Z(n4736) );
  IV U4866 ( .A(n4738), .Z(n4758) );
  XOR U4867 ( .A(n4762), .B(n4763), .Z(n4741) );
  AND U4868 ( .A(n4764), .B(n4765), .Z(n4763) );
  XOR U4869 ( .A(n4766), .B(n4767), .Z(n4765) );
  XOR U4870 ( .A(n4762), .B(n4768), .Z(n4767) );
  XOR U4871 ( .A(n4760), .B(n4769), .Z(n4764) );
  XOR U4872 ( .A(n4762), .B(n4761), .Z(n4769) );
  NANDN U4873 ( .B(n1020), .A(n2615), .Z(n4752) );
  XNOR U4874 ( .A(n4750), .B(n4770), .Z(n4751) );
  AND U4875 ( .A(n2491), .B(n1079), .Z(n4770) );
  XNOR U4876 ( .A(n4755), .B(n4775), .Z(n4756) );
  AND U4877 ( .A(n2254), .B(n1196), .Z(n4775) );
  XOR U4878 ( .A(n4779), .B(n4757), .Z(n4774) );
  NAND U4879 ( .A(n1138), .B(n2370), .Z(n4757) );
  IV U4880 ( .A(n4759), .Z(n4779) );
  XOR U4881 ( .A(n4783), .B(n4784), .Z(n4762) );
  AND U4882 ( .A(n4785), .B(n4786), .Z(n4784) );
  XOR U4883 ( .A(n4787), .B(n4788), .Z(n4786) );
  XOR U4884 ( .A(n4783), .B(n4789), .Z(n4788) );
  XOR U4885 ( .A(n4781), .B(n4790), .Z(n4785) );
  XOR U4886 ( .A(n4783), .B(n4782), .Z(n4790) );
  NANDN U4887 ( .B(n1020), .A(n2743), .Z(n4773) );
  XNOR U4888 ( .A(n4771), .B(n4791), .Z(n4772) );
  AND U4889 ( .A(n2615), .B(n1079), .Z(n4791) );
  XNOR U4890 ( .A(n4776), .B(n4796), .Z(n4777) );
  AND U4891 ( .A(n2370), .B(n1196), .Z(n4796) );
  XOR U4892 ( .A(n4800), .B(n4778), .Z(n4795) );
  NAND U4893 ( .A(n1138), .B(n2491), .Z(n4778) );
  IV U4894 ( .A(n4780), .Z(n4800) );
  XOR U4895 ( .A(n4804), .B(n4805), .Z(n4783) );
  AND U4896 ( .A(n4806), .B(n4807), .Z(n4805) );
  XOR U4897 ( .A(n4808), .B(n4809), .Z(n4807) );
  XOR U4898 ( .A(n4804), .B(n4810), .Z(n4809) );
  XOR U4899 ( .A(n4802), .B(n4811), .Z(n4806) );
  XOR U4900 ( .A(n4804), .B(n4803), .Z(n4811) );
  OR U4901 ( .A(n1020), .B(n2872), .Z(n4794) );
  XNOR U4902 ( .A(n4792), .B(n4812), .Z(n4793) );
  AND U4903 ( .A(n2743), .B(n1079), .Z(n4812) );
  XNOR U4904 ( .A(n4797), .B(n4817), .Z(n4798) );
  AND U4905 ( .A(n2491), .B(n1196), .Z(n4817) );
  XOR U4906 ( .A(n4821), .B(n4799), .Z(n4816) );
  NAND U4907 ( .A(n1138), .B(n2615), .Z(n4799) );
  IV U4908 ( .A(n4801), .Z(n4821) );
  XOR U4909 ( .A(n4825), .B(n4826), .Z(n4804) );
  AND U4910 ( .A(n4827), .B(n4828), .Z(n4826) );
  XOR U4911 ( .A(n4829), .B(n4830), .Z(n4828) );
  XOR U4912 ( .A(n4825), .B(n4831), .Z(n4830) );
  XOR U4913 ( .A(n4823), .B(n4832), .Z(n4827) );
  XOR U4914 ( .A(n4825), .B(n4824), .Z(n4832) );
  OR U4915 ( .A(n1020), .B(n3010), .Z(n4815) );
  XNOR U4916 ( .A(n4813), .B(n4833), .Z(n4814) );
  ANDN U4917 ( .A(n1079), .B(n2872), .Z(n4833) );
  XNOR U4918 ( .A(n4818), .B(n4838), .Z(n4819) );
  AND U4919 ( .A(n2615), .B(n1196), .Z(n4838) );
  XOR U4920 ( .A(n4842), .B(n4820), .Z(n4837) );
  NAND U4921 ( .A(n1138), .B(n2743), .Z(n4820) );
  IV U4922 ( .A(n4822), .Z(n4842) );
  XOR U4923 ( .A(n4846), .B(n4847), .Z(n4825) );
  AND U4924 ( .A(n4848), .B(n4849), .Z(n4847) );
  XOR U4925 ( .A(n4850), .B(n4851), .Z(n4849) );
  XOR U4926 ( .A(n4846), .B(n4852), .Z(n4851) );
  XOR U4927 ( .A(n4844), .B(n4853), .Z(n4848) );
  XOR U4928 ( .A(n4846), .B(n4845), .Z(n4853) );
  NANDN U4929 ( .B(n1020), .A(n3146), .Z(n4836) );
  XNOR U4930 ( .A(n4834), .B(n4854), .Z(n4835) );
  ANDN U4931 ( .A(n1079), .B(n3010), .Z(n4854) );
  XNOR U4932 ( .A(n4839), .B(n4859), .Z(n4840) );
  AND U4933 ( .A(n2743), .B(n1196), .Z(n4859) );
  XOR U4934 ( .A(n4863), .B(n4841), .Z(n4858) );
  NANDN U4935 ( .B(n2872), .A(n1138), .Z(n4841) );
  IV U4936 ( .A(n4843), .Z(n4863) );
  XOR U4937 ( .A(n4868), .B(n4869), .Z(n4714) );
  XNOR U4938 ( .A(n4870), .B(n4867), .Z(n4868) );
  XNOR U4939 ( .A(n4860), .B(n4872), .Z(n4861) );
  ANDN U4940 ( .A(n1196), .B(n2872), .Z(n4872) );
  XOR U4941 ( .A(n4875), .B(n4873), .Z(n4874) );
  ANDN U4942 ( .A(n1196), .B(n3010), .Z(n4875) );
  AND U4943 ( .A(n3146), .B(n1138), .Z(n4876) );
  XOR U4944 ( .A(n4880), .B(n4862), .Z(n4871) );
  NANDN U4945 ( .B(n3010), .A(n1138), .Z(n4862) );
  IV U4946 ( .A(n4864), .Z(n4880) );
  NAND U4947 ( .A(n1138), .B(n3835), .Z(n4879) );
  XNOR U4948 ( .A(n4877), .B(n4881), .Z(n4878) );
  AND U4949 ( .A(n3146), .B(n1196), .Z(n4881) );
  AND U4950 ( .A(n4882), .B(g_input[0]), .Z(n4877) );
  NANDN U4951 ( .B(n1138), .A(n4883), .Z(n4882) );
  NAND U4952 ( .A(n3835), .B(n1196), .Z(n4883) );
  XNOR U4953 ( .A(n4856), .B(n4857), .Z(n4866) );
  NANDN U4954 ( .B(n1020), .A(n3835), .Z(n4857) );
  XNOR U4955 ( .A(n4855), .B(n4886), .Z(n4856) );
  AND U4956 ( .A(n3146), .B(n1079), .Z(n4886) );
  AND U4957 ( .A(n4887), .B(g_input[0]), .Z(n4855) );
  NAND U4958 ( .A(n4888), .B(n1020), .Z(n4887) );
  NAND U4959 ( .A(n3835), .B(n1079), .Z(n4888) );
  XOR U4960 ( .A(n4891), .B(n4892), .Z(n4867) );
  XNOR U4961 ( .A(n3113), .B(n4894), .Z(n3114) );
  AND U4962 ( .A(n1554), .B(n1522), .Z(n4894) );
  XNOR U4963 ( .A(n4525), .B(g_input[16]), .Z(n4524) );
  NOR U4964 ( .A(n4895), .B(n4896), .Z(n4525) );
  XOR U4965 ( .A(n4900), .B(n3115), .Z(n4893) );
  NAND U4966 ( .A(n1435), .B(n1646), .Z(n3115) );
  IV U4967 ( .A(n3117), .Z(n4900) );
  NAND U4968 ( .A(n1284), .B(n1931), .Z(n4719) );
  XNOR U4969 ( .A(n4717), .B(n4902), .Z(n4718) );
  AND U4970 ( .A(n1831), .B(n1352), .Z(n4902) );
  XNOR U4971 ( .A(n4897), .B(n4907), .Z(n4898) );
  AND U4972 ( .A(n1646), .B(n1522), .Z(n4907) );
  XOR U4973 ( .A(n4895), .B(g_input[15]), .Z(n4896) );
  NANDN U4974 ( .B(n4908), .A(n4909), .Z(n4895) );
  XOR U4975 ( .A(n4913), .B(n4899), .Z(n4906) );
  NAND U4976 ( .A(n1435), .B(n1737), .Z(n4899) );
  IV U4977 ( .A(n4901), .Z(n4913) );
  NAND U4978 ( .A(n1284), .B(n2036), .Z(n4905) );
  XNOR U4979 ( .A(n4903), .B(n4915), .Z(n4904) );
  AND U4980 ( .A(n1931), .B(n1352), .Z(n4915) );
  XNOR U4981 ( .A(n4910), .B(n4920), .Z(n4911) );
  AND U4982 ( .A(n1737), .B(n1522), .Z(n4920) );
  XNOR U4983 ( .A(n4909), .B(g_input[14]), .Z(n4908) );
  NOR U4984 ( .A(n4921), .B(n4922), .Z(n4909) );
  XOR U4985 ( .A(n4926), .B(n4912), .Z(n4919) );
  NAND U4986 ( .A(n1435), .B(n1831), .Z(n4912) );
  IV U4987 ( .A(n4914), .Z(n4926) );
  NAND U4988 ( .A(n1284), .B(n2141), .Z(n4918) );
  XNOR U4989 ( .A(n4916), .B(n4928), .Z(n4917) );
  AND U4990 ( .A(n2036), .B(n1352), .Z(n4928) );
  XNOR U4991 ( .A(n4923), .B(n4933), .Z(n4924) );
  AND U4992 ( .A(n1831), .B(n1522), .Z(n4933) );
  XOR U4993 ( .A(n4921), .B(g_input[13]), .Z(n4922) );
  NANDN U4994 ( .B(n4934), .A(n4935), .Z(n4921) );
  XOR U4995 ( .A(n4939), .B(n4925), .Z(n4932) );
  NAND U4996 ( .A(n1435), .B(n1931), .Z(n4925) );
  IV U4997 ( .A(n4927), .Z(n4939) );
  NAND U4998 ( .A(n1284), .B(n2254), .Z(n4931) );
  XNOR U4999 ( .A(n4929), .B(n4941), .Z(n4930) );
  AND U5000 ( .A(n2141), .B(n1352), .Z(n4941) );
  XNOR U5001 ( .A(n4936), .B(n4946), .Z(n4937) );
  AND U5002 ( .A(n1931), .B(n1522), .Z(n4946) );
  XNOR U5003 ( .A(n4935), .B(g_input[12]), .Z(n4934) );
  NOR U5004 ( .A(n4947), .B(n4948), .Z(n4935) );
  XOR U5005 ( .A(n4952), .B(n4938), .Z(n4945) );
  NAND U5006 ( .A(n1435), .B(n2036), .Z(n4938) );
  IV U5007 ( .A(n4940), .Z(n4952) );
  NAND U5008 ( .A(n1284), .B(n2370), .Z(n4944) );
  XNOR U5009 ( .A(n4942), .B(n4954), .Z(n4943) );
  AND U5010 ( .A(n2254), .B(n1352), .Z(n4954) );
  XNOR U5011 ( .A(n4949), .B(n4959), .Z(n4950) );
  AND U5012 ( .A(n2036), .B(n1522), .Z(n4959) );
  XOR U5013 ( .A(n4947), .B(g_input[11]), .Z(n4948) );
  NANDN U5014 ( .B(n4960), .A(n4961), .Z(n4947) );
  XOR U5015 ( .A(n4965), .B(n4951), .Z(n4958) );
  NAND U5016 ( .A(n1435), .B(n2141), .Z(n4951) );
  IV U5017 ( .A(n4953), .Z(n4965) );
  NAND U5018 ( .A(n1284), .B(n2491), .Z(n4957) );
  XNOR U5019 ( .A(n4955), .B(n4967), .Z(n4956) );
  AND U5020 ( .A(n2370), .B(n1352), .Z(n4967) );
  XNOR U5021 ( .A(n4962), .B(n4972), .Z(n4963) );
  AND U5022 ( .A(n2141), .B(n1522), .Z(n4972) );
  XNOR U5023 ( .A(n4961), .B(g_input[10]), .Z(n4960) );
  NOR U5024 ( .A(n4973), .B(n4974), .Z(n4961) );
  XOR U5025 ( .A(n4978), .B(n4964), .Z(n4971) );
  NAND U5026 ( .A(n1435), .B(n2254), .Z(n4964) );
  IV U5027 ( .A(n4966), .Z(n4978) );
  NAND U5028 ( .A(n1284), .B(n2615), .Z(n4970) );
  XNOR U5029 ( .A(n4968), .B(n4980), .Z(n4969) );
  AND U5030 ( .A(n2491), .B(n1352), .Z(n4980) );
  XNOR U5031 ( .A(n4975), .B(n4985), .Z(n4976) );
  AND U5032 ( .A(n2254), .B(n1522), .Z(n4985) );
  XOR U5033 ( .A(n4973), .B(g_input[9]), .Z(n4974) );
  NANDN U5034 ( .B(n4986), .A(n4987), .Z(n4973) );
  XOR U5035 ( .A(n4991), .B(n4977), .Z(n4984) );
  NAND U5036 ( .A(n1435), .B(n2370), .Z(n4977) );
  IV U5037 ( .A(n4979), .Z(n4991) );
  NAND U5038 ( .A(n1284), .B(n2743), .Z(n4983) );
  XNOR U5039 ( .A(n4981), .B(n4993), .Z(n4982) );
  AND U5040 ( .A(n2615), .B(n1352), .Z(n4993) );
  XNOR U5041 ( .A(n4997), .B(n4994), .Z(n4996) );
  XNOR U5042 ( .A(n4988), .B(n4999), .Z(n4989) );
  AND U5043 ( .A(n2370), .B(n1522), .Z(n4999) );
  XNOR U5044 ( .A(n5003), .B(n5000), .Z(n5002) );
  XOR U5045 ( .A(n5004), .B(n4990), .Z(n4998) );
  NAND U5046 ( .A(n1435), .B(n2491), .Z(n4990) );
  IV U5047 ( .A(n4992), .Z(n5004) );
  XNOR U5048 ( .A(n5005), .B(n5006), .Z(n4992) );
  AND U5049 ( .A(n5007), .B(n5008), .Z(n5006) );
  XOR U5050 ( .A(n5001), .B(n5009), .Z(n5008) );
  XNOR U5051 ( .A(n5003), .B(n5005), .Z(n5009) );
  NAND U5052 ( .A(n1435), .B(n2615), .Z(n5003) );
  XOR U5053 ( .A(n5000), .B(n5010), .Z(n5001) );
  AND U5054 ( .A(n2491), .B(n1522), .Z(n5010) );
  XNOR U5055 ( .A(n5014), .B(n5011), .Z(n5013) );
  XOR U5056 ( .A(n4995), .B(n5015), .Z(n5007) );
  XNOR U5057 ( .A(n4997), .B(n5005), .Z(n5015) );
  NANDN U5058 ( .B(n2872), .A(n1284), .Z(n4997) );
  XOR U5059 ( .A(n4994), .B(n5016), .Z(n4995) );
  AND U5060 ( .A(n2743), .B(n1352), .Z(n5016) );
  XNOR U5061 ( .A(n5020), .B(n5017), .Z(n5019) );
  XOR U5062 ( .A(n5021), .B(n5022), .Z(n5005) );
  AND U5063 ( .A(n5023), .B(n5024), .Z(n5022) );
  XOR U5064 ( .A(n5012), .B(n5025), .Z(n5024) );
  XNOR U5065 ( .A(n5014), .B(n5021), .Z(n5025) );
  NAND U5066 ( .A(n1435), .B(n2743), .Z(n5014) );
  XOR U5067 ( .A(n5011), .B(n5026), .Z(n5012) );
  AND U5068 ( .A(n2615), .B(n1522), .Z(n5026) );
  XNOR U5069 ( .A(n5030), .B(n5027), .Z(n5029) );
  XOR U5070 ( .A(n5018), .B(n5031), .Z(n5023) );
  XNOR U5071 ( .A(n5020), .B(n5021), .Z(n5031) );
  NANDN U5072 ( .B(n3010), .A(n1284), .Z(n5020) );
  XOR U5073 ( .A(n5017), .B(n5032), .Z(n5018) );
  ANDN U5074 ( .A(n1352), .B(n2872), .Z(n5032) );
  XNOR U5075 ( .A(n5036), .B(n5033), .Z(n5035) );
  XOR U5076 ( .A(n5037), .B(n5038), .Z(n5021) );
  AND U5077 ( .A(n5039), .B(n5040), .Z(n5038) );
  XOR U5078 ( .A(n5028), .B(n5041), .Z(n5040) );
  XNOR U5079 ( .A(n5030), .B(n5037), .Z(n5041) );
  NANDN U5080 ( .B(n2872), .A(n1435), .Z(n5030) );
  XOR U5081 ( .A(n5027), .B(n5042), .Z(n5028) );
  AND U5082 ( .A(n2743), .B(n1522), .Z(n5042) );
  XOR U5083 ( .A(n5034), .B(n5046), .Z(n5039) );
  XNOR U5084 ( .A(n5036), .B(n5037), .Z(n5046) );
  NAND U5085 ( .A(n1284), .B(n3146), .Z(n5036) );
  XOR U5086 ( .A(n5033), .B(n5047), .Z(n5034) );
  ANDN U5087 ( .A(n1352), .B(n3010), .Z(n5047) );
  NAND U5088 ( .A(n1284), .B(n3835), .Z(n5050) );
  XNOR U5089 ( .A(n5048), .B(n5052), .Z(n5049) );
  AND U5090 ( .A(n3146), .B(n1352), .Z(n5052) );
  AND U5091 ( .A(n5053), .B(g_input[0]), .Z(n5048) );
  NANDN U5092 ( .B(n1284), .A(n5054), .Z(n5053) );
  NAND U5093 ( .A(n3835), .B(n1352), .Z(n5054) );
  XNOR U5094 ( .A(n5043), .B(n5058), .Z(n5044) );
  ANDN U5095 ( .A(n1522), .B(n2872), .Z(n5058) );
  XOR U5096 ( .A(n5061), .B(n5059), .Z(n5060) );
  ANDN U5097 ( .A(n1522), .B(n3010), .Z(n5061) );
  AND U5098 ( .A(n3146), .B(n1435), .Z(n5062) );
  XOR U5099 ( .A(n5066), .B(n5045), .Z(n5057) );
  NANDN U5100 ( .B(n3010), .A(n1435), .Z(n5045) );
  IV U5101 ( .A(n5051), .Z(n5066) );
  NAND U5102 ( .A(n1435), .B(n3835), .Z(n5065) );
  XNOR U5103 ( .A(n5063), .B(n5067), .Z(n5064) );
  AND U5104 ( .A(n3146), .B(n1522), .Z(n5067) );
  AND U5105 ( .A(n5068), .B(g_input[0]), .Z(n5063) );
  NANDN U5106 ( .B(n1435), .A(n5069), .Z(n5068) );
  NAND U5107 ( .A(n3835), .B(n1522), .Z(n5069) );
  XNOR U5108 ( .A(n5072), .B(n3136), .Z(n3126) );
  XNOR U5109 ( .A(n3123), .B(n3124), .Z(n3136) );
  NANDN U5110 ( .B(n834), .A(n2743), .Z(n3124) );
  XNOR U5111 ( .A(n3122), .B(n5073), .Z(n3123) );
  AND U5112 ( .A(n2615), .B(n872), .Z(n5073) );
  XNOR U5113 ( .A(n5077), .B(n5074), .Z(n5076) );
  XNOR U5114 ( .A(n3135), .B(n3125), .Z(n5072) );
  XOR U5115 ( .A(n5078), .B(n5079), .Z(n3125) );
  XNOR U5116 ( .A(n3130), .B(n5081), .Z(n3131) );
  AND U5117 ( .A(n2370), .B(n984), .Z(n5081) );
  XNOR U5118 ( .A(n4987), .B(g_input[8]), .Z(n4986) );
  NOR U5119 ( .A(n5082), .B(n5083), .Z(n4987) );
  XNOR U5120 ( .A(n5087), .B(n5084), .Z(n5086) );
  XOR U5121 ( .A(n5088), .B(n3132), .Z(n5080) );
  NAND U5122 ( .A(n928), .B(n2491), .Z(n3132) );
  IV U5123 ( .A(n3134), .Z(n5088) );
  XNOR U5124 ( .A(n5089), .B(n5090), .Z(n3134) );
  AND U5125 ( .A(n5091), .B(n5092), .Z(n5090) );
  XOR U5126 ( .A(n5085), .B(n5093), .Z(n5092) );
  XNOR U5127 ( .A(n5087), .B(n5089), .Z(n5093) );
  NAND U5128 ( .A(n928), .B(n2615), .Z(n5087) );
  XOR U5129 ( .A(n5084), .B(n5094), .Z(n5085) );
  AND U5130 ( .A(n2491), .B(n984), .Z(n5094) );
  XOR U5131 ( .A(n5082), .B(g_input[7]), .Z(n5083) );
  NANDN U5132 ( .B(n5095), .A(n5096), .Z(n5082) );
  XNOR U5133 ( .A(n5100), .B(n5097), .Z(n5099) );
  XOR U5134 ( .A(n5075), .B(n5101), .Z(n5091) );
  XNOR U5135 ( .A(n5077), .B(n5089), .Z(n5101) );
  OR U5136 ( .A(n834), .B(n2872), .Z(n5077) );
  XOR U5137 ( .A(n5074), .B(n5102), .Z(n5075) );
  AND U5138 ( .A(n2743), .B(n872), .Z(n5102) );
  XNOR U5139 ( .A(n5106), .B(n5103), .Z(n5105) );
  XOR U5140 ( .A(n5107), .B(n5108), .Z(n5089) );
  AND U5141 ( .A(n5109), .B(n5110), .Z(n5108) );
  XOR U5142 ( .A(n5098), .B(n5111), .Z(n5110) );
  XNOR U5143 ( .A(n5100), .B(n5107), .Z(n5111) );
  NAND U5144 ( .A(n928), .B(n2743), .Z(n5100) );
  XOR U5145 ( .A(n5097), .B(n5112), .Z(n5098) );
  AND U5146 ( .A(n2615), .B(n984), .Z(n5112) );
  XNOR U5147 ( .A(n5096), .B(g_input[6]), .Z(n5095) );
  NOR U5148 ( .A(n5113), .B(n5114), .Z(n5096) );
  XNOR U5149 ( .A(n5118), .B(n5115), .Z(n5117) );
  XOR U5150 ( .A(n5104), .B(n5119), .Z(n5109) );
  XNOR U5151 ( .A(n5106), .B(n5107), .Z(n5119) );
  OR U5152 ( .A(n834), .B(n3010), .Z(n5106) );
  XOR U5153 ( .A(n5103), .B(n5120), .Z(n5104) );
  ANDN U5154 ( .A(n872), .B(n2872), .Z(n5120) );
  XNOR U5155 ( .A(n5124), .B(n5121), .Z(n5123) );
  XOR U5156 ( .A(n5125), .B(n5126), .Z(n5107) );
  AND U5157 ( .A(n5127), .B(n5128), .Z(n5126) );
  XOR U5158 ( .A(n5116), .B(n5129), .Z(n5128) );
  XNOR U5159 ( .A(n5118), .B(n5125), .Z(n5129) );
  NANDN U5160 ( .B(n2872), .A(n928), .Z(n5118) );
  XOR U5161 ( .A(n5115), .B(n5130), .Z(n5116) );
  AND U5162 ( .A(n2743), .B(n984), .Z(n5130) );
  XOR U5163 ( .A(n5113), .B(g_input[5]), .Z(n5114) );
  NANDN U5164 ( .B(n5131), .A(n5132), .Z(n5113) );
  XOR U5165 ( .A(n5122), .B(n5136), .Z(n5127) );
  XNOR U5166 ( .A(n5124), .B(n5125), .Z(n5136) );
  NANDN U5167 ( .B(n834), .A(n3146), .Z(n5124) );
  XOR U5168 ( .A(n5121), .B(n5137), .Z(n5122) );
  ANDN U5169 ( .A(n872), .B(n3010), .Z(n5137) );
  NANDN U5170 ( .B(n834), .A(n3835), .Z(n5140) );
  XNOR U5171 ( .A(n5138), .B(n5142), .Z(n5139) );
  AND U5172 ( .A(n3146), .B(n872), .Z(n5142) );
  AND U5173 ( .A(n5143), .B(g_input[0]), .Z(n5138) );
  NAND U5174 ( .A(n5144), .B(n834), .Z(n5143) );
  NAND U5175 ( .A(n3835), .B(n872), .Z(n5144) );
  XNOR U5176 ( .A(n5133), .B(n5148), .Z(n5134) );
  ANDN U5177 ( .A(n984), .B(n2872), .Z(n5148) );
  XOR U5178 ( .A(n5151), .B(n5149), .Z(n5150) );
  ANDN U5179 ( .A(n984), .B(n3010), .Z(n5151) );
  AND U5180 ( .A(n3146), .B(n928), .Z(n5152) );
  XOR U5181 ( .A(n5156), .B(n5135), .Z(n5147) );
  NANDN U5182 ( .B(n3010), .A(n928), .Z(n5135) );
  IV U5183 ( .A(n5141), .Z(n5156) );
  NAND U5184 ( .A(n928), .B(n3835), .Z(n5155) );
  XNOR U5185 ( .A(n5153), .B(n5157), .Z(n5154) );
  AND U5186 ( .A(n3146), .B(n984), .Z(n5157) );
  AND U5187 ( .A(n5158), .B(g_input[0]), .Z(n5153) );
  NANDN U5188 ( .B(n928), .A(n5159), .Z(n5158) );
  NAND U5189 ( .A(n3835), .B(n984), .Z(n5159) );
  XNOR U5190 ( .A(n3139), .B(n5163), .Z(n3140) );
  ANDN U5191 ( .A(n806), .B(n2872), .Z(n5163) );
  XNOR U5192 ( .A(n5132), .B(g_input[4]), .Z(n5131) );
  NOR U5193 ( .A(n5164), .B(n5165), .Z(n5132) );
  XOR U5194 ( .A(n5168), .B(n5166), .Z(n5167) );
  ANDN U5195 ( .A(n806), .B(n3010), .Z(n5168) );
  AND U5196 ( .A(n3146), .B(n771), .Z(n5169) );
  XOR U5197 ( .A(n5173), .B(n3141), .Z(n5162) );
  NANDN U5198 ( .B(n3010), .A(n771), .Z(n3141) );
  NANDN U5199 ( .B(n5174), .A(n5175), .Z(n5164) );
  IV U5200 ( .A(n3143), .Z(n5173) );
  NAND U5201 ( .A(n771), .B(n3835), .Z(n5172) );
  XNOR U5202 ( .A(n5170), .B(n5176), .Z(n5171) );
  AND U5203 ( .A(n3146), .B(n806), .Z(n5176) );
  AND U5204 ( .A(n5177), .B(g_input[0]), .Z(n5170) );
  NANDN U5205 ( .B(n771), .A(n5178), .Z(n5177) );
  NAND U5206 ( .A(n3835), .B(n806), .Z(n5178) );
  XNOR U5207 ( .A(n3150), .B(n3151), .Z(n3145) );
  NANDN U5208 ( .B(n716), .A(n3835), .Z(n3151) );
  XNOR U5209 ( .A(n3149), .B(n5181), .Z(n3150) );
  AND U5210 ( .A(n3146), .B(n746), .Z(n5181) );
  XNOR U5211 ( .A(n5175), .B(g_input[2]), .Z(n5174) );
  AND U5212 ( .A(n5183), .B(g_input[0]), .Z(n3149) );
  NAND U5213 ( .A(n5184), .B(n716), .Z(n5183) );
  NANDN U5214 ( .B(n5185), .A(n5186), .Z(n716) );
  ANDN U5215 ( .A(e_input[31]), .B(n5187), .Z(n5186) );
  NAND U5216 ( .A(n3835), .B(n746), .Z(n5184) );
  XOR U5217 ( .A(n5187), .B(e_input[30]), .Z(n5185) );
  OR U5218 ( .A(n5180), .B(n5188), .Z(n5187) );
  XOR U5219 ( .A(n5188), .B(e_input[29]), .Z(n5180) );
  OR U5220 ( .A(n5179), .B(n5189), .Z(n5188) );
  XOR U5221 ( .A(n5189), .B(e_input[28]), .Z(n5179) );
  OR U5222 ( .A(n5145), .B(n5190), .Z(n5189) );
  XOR U5223 ( .A(n5190), .B(e_input[27]), .Z(n5145) );
  OR U5224 ( .A(n5146), .B(n5191), .Z(n5190) );
  XOR U5225 ( .A(n5191), .B(e_input[26]), .Z(n5146) );
  OR U5226 ( .A(n5161), .B(n5192), .Z(n5191) );
  XOR U5227 ( .A(n5192), .B(e_input[25]), .Z(n5161) );
  OR U5228 ( .A(n5160), .B(n5193), .Z(n5192) );
  XOR U5229 ( .A(n5193), .B(e_input[24]), .Z(n5160) );
  OR U5230 ( .A(n4889), .B(n5194), .Z(n5193) );
  XOR U5231 ( .A(n5194), .B(e_input[23]), .Z(n4889) );
  OR U5232 ( .A(n4890), .B(n5195), .Z(n5194) );
  XOR U5233 ( .A(n5195), .B(e_input[22]), .Z(n4890) );
  OR U5234 ( .A(n4885), .B(n5196), .Z(n5195) );
  XOR U5235 ( .A(n5196), .B(e_input[21]), .Z(n4885) );
  OR U5236 ( .A(n4884), .B(n5197), .Z(n5196) );
  XOR U5237 ( .A(n5197), .B(e_input[20]), .Z(n4884) );
  OR U5238 ( .A(n5056), .B(n5198), .Z(n5197) );
  XOR U5239 ( .A(n5198), .B(e_input[19]), .Z(n5056) );
  OR U5240 ( .A(n5055), .B(n5199), .Z(n5198) );
  XOR U5241 ( .A(n5199), .B(e_input[18]), .Z(n5055) );
  OR U5242 ( .A(n5071), .B(n5200), .Z(n5199) );
  XOR U5243 ( .A(n5200), .B(e_input[17]), .Z(n5071) );
  OR U5244 ( .A(n5070), .B(n5201), .Z(n5200) );
  XOR U5245 ( .A(n5201), .B(e_input[16]), .Z(n5070) );
  OR U5246 ( .A(n3875), .B(n5202), .Z(n5201) );
  XOR U5247 ( .A(n5202), .B(e_input[15]), .Z(n3875) );
  OR U5248 ( .A(n3874), .B(n5203), .Z(n5202) );
  XOR U5249 ( .A(n5203), .B(e_input[14]), .Z(n3874) );
  OR U5250 ( .A(n3870), .B(n5204), .Z(n5203) );
  XOR U5251 ( .A(n5204), .B(e_input[13]), .Z(n3870) );
  OR U5252 ( .A(n3869), .B(n5205), .Z(n5204) );
  XOR U5253 ( .A(n5205), .B(e_input[12]), .Z(n3869) );
  OR U5254 ( .A(n3840), .B(n5206), .Z(n5205) );
  XOR U5255 ( .A(n5206), .B(e_input[11]), .Z(n3840) );
  OR U5256 ( .A(n3839), .B(n5207), .Z(n5206) );
  XOR U5257 ( .A(n5207), .B(e_input[10]), .Z(n3839) );
  OR U5258 ( .A(n3855), .B(n5208), .Z(n5207) );
  XOR U5259 ( .A(n5208), .B(e_input[9]), .Z(n3855) );
  OR U5260 ( .A(n3854), .B(n5209), .Z(n5208) );
  XOR U5261 ( .A(n5209), .B(e_input[8]), .Z(n3854) );
  OR U5262 ( .A(n4325), .B(n5210), .Z(n5209) );
  XOR U5263 ( .A(n5210), .B(e_input[7]), .Z(n4325) );
  OR U5264 ( .A(n4324), .B(n5211), .Z(n5210) );
  XOR U5265 ( .A(n5211), .B(e_input[6]), .Z(n4324) );
  OR U5266 ( .A(n4320), .B(n5212), .Z(n5211) );
  XOR U5267 ( .A(n5212), .B(e_input[5]), .Z(n4320) );
  OR U5268 ( .A(n4319), .B(n5213), .Z(n5212) );
  XOR U5269 ( .A(n5213), .B(e_input[4]), .Z(n4319) );
  OR U5270 ( .A(n4684), .B(n5214), .Z(n5213) );
  XOR U5271 ( .A(n5214), .B(e_input[3]), .Z(n4684) );
  OR U5272 ( .A(n4683), .B(n5215), .Z(n5214) );
  XOR U5273 ( .A(n5215), .B(e_input[2]), .Z(n4683) );
  NANDN U5274 ( .B(e_input[0]), .A(n4698), .Z(n5215) );
  XNOR U5275 ( .A(e_input[0]), .B(e_input[1]), .Z(n4698) );
  XOR U5276 ( .A(g_input[0]), .B(g_input[1]), .Z(n5182) );
  AND U5277 ( .A(n5216), .B(n5217), .Z(\_MxM/N31 ) );
  XOR U5278 ( .A(\_MxM/n[13] ), .B(\_MxM/add_43/carry[13] ), .Z(n5217) );
  AND U5279 ( .A(\_MxM/N16 ), .B(n5216), .Z(\_MxM/N30 ) );
  AND U5280 ( .A(\_MxM/N15 ), .B(n5216), .Z(\_MxM/N29 ) );
  AND U5281 ( .A(\_MxM/N14 ), .B(n5216), .Z(\_MxM/N28 ) );
  AND U5282 ( .A(\_MxM/N13 ), .B(n5216), .Z(\_MxM/N27 ) );
  AND U5283 ( .A(\_MxM/N12 ), .B(n5216), .Z(\_MxM/N26 ) );
  AND U5284 ( .A(\_MxM/N11 ), .B(n5216), .Z(\_MxM/N25 ) );
  AND U5285 ( .A(\_MxM/N10 ), .B(n5216), .Z(\_MxM/N24 ) );
  AND U5286 ( .A(\_MxM/N9 ), .B(n5216), .Z(\_MxM/N23 ) );
  AND U5287 ( .A(\_MxM/N8 ), .B(n5216), .Z(\_MxM/N22 ) );
  AND U5288 ( .A(\_MxM/N7 ), .B(n5216), .Z(\_MxM/N21 ) );
  AND U5289 ( .A(\_MxM/N6 ), .B(n5216), .Z(\_MxM/N20 ) );
  AND U5290 ( .A(\_MxM/N5 ), .B(n5216), .Z(\_MxM/N19 ) );
  NAND U5291 ( .A(n5218), .B(n5219), .Z(n5216) );
  AND U5292 ( .A(n5220), .B(n5221), .Z(n5219) );
  ANDN U5293 ( .A(n654), .B(\_MxM/N18 ), .Z(n5221) );
  NOR U5294 ( .A(\_MxM/n[12] ), .B(\_MxM/n[11] ), .Z(n654) );
  AND U5295 ( .A(\_MxM/n[10] ), .B(n5222), .Z(n5220) );
  NOR U5296 ( .A(n656), .B(n657), .Z(n5222) );
  OR U5297 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n657) );
  OR U5298 ( .A(\_MxM/n[5] ), .B(\_MxM/n[4] ), .Z(n656) );
  AND U5299 ( .A(n5223), .B(n5224), .Z(n5218) );
  AND U5300 ( .A(\_MxM/n[2] ), .B(n5225), .Z(n5224) );
  AND U5301 ( .A(\_MxM/n[1] ), .B(\_MxM/n[13] ), .Z(n5225) );
  AND U5302 ( .A(\_MxM/n[9] ), .B(n5226), .Z(n5223) );
  AND U5303 ( .A(\_MxM/n[8] ), .B(\_MxM/n[3] ), .Z(n5226) );
  IV U5304 ( .A(\_MxM/n[0] ), .Z(\_MxM/N18 ) );
endmodule

