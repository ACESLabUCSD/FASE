
module MxM_TG_W8_N1000 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n117 , \_MxM/n116 , \_MxM/n115 , \_MxM/n114 , \_MxM/n113 ,
         \_MxM/n112 , \_MxM/n111 , \_MxM/n110 , \_MxM/n109 , \_MxM/n108 ,
         \_MxM/n107 , \_MxM/n106 , \_MxM/n105 , \_MxM/n104 , \_MxM/n103 ,
         \_MxM/n102 , \_MxM/N24 , \_MxM/N23 , \_MxM/N22 , \_MxM/N21 ,
         \_MxM/N20 , \_MxM/N19 , \_MxM/N18 , \_MxM/N17 , \_MxM/N16 ,
         \_MxM/N15 , \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 ,
         \_MxM/N8 , \_MxM/N7 , \_MxM/N6 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/Y0[0] , \_MxM/Y0[1] ,
         \_MxM/Y0[2] , \_MxM/Y0[3] , \_MxM/Y0[4] , \_MxM/Y0[5] , \_MxM/Y0[6] ,
         \_MxM/Y0[7] , \_MxM/add_39/carry[9] , \_MxM/add_39/carry[8] ,
         \_MxM/add_39/carry[7] , \_MxM/add_39/carry[6] ,
         \_MxM/add_39/carry[5] , \_MxM/add_39/carry[4] ,
         \_MxM/add_39/carry[3] , \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n102 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n103 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n104 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n105 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n106 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n107 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n108 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n109 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n110 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n111 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n112 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n113 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n114 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n115 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n116 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n117 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N24 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N18 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N13 ) );
  MUX U1 ( .IN0(n311), .IN1(n327), .SEL(n313), .F(n292) );
  MUX U2 ( .IN0(g_input[3]), .IN1(n376), .SEL(g_input[7]), .F(n1) );
  IV U3 ( .A(n1), .Z(n221) );
  MUX U4 ( .IN0(n261), .IN1(n259), .SEL(n260), .F(n216) );
  NAND U5 ( .A(n134), .B(n168), .Z(n167) );
  MUX U6 ( .IN0(n244), .IN1(n2), .SEL(n243), .F(n199) );
  IV U7 ( .A(n242), .Z(n2) );
  MUX U8 ( .IN0(n3), .IN1(n144), .SEL(n145), .F(n112) );
  IV U9 ( .A(\_MxM/Y0[3] ), .Z(n3) );
  XOR U10 ( .A(n375), .B(g_input[3]), .Z(n376) );
  XNOR U11 ( .A(n363), .B(n364), .Z(n342) );
  MUX U12 ( .IN0(e_input[6]), .IN1(n401), .SEL(e_input[7]), .F(n110) );
  MUX U13 ( .IN0(e_input[3]), .IN1(n351), .SEL(e_input[7]), .F(n202) );
  MUX U14 ( .IN0(n205), .IN1(n4), .SEL(n206), .F(n157) );
  IV U15 ( .A(n207), .Z(n4) );
  XNOR U16 ( .A(n208), .B(n173), .Z(n165) );
  MUX U17 ( .IN0(n5), .IN1(n227), .SEL(n228), .F(n182) );
  IV U18 ( .A(\_MxM/Y0[1] ), .Z(n5) );
  XOR U19 ( .A(n80), .B(n90), .Z(n88) );
  MUX U20 ( .IN0(n6), .IN1(n381), .SEL(n382), .F(n377) );
  IV U21 ( .A(n383), .Z(n6) );
  MUX U22 ( .IN0(g_input[4]), .IN1(n328), .SEL(g_input[7]), .F(n7) );
  IV U23 ( .A(n7), .Z(n175) );
  MUX U24 ( .IN0(g_input[5]), .IN1(n310), .SEL(g_input[7]), .F(n138) );
  XOR U25 ( .A(n224), .B(n263), .Z(n225) );
  MUX U26 ( .IN0(g_input[6]), .IN1(n282), .SEL(g_input[7]), .F(n111) );
  MUX U27 ( .IN0(n245), .IN1(n8), .SEL(n246), .F(n205) );
  IV U28 ( .A(n247), .Z(n8) );
  XNOR U29 ( .A(n127), .B(n128), .Z(n151) );
  XOR U30 ( .A(n112), .B(n122), .Z(n120) );
  NOR U31 ( .A(g_input[0]), .B(n398), .Z(n386) );
  MUX U32 ( .IN0(n9), .IN1(n275), .SEL(n276), .F(n322) );
  IV U33 ( .A(n342), .Z(n9) );
  MUX U34 ( .IN0(n377), .IN1(n380), .SEL(n378), .F(n253) );
  MUX U35 ( .IN0(n292), .IN1(n308), .SEL(n294), .F(n286) );
  MUX U36 ( .IN0(n137), .IN1(n161), .SEL(n136), .F(n99) );
  NAND U37 ( .A(n199), .B(n240), .Z(n239) );
  XNOR U38 ( .A(n261), .B(n260), .Z(n247) );
  XNOR U39 ( .A(n166), .B(n165), .Z(n159) );
  XNOR U40 ( .A(n220), .B(n219), .Z(n207) );
  MUX U41 ( .IN0(\_MxM/Y0[6] ), .IN1(n62), .SEL(n57), .F(n50) );
  XOR U42 ( .A(n144), .B(n152), .Z(n150) );
  MUX U43 ( .IN0(g_input[2]), .IN1(n385), .SEL(g_input[7]), .F(n262) );
  XOR U44 ( .A(n352), .B(n333), .Z(n276) );
  XNOR U45 ( .A(n251), .B(n213), .Z(n219) );
  MUX U46 ( .IN0(n250), .IN1(n248), .SEL(n249), .F(n10) );
  IV U47 ( .A(n10), .Z(n204) );
  AND U48 ( .A(n105), .B(n71), .Z(n104) );
  MUX U49 ( .IN0(n11), .IN1(n159), .SEL(n158), .F(n128) );
  IV U50 ( .A(n157), .Z(n11) );
  MUX U51 ( .IN0(n12), .IN1(n182), .SEL(n183), .F(n144) );
  IV U52 ( .A(\_MxM/Y0[2] ), .Z(n12) );
  MUX U53 ( .IN0(\_MxM/Y0[7] ), .IN1(n50), .SEL(n51), .F(n13) );
  IV U54 ( .A(n13), .Z(n47) );
  XOR U55 ( .A(n228), .B(\_MxM/Y0[1] ), .Z(n16) );
  NAND U56 ( .A(n14), .B(n15), .Z(\_MxM/n117 ) );
  OR U57 ( .A(n16), .B(n17), .Z(n15) );
  NANDN U58 ( .B(n18), .A(\_MxM/Y0[0] ), .Z(n14) );
  NAND U59 ( .A(n19), .B(n20), .Z(\_MxM/n116 ) );
  NANDN U60 ( .B(n17), .A(n21), .Z(n20) );
  NANDN U61 ( .B(n22), .A(rst), .Z(n19) );
  NAND U62 ( .A(n23), .B(n24), .Z(\_MxM/n115 ) );
  NANDN U63 ( .B(n17), .A(n25), .Z(n24) );
  NANDN U64 ( .B(n18), .A(\_MxM/Y0[2] ), .Z(n23) );
  NAND U65 ( .A(n26), .B(n27), .Z(\_MxM/n114 ) );
  NANDN U66 ( .B(n17), .A(n28), .Z(n27) );
  NANDN U67 ( .B(n18), .A(\_MxM/Y0[3] ), .Z(n26) );
  NAND U68 ( .A(n29), .B(n30), .Z(\_MxM/n113 ) );
  NANDN U69 ( .B(n17), .A(n31), .Z(n30) );
  NANDN U70 ( .B(n18), .A(\_MxM/Y0[4] ), .Z(n29) );
  NAND U71 ( .A(n32), .B(n33), .Z(\_MxM/n112 ) );
  NANDN U72 ( .B(n17), .A(n34), .Z(n33) );
  NANDN U73 ( .B(n18), .A(\_MxM/Y0[5] ), .Z(n32) );
  NAND U74 ( .A(n35), .B(n36), .Z(\_MxM/n111 ) );
  OR U75 ( .A(n37), .B(n17), .Z(n36) );
  NANDN U76 ( .B(n18), .A(\_MxM/Y0[6] ), .Z(n35) );
  NAND U77 ( .A(n38), .B(n39), .Z(\_MxM/n110 ) );
  OR U78 ( .A(n17), .B(n40), .Z(n39) );
  NANDN U79 ( .B(n41), .A(n18), .Z(n17) );
  NANDN U80 ( .B(n18), .A(\_MxM/Y0[7] ), .Z(n38) );
  NAND U81 ( .A(n42), .B(n43), .Z(\_MxM/n109 ) );
  NANDN U82 ( .B(n18), .A(o[7]), .Z(n43) );
  AND U83 ( .A(n44), .B(n45), .Z(n42) );
  NANDN U84 ( .B(n41), .A(o[7]), .Z(n45) );
  OR U85 ( .A(n40), .B(n46), .Z(n44) );
  XOR U86 ( .A(n47), .B(n48), .Z(n40) );
  XNOR U87 ( .A(\_MxM/Y0[7] ), .B(n49), .Z(n48) );
  NAND U88 ( .A(n52), .B(n53), .Z(\_MxM/n108 ) );
  NANDN U89 ( .B(n18), .A(o[6]), .Z(n53) );
  AND U90 ( .A(n54), .B(n55), .Z(n52) );
  NANDN U91 ( .B(n41), .A(o[6]), .Z(n55) );
  OR U92 ( .A(n37), .B(n46), .Z(n54) );
  XOR U93 ( .A(n51), .B(\_MxM/Y0[7] ), .Z(n37) );
  XOR U94 ( .A(n50), .B(n49), .Z(n51) );
  NAND U95 ( .A(n58), .B(n59), .Z(\_MxM/n107 ) );
  NANDN U96 ( .B(n18), .A(o[5]), .Z(n59) );
  AND U97 ( .A(n60), .B(n61), .Z(n58) );
  NANDN U98 ( .B(n41), .A(o[5]), .Z(n61) );
  NANDN U99 ( .B(n46), .A(n34), .Z(n60) );
  XNOR U100 ( .A(n57), .B(\_MxM/Y0[6] ), .Z(n34) );
  XOR U101 ( .A(n62), .B(n63), .Z(n57) );
  ANDN U102 ( .A(n49), .B(n64), .Z(n63) );
  NANDN U103 ( .B(n65), .A(n66), .Z(n49) );
  ANDN U104 ( .A(n67), .B(n64), .Z(n65) );
  NAND U105 ( .A(n68), .B(n69), .Z(n64) );
  OR U106 ( .A(n70), .B(n71), .Z(n69) );
  AND U107 ( .A(n72), .B(n73), .Z(n68) );
  OR U108 ( .A(n74), .B(n75), .Z(n73) );
  OR U109 ( .A(n76), .B(n77), .Z(n72) );
  NOR U110 ( .A(n78), .B(n79), .Z(n67) );
  IV U111 ( .A(n56), .Z(n62) );
  XOR U112 ( .A(n80), .B(n81), .Z(n56) );
  ANDN U113 ( .A(n82), .B(n83), .Z(n81) );
  XNOR U114 ( .A(\_MxM/Y0[5] ), .B(n80), .Z(n82) );
  NAND U115 ( .A(n84), .B(n85), .Z(\_MxM/n106 ) );
  NANDN U116 ( .B(n18), .A(o[4]), .Z(n85) );
  AND U117 ( .A(n86), .B(n87), .Z(n84) );
  NANDN U118 ( .B(n41), .A(o[4]), .Z(n87) );
  NANDN U119 ( .B(n46), .A(n31), .Z(n86) );
  XNOR U120 ( .A(n83), .B(\_MxM/Y0[5] ), .Z(n31) );
  XNOR U121 ( .A(n88), .B(n89), .Z(n83) );
  AND U122 ( .A(n66), .B(n91), .Z(n90) );
  XOR U123 ( .A(n78), .B(n92), .Z(n91) );
  XOR U124 ( .A(n92), .B(n79), .Z(n78) );
  OR U125 ( .A(n93), .B(n94), .Z(n79) );
  IV U126 ( .A(n89), .Z(n92) );
  XNOR U127 ( .A(n77), .B(n76), .Z(n89) );
  OR U128 ( .A(n95), .B(n96), .Z(n76) );
  AND U129 ( .A(n97), .B(n98), .Z(n77) );
  XNOR U130 ( .A(n99), .B(n100), .Z(n98) );
  ANDN U131 ( .A(n101), .B(n102), .Z(n100) );
  XOR U132 ( .A(n99), .B(n103), .Z(n101) );
  XNOR U133 ( .A(n70), .B(n104), .Z(n97) );
  NAND U134 ( .A(n106), .B(n107), .Z(n71) );
  NANDN U135 ( .B(n108), .A(n109), .Z(n106) );
  NANDN U136 ( .B(n74), .A(n110), .Z(n105) );
  NANDN U137 ( .B(n75), .A(n111), .Z(n70) );
  XOR U138 ( .A(n112), .B(n113), .Z(n80) );
  ANDN U139 ( .A(n114), .B(n115), .Z(n113) );
  XNOR U140 ( .A(\_MxM/Y0[4] ), .B(n112), .Z(n114) );
  NAND U141 ( .A(n116), .B(n117), .Z(\_MxM/n105 ) );
  NANDN U142 ( .B(n18), .A(o[3]), .Z(n117) );
  AND U143 ( .A(n118), .B(n119), .Z(n116) );
  NANDN U144 ( .B(n41), .A(o[3]), .Z(n119) );
  NANDN U145 ( .B(n46), .A(n28), .Z(n118) );
  XNOR U146 ( .A(n115), .B(\_MxM/Y0[4] ), .Z(n28) );
  XNOR U147 ( .A(n120), .B(n121), .Z(n115) );
  AND U148 ( .A(n66), .B(n123), .Z(n122) );
  XOR U149 ( .A(n93), .B(n124), .Z(n123) );
  XOR U150 ( .A(n124), .B(n94), .Z(n93) );
  OR U151 ( .A(n125), .B(n126), .Z(n94) );
  IV U152 ( .A(n121), .Z(n124) );
  XNOR U153 ( .A(n96), .B(n95), .Z(n121) );
  OR U154 ( .A(n127), .B(n128), .Z(n95) );
  XOR U155 ( .A(n103), .B(n102), .Z(n96) );
  XOR U156 ( .A(n99), .B(n129), .Z(n102) );
  AND U157 ( .A(n130), .B(n131), .Z(n129) );
  NANDN U158 ( .B(n74), .A(n132), .Z(n131) );
  OR U159 ( .A(n133), .B(n134), .Z(n130) );
  XOR U160 ( .A(n108), .B(n109), .Z(n103) );
  NANDN U161 ( .B(n75), .A(n138), .Z(n109) );
  XNOR U162 ( .A(n107), .B(n139), .Z(n108) );
  AND U163 ( .A(n111), .B(n110), .Z(n139) );
  ANDN U164 ( .A(n140), .B(n141), .Z(n107) );
  NANDN U165 ( .B(n142), .A(n143), .Z(n140) );
  NAND U166 ( .A(n146), .B(n147), .Z(\_MxM/n104 ) );
  NANDN U167 ( .B(n18), .A(o[2]), .Z(n147) );
  AND U168 ( .A(n148), .B(n149), .Z(n146) );
  NANDN U169 ( .B(n41), .A(o[2]), .Z(n149) );
  NANDN U170 ( .B(n46), .A(n25), .Z(n148) );
  XNOR U171 ( .A(n145), .B(\_MxM/Y0[3] ), .Z(n25) );
  XNOR U172 ( .A(n150), .B(n151), .Z(n145) );
  AND U173 ( .A(n66), .B(n153), .Z(n152) );
  XOR U174 ( .A(n125), .B(n154), .Z(n153) );
  XOR U175 ( .A(n154), .B(n126), .Z(n125) );
  OR U176 ( .A(n155), .B(n156), .Z(n126) );
  IV U177 ( .A(n151), .Z(n154) );
  XOR U178 ( .A(n137), .B(n136), .Z(n127) );
  XNOR U179 ( .A(n160), .B(n161), .Z(n136) );
  IV U180 ( .A(n135), .Z(n161) );
  XOR U181 ( .A(n162), .B(n163), .Z(n135) );
  ANDN U182 ( .A(n164), .B(n165), .Z(n163) );
  XOR U183 ( .A(n162), .B(n166), .Z(n164) );
  XNOR U184 ( .A(n167), .B(n133), .Z(n160) );
  NAND U185 ( .A(n132), .B(n111), .Z(n133) );
  NANDN U186 ( .B(n74), .A(n169), .Z(n168) );
  XNOR U187 ( .A(n170), .B(n171), .Z(n134) );
  ANDN U188 ( .A(n172), .B(n173), .Z(n171) );
  XNOR U189 ( .A(n174), .B(n170), .Z(n172) );
  XOR U190 ( .A(n142), .B(n143), .Z(n137) );
  OR U191 ( .A(n175), .B(n75), .Z(n143) );
  XNOR U192 ( .A(n176), .B(n177), .Z(n142) );
  AND U193 ( .A(n138), .B(n110), .Z(n177) );
  IV U194 ( .A(n141), .Z(n176) );
  NAND U195 ( .A(n178), .B(n179), .Z(n141) );
  NANDN U196 ( .B(n180), .A(n181), .Z(n178) );
  NAND U197 ( .A(n184), .B(n185), .Z(\_MxM/n103 ) );
  NANDN U198 ( .B(n18), .A(o[1]), .Z(n185) );
  AND U199 ( .A(n186), .B(n187), .Z(n184) );
  NANDN U200 ( .B(n41), .A(o[1]), .Z(n187) );
  NANDN U201 ( .B(n46), .A(n21), .Z(n186) );
  XNOR U202 ( .A(n183), .B(\_MxM/Y0[2] ), .Z(n21) );
  XNOR U203 ( .A(n188), .B(n189), .Z(n183) );
  XOR U204 ( .A(n182), .B(n190), .Z(n188) );
  AND U205 ( .A(n66), .B(n191), .Z(n190) );
  XOR U206 ( .A(n155), .B(n192), .Z(n191) );
  XOR U207 ( .A(n192), .B(n156), .Z(n155) );
  NANDN U208 ( .B(n193), .A(n194), .Z(n156) );
  IV U209 ( .A(n189), .Z(n192) );
  XOR U210 ( .A(n159), .B(n158), .Z(n189) );
  XNOR U211 ( .A(n157), .B(n195), .Z(n158) );
  AND U212 ( .A(n196), .B(n197), .Z(n195) );
  OR U213 ( .A(n198), .B(n199), .Z(n197) );
  AND U214 ( .A(n200), .B(n201), .Z(n196) );
  NANDN U215 ( .B(n74), .A(n202), .Z(n201) );
  NAND U216 ( .A(n203), .B(n204), .Z(n200) );
  XNOR U217 ( .A(n170), .B(n209), .Z(n173) );
  AND U218 ( .A(n111), .B(n169), .Z(n209) );
  XOR U219 ( .A(n210), .B(n211), .Z(n170) );
  ANDN U220 ( .A(n212), .B(n213), .Z(n211) );
  XNOR U221 ( .A(n214), .B(n210), .Z(n212) );
  XOR U222 ( .A(n215), .B(n174), .Z(n208) );
  NAND U223 ( .A(n132), .B(n138), .Z(n174) );
  IV U224 ( .A(n162), .Z(n215) );
  XOR U225 ( .A(n216), .B(n217), .Z(n162) );
  ANDN U226 ( .A(n218), .B(n219), .Z(n217) );
  XOR U227 ( .A(n216), .B(n220), .Z(n218) );
  XNOR U228 ( .A(n180), .B(n181), .Z(n166) );
  OR U229 ( .A(n221), .B(n75), .Z(n181) );
  XNOR U230 ( .A(n179), .B(n222), .Z(n180) );
  ANDN U231 ( .A(n110), .B(n175), .Z(n222) );
  ANDN U232 ( .A(n223), .B(n224), .Z(n179) );
  NANDN U233 ( .B(n225), .A(n226), .Z(n223) );
  NAND U234 ( .A(n229), .B(n230), .Z(\_MxM/n102 ) );
  NANDN U235 ( .B(n18), .A(o[0]), .Z(n230) );
  AND U236 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U237 ( .B(n41), .A(o[0]), .Z(n232) );
  IV U238 ( .A(n233), .Z(n41) );
  OR U239 ( .A(n46), .B(n16), .Z(n231) );
  IV U240 ( .A(\_MxM/Y0[1] ), .Z(n22) );
  XOR U241 ( .A(n234), .B(n235), .Z(n228) );
  XNOR U242 ( .A(n236), .B(n227), .Z(n234) );
  NAND U243 ( .A(\_MxM/Y0[0] ), .B(n193), .Z(n227) );
  NAND U244 ( .A(n237), .B(n66), .Z(n236) );
  XOR U245 ( .A(e_input[7]), .B(g_input[7]), .Z(n66) );
  XNOR U246 ( .A(n194), .B(n235), .Z(n237) );
  XNOR U247 ( .A(n193), .B(n235), .Z(n194) );
  XNOR U248 ( .A(n207), .B(n206), .Z(n235) );
  XNOR U249 ( .A(n238), .B(n203), .Z(n206) );
  XNOR U250 ( .A(n239), .B(n198), .Z(n203) );
  NAND U251 ( .A(n111), .B(n202), .Z(n198) );
  NANDN U252 ( .B(n74), .A(n241), .Z(n240) );
  XNOR U253 ( .A(n204), .B(n205), .Z(n238) );
  XNOR U254 ( .A(n210), .B(n252), .Z(n213) );
  AND U255 ( .A(n138), .B(n169), .Z(n252) );
  XOR U256 ( .A(n253), .B(n254), .Z(n210) );
  ANDN U257 ( .A(n255), .B(n256), .Z(n254) );
  XNOR U258 ( .A(n257), .B(n253), .Z(n255) );
  XOR U259 ( .A(n258), .B(n214), .Z(n251) );
  NANDN U260 ( .B(n175), .A(n132), .Z(n214) );
  IV U261 ( .A(n216), .Z(n258) );
  XNOR U262 ( .A(n225), .B(n226), .Z(n220) );
  NANDN U263 ( .B(n75), .A(n262), .Z(n226) );
  ANDN U264 ( .A(n110), .B(n221), .Z(n263) );
  NAND U265 ( .A(n264), .B(n265), .Z(n224) );
  NANDN U266 ( .B(n266), .A(n267), .Z(n264) );
  XNOR U267 ( .A(n247), .B(n246), .Z(n193) );
  XNOR U268 ( .A(n268), .B(n250), .Z(n246) );
  XNOR U269 ( .A(n243), .B(n244), .Z(n250) );
  NAND U270 ( .A(n138), .B(n202), .Z(n244) );
  XNOR U271 ( .A(n242), .B(n269), .Z(n243) );
  AND U272 ( .A(n241), .B(n111), .Z(n269) );
  XOR U273 ( .A(n270), .B(n271), .Z(n242) );
  AND U274 ( .A(n272), .B(n273), .Z(n271) );
  XNOR U275 ( .A(n274), .B(n270), .Z(n273) );
  XNOR U276 ( .A(n249), .B(n245), .Z(n268) );
  XOR U277 ( .A(n275), .B(n276), .Z(n245) );
  XOR U278 ( .A(n277), .B(n278), .Z(n249) );
  AND U279 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U280 ( .B(n74), .A(n281), .Z(n280) );
  NANDN U281 ( .B(n282), .A(n283), .Z(n74) );
  AND U282 ( .A(n284), .B(g_input[7]), .Z(n283) );
  NANDN U283 ( .B(n285), .A(n286), .Z(n279) );
  IV U284 ( .A(n248), .Z(n277) );
  XNOR U285 ( .A(n287), .B(n288), .Z(n248) );
  AND U286 ( .A(n289), .B(n290), .Z(n288) );
  XOR U287 ( .A(n286), .B(n291), .Z(n290) );
  XNOR U288 ( .A(n285), .B(n287), .Z(n291) );
  NAND U289 ( .A(n111), .B(n281), .Z(n285) );
  XNOR U290 ( .A(n295), .B(n292), .Z(n294) );
  XOR U291 ( .A(n272), .B(n296), .Z(n289) );
  XNOR U292 ( .A(n274), .B(n287), .Z(n296) );
  NANDN U293 ( .B(n175), .A(n202), .Z(n274) );
  XOR U294 ( .A(n270), .B(n297), .Z(n272) );
  AND U295 ( .A(n241), .B(n138), .Z(n297) );
  XOR U296 ( .A(n298), .B(n299), .Z(n270) );
  AND U297 ( .A(n300), .B(n301), .Z(n299) );
  XNOR U298 ( .A(n302), .B(n298), .Z(n301) );
  XOR U299 ( .A(n303), .B(n304), .Z(n287) );
  AND U300 ( .A(n305), .B(n306), .Z(n304) );
  XOR U301 ( .A(n293), .B(n307), .Z(n306) );
  XNOR U302 ( .A(n295), .B(n303), .Z(n307) );
  NAND U303 ( .A(n138), .B(n281), .Z(n295) );
  XOR U304 ( .A(n292), .B(n308), .Z(n293) );
  AND U305 ( .A(n111), .B(e_input[0]), .Z(n308) );
  XNOR U306 ( .A(n284), .B(g_input[6]), .Z(n282) );
  NOR U307 ( .A(n309), .B(n310), .Z(n284) );
  XNOR U308 ( .A(n314), .B(n311), .Z(n313) );
  XOR U309 ( .A(n300), .B(n315), .Z(n305) );
  XNOR U310 ( .A(n302), .B(n303), .Z(n315) );
  NANDN U311 ( .B(n221), .A(n202), .Z(n302) );
  XOR U312 ( .A(n298), .B(n316), .Z(n300) );
  ANDN U313 ( .A(n241), .B(n175), .Z(n316) );
  XOR U314 ( .A(n317), .B(n318), .Z(n298) );
  AND U315 ( .A(n319), .B(n320), .Z(n318) );
  XNOR U316 ( .A(n321), .B(n317), .Z(n320) );
  XOR U317 ( .A(n322), .B(n323), .Z(n303) );
  AND U318 ( .A(n324), .B(n325), .Z(n323) );
  XOR U319 ( .A(n312), .B(n326), .Z(n325) );
  XNOR U320 ( .A(n314), .B(n322), .Z(n326) );
  NANDN U321 ( .B(n175), .A(n281), .Z(n314) );
  XOR U322 ( .A(n311), .B(n327), .Z(n312) );
  AND U323 ( .A(n138), .B(e_input[0]), .Z(n327) );
  XOR U324 ( .A(n309), .B(g_input[5]), .Z(n310) );
  NANDN U325 ( .B(n328), .A(n329), .Z(n309) );
  XOR U326 ( .A(n330), .B(n331), .Z(n311) );
  ANDN U327 ( .A(n332), .B(n333), .Z(n331) );
  XNOR U328 ( .A(n334), .B(n330), .Z(n332) );
  XOR U329 ( .A(n319), .B(n335), .Z(n324) );
  XNOR U330 ( .A(n321), .B(n322), .Z(n335) );
  NAND U331 ( .A(n202), .B(n262), .Z(n321) );
  XOR U332 ( .A(n317), .B(n336), .Z(n319) );
  ANDN U333 ( .A(n241), .B(n221), .Z(n336) );
  XOR U334 ( .A(n337), .B(n338), .Z(n317) );
  ANDN U335 ( .A(n339), .B(n340), .Z(n338) );
  XNOR U336 ( .A(n341), .B(n337), .Z(n339) );
  XNOR U337 ( .A(n343), .B(n341), .Z(n275) );
  NAND U338 ( .A(n202), .B(n344), .Z(n341) );
  IV U339 ( .A(n340), .Z(n343) );
  XNOR U340 ( .A(n337), .B(n345), .Z(n340) );
  AND U341 ( .A(n262), .B(n241), .Z(n345) );
  AND U342 ( .A(n346), .B(g_input[0]), .Z(n337) );
  NANDN U343 ( .B(n202), .A(n347), .Z(n346) );
  NAND U344 ( .A(n344), .B(n241), .Z(n347) );
  XNOR U345 ( .A(n348), .B(e_input[2]), .Z(n241) );
  NAND U346 ( .A(n349), .B(e_input[7]), .Z(n348) );
  XOR U347 ( .A(n350), .B(e_input[2]), .Z(n349) );
  XNOR U348 ( .A(n330), .B(n353), .Z(n333) );
  ANDN U349 ( .A(e_input[0]), .B(n175), .Z(n353) );
  XOR U350 ( .A(n354), .B(n355), .Z(n330) );
  AND U351 ( .A(n356), .B(n357), .Z(n355) );
  XOR U352 ( .A(n358), .B(n354), .Z(n357) );
  ANDN U353 ( .A(e_input[0]), .B(n221), .Z(n358) );
  XOR U354 ( .A(n359), .B(n354), .Z(n356) );
  AND U355 ( .A(n281), .B(n262), .Z(n359) );
  XOR U356 ( .A(n360), .B(n361), .Z(n354) );
  ANDN U357 ( .A(n362), .B(n363), .Z(n361) );
  XNOR U358 ( .A(n364), .B(n360), .Z(n362) );
  XOR U359 ( .A(n365), .B(n334), .Z(n352) );
  NANDN U360 ( .B(n221), .A(n281), .Z(n334) );
  IV U361 ( .A(n342), .Z(n365) );
  NAND U362 ( .A(n281), .B(n344), .Z(n364) );
  XNOR U363 ( .A(n360), .B(n366), .Z(n363) );
  AND U364 ( .A(n262), .B(e_input[0]), .Z(n366) );
  AND U365 ( .A(n367), .B(g_input[0]), .Z(n360) );
  NANDN U366 ( .B(n281), .A(n368), .Z(n367) );
  NAND U367 ( .A(n344), .B(e_input[0]), .Z(n368) );
  XNOR U368 ( .A(n369), .B(e_input[1]), .Z(n281) );
  NAND U369 ( .A(n370), .B(e_input[7]), .Z(n369) );
  XNOR U370 ( .A(e_input[1]), .B(n371), .Z(n370) );
  XOR U371 ( .A(n372), .B(n373), .Z(n260) );
  IV U372 ( .A(n256), .Z(n373) );
  XNOR U373 ( .A(n253), .B(n374), .Z(n256) );
  ANDN U374 ( .A(n169), .B(n175), .Z(n374) );
  XNOR U375 ( .A(n329), .B(g_input[4]), .Z(n328) );
  NOR U376 ( .A(n375), .B(n376), .Z(n329) );
  XOR U377 ( .A(n379), .B(n377), .Z(n378) );
  ANDN U378 ( .A(n169), .B(n221), .Z(n379) );
  AND U379 ( .A(n262), .B(n132), .Z(n380) );
  XOR U380 ( .A(n384), .B(n257), .Z(n372) );
  NANDN U381 ( .B(n221), .A(n132), .Z(n257) );
  NANDN U382 ( .B(n385), .A(n386), .Z(n375) );
  IV U383 ( .A(n259), .Z(n384) );
  XOR U384 ( .A(n387), .B(n383), .Z(n259) );
  NAND U385 ( .A(n132), .B(n344), .Z(n383) );
  IV U386 ( .A(n382), .Z(n387) );
  XNOR U387 ( .A(n381), .B(n388), .Z(n382) );
  AND U388 ( .A(n262), .B(n169), .Z(n388) );
  AND U389 ( .A(n389), .B(g_input[0]), .Z(n381) );
  NANDN U390 ( .B(n132), .A(n390), .Z(n389) );
  NAND U391 ( .A(n344), .B(n169), .Z(n390) );
  XNOR U392 ( .A(n391), .B(e_input[4]), .Z(n169) );
  NAND U393 ( .A(n392), .B(e_input[7]), .Z(n391) );
  XOR U394 ( .A(n393), .B(e_input[4]), .Z(n392) );
  XNOR U395 ( .A(n394), .B(e_input[5]), .Z(n132) );
  NAND U396 ( .A(n395), .B(e_input[7]), .Z(n394) );
  XOR U397 ( .A(n396), .B(e_input[5]), .Z(n395) );
  XNOR U398 ( .A(n266), .B(n267), .Z(n261) );
  NANDN U399 ( .B(n75), .A(n344), .Z(n267) );
  XNOR U400 ( .A(n265), .B(n397), .Z(n266) );
  AND U401 ( .A(n262), .B(n110), .Z(n397) );
  XNOR U402 ( .A(n386), .B(g_input[2]), .Z(n385) );
  AND U403 ( .A(n399), .B(g_input[0]), .Z(n265) );
  NAND U404 ( .A(n400), .B(n75), .Z(n399) );
  NANDN U405 ( .B(n401), .A(n402), .Z(n75) );
  ANDN U406 ( .A(e_input[7]), .B(n403), .Z(n402) );
  NAND U407 ( .A(n344), .B(n110), .Z(n400) );
  XOR U408 ( .A(n403), .B(e_input[6]), .Z(n401) );
  OR U409 ( .A(n396), .B(n404), .Z(n403) );
  XOR U410 ( .A(n404), .B(e_input[5]), .Z(n396) );
  OR U411 ( .A(n393), .B(n405), .Z(n404) );
  XOR U412 ( .A(n405), .B(e_input[4]), .Z(n393) );
  OR U413 ( .A(n351), .B(n406), .Z(n405) );
  XOR U414 ( .A(n406), .B(e_input[3]), .Z(n351) );
  OR U415 ( .A(n350), .B(n407), .Z(n406) );
  XOR U416 ( .A(n407), .B(e_input[2]), .Z(n350) );
  NANDN U417 ( .B(e_input[0]), .A(n371), .Z(n407) );
  XNOR U418 ( .A(e_input[0]), .B(e_input[1]), .Z(n371) );
  XNOR U419 ( .A(n408), .B(g_input[1]), .Z(n344) );
  NAND U420 ( .A(n409), .B(g_input[7]), .Z(n408) );
  XOR U421 ( .A(g_input[1]), .B(n398), .Z(n409) );
  XOR U422 ( .A(g_input[0]), .B(g_input[1]), .Z(n398) );
  NANDN U423 ( .B(n233), .A(n18), .Z(n46) );
  IV U424 ( .A(rst), .Z(n18) );
  NAND U425 ( .A(n410), .B(n411), .Z(n233) );
  AND U426 ( .A(n412), .B(n413), .Z(n411) );
  ANDN U427 ( .A(n414), .B(\_MxM/n[7] ), .Z(n413) );
  NOR U428 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n414) );
  NOR U429 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n412) );
  AND U430 ( .A(n415), .B(n416), .Z(n410) );
  NOR U431 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n416) );
  NOR U432 ( .A(\_MxM/n[0] ), .B(n417), .Z(n415) );
  AND U433 ( .A(n418), .B(n419), .Z(\_MxM/N24 ) );
  XOR U434 ( .A(\_MxM/n[9] ), .B(\_MxM/add_39/carry[9] ), .Z(n419) );
  AND U435 ( .A(\_MxM/N13 ), .B(n418), .Z(\_MxM/N23 ) );
  AND U436 ( .A(\_MxM/N12 ), .B(n418), .Z(\_MxM/N22 ) );
  AND U437 ( .A(\_MxM/N11 ), .B(n418), .Z(\_MxM/N21 ) );
  AND U438 ( .A(\_MxM/N10 ), .B(n418), .Z(\_MxM/N20 ) );
  AND U439 ( .A(\_MxM/N9 ), .B(n418), .Z(\_MxM/N19 ) );
  AND U440 ( .A(\_MxM/N8 ), .B(n418), .Z(\_MxM/N18 ) );
  AND U441 ( .A(\_MxM/N7 ), .B(n418), .Z(\_MxM/N17 ) );
  AND U442 ( .A(\_MxM/N6 ), .B(n418), .Z(\_MxM/N16 ) );
  NAND U443 ( .A(n420), .B(n421), .Z(n418) );
  AND U444 ( .A(n422), .B(n423), .Z(n421) );
  AND U445 ( .A(\_MxM/n[1] ), .B(n424), .Z(n423) );
  NOR U446 ( .A(\_MxM/N15 ), .B(n417), .Z(n424) );
  OR U447 ( .A(\_MxM/n[3] ), .B(\_MxM/n[4] ), .Z(n417) );
  AND U448 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n422) );
  AND U449 ( .A(n425), .B(n426), .Z(n420) );
  AND U450 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n426) );
  AND U451 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n425) );
  IV U452 ( .A(\_MxM/n[0] ), .Z(\_MxM/N15 ) );
endmodule

