
module MxM_TG_W16_N10000 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MxM/n219 , \_MxM/n218 , \_MxM/n217 , \_MxM/n216 , \_MxM/n215 ,
         \_MxM/n214 , \_MxM/n213 , \_MxM/n212 , \_MxM/n211 , \_MxM/n210 ,
         \_MxM/n209 , \_MxM/n208 , \_MxM/n207 , \_MxM/n206 , \_MxM/n205 ,
         \_MxM/n204 , \_MxM/n203 , \_MxM/n202 , \_MxM/n201 , \_MxM/n200 ,
         \_MxM/n199 , \_MxM/n198 , \_MxM/n197 , \_MxM/n196 , \_MxM/n195 ,
         \_MxM/n194 , \_MxM/n193 , \_MxM/n192 , \_MxM/n191 , \_MxM/n190 ,
         \_MxM/n189 , \_MxM/n188 , \_MxM/N32 , \_MxM/N31 , \_MxM/N30 ,
         \_MxM/N29 , \_MxM/N28 , \_MxM/N27 , \_MxM/N26 , \_MxM/N25 ,
         \_MxM/N24 , \_MxM/N23 , \_MxM/N22 , \_MxM/N21 , \_MxM/N20 ,
         \_MxM/N19 , \_MxM/N17 , \_MxM/N16 , \_MxM/N15 , \_MxM/N14 ,
         \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 ,
         \_MxM/N7 , \_MxM/N6 , \_MxM/n[0] , \_MxM/n[1] , \_MxM/n[2] ,
         \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] , \_MxM/n[7] ,
         \_MxM/n[8] , \_MxM/n[9] , \_MxM/n[10] , \_MxM/n[11] , \_MxM/n[12] ,
         \_MxM/n[13] , \_MxM/Y0[0] , \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] ,
         \_MxM/Y0[4] , \_MxM/Y0[5] , \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/Y0[8] ,
         \_MxM/Y0[9] , \_MxM/Y0[10] , \_MxM/Y0[11] , \_MxM/Y0[12] ,
         \_MxM/Y0[13] , \_MxM/Y0[14] , \_MxM/Y0[15] , \_MxM/add_39/carry[13] ,
         \_MxM/add_39/carry[12] , \_MxM/add_39/carry[11] ,
         \_MxM/add_39/carry[10] , \_MxM/add_39/carry[9] ,
         \_MxM/add_39/carry[8] , \_MxM/add_39/carry[7] ,
         \_MxM/add_39/carry[6] , \_MxM/add_39/carry[5] ,
         \_MxM/add_39/carry[4] , \_MxM/add_39/carry[3] ,
         \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n188 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n189 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n190 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n191 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n192 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n193 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n194 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n195 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n196 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n197 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n198 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n199 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n200 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n201 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n202 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n203 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/n204 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/n205 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/n206 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/n207 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/n208 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/n209 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/n210 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/n211 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n212 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n213 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n214 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n215 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n216 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n217 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n218 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n219 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[13]  ( .D(\_MxM/N32 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[13] ) );
  DFF \_MxM/n_reg[12]  ( .D(\_MxM/N31 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[12] ) );
  DFF \_MxM/n_reg[11]  ( .D(\_MxM/N30 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[11] ) );
  DFF \_MxM/n_reg[10]  ( .D(\_MxM/N29 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[10] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/N28 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/N27 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/N26 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N25 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N24 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N23 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N22 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N21 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N20 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N19 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_39/U1_1_9  ( .IN0(\_MxM/n[9] ), .IN1(\_MxM/add_39/carry[9] ), .COUT(\_MxM/add_39/carry[10] ), .SUM(\_MxM/N14 ) );
  HADDER \_MxM/add_39/U1_1_10  ( .IN0(\_MxM/n[10] ), .IN1(
        \_MxM/add_39/carry[10] ), .COUT(\_MxM/add_39/carry[11] ), .SUM(
        \_MxM/N15 ) );
  HADDER \_MxM/add_39/U1_1_11  ( .IN0(\_MxM/n[11] ), .IN1(
        \_MxM/add_39/carry[11] ), .COUT(\_MxM/add_39/carry[12] ), .SUM(
        \_MxM/N16 ) );
  HADDER \_MxM/add_39/U1_1_12  ( .IN0(\_MxM/n[12] ), .IN1(
        \_MxM/add_39/carry[12] ), .COUT(\_MxM/add_39/carry[13] ), .SUM(
        \_MxM/N17 ) );
  MUX U1 ( .IN0(n1), .IN1(n1306), .SEL(n1307), .F(n1290) );
  IV U2 ( .A(n1308), .Z(n1) );
  MUX U3 ( .IN0(n2), .IN1(n973), .SEL(n974), .F(n950) );
  IV U4 ( .A(n975), .Z(n2) );
  MUX U5 ( .IN0(n1381), .IN1(n1399), .SEL(n1383), .F(n1362) );
  XOR U6 ( .A(n1164), .B(n1154), .Z(n970) );
  XOR U7 ( .A(n976), .B(n958), .Z(n962) );
  MUX U8 ( .IN0(n3), .IN1(n723), .SEL(n724), .F(n653) );
  IV U9 ( .A(n725), .Z(n3) );
  MUX U10 ( .IN0(n4), .IN1(n884), .SEL(n885), .F(n809) );
  IV U11 ( .A(n886), .Z(n4) );
  MUX U12 ( .IN0(n5), .IN1(n950), .SEL(n951), .F(n927) );
  IV U13 ( .A(n952), .Z(n5) );
  MUX U14 ( .IN0(n6), .IN1(n1146), .SEL(n1147), .F(n1136) );
  IV U15 ( .A(n1148), .Z(n6) );
  XOR U16 ( .A(n1149), .B(n1141), .Z(n947) );
  MUX U17 ( .IN0(n1101), .IN1(n1104), .SEL(n1102), .F(n1086) );
  MUX U18 ( .IN0(n7), .IN1(n448), .SEL(n449), .F(n397) );
  IV U19 ( .A(n450), .Z(n7) );
  MUX U20 ( .IN0(n8), .IN1(n800), .SEL(n801), .F(n723) );
  IV U21 ( .A(n802), .Z(n8) );
  XNOR U22 ( .A(n1444), .B(n1445), .Z(n888) );
  XOR U23 ( .A(n951), .B(n952), .Z(n963) );
  MUX U24 ( .IN0(n9), .IN1(n900), .SEL(n901), .F(n838) );
  IV U25 ( .A(n902), .Z(n9) );
  XOR U26 ( .A(n1137), .B(n1138), .Z(n945) );
  MUX U27 ( .IN0(n10), .IN1(n577), .SEL(n578), .F(n512) );
  IV U28 ( .A(n579), .Z(n10) );
  MUX U29 ( .IN0(e_input[8]), .IN1(n1429), .SEL(e_input[15]), .F(n460) );
  MUX U30 ( .IN0(n1142), .IN1(n11), .SEL(n1141), .F(n1133) );
  IV U31 ( .A(n1140), .Z(n11) );
  MUX U32 ( .IN0(e_input[13]), .IN1(n1455), .SEL(e_input[15]), .F(n242) );
  MUX U33 ( .IN0(n1317), .IN1(n1320), .SEL(n1318), .F(n1301) );
  MUX U34 ( .IN0(n12), .IN1(n927), .SEL(n928), .F(n908) );
  IV U35 ( .A(n929), .Z(n12) );
  MUX U36 ( .IN0(n13), .IN1(n1136), .SEL(n1137), .F(n915) );
  IV U37 ( .A(n1138), .Z(n13) );
  XOR U38 ( .A(n953), .B(n935), .Z(n939) );
  MUX U39 ( .IN0(e_input[9]), .IN1(n1430), .SEL(e_input[15]), .F(n406) );
  MUX U40 ( .IN0(n283), .IN1(n14), .SEL(n282), .F(n244) );
  IV U41 ( .A(n281), .Z(n14) );
  MUX U42 ( .IN0(e_input[11]), .IN1(n1410), .SEL(e_input[15]), .F(n312) );
  MUX U43 ( .IN0(n373), .IN1(n371), .SEL(n372), .F(n326) );
  MUX U44 ( .IN0(n15), .IN1(n166), .SEL(n165), .F(n174) );
  IV U45 ( .A(n177), .Z(n15) );
  MUX U46 ( .IN0(n16), .IN1(n1321), .SEL(n1322), .F(n1317) );
  IV U47 ( .A(n1323), .Z(n16) );
  XOR U48 ( .A(n1147), .B(n1148), .Z(n968) );
  MUX U49 ( .IN0(n17), .IN1(n704), .SEL(n705), .F(n635) );
  IV U50 ( .A(n706), .Z(n17) );
  MUX U51 ( .IN0(n18), .IN1(n763), .SEL(n764), .F(n700) );
  IV U52 ( .A(n765), .Z(n18) );
  MUX U53 ( .IN0(e_input[10]), .IN1(n1409), .SEL(e_input[15]), .F(n353) );
  MUX U54 ( .IN0(n463), .IN1(n19), .SEL(n462), .F(n408) );
  IV U55 ( .A(n461), .Z(n19) );
  MUX U56 ( .IN0(n539), .IN1(n537), .SEL(n538), .F(n472) );
  XNOR U57 ( .A(n1431), .B(n885), .Z(n889) );
  XOR U58 ( .A(n175), .B(n196), .Z(n194) );
  MUX U59 ( .IN0(n1362), .IN1(n1380), .SEL(n1364), .F(n1331) );
  MUX U60 ( .IN0(n1250), .IN1(n1272), .SEL(n1252), .F(n1232) );
  MUX U61 ( .IN0(n20), .IN1(n908), .SEL(n909), .F(n846) );
  IV U62 ( .A(n910), .Z(n20) );
  MUX U63 ( .IN0(n21), .IN1(n1153), .SEL(n1154), .F(n1140) );
  IV U64 ( .A(n1155), .Z(n21) );
  MUX U65 ( .IN0(n22), .IN1(n875), .SEL(n876), .F(n800) );
  IV U66 ( .A(n877), .Z(n22) );
  MUX U67 ( .IN0(g_input[11]), .IN1(n1184), .SEL(g_input[15]), .F(n329) );
  MUX U68 ( .IN0(n411), .IN1(n27), .SEL(n410), .F(n360) );
  MUX U69 ( .IN0(n672), .IN1(n670), .SEL(n671), .F(n602) );
  MUX U70 ( .IN0(n702), .IN1(n23), .SEL(n701), .F(n630) );
  IV U71 ( .A(n700), .Z(n23) );
  NAND U72 ( .A(n244), .B(n279), .Z(n278) );
  XOR U73 ( .A(n222), .B(n230), .Z(n228) );
  MUX U74 ( .IN0(n24), .IN1(n1168), .SEL(n1169), .F(n1153) );
  IV U75 ( .A(n1170), .Z(n24) );
  MUX U76 ( .IN0(n25), .IN1(n715), .SEL(n716), .F(n645) );
  IV U77 ( .A(n717), .Z(n25) );
  MUX U78 ( .IN0(n26), .IN1(n771), .SEL(n772), .F(n704) );
  IV U79 ( .A(n773), .Z(n26) );
  MUX U80 ( .IN0(e_input[4]), .IN1(n1115), .SEL(e_input[15]), .F(n699) );
  XOR U81 ( .A(n1411), .B(n1396), .Z(n1336) );
  MUX U82 ( .IN0(n455), .IN1(n457), .SEL(n456), .F(n27) );
  IV U83 ( .A(n27), .Z(n409) );
  MUX U84 ( .IN0(n633), .IN1(n28), .SEL(n632), .F(n560) );
  IV U85 ( .A(n631), .Z(n28) );
  MUX U86 ( .IN0(n740), .IN1(n738), .SEL(n739), .F(n670) );
  MUX U87 ( .IN0(n858), .IN1(n29), .SEL(n857), .F(n781) );
  IV U88 ( .A(n856), .Z(n29) );
  XNOR U89 ( .A(n363), .B(n323), .Z(n327) );
  XOR U90 ( .A(n253), .B(n261), .Z(n259) );
  XOR U91 ( .A(n928), .B(n929), .Z(n940) );
  MUX U92 ( .IN0(n1256), .IN1(n1266), .SEL(n1258), .F(n1242) );
  MUX U93 ( .IN0(n1331), .IN1(n1361), .SEL(n1333), .F(n867) );
  XNOR U94 ( .A(n1108), .B(n1109), .Z(n1092) );
  MUX U95 ( .IN0(g_input[9]), .IN1(n1222), .SEL(g_input[15]), .F(n423) );
  MUX U96 ( .IN0(g_input[12]), .IN1(n1166), .SEL(g_input[15]), .F(n284) );
  XOR U97 ( .A(n332), .B(n375), .Z(n333) );
  MUX U98 ( .IN0(n727), .IN1(n729), .SEL(n728), .F(n659) );
  MUX U99 ( .IN0(n769), .IN1(n767), .SEL(n768), .F(n694) );
  XOR U100 ( .A(n857), .B(n858), .Z(n864) );
  XNOR U101 ( .A(n360), .B(n403), .Z(n361) );
  XNOR U102 ( .A(n464), .B(n417), .Z(n421) );
  MUX U103 ( .IN0(n30), .IN1(n648), .SEL(n649), .F(n580) );
  IV U104 ( .A(n650), .Z(n30) );
  MUX U105 ( .IN0(n507), .IN1(n509), .SEL(n508), .F(n31) );
  IV U106 ( .A(n31), .Z(n443) );
  XOR U107 ( .A(n290), .B(n298), .Z(n296) );
  MUX U108 ( .IN0(n1248), .IN1(n32), .SEL(n1098), .F(n1229) );
  IV U109 ( .A(n1097), .Z(n32) );
  MUX U110 ( .IN0(n1094), .IN1(n1092), .SEL(n1093), .F(n1065) );
  XOR U111 ( .A(n1139), .B(n1133), .Z(n924) );
  MUX U112 ( .IN0(n33), .IN1(n867), .SEL(n868), .F(n792) );
  IV U113 ( .A(n869), .Z(n33) );
  MUX U114 ( .IN0(n34), .IN1(n915), .SEL(n916), .F(n856) );
  IV U115 ( .A(n917), .Z(n34) );
  XOR U116 ( .A(n930), .B(n901), .Z(n905) );
  MUX U117 ( .IN0(n591), .IN1(n593), .SEL(n592), .F(n526) );
  MUX U118 ( .IN0(n817), .IN1(n815), .SEL(n816), .F(n738) );
  XOR U119 ( .A(n1337), .B(n876), .Z(n880) );
  XNOR U120 ( .A(n412), .B(n368), .Z(n372) );
  MUX U121 ( .IN0(n35), .IN1(n451), .SEL(n452), .F(n400) );
  IV U122 ( .A(n453), .Z(n35) );
  MUX U123 ( .IN0(n36), .IN1(n566), .SEL(n567), .F(n506) );
  IV U124 ( .A(n568), .Z(n36) );
  NAND U125 ( .A(n630), .B(n698), .Z(n697) );
  MUX U126 ( .IN0(n572), .IN1(n574), .SEL(n573), .F(n507) );
  MUX U127 ( .IN0(n37), .IN1(n546), .SEL(n547), .F(n481) );
  IV U128 ( .A(\_MxM/Y0[5] ), .Z(n37) );
  XOR U129 ( .A(n335), .B(n343), .Z(n341) );
  MUX U130 ( .IN0(n38), .IN1(n1301), .SEL(n1302), .F(n1284) );
  IV U131 ( .A(n1303), .Z(n38) );
  MUX U132 ( .IN0(g_input[1]), .IN1(n1457), .SEL(g_input[15]), .F(n1111) );
  MUX U133 ( .IN0(n39), .IN1(n512), .SEL(n513), .F(n448) );
  IV U134 ( .A(n514), .Z(n39) );
  MUX U135 ( .IN0(g_input[6]), .IN1(n1353), .SEL(g_input[15]), .F(n605) );
  MUX U136 ( .IN0(g_input[7]), .IN1(n1340), .SEL(g_input[15]), .F(n540) );
  MUX U137 ( .IN0(g_input[5]), .IN1(n1373), .SEL(g_input[15]), .F(n673) );
  MUX U138 ( .IN0(n40), .IN1(n846), .SEL(n847), .F(n771) );
  IV U139 ( .A(n848), .Z(n40) );
  XOR U140 ( .A(n916), .B(n917), .Z(n922) );
  MUX U141 ( .IN0(n659), .IN1(n661), .SEL(n660), .F(n591) );
  XNOR U142 ( .A(n898), .B(n839), .Z(n843) );
  XOR U143 ( .A(n250), .B(n285), .Z(n251) );
  MUX U144 ( .IN0(n41), .IN1(n315), .SEL(n316), .F(n268) );
  IV U145 ( .A(n317), .Z(n41) );
  NAND U146 ( .A(n408), .B(n459), .Z(n458) );
  MUX U147 ( .IN0(n562), .IN1(n560), .SEL(n561), .F(n504) );
  XNOR U148 ( .A(n594), .B(n534), .Z(n538) );
  MUX U149 ( .IN0(n42), .IN1(n795), .SEL(n796), .F(n718) );
  IV U150 ( .A(n797), .Z(n42) );
  MUX U151 ( .IN0(n43), .IN1(n642), .SEL(n641), .F(n572) );
  IV U152 ( .A(n640), .Z(n43) );
  MUX U153 ( .IN0(n44), .IN1(n611), .SEL(n612), .F(n546) );
  IV U154 ( .A(\_MxM/Y0[4] ), .Z(n44) );
  XOR U155 ( .A(n380), .B(n388), .Z(n386) );
  MUX U156 ( .IN0(n1065), .IN1(n45), .SEL(n1066), .F(n1038) );
  IV U157 ( .A(n1067), .Z(n45) );
  MUX U158 ( .IN0(n1157), .IN1(n46), .SEL(n970), .F(n1144) );
  IV U159 ( .A(n968), .Z(n46) );
  XNOR U160 ( .A(n1322), .B(n1323), .Z(n1309) );
  MUX U161 ( .IN0(n47), .IN1(n645), .SEL(n646), .F(n577) );
  IV U162 ( .A(n647), .Z(n47) );
  MUX U163 ( .IN0(g_input[3]), .IN1(n1434), .SEL(g_input[15]), .F(n48) );
  IV U164 ( .A(n48), .Z(n818) );
  MUX U165 ( .IN0(g_input[4]), .IN1(n1391), .SEL(g_input[15]), .F(n49) );
  IV U166 ( .A(n49), .Z(n741) );
  MUX U167 ( .IN0(n904), .IN1(n50), .SEL(n905), .F(n842) );
  IV U168 ( .A(n906), .Z(n50) );
  XOR U169 ( .A(n1235), .B(n1236), .Z(n1097) );
  MUX U170 ( .IN0(n328), .IN1(n326), .SEL(n327), .F(n273) );
  MUX U171 ( .IN0(n51), .IN1(n635), .SEL(n636), .F(n566) );
  IV U172 ( .A(n637), .Z(n51) );
  XOR U173 ( .A(n543), .B(n606), .Z(n544) );
  MUX U174 ( .IN0(n804), .IN1(n806), .SEL(n805), .F(n727) );
  MUX U175 ( .IN0(n890), .IN1(n888), .SEL(n889), .F(n815) );
  MUX U176 ( .IN0(n52), .IN1(n357), .SEL(n358), .F(n315) );
  IV U177 ( .A(n359), .Z(n52) );
  XOR U178 ( .A(n518), .B(n462), .Z(n456) );
  XNOR U179 ( .A(n529), .B(n469), .Z(n473) );
  MUX U180 ( .IN0(n53), .IN1(n580), .SEL(n581), .F(n515) );
  IV U181 ( .A(n582), .Z(n53) );
  XOR U182 ( .A(n693), .B(n631), .Z(n632) );
  MUX U183 ( .IN0(n789), .IN1(n54), .SEL(n788), .F(n710) );
  IV U184 ( .A(n787), .Z(n54) );
  MUX U185 ( .IN0(n707), .IN1(n55), .SEL(n708), .F(n640) );
  IV U186 ( .A(n709), .Z(n55) );
  MUX U187 ( .IN0(n56), .IN1(n679), .SEL(n680), .F(n611) );
  IV U188 ( .A(\_MxM/Y0[3] ), .Z(n56) );
  XOR U189 ( .A(n435), .B(n441), .Z(n430) );
  MUX U190 ( .IN0(n57), .IN1(n1095), .SEL(n912), .F(n1068) );
  IV U191 ( .A(n911), .Z(n57) );
  MUX U192 ( .IN0(n1011), .IN1(n58), .SEL(n1012), .F(n984) );
  IV U193 ( .A(n1013), .Z(n58) );
  MUX U194 ( .IN0(e_input[1]), .IN1(n59), .SEL(e_input[15]), .F(n1128) );
  IV U195 ( .A(n1328), .Z(n59) );
  MUX U196 ( .IN0(e_input[6]), .IN1(n1120), .SEL(e_input[15]), .F(n565) );
  MUX U197 ( .IN0(e_input[3]), .IN1(n1314), .SEL(e_input[15]), .F(n784) );
  MUX U198 ( .IN0(n879), .IN1(n881), .SEL(n880), .F(n804) );
  MUX U199 ( .IN0(e_input[14]), .IN1(n1460), .SEL(e_input[15]), .F(n211) );
  NAND U200 ( .A(n309), .B(n352), .Z(n351) );
  XOR U201 ( .A(n583), .B(n523), .Z(n527) );
  XNOR U202 ( .A(n662), .B(n599), .Z(n603) );
  MUX U203 ( .IN0(n60), .IN1(n718), .SEL(n719), .F(n648) );
  IV U204 ( .A(n720), .Z(n60) );
  XNOR U205 ( .A(n761), .B(n701), .Z(n695) );
  MUX U206 ( .IN0(n774), .IN1(n61), .SEL(n775), .F(n707) );
  IV U207 ( .A(n776), .Z(n61) );
  MUX U208 ( .IN0(n62), .IN1(n253), .SEL(n254), .F(n222) );
  IV U209 ( .A(\_MxM/Y0[11] ), .Z(n62) );
  XOR U210 ( .A(n481), .B(n489), .Z(n487) );
  MUX U211 ( .IN0(n1229), .IN1(n63), .SEL(n1074), .F(n1210) );
  IV U212 ( .A(n1072), .Z(n63) );
  MUX U213 ( .IN0(n1284), .IN1(n1300), .SEL(n1286), .F(n1267) );
  MUX U214 ( .IN0(n961), .IN1(n64), .SEL(n962), .F(n938) );
  IV U215 ( .A(n963), .Z(n64) );
  XOR U216 ( .A(n909), .B(n910), .Z(n906) );
  XOR U217 ( .A(n1307), .B(n1308), .Z(n1122) );
  MUX U218 ( .IN0(n65), .IN1(n792), .SEL(n793), .F(n715) );
  IV U219 ( .A(n794), .Z(n65) );
  MUX U220 ( .IN0(g_input[10]), .IN1(n1202), .SEL(g_input[15]), .F(n374) );
  XNOR U221 ( .A(n1099), .B(n1089), .Z(n1093) );
  XOR U222 ( .A(n426), .B(n476), .Z(n427) );
  MUX U223 ( .IN0(n474), .IN1(n472), .SEL(n473), .F(n420) );
  MUX U224 ( .IN0(n696), .IN1(n694), .SEL(n695), .F(n631) );
  MUX U225 ( .IN0(g_input[13]), .IN1(n1152), .SEL(g_input[15]), .F(n247) );
  MUX U226 ( .IN0(n66), .IN1(n515), .SEL(n516), .F(n451) );
  IV U227 ( .A(n517), .Z(n66) );
  XOR U228 ( .A(n651), .B(n588), .Z(n592) );
  XNOR U229 ( .A(n807), .B(n735), .Z(n739) );
  MUX U230 ( .IN0(n67), .IN1(n870), .SEL(n871), .F(n795) );
  IV U231 ( .A(n872), .Z(n67) );
  MUX U232 ( .IN0(n68), .IN1(n859), .SEL(n860), .F(n787) );
  IV U233 ( .A(n861), .Z(n68) );
  MUX U234 ( .IN0(g_input[14]), .IN1(n1129), .SEL(g_input[15]), .F(n212) );
  MUX U235 ( .IN0(n270), .IN1(n69), .SEL(n269), .F(n238) );
  IV U236 ( .A(n268), .Z(n69) );
  XNOR U237 ( .A(n572), .B(n571), .Z(n624) );
  MUX U238 ( .IN0(\_MxM/Y0[13] ), .IN1(n70), .SEL(n176), .F(n168) );
  IV U239 ( .A(n175), .Z(n70) );
  MUX U240 ( .IN0(n71), .IN1(n335), .SEL(n336), .F(n290) );
  IV U241 ( .A(\_MxM/Y0[9] ), .Z(n71) );
  MUX U242 ( .IN0(n72), .IN1(n824), .SEL(n825), .F(n747) );
  IV U243 ( .A(\_MxM/Y0[1] ), .Z(n72) );
  XOR U244 ( .A(n546), .B(n554), .Z(n552) );
  MUX U245 ( .IN0(n1210), .IN1(n73), .SEL(n1047), .F(n1191) );
  IV U246 ( .A(n1045), .Z(n73) );
  MUX U247 ( .IN0(n984), .IN1(n74), .SEL(n985), .F(n961) );
  IV U248 ( .A(n986), .Z(n74) );
  MUX U249 ( .IN0(n1267), .IN1(n1283), .SEL(n1269), .F(n1256) );
  MUX U250 ( .IN0(n1144), .IN1(n75), .SEL(n947), .F(n1134) );
  IV U251 ( .A(n945), .Z(n75) );
  MUX U252 ( .IN0(g_input[8]), .IN1(n1240), .SEL(g_input[15]), .F(n475) );
  MUX U253 ( .IN0(g_input[2]), .IN1(n1447), .SEL(g_input[15]), .F(n891) );
  MUX U254 ( .IN0(n76), .IN1(n838), .SEL(n839), .F(n763) );
  IV U255 ( .A(n840), .Z(n76) );
  MUX U256 ( .IN0(n77), .IN1(n397), .SEL(n398), .F(n354) );
  IV U257 ( .A(n399), .Z(n77) );
  MUX U258 ( .IN0(n526), .IN1(n528), .SEL(n527), .F(n455) );
  MUX U259 ( .IN0(n604), .IN1(n602), .SEL(n603), .F(n537) );
  XOR U260 ( .A(n821), .B(n892), .Z(n822) );
  MUX U261 ( .IN0(n844), .IN1(n842), .SEL(n843), .F(n767) );
  XNOR U262 ( .A(n273), .B(n274), .Z(n272) );
  MUX U263 ( .IN0(n78), .IN1(n400), .SEL(n401), .F(n357) );
  IV U264 ( .A(n402), .Z(n78) );
  XOR U265 ( .A(n567), .B(n568), .Z(n562) );
  XOR U266 ( .A(n798), .B(n724), .Z(n728) );
  XNOR U267 ( .A(n882), .B(n812), .Z(n816) );
  NAND U268 ( .A(n781), .B(n854), .Z(n853) );
  XNOR U269 ( .A(n277), .B(n276), .Z(n270) );
  XNOR U270 ( .A(n672), .B(n671), .Z(n650) );
  MUX U271 ( .IN0(n712), .IN1(n710), .SEL(n711), .F(n79) );
  IV U272 ( .A(n79), .Z(n639) );
  MUX U273 ( .IN0(n849), .IN1(n80), .SEL(n850), .F(n774) );
  IV U274 ( .A(n851), .Z(n80) );
  MUX U275 ( .IN0(n443), .IN1(n81), .SEL(n444), .F(n394) );
  IV U276 ( .A(n445), .Z(n81) );
  MUX U277 ( .IN0(n82), .IN1(n222), .SEL(n223), .F(n175) );
  IV U278 ( .A(\_MxM/Y0[12] ), .Z(n82) );
  MUX U279 ( .IN0(n83), .IN1(n380), .SEL(n381), .F(n335) );
  IV U280 ( .A(\_MxM/Y0[8] ), .Z(n83) );
  XOR U281 ( .A(n611), .B(n619), .Z(n617) );
  MUX U282 ( .IN0(n1191), .IN1(n84), .SEL(n1020), .F(n1172) );
  IV U283 ( .A(n1018), .Z(n84) );
  MUX U284 ( .IN0(n85), .IN1(n1335), .SEL(n1336), .F(n1385) );
  IV U285 ( .A(n1405), .Z(n85) );
  NOR U286 ( .A(g_input[0]), .B(n1457), .Z(n1448) );
  XOR U287 ( .A(n1315), .B(n1302), .Z(n1123) );
  MUX U288 ( .IN0(n1134), .IN1(n86), .SEL(n924), .F(n862) );
  IV U289 ( .A(n922), .Z(n86) );
  MUX U290 ( .IN0(n422), .IN1(n420), .SEL(n421), .F(n371) );
  XOR U291 ( .A(n676), .B(n742), .Z(n677) );
  MUX U292 ( .IN0(n356), .IN1(n87), .SEL(n355), .F(n309) );
  IV U293 ( .A(n354), .Z(n87) );
  MUX U294 ( .IN0(e_input[7]), .IN1(n1121), .SEL(e_input[15]), .F(n498) );
  XNOR U295 ( .A(n730), .B(n667), .Z(n671) );
  XOR U296 ( .A(n721), .B(n656), .Z(n660) );
  XNOR U297 ( .A(n836), .B(n764), .Z(n768) );
  XNOR U298 ( .A(n890), .B(n889), .Z(n872) );
  MUX U299 ( .IN0(n246), .IN1(n272), .SEL(n245), .F(n217) );
  XNOR U300 ( .A(n328), .B(n327), .Z(n317) );
  XNOR U301 ( .A(n539), .B(n538), .Z(n517) );
  XNOR U302 ( .A(n604), .B(n603), .Z(n582) );
  XNOR U303 ( .A(n710), .B(n777), .Z(n711) );
  XNOR U304 ( .A(n453), .B(n452), .Z(n445) );
  XOR U305 ( .A(n559), .B(n500), .Z(n508) );
  XNOR U306 ( .A(n720), .B(n719), .Z(n709) );
  XNOR U307 ( .A(n797), .B(n796), .Z(n776) );
  XNOR U308 ( .A(n236), .B(n235), .Z(n260) );
  MUX U309 ( .IN0(n88), .IN1(n429), .SEL(n430), .F(n380) );
  IV U310 ( .A(\_MxM/Y0[7] ), .Z(n88) );
  MUX U311 ( .IN0(\_MxM/Y0[14] ), .IN1(n168), .SEL(n169), .F(n158) );
  XOR U312 ( .A(n679), .B(n687), .Z(n685) );
  MUX U313 ( .IN0(n1038), .IN1(n89), .SEL(n1039), .F(n1011) );
  IV U314 ( .A(n1040), .Z(n89) );
  MUX U315 ( .IN0(n90), .IN1(n1122), .SEL(n1123), .F(n1295) );
  IV U316 ( .A(n1309), .Z(n90) );
  MUX U317 ( .IN0(n1172), .IN1(n91), .SEL(n993), .F(n1157) );
  IV U318 ( .A(n991), .Z(n91) );
  XOR U319 ( .A(n1433), .B(g_input[3]), .Z(n1434) );
  MUX U320 ( .IN0(n938), .IN1(n92), .SEL(n939), .F(n904) );
  IV U321 ( .A(n940), .Z(n92) );
  XOR U322 ( .A(n1403), .B(n1404), .Z(n1335) );
  XOR U323 ( .A(n1254), .B(n1245), .Z(n1098) );
  MUX U324 ( .IN0(e_input[5]), .IN1(n1116), .SEL(e_input[15]), .F(n628) );
  MUX U325 ( .IN0(e_input[2]), .IN1(n1313), .SEL(e_input[15]), .F(n855) );
  XNOR U326 ( .A(n1094), .B(n1093), .Z(n911) );
  XNOR U327 ( .A(n318), .B(n282), .Z(n276) );
  MUX U328 ( .IN0(n362), .IN1(n360), .SEL(n361), .F(n93) );
  IV U329 ( .A(n93), .Z(n314) );
  XOR U330 ( .A(n636), .B(n637), .Z(n633) );
  XOR U331 ( .A(n873), .B(n801), .Z(n805) );
  MUX U332 ( .IN0(n864), .IN1(n1124), .SEL(n863), .F(n786) );
  XNOR U333 ( .A(n844), .B(n843), .Z(n861) );
  AND U334 ( .A(n206), .B(n183), .Z(n205) );
  XNOR U335 ( .A(n373), .B(n372), .Z(n359) );
  XNOR U336 ( .A(n422), .B(n421), .Z(n402) );
  XNOR U337 ( .A(n474), .B(n473), .Z(n453) );
  XNOR U338 ( .A(n696), .B(n695), .Z(n712) );
  XNOR U339 ( .A(n740), .B(n739), .Z(n720) );
  XNOR U340 ( .A(n817), .B(n816), .Z(n797) );
  XNOR U341 ( .A(n769), .B(n768), .Z(n789) );
  XNOR U342 ( .A(n872), .B(n871), .Z(n851) );
  XNOR U343 ( .A(n237), .B(n238), .Z(n236) );
  XNOR U344 ( .A(n517), .B(n516), .Z(n509) );
  XNOR U345 ( .A(n582), .B(n581), .Z(n574) );
  XNOR U346 ( .A(n650), .B(n649), .Z(n642) );
  MUX U347 ( .IN0(n94), .IN1(n290), .SEL(n291), .F(n253) );
  IV U348 ( .A(\_MxM/Y0[10] ), .Z(n94) );
  MUX U349 ( .IN0(n95), .IN1(n481), .SEL(n482), .F(n429) );
  IV U350 ( .A(\_MxM/Y0[6] ), .Z(n95) );
  MUX U351 ( .IN0(n96), .IN1(n747), .SEL(n748), .F(n679) );
  IV U352 ( .A(\_MxM/Y0[2] ), .Z(n96) );
  MUX U353 ( .IN0(\_MxM/Y0[15] ), .IN1(n158), .SEL(n159), .F(n97) );
  IV U354 ( .A(n97), .Z(n155) );
  XOR U355 ( .A(n825), .B(\_MxM/Y0[1] ), .Z(n100) );
  NAND U356 ( .A(n98), .B(n99), .Z(\_MxM/n219 ) );
  OR U357 ( .A(n100), .B(n101), .Z(n99) );
  NANDN U358 ( .B(n102), .A(\_MxM/Y0[0] ), .Z(n98) );
  NAND U359 ( .A(n103), .B(n104), .Z(\_MxM/n218 ) );
  NANDN U360 ( .B(n101), .A(n105), .Z(n104) );
  NANDN U361 ( .B(n106), .A(rst), .Z(n103) );
  NAND U362 ( .A(n107), .B(n108), .Z(\_MxM/n217 ) );
  NANDN U363 ( .B(n101), .A(n109), .Z(n108) );
  NANDN U364 ( .B(n102), .A(\_MxM/Y0[2] ), .Z(n107) );
  NAND U365 ( .A(n110), .B(n111), .Z(\_MxM/n216 ) );
  NANDN U366 ( .B(n101), .A(n112), .Z(n111) );
  NANDN U367 ( .B(n102), .A(\_MxM/Y0[3] ), .Z(n110) );
  NAND U368 ( .A(n113), .B(n114), .Z(\_MxM/n215 ) );
  NANDN U369 ( .B(n101), .A(n115), .Z(n114) );
  NANDN U370 ( .B(n102), .A(\_MxM/Y0[4] ), .Z(n113) );
  NAND U371 ( .A(n116), .B(n117), .Z(\_MxM/n214 ) );
  NANDN U372 ( .B(n101), .A(n118), .Z(n117) );
  NANDN U373 ( .B(n102), .A(\_MxM/Y0[5] ), .Z(n116) );
  NAND U374 ( .A(n119), .B(n120), .Z(\_MxM/n213 ) );
  NANDN U375 ( .B(n101), .A(n121), .Z(n120) );
  NANDN U376 ( .B(n102), .A(\_MxM/Y0[6] ), .Z(n119) );
  NAND U377 ( .A(n122), .B(n123), .Z(\_MxM/n212 ) );
  NANDN U378 ( .B(n101), .A(n124), .Z(n123) );
  NANDN U379 ( .B(n102), .A(\_MxM/Y0[7] ), .Z(n122) );
  NAND U380 ( .A(n125), .B(n126), .Z(\_MxM/n211 ) );
  NANDN U381 ( .B(n101), .A(n127), .Z(n126) );
  NANDN U382 ( .B(n102), .A(\_MxM/Y0[8] ), .Z(n125) );
  NAND U383 ( .A(n128), .B(n129), .Z(\_MxM/n210 ) );
  NANDN U384 ( .B(n101), .A(n130), .Z(n129) );
  NANDN U385 ( .B(n102), .A(\_MxM/Y0[9] ), .Z(n128) );
  NAND U386 ( .A(n131), .B(n132), .Z(\_MxM/n209 ) );
  NANDN U387 ( .B(n101), .A(n133), .Z(n132) );
  NANDN U388 ( .B(n102), .A(\_MxM/Y0[10] ), .Z(n131) );
  NAND U389 ( .A(n134), .B(n135), .Z(\_MxM/n208 ) );
  NANDN U390 ( .B(n101), .A(n136), .Z(n135) );
  NANDN U391 ( .B(n102), .A(\_MxM/Y0[11] ), .Z(n134) );
  NAND U392 ( .A(n137), .B(n138), .Z(\_MxM/n207 ) );
  NANDN U393 ( .B(n101), .A(n139), .Z(n138) );
  NANDN U394 ( .B(n102), .A(\_MxM/Y0[12] ), .Z(n137) );
  NAND U395 ( .A(n140), .B(n141), .Z(\_MxM/n206 ) );
  NANDN U396 ( .B(n101), .A(n142), .Z(n141) );
  NANDN U397 ( .B(n102), .A(\_MxM/Y0[13] ), .Z(n140) );
  NAND U398 ( .A(n143), .B(n144), .Z(\_MxM/n205 ) );
  OR U399 ( .A(n145), .B(n101), .Z(n144) );
  NANDN U400 ( .B(n102), .A(\_MxM/Y0[14] ), .Z(n143) );
  NAND U401 ( .A(n146), .B(n147), .Z(\_MxM/n204 ) );
  OR U402 ( .A(n101), .B(n148), .Z(n147) );
  NANDN U403 ( .B(n149), .A(n102), .Z(n101) );
  NANDN U404 ( .B(n102), .A(\_MxM/Y0[15] ), .Z(n146) );
  NAND U405 ( .A(n150), .B(n151), .Z(\_MxM/n203 ) );
  NANDN U406 ( .B(n102), .A(o[15]), .Z(n151) );
  AND U407 ( .A(n152), .B(n153), .Z(n150) );
  NANDN U408 ( .B(n149), .A(o[15]), .Z(n153) );
  OR U409 ( .A(n148), .B(n154), .Z(n152) );
  XOR U410 ( .A(n155), .B(n156), .Z(n148) );
  XNOR U411 ( .A(\_MxM/Y0[15] ), .B(n157), .Z(n156) );
  NAND U412 ( .A(n160), .B(n161), .Z(\_MxM/n202 ) );
  NANDN U413 ( .B(n102), .A(o[14]), .Z(n161) );
  AND U414 ( .A(n162), .B(n163), .Z(n160) );
  NANDN U415 ( .B(n149), .A(o[14]), .Z(n163) );
  OR U416 ( .A(n145), .B(n154), .Z(n162) );
  XOR U417 ( .A(n159), .B(\_MxM/Y0[15] ), .Z(n145) );
  XOR U418 ( .A(n158), .B(n157), .Z(n159) );
  NAND U419 ( .A(n164), .B(n165), .Z(n157) );
  OR U420 ( .A(n166), .B(n167), .Z(n164) );
  NAND U421 ( .A(n170), .B(n171), .Z(\_MxM/n201 ) );
  NANDN U422 ( .B(n102), .A(o[13]), .Z(n171) );
  AND U423 ( .A(n172), .B(n173), .Z(n170) );
  NANDN U424 ( .B(n149), .A(o[13]), .Z(n173) );
  NANDN U425 ( .B(n154), .A(n142), .Z(n172) );
  XNOR U426 ( .A(n169), .B(\_MxM/Y0[14] ), .Z(n142) );
  XNOR U427 ( .A(n174), .B(n168), .Z(n169) );
  XNOR U428 ( .A(n167), .B(n177), .Z(n166) );
  OR U429 ( .A(n178), .B(n179), .Z(n167) );
  AND U430 ( .A(n180), .B(n181), .Z(n177) );
  OR U431 ( .A(n182), .B(n183), .Z(n181) );
  AND U432 ( .A(n184), .B(n185), .Z(n180) );
  OR U433 ( .A(n186), .B(n187), .Z(n185) );
  OR U434 ( .A(n188), .B(n189), .Z(n184) );
  NAND U435 ( .A(n190), .B(n191), .Z(\_MxM/n200 ) );
  NANDN U436 ( .B(n102), .A(o[12]), .Z(n191) );
  AND U437 ( .A(n192), .B(n193), .Z(n190) );
  NANDN U438 ( .B(n149), .A(o[12]), .Z(n193) );
  NANDN U439 ( .B(n154), .A(n139), .Z(n192) );
  XNOR U440 ( .A(n176), .B(\_MxM/Y0[13] ), .Z(n139) );
  XNOR U441 ( .A(n194), .B(n195), .Z(n176) );
  AND U442 ( .A(n165), .B(n197), .Z(n196) );
  XOR U443 ( .A(n178), .B(n198), .Z(n197) );
  XOR U444 ( .A(n198), .B(n179), .Z(n178) );
  OR U445 ( .A(n199), .B(n200), .Z(n179) );
  IV U446 ( .A(n195), .Z(n198) );
  XNOR U447 ( .A(n189), .B(n188), .Z(n195) );
  OR U448 ( .A(n201), .B(n202), .Z(n188) );
  AND U449 ( .A(n203), .B(n204), .Z(n189) );
  XNOR U450 ( .A(n182), .B(n205), .Z(n204) );
  NAND U451 ( .A(n207), .B(n208), .Z(n183) );
  NANDN U452 ( .B(n209), .A(n210), .Z(n207) );
  NANDN U453 ( .B(n186), .A(n211), .Z(n206) );
  NANDN U454 ( .B(n187), .A(n212), .Z(n182) );
  AND U455 ( .A(n213), .B(n214), .Z(n203) );
  OR U456 ( .A(n215), .B(n216), .Z(n214) );
  XNOR U457 ( .A(n217), .B(n218), .Z(n213) );
  ANDN U458 ( .A(n219), .B(n220), .Z(n218) );
  XOR U459 ( .A(n217), .B(n221), .Z(n219) );
  NAND U460 ( .A(n224), .B(n225), .Z(\_MxM/n199 ) );
  NANDN U461 ( .B(n102), .A(o[11]), .Z(n225) );
  AND U462 ( .A(n226), .B(n227), .Z(n224) );
  NANDN U463 ( .B(n149), .A(o[11]), .Z(n227) );
  NANDN U464 ( .B(n154), .A(n136), .Z(n226) );
  XNOR U465 ( .A(n223), .B(\_MxM/Y0[12] ), .Z(n136) );
  XNOR U466 ( .A(n228), .B(n229), .Z(n223) );
  AND U467 ( .A(n165), .B(n231), .Z(n230) );
  XOR U468 ( .A(n199), .B(n232), .Z(n231) );
  XOR U469 ( .A(n232), .B(n200), .Z(n199) );
  OR U470 ( .A(n233), .B(n234), .Z(n200) );
  IV U471 ( .A(n229), .Z(n232) );
  XNOR U472 ( .A(n202), .B(n201), .Z(n229) );
  OR U473 ( .A(n235), .B(n236), .Z(n201) );
  XNOR U474 ( .A(n216), .B(n215), .Z(n202) );
  OR U475 ( .A(n237), .B(n238), .Z(n215) );
  XOR U476 ( .A(n221), .B(n220), .Z(n216) );
  XOR U477 ( .A(n217), .B(n239), .Z(n220) );
  AND U478 ( .A(n240), .B(n241), .Z(n239) );
  NANDN U479 ( .B(n186), .A(n242), .Z(n241) );
  OR U480 ( .A(n243), .B(n244), .Z(n240) );
  XOR U481 ( .A(n209), .B(n210), .Z(n221) );
  NANDN U482 ( .B(n187), .A(n247), .Z(n210) );
  XNOR U483 ( .A(n208), .B(n248), .Z(n209) );
  AND U484 ( .A(n212), .B(n211), .Z(n248) );
  ANDN U485 ( .A(n249), .B(n250), .Z(n208) );
  NANDN U486 ( .B(n251), .A(n252), .Z(n249) );
  NAND U487 ( .A(n255), .B(n256), .Z(\_MxM/n198 ) );
  NANDN U488 ( .B(n102), .A(o[10]), .Z(n256) );
  AND U489 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U490 ( .B(n149), .A(o[10]), .Z(n258) );
  NANDN U491 ( .B(n154), .A(n133), .Z(n257) );
  XNOR U492 ( .A(n254), .B(\_MxM/Y0[11] ), .Z(n133) );
  XNOR U493 ( .A(n259), .B(n260), .Z(n254) );
  AND U494 ( .A(n165), .B(n262), .Z(n261) );
  XOR U495 ( .A(n233), .B(n263), .Z(n262) );
  XOR U496 ( .A(n263), .B(n234), .Z(n233) );
  OR U497 ( .A(n264), .B(n265), .Z(n234) );
  IV U498 ( .A(n260), .Z(n263) );
  OR U499 ( .A(n266), .B(n267), .Z(n235) );
  XOR U500 ( .A(n246), .B(n245), .Z(n237) );
  XNOR U501 ( .A(n271), .B(n272), .Z(n245) );
  ANDN U502 ( .A(n275), .B(n276), .Z(n274) );
  XOR U503 ( .A(n273), .B(n277), .Z(n275) );
  XNOR U504 ( .A(n278), .B(n243), .Z(n271) );
  NAND U505 ( .A(n242), .B(n212), .Z(n243) );
  NANDN U506 ( .B(n186), .A(n280), .Z(n279) );
  XOR U507 ( .A(n251), .B(n252), .Z(n246) );
  NANDN U508 ( .B(n187), .A(n284), .Z(n252) );
  AND U509 ( .A(n247), .B(n211), .Z(n285) );
  NAND U510 ( .A(n286), .B(n287), .Z(n250) );
  NANDN U511 ( .B(n288), .A(n289), .Z(n286) );
  NAND U512 ( .A(n292), .B(n293), .Z(\_MxM/n197 ) );
  NANDN U513 ( .B(n102), .A(o[9]), .Z(n293) );
  AND U514 ( .A(n294), .B(n295), .Z(n292) );
  NANDN U515 ( .B(n149), .A(o[9]), .Z(n295) );
  NANDN U516 ( .B(n154), .A(n130), .Z(n294) );
  XNOR U517 ( .A(n291), .B(\_MxM/Y0[10] ), .Z(n130) );
  XNOR U518 ( .A(n296), .B(n297), .Z(n291) );
  AND U519 ( .A(n165), .B(n299), .Z(n298) );
  XOR U520 ( .A(n264), .B(n300), .Z(n299) );
  XOR U521 ( .A(n300), .B(n265), .Z(n264) );
  OR U522 ( .A(n301), .B(n302), .Z(n265) );
  IV U523 ( .A(n297), .Z(n300) );
  XNOR U524 ( .A(n267), .B(n266), .Z(n297) );
  OR U525 ( .A(n303), .B(n304), .Z(n266) );
  XNOR U526 ( .A(n270), .B(n269), .Z(n267) );
  XOR U527 ( .A(n268), .B(n305), .Z(n269) );
  AND U528 ( .A(n306), .B(n307), .Z(n305) );
  OR U529 ( .A(n308), .B(n309), .Z(n307) );
  AND U530 ( .A(n310), .B(n311), .Z(n306) );
  NANDN U531 ( .B(n186), .A(n312), .Z(n311) );
  NAND U532 ( .A(n313), .B(n314), .Z(n310) );
  XNOR U533 ( .A(n281), .B(n319), .Z(n282) );
  AND U534 ( .A(n212), .B(n280), .Z(n319) );
  XOR U535 ( .A(n320), .B(n321), .Z(n281) );
  ANDN U536 ( .A(n322), .B(n323), .Z(n321) );
  XNOR U537 ( .A(n324), .B(n320), .Z(n322) );
  XOR U538 ( .A(n325), .B(n283), .Z(n318) );
  NAND U539 ( .A(n242), .B(n247), .Z(n283) );
  IV U540 ( .A(n273), .Z(n325) );
  XNOR U541 ( .A(n288), .B(n289), .Z(n277) );
  NANDN U542 ( .B(n187), .A(n329), .Z(n289) );
  XNOR U543 ( .A(n287), .B(n330), .Z(n288) );
  AND U544 ( .A(n284), .B(n211), .Z(n330) );
  ANDN U545 ( .A(n331), .B(n332), .Z(n287) );
  NANDN U546 ( .B(n333), .A(n334), .Z(n331) );
  NAND U547 ( .A(n337), .B(n338), .Z(\_MxM/n196 ) );
  NANDN U548 ( .B(n102), .A(o[8]), .Z(n338) );
  AND U549 ( .A(n339), .B(n340), .Z(n337) );
  NANDN U550 ( .B(n149), .A(o[8]), .Z(n340) );
  NANDN U551 ( .B(n154), .A(n127), .Z(n339) );
  XNOR U552 ( .A(n336), .B(\_MxM/Y0[9] ), .Z(n127) );
  XNOR U553 ( .A(n341), .B(n342), .Z(n336) );
  AND U554 ( .A(n165), .B(n344), .Z(n343) );
  XOR U555 ( .A(n301), .B(n345), .Z(n344) );
  XOR U556 ( .A(n345), .B(n302), .Z(n301) );
  OR U557 ( .A(n346), .B(n347), .Z(n302) );
  IV U558 ( .A(n342), .Z(n345) );
  XNOR U559 ( .A(n304), .B(n303), .Z(n342) );
  OR U560 ( .A(n348), .B(n349), .Z(n303) );
  XNOR U561 ( .A(n317), .B(n316), .Z(n304) );
  XOR U562 ( .A(n350), .B(n313), .Z(n316) );
  XNOR U563 ( .A(n351), .B(n308), .Z(n313) );
  NAND U564 ( .A(n312), .B(n212), .Z(n308) );
  NANDN U565 ( .B(n186), .A(n353), .Z(n352) );
  XNOR U566 ( .A(n314), .B(n315), .Z(n350) );
  XNOR U567 ( .A(n320), .B(n364), .Z(n323) );
  AND U568 ( .A(n247), .B(n280), .Z(n364) );
  XOR U569 ( .A(n365), .B(n366), .Z(n320) );
  ANDN U570 ( .A(n367), .B(n368), .Z(n366) );
  XNOR U571 ( .A(n369), .B(n365), .Z(n367) );
  XOR U572 ( .A(n370), .B(n324), .Z(n363) );
  NAND U573 ( .A(n242), .B(n284), .Z(n324) );
  IV U574 ( .A(n326), .Z(n370) );
  XNOR U575 ( .A(n333), .B(n334), .Z(n328) );
  NANDN U576 ( .B(n187), .A(n374), .Z(n334) );
  AND U577 ( .A(n329), .B(n211), .Z(n375) );
  NAND U578 ( .A(n376), .B(n377), .Z(n332) );
  NANDN U579 ( .B(n378), .A(n379), .Z(n376) );
  NAND U580 ( .A(n382), .B(n383), .Z(\_MxM/n195 ) );
  NANDN U581 ( .B(n102), .A(o[7]), .Z(n383) );
  AND U582 ( .A(n384), .B(n385), .Z(n382) );
  NANDN U583 ( .B(n149), .A(o[7]), .Z(n385) );
  NANDN U584 ( .B(n154), .A(n124), .Z(n384) );
  XNOR U585 ( .A(n381), .B(\_MxM/Y0[8] ), .Z(n124) );
  XNOR U586 ( .A(n386), .B(n387), .Z(n381) );
  AND U587 ( .A(n165), .B(n389), .Z(n388) );
  XOR U588 ( .A(n346), .B(n390), .Z(n389) );
  XOR U589 ( .A(n390), .B(n347), .Z(n346) );
  OR U590 ( .A(n391), .B(n392), .Z(n347) );
  IV U591 ( .A(n387), .Z(n390) );
  XNOR U592 ( .A(n349), .B(n348), .Z(n387) );
  NANDN U593 ( .B(n393), .A(n394), .Z(n348) );
  XNOR U594 ( .A(n359), .B(n358), .Z(n349) );
  XOR U595 ( .A(n395), .B(n362), .Z(n358) );
  XNOR U596 ( .A(n355), .B(n356), .Z(n362) );
  NAND U597 ( .A(n312), .B(n247), .Z(n356) );
  XNOR U598 ( .A(n354), .B(n396), .Z(n355) );
  AND U599 ( .A(n212), .B(n353), .Z(n396) );
  XNOR U600 ( .A(n361), .B(n357), .Z(n395) );
  AND U601 ( .A(n404), .B(n405), .Z(n403) );
  NANDN U602 ( .B(n186), .A(n406), .Z(n405) );
  OR U603 ( .A(n407), .B(n408), .Z(n404) );
  XNOR U604 ( .A(n365), .B(n413), .Z(n368) );
  AND U605 ( .A(n284), .B(n280), .Z(n413) );
  XOR U606 ( .A(n414), .B(n415), .Z(n365) );
  ANDN U607 ( .A(n416), .B(n417), .Z(n415) );
  XNOR U608 ( .A(n418), .B(n414), .Z(n416) );
  XOR U609 ( .A(n419), .B(n369), .Z(n412) );
  NAND U610 ( .A(n242), .B(n329), .Z(n369) );
  IV U611 ( .A(n371), .Z(n419) );
  XNOR U612 ( .A(n378), .B(n379), .Z(n373) );
  NANDN U613 ( .B(n187), .A(n423), .Z(n379) );
  XNOR U614 ( .A(n377), .B(n424), .Z(n378) );
  AND U615 ( .A(n374), .B(n211), .Z(n424) );
  ANDN U616 ( .A(n425), .B(n426), .Z(n377) );
  NANDN U617 ( .B(n427), .A(n428), .Z(n425) );
  NAND U618 ( .A(n431), .B(n432), .Z(\_MxM/n194 ) );
  NANDN U619 ( .B(n102), .A(o[6]), .Z(n432) );
  AND U620 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U621 ( .B(n149), .A(o[6]), .Z(n434) );
  NANDN U622 ( .B(n154), .A(n121), .Z(n433) );
  XNOR U623 ( .A(n430), .B(\_MxM/Y0[7] ), .Z(n121) );
  XNOR U624 ( .A(n436), .B(n437), .Z(n435) );
  AND U625 ( .A(n165), .B(n438), .Z(n437) );
  XOR U626 ( .A(n391), .B(n441), .Z(n438) );
  XOR U627 ( .A(n441), .B(n392), .Z(n391) );
  OR U628 ( .A(n439), .B(n440), .Z(n392) );
  XNOR U629 ( .A(n393), .B(n394), .Z(n441) );
  XNOR U630 ( .A(n402), .B(n401), .Z(n393) );
  XOR U631 ( .A(n446), .B(n411), .Z(n401) );
  XNOR U632 ( .A(n398), .B(n399), .Z(n411) );
  NAND U633 ( .A(n312), .B(n284), .Z(n399) );
  XNOR U634 ( .A(n397), .B(n447), .Z(n398) );
  AND U635 ( .A(n247), .B(n353), .Z(n447) );
  XNOR U636 ( .A(n410), .B(n400), .Z(n446) );
  XNOR U637 ( .A(n454), .B(n409), .Z(n410) );
  XNOR U638 ( .A(n458), .B(n407), .Z(n454) );
  NAND U639 ( .A(n406), .B(n212), .Z(n407) );
  NANDN U640 ( .B(n186), .A(n460), .Z(n459) );
  XNOR U641 ( .A(n414), .B(n465), .Z(n417) );
  AND U642 ( .A(n329), .B(n280), .Z(n465) );
  XOR U643 ( .A(n466), .B(n467), .Z(n414) );
  ANDN U644 ( .A(n468), .B(n469), .Z(n467) );
  XNOR U645 ( .A(n470), .B(n466), .Z(n468) );
  XOR U646 ( .A(n471), .B(n418), .Z(n464) );
  NAND U647 ( .A(n242), .B(n374), .Z(n418) );
  IV U648 ( .A(n420), .Z(n471) );
  XNOR U649 ( .A(n427), .B(n428), .Z(n422) );
  NANDN U650 ( .B(n187), .A(n475), .Z(n428) );
  AND U651 ( .A(n423), .B(n211), .Z(n476) );
  NAND U652 ( .A(n477), .B(n478), .Z(n426) );
  NANDN U653 ( .B(n479), .A(n480), .Z(n477) );
  IV U654 ( .A(n429), .Z(n436) );
  NAND U655 ( .A(n483), .B(n484), .Z(\_MxM/n193 ) );
  NANDN U656 ( .B(n102), .A(o[5]), .Z(n484) );
  AND U657 ( .A(n485), .B(n486), .Z(n483) );
  NANDN U658 ( .B(n149), .A(o[5]), .Z(n486) );
  NANDN U659 ( .B(n154), .A(n118), .Z(n485) );
  XNOR U660 ( .A(n482), .B(\_MxM/Y0[6] ), .Z(n118) );
  XNOR U661 ( .A(n487), .B(n488), .Z(n482) );
  AND U662 ( .A(n165), .B(n490), .Z(n489) );
  XOR U663 ( .A(n439), .B(n491), .Z(n490) );
  XOR U664 ( .A(n491), .B(n440), .Z(n439) );
  OR U665 ( .A(n492), .B(n493), .Z(n440) );
  IV U666 ( .A(n488), .Z(n491) );
  XOR U667 ( .A(n445), .B(n444), .Z(n488) );
  XNOR U668 ( .A(n443), .B(n494), .Z(n444) );
  AND U669 ( .A(n442), .B(n495), .Z(n494) );
  AND U670 ( .A(n496), .B(n497), .Z(n495) );
  NANDN U671 ( .B(n186), .A(n498), .Z(n497) );
  OR U672 ( .A(n499), .B(n500), .Z(n496) );
  AND U673 ( .A(n501), .B(n502), .Z(n442) );
  NANDN U674 ( .B(n503), .A(n504), .Z(n502) );
  NANDN U675 ( .B(n505), .A(n506), .Z(n501) );
  XNOR U676 ( .A(n510), .B(n457), .Z(n452) );
  XNOR U677 ( .A(n449), .B(n450), .Z(n457) );
  NAND U678 ( .A(n312), .B(n329), .Z(n450) );
  XNOR U679 ( .A(n448), .B(n511), .Z(n449) );
  AND U680 ( .A(n284), .B(n353), .Z(n511) );
  XNOR U681 ( .A(n456), .B(n451), .Z(n510) );
  XNOR U682 ( .A(n461), .B(n519), .Z(n462) );
  AND U683 ( .A(n212), .B(n460), .Z(n519) );
  XOR U684 ( .A(n520), .B(n521), .Z(n461) );
  ANDN U685 ( .A(n522), .B(n523), .Z(n521) );
  XNOR U686 ( .A(n524), .B(n520), .Z(n522) );
  XOR U687 ( .A(n525), .B(n463), .Z(n518) );
  NAND U688 ( .A(n406), .B(n247), .Z(n463) );
  IV U689 ( .A(n455), .Z(n525) );
  XNOR U690 ( .A(n466), .B(n530), .Z(n469) );
  AND U691 ( .A(n374), .B(n280), .Z(n530) );
  XOR U692 ( .A(n531), .B(n532), .Z(n466) );
  ANDN U693 ( .A(n533), .B(n534), .Z(n532) );
  XNOR U694 ( .A(n535), .B(n531), .Z(n533) );
  XOR U695 ( .A(n536), .B(n470), .Z(n529) );
  NAND U696 ( .A(n242), .B(n423), .Z(n470) );
  IV U697 ( .A(n472), .Z(n536) );
  XNOR U698 ( .A(n479), .B(n480), .Z(n474) );
  NANDN U699 ( .B(n187), .A(n540), .Z(n480) );
  XNOR U700 ( .A(n478), .B(n541), .Z(n479) );
  AND U701 ( .A(n475), .B(n211), .Z(n541) );
  ANDN U702 ( .A(n542), .B(n543), .Z(n478) );
  NANDN U703 ( .B(n544), .A(n545), .Z(n542) );
  NAND U704 ( .A(n548), .B(n549), .Z(\_MxM/n192 ) );
  NANDN U705 ( .B(n102), .A(o[4]), .Z(n549) );
  AND U706 ( .A(n550), .B(n551), .Z(n548) );
  NANDN U707 ( .B(n149), .A(o[4]), .Z(n551) );
  NANDN U708 ( .B(n154), .A(n115), .Z(n550) );
  XNOR U709 ( .A(n547), .B(\_MxM/Y0[5] ), .Z(n115) );
  XNOR U710 ( .A(n552), .B(n553), .Z(n547) );
  AND U711 ( .A(n165), .B(n555), .Z(n554) );
  XOR U712 ( .A(n492), .B(n556), .Z(n555) );
  XOR U713 ( .A(n556), .B(n493), .Z(n492) );
  OR U714 ( .A(n557), .B(n558), .Z(n493) );
  IV U715 ( .A(n553), .Z(n556) );
  XOR U716 ( .A(n509), .B(n508), .Z(n553) );
  XOR U717 ( .A(n503), .B(n504), .Z(n500) );
  XOR U718 ( .A(n563), .B(n505), .Z(n503) );
  NAND U719 ( .A(n212), .B(n498), .Z(n505) );
  NANDN U720 ( .B(n506), .A(n564), .Z(n563) );
  NANDN U721 ( .B(n186), .A(n565), .Z(n564) );
  XOR U722 ( .A(n569), .B(n499), .Z(n559) );
  OR U723 ( .A(n570), .B(n571), .Z(n499) );
  IV U724 ( .A(n507), .Z(n569) );
  XNOR U725 ( .A(n575), .B(n528), .Z(n516) );
  XNOR U726 ( .A(n513), .B(n514), .Z(n528) );
  NAND U727 ( .A(n312), .B(n374), .Z(n514) );
  XNOR U728 ( .A(n512), .B(n576), .Z(n513) );
  AND U729 ( .A(n329), .B(n353), .Z(n576) );
  XNOR U730 ( .A(n527), .B(n515), .Z(n575) );
  XNOR U731 ( .A(n520), .B(n584), .Z(n523) );
  AND U732 ( .A(n247), .B(n460), .Z(n584) );
  XOR U733 ( .A(n585), .B(n586), .Z(n520) );
  ANDN U734 ( .A(n587), .B(n588), .Z(n586) );
  XNOR U735 ( .A(n589), .B(n585), .Z(n587) );
  XOR U736 ( .A(n590), .B(n524), .Z(n583) );
  NAND U737 ( .A(n406), .B(n284), .Z(n524) );
  IV U738 ( .A(n526), .Z(n590) );
  XNOR U739 ( .A(n531), .B(n595), .Z(n534) );
  AND U740 ( .A(n423), .B(n280), .Z(n595) );
  XOR U741 ( .A(n596), .B(n597), .Z(n531) );
  ANDN U742 ( .A(n598), .B(n599), .Z(n597) );
  XNOR U743 ( .A(n600), .B(n596), .Z(n598) );
  XOR U744 ( .A(n601), .B(n535), .Z(n594) );
  NAND U745 ( .A(n242), .B(n475), .Z(n535) );
  IV U746 ( .A(n537), .Z(n601) );
  XNOR U747 ( .A(n544), .B(n545), .Z(n539) );
  NANDN U748 ( .B(n187), .A(n605), .Z(n545) );
  AND U749 ( .A(n540), .B(n211), .Z(n606) );
  NAND U750 ( .A(n607), .B(n608), .Z(n543) );
  NANDN U751 ( .B(n609), .A(n610), .Z(n607) );
  NAND U752 ( .A(n613), .B(n614), .Z(\_MxM/n191 ) );
  NANDN U753 ( .B(n102), .A(o[3]), .Z(n614) );
  AND U754 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U755 ( .B(n149), .A(o[3]), .Z(n616) );
  NANDN U756 ( .B(n154), .A(n112), .Z(n615) );
  XNOR U757 ( .A(n612), .B(\_MxM/Y0[4] ), .Z(n112) );
  XNOR U758 ( .A(n617), .B(n618), .Z(n612) );
  AND U759 ( .A(n165), .B(n620), .Z(n619) );
  XOR U760 ( .A(n557), .B(n621), .Z(n620) );
  XOR U761 ( .A(n621), .B(n558), .Z(n557) );
  OR U762 ( .A(n622), .B(n623), .Z(n558) );
  IV U763 ( .A(n618), .Z(n621) );
  XOR U764 ( .A(n574), .B(n573), .Z(n618) );
  XOR U765 ( .A(n624), .B(n570), .Z(n573) );
  XOR U766 ( .A(n562), .B(n561), .Z(n570) );
  XOR U767 ( .A(n560), .B(n625), .Z(n561) );
  AND U768 ( .A(n626), .B(n627), .Z(n625) );
  NANDN U769 ( .B(n186), .A(n628), .Z(n627) );
  OR U770 ( .A(n629), .B(n630), .Z(n626) );
  NAND U771 ( .A(n247), .B(n498), .Z(n568) );
  XNOR U772 ( .A(n566), .B(n634), .Z(n567) );
  AND U773 ( .A(n565), .B(n212), .Z(n634) );
  NANDN U774 ( .B(n638), .A(n639), .Z(n571) );
  XNOR U775 ( .A(n643), .B(n593), .Z(n581) );
  XNOR U776 ( .A(n578), .B(n579), .Z(n593) );
  NAND U777 ( .A(n312), .B(n423), .Z(n579) );
  XNOR U778 ( .A(n577), .B(n644), .Z(n578) );
  AND U779 ( .A(n374), .B(n353), .Z(n644) );
  XNOR U780 ( .A(n592), .B(n580), .Z(n643) );
  XNOR U781 ( .A(n585), .B(n652), .Z(n588) );
  AND U782 ( .A(n284), .B(n460), .Z(n652) );
  XOR U783 ( .A(n653), .B(n654), .Z(n585) );
  ANDN U784 ( .A(n655), .B(n656), .Z(n654) );
  XNOR U785 ( .A(n657), .B(n653), .Z(n655) );
  XOR U786 ( .A(n658), .B(n589), .Z(n651) );
  NAND U787 ( .A(n406), .B(n329), .Z(n589) );
  IV U788 ( .A(n591), .Z(n658) );
  XNOR U789 ( .A(n596), .B(n663), .Z(n599) );
  AND U790 ( .A(n475), .B(n280), .Z(n663) );
  XOR U791 ( .A(n664), .B(n665), .Z(n596) );
  ANDN U792 ( .A(n666), .B(n667), .Z(n665) );
  XNOR U793 ( .A(n668), .B(n664), .Z(n666) );
  XOR U794 ( .A(n669), .B(n600), .Z(n662) );
  NAND U795 ( .A(n242), .B(n540), .Z(n600) );
  IV U796 ( .A(n602), .Z(n669) );
  XNOR U797 ( .A(n609), .B(n610), .Z(n604) );
  NANDN U798 ( .B(n187), .A(n673), .Z(n610) );
  XNOR U799 ( .A(n608), .B(n674), .Z(n609) );
  AND U800 ( .A(n605), .B(n211), .Z(n674) );
  ANDN U801 ( .A(n675), .B(n676), .Z(n608) );
  NANDN U802 ( .B(n677), .A(n678), .Z(n675) );
  NAND U803 ( .A(n681), .B(n682), .Z(\_MxM/n190 ) );
  NANDN U804 ( .B(n102), .A(o[2]), .Z(n682) );
  AND U805 ( .A(n683), .B(n684), .Z(n681) );
  NANDN U806 ( .B(n149), .A(o[2]), .Z(n684) );
  NANDN U807 ( .B(n154), .A(n109), .Z(n683) );
  XNOR U808 ( .A(n680), .B(\_MxM/Y0[3] ), .Z(n109) );
  XNOR U809 ( .A(n685), .B(n686), .Z(n680) );
  AND U810 ( .A(n165), .B(n688), .Z(n687) );
  XOR U811 ( .A(n622), .B(n689), .Z(n688) );
  XOR U812 ( .A(n689), .B(n623), .Z(n622) );
  OR U813 ( .A(n690), .B(n691), .Z(n623) );
  IV U814 ( .A(n686), .Z(n689) );
  XOR U815 ( .A(n642), .B(n641), .Z(n686) );
  XOR U816 ( .A(n692), .B(n638), .Z(n641) );
  XOR U817 ( .A(n633), .B(n632), .Z(n638) );
  XNOR U818 ( .A(n697), .B(n629), .Z(n693) );
  NAND U819 ( .A(n212), .B(n628), .Z(n629) );
  NANDN U820 ( .B(n186), .A(n699), .Z(n698) );
  NAND U821 ( .A(n284), .B(n498), .Z(n637) );
  XNOR U822 ( .A(n635), .B(n703), .Z(n636) );
  AND U823 ( .A(n565), .B(n247), .Z(n703) );
  XNOR U824 ( .A(n639), .B(n640), .Z(n692) );
  XNOR U825 ( .A(n713), .B(n661), .Z(n649) );
  XNOR U826 ( .A(n646), .B(n647), .Z(n661) );
  NAND U827 ( .A(n312), .B(n475), .Z(n647) );
  XNOR U828 ( .A(n645), .B(n714), .Z(n646) );
  AND U829 ( .A(n423), .B(n353), .Z(n714) );
  XNOR U830 ( .A(n660), .B(n648), .Z(n713) );
  XNOR U831 ( .A(n653), .B(n722), .Z(n656) );
  AND U832 ( .A(n329), .B(n460), .Z(n722) );
  XOR U833 ( .A(n726), .B(n657), .Z(n721) );
  NAND U834 ( .A(n406), .B(n374), .Z(n657) );
  IV U835 ( .A(n659), .Z(n726) );
  XNOR U836 ( .A(n664), .B(n731), .Z(n667) );
  AND U837 ( .A(n540), .B(n280), .Z(n731) );
  XOR U838 ( .A(n732), .B(n733), .Z(n664) );
  ANDN U839 ( .A(n734), .B(n735), .Z(n733) );
  XNOR U840 ( .A(n736), .B(n732), .Z(n734) );
  XOR U841 ( .A(n737), .B(n668), .Z(n730) );
  NAND U842 ( .A(n242), .B(n605), .Z(n668) );
  IV U843 ( .A(n670), .Z(n737) );
  XNOR U844 ( .A(n677), .B(n678), .Z(n672) );
  OR U845 ( .A(n741), .B(n187), .Z(n678) );
  AND U846 ( .A(n673), .B(n211), .Z(n742) );
  NAND U847 ( .A(n743), .B(n744), .Z(n676) );
  NANDN U848 ( .B(n745), .A(n746), .Z(n743) );
  NAND U849 ( .A(n749), .B(n750), .Z(\_MxM/n189 ) );
  NANDN U850 ( .B(n102), .A(o[1]), .Z(n750) );
  AND U851 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U852 ( .B(n149), .A(o[1]), .Z(n752) );
  NANDN U853 ( .B(n154), .A(n105), .Z(n751) );
  XNOR U854 ( .A(n748), .B(\_MxM/Y0[2] ), .Z(n105) );
  XNOR U855 ( .A(n753), .B(n754), .Z(n748) );
  XOR U856 ( .A(n747), .B(n755), .Z(n753) );
  AND U857 ( .A(n165), .B(n756), .Z(n755) );
  XOR U858 ( .A(n690), .B(n757), .Z(n756) );
  XOR U859 ( .A(n757), .B(n691), .Z(n690) );
  NANDN U860 ( .B(n758), .A(n759), .Z(n691) );
  IV U861 ( .A(n754), .Z(n757) );
  XOR U862 ( .A(n709), .B(n708), .Z(n754) );
  XNOR U863 ( .A(n760), .B(n712), .Z(n708) );
  XNOR U864 ( .A(n700), .B(n762), .Z(n701) );
  AND U865 ( .A(n699), .B(n212), .Z(n762) );
  XOR U866 ( .A(n766), .B(n702), .Z(n761) );
  NAND U867 ( .A(n247), .B(n628), .Z(n702) );
  IV U868 ( .A(n694), .Z(n766) );
  XNOR U869 ( .A(n705), .B(n706), .Z(n696) );
  NAND U870 ( .A(n329), .B(n498), .Z(n706) );
  XNOR U871 ( .A(n704), .B(n770), .Z(n705) );
  AND U872 ( .A(n565), .B(n284), .Z(n770) );
  XNOR U873 ( .A(n711), .B(n707), .Z(n760) );
  AND U874 ( .A(n778), .B(n779), .Z(n777) );
  OR U875 ( .A(n780), .B(n781), .Z(n779) );
  AND U876 ( .A(n782), .B(n783), .Z(n778) );
  NANDN U877 ( .B(n186), .A(n784), .Z(n783) );
  NANDN U878 ( .B(n785), .A(n786), .Z(n782) );
  XNOR U879 ( .A(n790), .B(n729), .Z(n719) );
  XNOR U880 ( .A(n716), .B(n717), .Z(n729) );
  NAND U881 ( .A(n312), .B(n540), .Z(n717) );
  XNOR U882 ( .A(n715), .B(n791), .Z(n716) );
  AND U883 ( .A(n475), .B(n353), .Z(n791) );
  XNOR U884 ( .A(n728), .B(n718), .Z(n790) );
  XNOR U885 ( .A(n723), .B(n799), .Z(n724) );
  AND U886 ( .A(n374), .B(n460), .Z(n799) );
  XOR U887 ( .A(n803), .B(n725), .Z(n798) );
  NAND U888 ( .A(n406), .B(n423), .Z(n725) );
  IV U889 ( .A(n727), .Z(n803) );
  XNOR U890 ( .A(n732), .B(n808), .Z(n735) );
  AND U891 ( .A(n605), .B(n280), .Z(n808) );
  XOR U892 ( .A(n809), .B(n810), .Z(n732) );
  ANDN U893 ( .A(n811), .B(n812), .Z(n810) );
  XNOR U894 ( .A(n813), .B(n809), .Z(n811) );
  XOR U895 ( .A(n814), .B(n736), .Z(n807) );
  NAND U896 ( .A(n242), .B(n673), .Z(n736) );
  IV U897 ( .A(n738), .Z(n814) );
  XNOR U898 ( .A(n745), .B(n746), .Z(n740) );
  OR U899 ( .A(n818), .B(n187), .Z(n746) );
  XNOR U900 ( .A(n744), .B(n819), .Z(n745) );
  ANDN U901 ( .A(n211), .B(n741), .Z(n819) );
  ANDN U902 ( .A(n820), .B(n821), .Z(n744) );
  NANDN U903 ( .B(n822), .A(n823), .Z(n820) );
  NAND U904 ( .A(n826), .B(n827), .Z(\_MxM/n188 ) );
  NANDN U905 ( .B(n102), .A(o[0]), .Z(n827) );
  AND U906 ( .A(n828), .B(n829), .Z(n826) );
  NANDN U907 ( .B(n149), .A(o[0]), .Z(n829) );
  IV U908 ( .A(n830), .Z(n149) );
  OR U909 ( .A(n154), .B(n100), .Z(n828) );
  IV U910 ( .A(\_MxM/Y0[1] ), .Z(n106) );
  XOR U911 ( .A(n831), .B(n832), .Z(n825) );
  XNOR U912 ( .A(n833), .B(n824), .Z(n831) );
  NAND U913 ( .A(\_MxM/Y0[0] ), .B(n758), .Z(n824) );
  NAND U914 ( .A(n834), .B(n165), .Z(n833) );
  XOR U915 ( .A(e_input[15]), .B(g_input[15]), .Z(n165) );
  XNOR U916 ( .A(n759), .B(n832), .Z(n834) );
  XNOR U917 ( .A(n758), .B(n832), .Z(n759) );
  XNOR U918 ( .A(n776), .B(n775), .Z(n832) );
  XNOR U919 ( .A(n835), .B(n789), .Z(n775) );
  XNOR U920 ( .A(n763), .B(n837), .Z(n764) );
  AND U921 ( .A(n699), .B(n247), .Z(n837) );
  XOR U922 ( .A(n841), .B(n765), .Z(n836) );
  NAND U923 ( .A(n284), .B(n628), .Z(n765) );
  IV U924 ( .A(n767), .Z(n841) );
  XNOR U925 ( .A(n772), .B(n773), .Z(n769) );
  NAND U926 ( .A(n374), .B(n498), .Z(n773) );
  XNOR U927 ( .A(n771), .B(n845), .Z(n772) );
  AND U928 ( .A(n565), .B(n329), .Z(n845) );
  XNOR U929 ( .A(n788), .B(n774), .Z(n835) );
  XNOR U930 ( .A(n852), .B(n785), .Z(n788) );
  XOR U931 ( .A(n853), .B(n780), .Z(n785) );
  NAND U932 ( .A(n212), .B(n784), .Z(n780) );
  NANDN U933 ( .B(n186), .A(n855), .Z(n854) );
  XNOR U934 ( .A(n786), .B(n787), .Z(n852) );
  XNOR U935 ( .A(n865), .B(n806), .Z(n796) );
  XNOR U936 ( .A(n793), .B(n794), .Z(n806) );
  NAND U937 ( .A(n312), .B(n605), .Z(n794) );
  XNOR U938 ( .A(n792), .B(n866), .Z(n793) );
  AND U939 ( .A(n540), .B(n353), .Z(n866) );
  XNOR U940 ( .A(n805), .B(n795), .Z(n865) );
  XNOR U941 ( .A(n800), .B(n874), .Z(n801) );
  AND U942 ( .A(n423), .B(n460), .Z(n874) );
  XOR U943 ( .A(n878), .B(n802), .Z(n873) );
  NAND U944 ( .A(n406), .B(n475), .Z(n802) );
  IV U945 ( .A(n804), .Z(n878) );
  XNOR U946 ( .A(n809), .B(n883), .Z(n812) );
  AND U947 ( .A(n673), .B(n280), .Z(n883) );
  XOR U948 ( .A(n887), .B(n813), .Z(n882) );
  NANDN U949 ( .B(n741), .A(n242), .Z(n813) );
  IV U950 ( .A(n815), .Z(n887) );
  XNOR U951 ( .A(n822), .B(n823), .Z(n817) );
  NANDN U952 ( .B(n187), .A(n891), .Z(n823) );
  ANDN U953 ( .A(n211), .B(n818), .Z(n892) );
  NAND U954 ( .A(n893), .B(n894), .Z(n821) );
  NANDN U955 ( .B(n895), .A(n896), .Z(n893) );
  XNOR U956 ( .A(n851), .B(n850), .Z(n758) );
  XNOR U957 ( .A(n897), .B(n861), .Z(n850) );
  XNOR U958 ( .A(n838), .B(n899), .Z(n839) );
  AND U959 ( .A(n699), .B(n284), .Z(n899) );
  XOR U960 ( .A(n903), .B(n840), .Z(n898) );
  NAND U961 ( .A(n329), .B(n628), .Z(n840) );
  IV U962 ( .A(n842), .Z(n903) );
  XNOR U963 ( .A(n847), .B(n848), .Z(n844) );
  NAND U964 ( .A(n423), .B(n498), .Z(n848) );
  XNOR U965 ( .A(n846), .B(n907), .Z(n847) );
  AND U966 ( .A(n565), .B(n374), .Z(n907) );
  XNOR U967 ( .A(n860), .B(n849), .Z(n897) );
  XOR U968 ( .A(n911), .B(n912), .Z(n849) );
  XNOR U969 ( .A(n913), .B(n864), .Z(n860) );
  NAND U970 ( .A(n247), .B(n784), .Z(n858) );
  XNOR U971 ( .A(n856), .B(n914), .Z(n857) );
  AND U972 ( .A(n855), .B(n212), .Z(n914) );
  XNOR U973 ( .A(n863), .B(n859), .Z(n913) );
  XOR U974 ( .A(n918), .B(n919), .Z(n859) );
  AND U975 ( .A(n920), .B(n921), .Z(n919) );
  XOR U976 ( .A(n922), .B(n923), .Z(n921) );
  XOR U977 ( .A(n918), .B(n924), .Z(n923) );
  XOR U978 ( .A(n905), .B(n925), .Z(n920) );
  XOR U979 ( .A(n918), .B(n906), .Z(n925) );
  NAND U980 ( .A(n498), .B(n475), .Z(n910) );
  XNOR U981 ( .A(n908), .B(n926), .Z(n909) );
  AND U982 ( .A(n565), .B(n423), .Z(n926) );
  XNOR U983 ( .A(n900), .B(n931), .Z(n901) );
  AND U984 ( .A(n699), .B(n329), .Z(n931) );
  XOR U985 ( .A(n932), .B(n933), .Z(n900) );
  ANDN U986 ( .A(n934), .B(n935), .Z(n933) );
  XNOR U987 ( .A(n936), .B(n932), .Z(n934) );
  XOR U988 ( .A(n937), .B(n902), .Z(n930) );
  NAND U989 ( .A(n374), .B(n628), .Z(n902) );
  IV U990 ( .A(n904), .Z(n937) );
  XOR U991 ( .A(n941), .B(n942), .Z(n918) );
  AND U992 ( .A(n943), .B(n944), .Z(n942) );
  XOR U993 ( .A(n945), .B(n946), .Z(n944) );
  XOR U994 ( .A(n941), .B(n947), .Z(n946) );
  XOR U995 ( .A(n939), .B(n948), .Z(n943) );
  XOR U996 ( .A(n941), .B(n940), .Z(n948) );
  NAND U997 ( .A(n498), .B(n540), .Z(n929) );
  XNOR U998 ( .A(n927), .B(n949), .Z(n928) );
  AND U999 ( .A(n475), .B(n565), .Z(n949) );
  XNOR U1000 ( .A(n932), .B(n954), .Z(n935) );
  AND U1001 ( .A(n699), .B(n374), .Z(n954) );
  XOR U1002 ( .A(n955), .B(n956), .Z(n932) );
  ANDN U1003 ( .A(n957), .B(n958), .Z(n956) );
  XNOR U1004 ( .A(n959), .B(n955), .Z(n957) );
  XOR U1005 ( .A(n960), .B(n936), .Z(n953) );
  NAND U1006 ( .A(n423), .B(n628), .Z(n936) );
  IV U1007 ( .A(n938), .Z(n960) );
  XOR U1008 ( .A(n964), .B(n965), .Z(n941) );
  AND U1009 ( .A(n966), .B(n967), .Z(n965) );
  XOR U1010 ( .A(n968), .B(n969), .Z(n967) );
  XOR U1011 ( .A(n964), .B(n970), .Z(n969) );
  XOR U1012 ( .A(n962), .B(n971), .Z(n966) );
  XOR U1013 ( .A(n964), .B(n963), .Z(n971) );
  NAND U1014 ( .A(n498), .B(n605), .Z(n952) );
  XNOR U1015 ( .A(n950), .B(n972), .Z(n951) );
  AND U1016 ( .A(n540), .B(n565), .Z(n972) );
  XNOR U1017 ( .A(n955), .B(n977), .Z(n958) );
  AND U1018 ( .A(n699), .B(n423), .Z(n977) );
  XOR U1019 ( .A(n978), .B(n979), .Z(n955) );
  ANDN U1020 ( .A(n980), .B(n981), .Z(n979) );
  XNOR U1021 ( .A(n982), .B(n978), .Z(n980) );
  XOR U1022 ( .A(n983), .B(n959), .Z(n976) );
  NAND U1023 ( .A(n628), .B(n475), .Z(n959) );
  IV U1024 ( .A(n961), .Z(n983) );
  XOR U1025 ( .A(n987), .B(n988), .Z(n964) );
  AND U1026 ( .A(n989), .B(n990), .Z(n988) );
  XOR U1027 ( .A(n991), .B(n992), .Z(n990) );
  XOR U1028 ( .A(n987), .B(n993), .Z(n992) );
  XOR U1029 ( .A(n985), .B(n994), .Z(n989) );
  XOR U1030 ( .A(n987), .B(n986), .Z(n994) );
  XNOR U1031 ( .A(n995), .B(n975), .Z(n986) );
  NAND U1032 ( .A(n498), .B(n673), .Z(n975) );
  IV U1033 ( .A(n974), .Z(n995) );
  XNOR U1034 ( .A(n973), .B(n996), .Z(n974) );
  AND U1035 ( .A(n605), .B(n565), .Z(n996) );
  XOR U1036 ( .A(n997), .B(n998), .Z(n973) );
  ANDN U1037 ( .A(n999), .B(n1000), .Z(n998) );
  XNOR U1038 ( .A(n1001), .B(n997), .Z(n999) );
  XNOR U1039 ( .A(n1002), .B(n1003), .Z(n985) );
  IV U1040 ( .A(n981), .Z(n1003) );
  XNOR U1041 ( .A(n978), .B(n1004), .Z(n981) );
  AND U1042 ( .A(n475), .B(n699), .Z(n1004) );
  XOR U1043 ( .A(n1005), .B(n1006), .Z(n978) );
  ANDN U1044 ( .A(n1007), .B(n1008), .Z(n1006) );
  XNOR U1045 ( .A(n1009), .B(n1005), .Z(n1007) );
  XOR U1046 ( .A(n1010), .B(n982), .Z(n1002) );
  NAND U1047 ( .A(n628), .B(n540), .Z(n982) );
  IV U1048 ( .A(n984), .Z(n1010) );
  XOR U1049 ( .A(n1014), .B(n1015), .Z(n987) );
  AND U1050 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR U1051 ( .A(n1018), .B(n1019), .Z(n1017) );
  XOR U1052 ( .A(n1014), .B(n1020), .Z(n1019) );
  XOR U1053 ( .A(n1012), .B(n1021), .Z(n1016) );
  XOR U1054 ( .A(n1014), .B(n1013), .Z(n1021) );
  XNOR U1055 ( .A(n1022), .B(n1001), .Z(n1013) );
  NANDN U1056 ( .B(n741), .A(n498), .Z(n1001) );
  IV U1057 ( .A(n1000), .Z(n1022) );
  XNOR U1058 ( .A(n997), .B(n1023), .Z(n1000) );
  AND U1059 ( .A(n673), .B(n565), .Z(n1023) );
  XOR U1060 ( .A(n1024), .B(n1025), .Z(n997) );
  ANDN U1061 ( .A(n1026), .B(n1027), .Z(n1025) );
  XNOR U1062 ( .A(n1028), .B(n1024), .Z(n1026) );
  XNOR U1063 ( .A(n1029), .B(n1030), .Z(n1012) );
  IV U1064 ( .A(n1008), .Z(n1030) );
  XNOR U1065 ( .A(n1005), .B(n1031), .Z(n1008) );
  AND U1066 ( .A(n540), .B(n699), .Z(n1031) );
  XOR U1067 ( .A(n1032), .B(n1033), .Z(n1005) );
  ANDN U1068 ( .A(n1034), .B(n1035), .Z(n1033) );
  XNOR U1069 ( .A(n1036), .B(n1032), .Z(n1034) );
  XOR U1070 ( .A(n1037), .B(n1009), .Z(n1029) );
  NAND U1071 ( .A(n628), .B(n605), .Z(n1009) );
  IV U1072 ( .A(n1011), .Z(n1037) );
  XOR U1073 ( .A(n1041), .B(n1042), .Z(n1014) );
  AND U1074 ( .A(n1043), .B(n1044), .Z(n1042) );
  XOR U1075 ( .A(n1045), .B(n1046), .Z(n1044) );
  XOR U1076 ( .A(n1041), .B(n1047), .Z(n1046) );
  XOR U1077 ( .A(n1039), .B(n1048), .Z(n1043) );
  XOR U1078 ( .A(n1041), .B(n1040), .Z(n1048) );
  XNOR U1079 ( .A(n1049), .B(n1028), .Z(n1040) );
  NANDN U1080 ( .B(n818), .A(n498), .Z(n1028) );
  IV U1081 ( .A(n1027), .Z(n1049) );
  XNOR U1082 ( .A(n1024), .B(n1050), .Z(n1027) );
  ANDN U1083 ( .A(n565), .B(n741), .Z(n1050) );
  XOR U1084 ( .A(n1051), .B(n1052), .Z(n1024) );
  ANDN U1085 ( .A(n1053), .B(n1054), .Z(n1052) );
  XNOR U1086 ( .A(n1055), .B(n1051), .Z(n1053) );
  XNOR U1087 ( .A(n1056), .B(n1057), .Z(n1039) );
  IV U1088 ( .A(n1035), .Z(n1057) );
  XNOR U1089 ( .A(n1032), .B(n1058), .Z(n1035) );
  AND U1090 ( .A(n605), .B(n699), .Z(n1058) );
  XOR U1091 ( .A(n1059), .B(n1060), .Z(n1032) );
  ANDN U1092 ( .A(n1061), .B(n1062), .Z(n1060) );
  XNOR U1093 ( .A(n1063), .B(n1059), .Z(n1061) );
  XOR U1094 ( .A(n1064), .B(n1036), .Z(n1056) );
  NAND U1095 ( .A(n628), .B(n673), .Z(n1036) );
  IV U1096 ( .A(n1038), .Z(n1064) );
  XOR U1097 ( .A(n1068), .B(n1069), .Z(n1041) );
  AND U1098 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U1099 ( .A(n1072), .B(n1073), .Z(n1071) );
  XOR U1100 ( .A(n1068), .B(n1074), .Z(n1073) );
  XOR U1101 ( .A(n1066), .B(n1075), .Z(n1070) );
  XOR U1102 ( .A(n1068), .B(n1067), .Z(n1075) );
  XNOR U1103 ( .A(n1076), .B(n1055), .Z(n1067) );
  NAND U1104 ( .A(n498), .B(n891), .Z(n1055) );
  IV U1105 ( .A(n1054), .Z(n1076) );
  XNOR U1106 ( .A(n1051), .B(n1077), .Z(n1054) );
  ANDN U1107 ( .A(n565), .B(n818), .Z(n1077) );
  XOR U1108 ( .A(n1078), .B(n1079), .Z(n1051) );
  ANDN U1109 ( .A(n1080), .B(n1081), .Z(n1079) );
  XNOR U1110 ( .A(n1082), .B(n1078), .Z(n1080) );
  XNOR U1111 ( .A(n1083), .B(n1084), .Z(n1066) );
  IV U1112 ( .A(n1062), .Z(n1084) );
  XNOR U1113 ( .A(n1059), .B(n1085), .Z(n1062) );
  AND U1114 ( .A(n673), .B(n699), .Z(n1085) );
  XOR U1115 ( .A(n1086), .B(n1087), .Z(n1059) );
  ANDN U1116 ( .A(n1088), .B(n1089), .Z(n1087) );
  XNOR U1117 ( .A(n1090), .B(n1086), .Z(n1088) );
  XOR U1118 ( .A(n1091), .B(n1063), .Z(n1083) );
  NANDN U1119 ( .B(n741), .A(n628), .Z(n1063) );
  IV U1120 ( .A(n1065), .Z(n1091) );
  XOR U1121 ( .A(n1096), .B(n1097), .Z(n912) );
  XNOR U1122 ( .A(n1098), .B(n1095), .Z(n1096) );
  XNOR U1123 ( .A(n1086), .B(n1100), .Z(n1089) );
  ANDN U1124 ( .A(n699), .B(n741), .Z(n1100) );
  XOR U1125 ( .A(n1103), .B(n1101), .Z(n1102) );
  ANDN U1126 ( .A(n699), .B(n818), .Z(n1103) );
  AND U1127 ( .A(n891), .B(n628), .Z(n1104) );
  XOR U1128 ( .A(n1105), .B(n1106), .Z(n1101) );
  ANDN U1129 ( .A(n1107), .B(n1108), .Z(n1106) );
  XNOR U1130 ( .A(n1109), .B(n1105), .Z(n1107) );
  XOR U1131 ( .A(n1110), .B(n1090), .Z(n1099) );
  NANDN U1132 ( .B(n818), .A(n628), .Z(n1090) );
  IV U1133 ( .A(n1092), .Z(n1110) );
  NAND U1134 ( .A(n628), .B(n1111), .Z(n1109) );
  XNOR U1135 ( .A(n1105), .B(n1112), .Z(n1108) );
  AND U1136 ( .A(n891), .B(n699), .Z(n1112) );
  AND U1137 ( .A(n1113), .B(g_input[0]), .Z(n1105) );
  NANDN U1138 ( .B(n628), .A(n1114), .Z(n1113) );
  NAND U1139 ( .A(n1111), .B(n699), .Z(n1114) );
  XNOR U1140 ( .A(n1081), .B(n1082), .Z(n1094) );
  NAND U1141 ( .A(n498), .B(n1111), .Z(n1082) );
  XNOR U1142 ( .A(n1078), .B(n1117), .Z(n1081) );
  AND U1143 ( .A(n891), .B(n565), .Z(n1117) );
  AND U1144 ( .A(n1118), .B(g_input[0]), .Z(n1078) );
  NANDN U1145 ( .B(n498), .A(n1119), .Z(n1118) );
  NAND U1146 ( .A(n1111), .B(n565), .Z(n1119) );
  XOR U1147 ( .A(n1122), .B(n1123), .Z(n1095) );
  XOR U1148 ( .A(n1124), .B(n1125), .Z(n863) );
  AND U1149 ( .A(n1126), .B(n1127), .Z(n1125) );
  NANDN U1150 ( .B(n186), .A(n1128), .Z(n1127) );
  NANDN U1151 ( .B(n1129), .A(n1130), .Z(n186) );
  AND U1152 ( .A(n1131), .B(g_input[15]), .Z(n1130) );
  OR U1153 ( .A(n1132), .B(n1133), .Z(n1126) );
  IV U1154 ( .A(n862), .Z(n1124) );
  NAND U1155 ( .A(n284), .B(n784), .Z(n917) );
  XNOR U1156 ( .A(n915), .B(n1135), .Z(n916) );
  AND U1157 ( .A(n855), .B(n247), .Z(n1135) );
  XOR U1158 ( .A(n1143), .B(n1132), .Z(n1139) );
  NAND U1159 ( .A(n212), .B(n1128), .Z(n1132) );
  IV U1160 ( .A(n1134), .Z(n1143) );
  NAND U1161 ( .A(n329), .B(n784), .Z(n1138) );
  XNOR U1162 ( .A(n1136), .B(n1145), .Z(n1137) );
  AND U1163 ( .A(n855), .B(n284), .Z(n1145) );
  XNOR U1164 ( .A(n1140), .B(n1150), .Z(n1141) );
  AND U1165 ( .A(n212), .B(e_input[0]), .Z(n1150) );
  XNOR U1166 ( .A(n1131), .B(g_input[14]), .Z(n1129) );
  NOR U1167 ( .A(n1151), .B(n1152), .Z(n1131) );
  XOR U1168 ( .A(n1156), .B(n1142), .Z(n1149) );
  NAND U1169 ( .A(n247), .B(n1128), .Z(n1142) );
  IV U1170 ( .A(n1144), .Z(n1156) );
  NAND U1171 ( .A(n374), .B(n784), .Z(n1148) );
  XNOR U1172 ( .A(n1146), .B(n1158), .Z(n1147) );
  AND U1173 ( .A(n855), .B(n329), .Z(n1158) );
  XOR U1174 ( .A(n1159), .B(n1160), .Z(n1146) );
  ANDN U1175 ( .A(n1161), .B(n1162), .Z(n1160) );
  XNOR U1176 ( .A(n1163), .B(n1159), .Z(n1161) );
  XNOR U1177 ( .A(n1153), .B(n1165), .Z(n1154) );
  AND U1178 ( .A(n247), .B(e_input[0]), .Z(n1165) );
  XOR U1179 ( .A(n1151), .B(g_input[13]), .Z(n1152) );
  NANDN U1180 ( .B(n1166), .A(n1167), .Z(n1151) );
  XOR U1181 ( .A(n1171), .B(n1155), .Z(n1164) );
  NAND U1182 ( .A(n284), .B(n1128), .Z(n1155) );
  IV U1183 ( .A(n1157), .Z(n1171) );
  XNOR U1184 ( .A(n1173), .B(n1163), .Z(n991) );
  NAND U1185 ( .A(n423), .B(n784), .Z(n1163) );
  IV U1186 ( .A(n1162), .Z(n1173) );
  XNOR U1187 ( .A(n1159), .B(n1174), .Z(n1162) );
  AND U1188 ( .A(n855), .B(n374), .Z(n1174) );
  XOR U1189 ( .A(n1175), .B(n1176), .Z(n1159) );
  ANDN U1190 ( .A(n1177), .B(n1178), .Z(n1176) );
  XNOR U1191 ( .A(n1179), .B(n1175), .Z(n1177) );
  XNOR U1192 ( .A(n1180), .B(n1181), .Z(n993) );
  IV U1193 ( .A(n1169), .Z(n1181) );
  XNOR U1194 ( .A(n1168), .B(n1182), .Z(n1169) );
  AND U1195 ( .A(n284), .B(e_input[0]), .Z(n1182) );
  XNOR U1196 ( .A(n1167), .B(g_input[12]), .Z(n1166) );
  NOR U1197 ( .A(n1183), .B(n1184), .Z(n1167) );
  XOR U1198 ( .A(n1185), .B(n1186), .Z(n1168) );
  ANDN U1199 ( .A(n1187), .B(n1188), .Z(n1186) );
  XNOR U1200 ( .A(n1189), .B(n1185), .Z(n1187) );
  XOR U1201 ( .A(n1190), .B(n1170), .Z(n1180) );
  NAND U1202 ( .A(n329), .B(n1128), .Z(n1170) );
  IV U1203 ( .A(n1172), .Z(n1190) );
  XNOR U1204 ( .A(n1192), .B(n1179), .Z(n1018) );
  NAND U1205 ( .A(n475), .B(n784), .Z(n1179) );
  IV U1206 ( .A(n1178), .Z(n1192) );
  XNOR U1207 ( .A(n1175), .B(n1193), .Z(n1178) );
  AND U1208 ( .A(n855), .B(n423), .Z(n1193) );
  XOR U1209 ( .A(n1194), .B(n1195), .Z(n1175) );
  ANDN U1210 ( .A(n1196), .B(n1197), .Z(n1195) );
  XNOR U1211 ( .A(n1198), .B(n1194), .Z(n1196) );
  XNOR U1212 ( .A(n1199), .B(n1200), .Z(n1020) );
  IV U1213 ( .A(n1188), .Z(n1200) );
  XNOR U1214 ( .A(n1185), .B(n1201), .Z(n1188) );
  AND U1215 ( .A(n329), .B(e_input[0]), .Z(n1201) );
  XOR U1216 ( .A(n1183), .B(g_input[11]), .Z(n1184) );
  NANDN U1217 ( .B(n1202), .A(n1203), .Z(n1183) );
  XOR U1218 ( .A(n1204), .B(n1205), .Z(n1185) );
  ANDN U1219 ( .A(n1206), .B(n1207), .Z(n1205) );
  XNOR U1220 ( .A(n1208), .B(n1204), .Z(n1206) );
  XOR U1221 ( .A(n1209), .B(n1189), .Z(n1199) );
  NAND U1222 ( .A(n374), .B(n1128), .Z(n1189) );
  IV U1223 ( .A(n1191), .Z(n1209) );
  XNOR U1224 ( .A(n1211), .B(n1198), .Z(n1045) );
  NAND U1225 ( .A(n540), .B(n784), .Z(n1198) );
  IV U1226 ( .A(n1197), .Z(n1211) );
  XNOR U1227 ( .A(n1194), .B(n1212), .Z(n1197) );
  AND U1228 ( .A(n855), .B(n475), .Z(n1212) );
  XOR U1229 ( .A(n1213), .B(n1214), .Z(n1194) );
  ANDN U1230 ( .A(n1215), .B(n1216), .Z(n1214) );
  XNOR U1231 ( .A(n1217), .B(n1213), .Z(n1215) );
  XNOR U1232 ( .A(n1218), .B(n1219), .Z(n1047) );
  IV U1233 ( .A(n1207), .Z(n1219) );
  XNOR U1234 ( .A(n1204), .B(n1220), .Z(n1207) );
  AND U1235 ( .A(n374), .B(e_input[0]), .Z(n1220) );
  XNOR U1236 ( .A(n1203), .B(g_input[10]), .Z(n1202) );
  NOR U1237 ( .A(n1221), .B(n1222), .Z(n1203) );
  XOR U1238 ( .A(n1223), .B(n1224), .Z(n1204) );
  ANDN U1239 ( .A(n1225), .B(n1226), .Z(n1224) );
  XNOR U1240 ( .A(n1227), .B(n1223), .Z(n1225) );
  XOR U1241 ( .A(n1228), .B(n1208), .Z(n1218) );
  NAND U1242 ( .A(n423), .B(n1128), .Z(n1208) );
  IV U1243 ( .A(n1210), .Z(n1228) );
  XNOR U1244 ( .A(n1230), .B(n1217), .Z(n1072) );
  NAND U1245 ( .A(n605), .B(n784), .Z(n1217) );
  IV U1246 ( .A(n1216), .Z(n1230) );
  XNOR U1247 ( .A(n1213), .B(n1231), .Z(n1216) );
  AND U1248 ( .A(n855), .B(n540), .Z(n1231) );
  XOR U1249 ( .A(n1232), .B(n1233), .Z(n1213) );
  ANDN U1250 ( .A(n1234), .B(n1235), .Z(n1233) );
  XNOR U1251 ( .A(n1236), .B(n1232), .Z(n1234) );
  XNOR U1252 ( .A(n1237), .B(n1238), .Z(n1074) );
  IV U1253 ( .A(n1226), .Z(n1238) );
  XNOR U1254 ( .A(n1223), .B(n1239), .Z(n1226) );
  AND U1255 ( .A(n423), .B(e_input[0]), .Z(n1239) );
  XOR U1256 ( .A(n1221), .B(g_input[9]), .Z(n1222) );
  NANDN U1257 ( .B(n1240), .A(n1241), .Z(n1221) );
  XOR U1258 ( .A(n1242), .B(n1243), .Z(n1223) );
  ANDN U1259 ( .A(n1244), .B(n1245), .Z(n1243) );
  XNOR U1260 ( .A(n1246), .B(n1242), .Z(n1244) );
  XOR U1261 ( .A(n1247), .B(n1227), .Z(n1237) );
  NAND U1262 ( .A(n475), .B(n1128), .Z(n1227) );
  IV U1263 ( .A(n1229), .Z(n1247) );
  NAND U1264 ( .A(n673), .B(n784), .Z(n1236) );
  XNOR U1265 ( .A(n1232), .B(n1249), .Z(n1235) );
  AND U1266 ( .A(n855), .B(n605), .Z(n1249) );
  XNOR U1267 ( .A(n1253), .B(n1250), .Z(n1252) );
  XNOR U1268 ( .A(n1242), .B(n1255), .Z(n1245) );
  AND U1269 ( .A(n475), .B(e_input[0]), .Z(n1255) );
  XNOR U1270 ( .A(n1259), .B(n1256), .Z(n1258) );
  XOR U1271 ( .A(n1260), .B(n1246), .Z(n1254) );
  NAND U1272 ( .A(n540), .B(n1128), .Z(n1246) );
  IV U1273 ( .A(n1248), .Z(n1260) );
  XNOR U1274 ( .A(n1261), .B(n1262), .Z(n1248) );
  AND U1275 ( .A(n1263), .B(n1264), .Z(n1262) );
  XOR U1276 ( .A(n1257), .B(n1265), .Z(n1264) );
  XNOR U1277 ( .A(n1259), .B(n1261), .Z(n1265) );
  NAND U1278 ( .A(n605), .B(n1128), .Z(n1259) );
  XOR U1279 ( .A(n1256), .B(n1266), .Z(n1257) );
  AND U1280 ( .A(n540), .B(e_input[0]), .Z(n1266) );
  XNOR U1281 ( .A(n1270), .B(n1267), .Z(n1269) );
  XOR U1282 ( .A(n1251), .B(n1271), .Z(n1263) );
  XNOR U1283 ( .A(n1253), .B(n1261), .Z(n1271) );
  NANDN U1284 ( .B(n741), .A(n784), .Z(n1253) );
  XOR U1285 ( .A(n1250), .B(n1272), .Z(n1251) );
  AND U1286 ( .A(n855), .B(n673), .Z(n1272) );
  XOR U1287 ( .A(n1273), .B(n1274), .Z(n1250) );
  AND U1288 ( .A(n1275), .B(n1276), .Z(n1274) );
  XNOR U1289 ( .A(n1277), .B(n1273), .Z(n1276) );
  XOR U1290 ( .A(n1278), .B(n1279), .Z(n1261) );
  AND U1291 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U1292 ( .A(n1268), .B(n1282), .Z(n1281) );
  XNOR U1293 ( .A(n1270), .B(n1278), .Z(n1282) );
  NAND U1294 ( .A(n673), .B(n1128), .Z(n1270) );
  XOR U1295 ( .A(n1267), .B(n1283), .Z(n1268) );
  AND U1296 ( .A(n605), .B(e_input[0]), .Z(n1283) );
  XNOR U1297 ( .A(n1287), .B(n1284), .Z(n1286) );
  XOR U1298 ( .A(n1275), .B(n1288), .Z(n1280) );
  XNOR U1299 ( .A(n1277), .B(n1278), .Z(n1288) );
  NANDN U1300 ( .B(n818), .A(n784), .Z(n1277) );
  XOR U1301 ( .A(n1273), .B(n1289), .Z(n1275) );
  ANDN U1302 ( .A(n855), .B(n741), .Z(n1289) );
  XOR U1303 ( .A(n1290), .B(n1291), .Z(n1273) );
  AND U1304 ( .A(n1292), .B(n1293), .Z(n1291) );
  XNOR U1305 ( .A(n1294), .B(n1290), .Z(n1293) );
  XOR U1306 ( .A(n1295), .B(n1296), .Z(n1278) );
  AND U1307 ( .A(n1297), .B(n1298), .Z(n1296) );
  XOR U1308 ( .A(n1285), .B(n1299), .Z(n1298) );
  XNOR U1309 ( .A(n1287), .B(n1295), .Z(n1299) );
  NANDN U1310 ( .B(n741), .A(n1128), .Z(n1287) );
  XOR U1311 ( .A(n1284), .B(n1300), .Z(n1285) );
  AND U1312 ( .A(n673), .B(e_input[0]), .Z(n1300) );
  XOR U1313 ( .A(n1292), .B(n1304), .Z(n1297) );
  XNOR U1314 ( .A(n1294), .B(n1295), .Z(n1304) );
  NAND U1315 ( .A(n784), .B(n891), .Z(n1294) );
  XOR U1316 ( .A(n1290), .B(n1305), .Z(n1292) );
  ANDN U1317 ( .A(n855), .B(n818), .Z(n1305) );
  NAND U1318 ( .A(n784), .B(n1111), .Z(n1308) );
  XNOR U1319 ( .A(n1306), .B(n1310), .Z(n1307) );
  AND U1320 ( .A(n891), .B(n855), .Z(n1310) );
  AND U1321 ( .A(n1311), .B(g_input[0]), .Z(n1306) );
  NANDN U1322 ( .B(n784), .A(n1312), .Z(n1311) );
  NAND U1323 ( .A(n1111), .B(n855), .Z(n1312) );
  XNOR U1324 ( .A(n1301), .B(n1316), .Z(n1302) );
  ANDN U1325 ( .A(e_input[0]), .B(n741), .Z(n1316) );
  XOR U1326 ( .A(n1319), .B(n1317), .Z(n1318) );
  ANDN U1327 ( .A(e_input[0]), .B(n818), .Z(n1319) );
  AND U1328 ( .A(n1128), .B(n891), .Z(n1320) );
  XOR U1329 ( .A(n1324), .B(n1303), .Z(n1315) );
  NANDN U1330 ( .B(n818), .A(n1128), .Z(n1303) );
  IV U1331 ( .A(n1309), .Z(n1324) );
  NAND U1332 ( .A(n1128), .B(n1111), .Z(n1323) );
  XNOR U1333 ( .A(n1321), .B(n1325), .Z(n1322) );
  AND U1334 ( .A(n891), .B(e_input[0]), .Z(n1325) );
  AND U1335 ( .A(n1326), .B(g_input[0]), .Z(n1321) );
  NANDN U1336 ( .B(n1128), .A(n1327), .Z(n1326) );
  NAND U1337 ( .A(n1111), .B(e_input[0]), .Z(n1327) );
  XNOR U1338 ( .A(n1329), .B(n881), .Z(n871) );
  XNOR U1339 ( .A(n868), .B(n869), .Z(n881) );
  NAND U1340 ( .A(n312), .B(n673), .Z(n869) );
  XNOR U1341 ( .A(n867), .B(n1330), .Z(n868) );
  AND U1342 ( .A(n605), .B(n353), .Z(n1330) );
  XNOR U1343 ( .A(n1334), .B(n1331), .Z(n1333) );
  XNOR U1344 ( .A(n880), .B(n870), .Z(n1329) );
  XOR U1345 ( .A(n1335), .B(n1336), .Z(n870) );
  XNOR U1346 ( .A(n875), .B(n1338), .Z(n876) );
  AND U1347 ( .A(n475), .B(n460), .Z(n1338) );
  XNOR U1348 ( .A(n1241), .B(g_input[8]), .Z(n1240) );
  NOR U1349 ( .A(n1339), .B(n1340), .Z(n1241) );
  XOR U1350 ( .A(n1341), .B(n1342), .Z(n875) );
  AND U1351 ( .A(n1343), .B(n1344), .Z(n1342) );
  XNOR U1352 ( .A(n1345), .B(n1341), .Z(n1344) );
  XOR U1353 ( .A(n1346), .B(n877), .Z(n1337) );
  NAND U1354 ( .A(n406), .B(n540), .Z(n877) );
  IV U1355 ( .A(n879), .Z(n1346) );
  XNOR U1356 ( .A(n1347), .B(n1348), .Z(n879) );
  AND U1357 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U1358 ( .A(n1343), .B(n1351), .Z(n1350) );
  XNOR U1359 ( .A(n1345), .B(n1347), .Z(n1351) );
  NAND U1360 ( .A(n406), .B(n605), .Z(n1345) );
  XOR U1361 ( .A(n1341), .B(n1352), .Z(n1343) );
  AND U1362 ( .A(n540), .B(n460), .Z(n1352) );
  XOR U1363 ( .A(n1339), .B(g_input[7]), .Z(n1340) );
  NANDN U1364 ( .B(n1353), .A(n1354), .Z(n1339) );
  XOR U1365 ( .A(n1355), .B(n1356), .Z(n1341) );
  AND U1366 ( .A(n1357), .B(n1358), .Z(n1356) );
  XNOR U1367 ( .A(n1359), .B(n1355), .Z(n1358) );
  XOR U1368 ( .A(n1332), .B(n1360), .Z(n1349) );
  XNOR U1369 ( .A(n1334), .B(n1347), .Z(n1360) );
  NANDN U1370 ( .B(n741), .A(n312), .Z(n1334) );
  XOR U1371 ( .A(n1331), .B(n1361), .Z(n1332) );
  AND U1372 ( .A(n673), .B(n353), .Z(n1361) );
  XNOR U1373 ( .A(n1365), .B(n1362), .Z(n1364) );
  XOR U1374 ( .A(n1366), .B(n1367), .Z(n1347) );
  AND U1375 ( .A(n1368), .B(n1369), .Z(n1367) );
  XOR U1376 ( .A(n1357), .B(n1370), .Z(n1369) );
  XNOR U1377 ( .A(n1359), .B(n1366), .Z(n1370) );
  NAND U1378 ( .A(n406), .B(n673), .Z(n1359) );
  XOR U1379 ( .A(n1355), .B(n1371), .Z(n1357) );
  AND U1380 ( .A(n605), .B(n460), .Z(n1371) );
  XNOR U1381 ( .A(n1354), .B(g_input[6]), .Z(n1353) );
  NOR U1382 ( .A(n1372), .B(n1373), .Z(n1354) );
  XOR U1383 ( .A(n1374), .B(n1375), .Z(n1355) );
  AND U1384 ( .A(n1376), .B(n1377), .Z(n1375) );
  XNOR U1385 ( .A(n1378), .B(n1374), .Z(n1377) );
  XOR U1386 ( .A(n1363), .B(n1379), .Z(n1368) );
  XNOR U1387 ( .A(n1365), .B(n1366), .Z(n1379) );
  NANDN U1388 ( .B(n818), .A(n312), .Z(n1365) );
  XOR U1389 ( .A(n1362), .B(n1380), .Z(n1363) );
  ANDN U1390 ( .A(n353), .B(n741), .Z(n1380) );
  XNOR U1391 ( .A(n1384), .B(n1381), .Z(n1383) );
  XOR U1392 ( .A(n1385), .B(n1386), .Z(n1366) );
  AND U1393 ( .A(n1387), .B(n1388), .Z(n1386) );
  XOR U1394 ( .A(n1376), .B(n1389), .Z(n1388) );
  XNOR U1395 ( .A(n1378), .B(n1385), .Z(n1389) );
  NANDN U1396 ( .B(n741), .A(n406), .Z(n1378) );
  XOR U1397 ( .A(n1374), .B(n1390), .Z(n1376) );
  AND U1398 ( .A(n673), .B(n460), .Z(n1390) );
  XOR U1399 ( .A(n1372), .B(g_input[5]), .Z(n1373) );
  NANDN U1400 ( .B(n1391), .A(n1392), .Z(n1372) );
  XOR U1401 ( .A(n1393), .B(n1394), .Z(n1374) );
  ANDN U1402 ( .A(n1395), .B(n1396), .Z(n1394) );
  XNOR U1403 ( .A(n1397), .B(n1393), .Z(n1395) );
  XOR U1404 ( .A(n1382), .B(n1398), .Z(n1387) );
  XNOR U1405 ( .A(n1384), .B(n1385), .Z(n1398) );
  NAND U1406 ( .A(n312), .B(n891), .Z(n1384) );
  XOR U1407 ( .A(n1381), .B(n1399), .Z(n1382) );
  ANDN U1408 ( .A(n353), .B(n818), .Z(n1399) );
  XOR U1409 ( .A(n1400), .B(n1401), .Z(n1381) );
  ANDN U1410 ( .A(n1402), .B(n1403), .Z(n1401) );
  XNOR U1411 ( .A(n1404), .B(n1400), .Z(n1402) );
  NAND U1412 ( .A(n312), .B(n1111), .Z(n1404) );
  XNOR U1413 ( .A(n1400), .B(n1406), .Z(n1403) );
  AND U1414 ( .A(n891), .B(n353), .Z(n1406) );
  AND U1415 ( .A(n1407), .B(g_input[0]), .Z(n1400) );
  NANDN U1416 ( .B(n312), .A(n1408), .Z(n1407) );
  NAND U1417 ( .A(n1111), .B(n353), .Z(n1408) );
  XNOR U1418 ( .A(n1393), .B(n1412), .Z(n1396) );
  ANDN U1419 ( .A(n460), .B(n741), .Z(n1412) );
  XOR U1420 ( .A(n1413), .B(n1414), .Z(n1393) );
  AND U1421 ( .A(n1415), .B(n1416), .Z(n1414) );
  XOR U1422 ( .A(n1417), .B(n1413), .Z(n1416) );
  ANDN U1423 ( .A(n460), .B(n818), .Z(n1417) );
  XOR U1424 ( .A(n1418), .B(n1413), .Z(n1415) );
  AND U1425 ( .A(n891), .B(n406), .Z(n1418) );
  XOR U1426 ( .A(n1419), .B(n1420), .Z(n1413) );
  ANDN U1427 ( .A(n1421), .B(n1422), .Z(n1420) );
  XNOR U1428 ( .A(n1423), .B(n1419), .Z(n1421) );
  XOR U1429 ( .A(n1424), .B(n1397), .Z(n1411) );
  NANDN U1430 ( .B(n818), .A(n406), .Z(n1397) );
  IV U1431 ( .A(n1405), .Z(n1424) );
  XOR U1432 ( .A(n1425), .B(n1423), .Z(n1405) );
  NAND U1433 ( .A(n406), .B(n1111), .Z(n1423) );
  IV U1434 ( .A(n1422), .Z(n1425) );
  XNOR U1435 ( .A(n1419), .B(n1426), .Z(n1422) );
  AND U1436 ( .A(n891), .B(n460), .Z(n1426) );
  AND U1437 ( .A(n1427), .B(g_input[0]), .Z(n1419) );
  NANDN U1438 ( .B(n406), .A(n1428), .Z(n1427) );
  NAND U1439 ( .A(n1111), .B(n460), .Z(n1428) );
  XNOR U1440 ( .A(n884), .B(n1432), .Z(n885) );
  ANDN U1441 ( .A(n280), .B(n741), .Z(n1432) );
  XNOR U1442 ( .A(n1392), .B(g_input[4]), .Z(n1391) );
  NOR U1443 ( .A(n1433), .B(n1434), .Z(n1392) );
  XOR U1444 ( .A(n1435), .B(n1436), .Z(n884) );
  AND U1445 ( .A(n1437), .B(n1438), .Z(n1436) );
  XOR U1446 ( .A(n1439), .B(n1435), .Z(n1438) );
  ANDN U1447 ( .A(n280), .B(n818), .Z(n1439) );
  XOR U1448 ( .A(n1440), .B(n1435), .Z(n1437) );
  AND U1449 ( .A(n891), .B(n242), .Z(n1440) );
  XOR U1450 ( .A(n1441), .B(n1442), .Z(n1435) );
  ANDN U1451 ( .A(n1443), .B(n1444), .Z(n1442) );
  XNOR U1452 ( .A(n1445), .B(n1441), .Z(n1443) );
  XOR U1453 ( .A(n1446), .B(n886), .Z(n1431) );
  NANDN U1454 ( .B(n818), .A(n242), .Z(n886) );
  NANDN U1455 ( .B(n1447), .A(n1448), .Z(n1433) );
  IV U1456 ( .A(n888), .Z(n1446) );
  NAND U1457 ( .A(n242), .B(n1111), .Z(n1445) );
  XNOR U1458 ( .A(n1441), .B(n1449), .Z(n1444) );
  AND U1459 ( .A(n891), .B(n280), .Z(n1449) );
  AND U1460 ( .A(n1450), .B(g_input[0]), .Z(n1441) );
  NANDN U1461 ( .B(n242), .A(n1451), .Z(n1450) );
  NAND U1462 ( .A(n1111), .B(n280), .Z(n1451) );
  XNOR U1463 ( .A(n1452), .B(e_input[12]), .Z(n280) );
  NAND U1464 ( .A(n1453), .B(e_input[15]), .Z(n1452) );
  XOR U1465 ( .A(n1454), .B(e_input[12]), .Z(n1453) );
  XNOR U1466 ( .A(n895), .B(n896), .Z(n890) );
  NANDN U1467 ( .B(n187), .A(n1111), .Z(n896) );
  XNOR U1468 ( .A(n894), .B(n1456), .Z(n895) );
  AND U1469 ( .A(n891), .B(n211), .Z(n1456) );
  XNOR U1470 ( .A(n1448), .B(g_input[2]), .Z(n1447) );
  AND U1471 ( .A(n1458), .B(g_input[0]), .Z(n894) );
  NAND U1472 ( .A(n1459), .B(n187), .Z(n1458) );
  NANDN U1473 ( .B(n1460), .A(n1461), .Z(n187) );
  ANDN U1474 ( .A(e_input[15]), .B(n1462), .Z(n1461) );
  NAND U1475 ( .A(n1111), .B(n211), .Z(n1459) );
  XOR U1476 ( .A(n1462), .B(e_input[14]), .Z(n1460) );
  OR U1477 ( .A(n1455), .B(n1463), .Z(n1462) );
  XOR U1478 ( .A(n1463), .B(e_input[13]), .Z(n1455) );
  OR U1479 ( .A(n1454), .B(n1464), .Z(n1463) );
  XOR U1480 ( .A(n1464), .B(e_input[12]), .Z(n1454) );
  OR U1481 ( .A(n1410), .B(n1465), .Z(n1464) );
  XOR U1482 ( .A(n1465), .B(e_input[11]), .Z(n1410) );
  OR U1483 ( .A(n1409), .B(n1466), .Z(n1465) );
  XOR U1484 ( .A(n1466), .B(e_input[10]), .Z(n1409) );
  OR U1485 ( .A(n1430), .B(n1467), .Z(n1466) );
  XOR U1486 ( .A(n1467), .B(e_input[9]), .Z(n1430) );
  OR U1487 ( .A(n1429), .B(n1468), .Z(n1467) );
  XOR U1488 ( .A(n1468), .B(e_input[8]), .Z(n1429) );
  OR U1489 ( .A(n1121), .B(n1469), .Z(n1468) );
  XOR U1490 ( .A(n1469), .B(e_input[7]), .Z(n1121) );
  OR U1491 ( .A(n1120), .B(n1470), .Z(n1469) );
  XOR U1492 ( .A(n1470), .B(e_input[6]), .Z(n1120) );
  OR U1493 ( .A(n1116), .B(n1471), .Z(n1470) );
  XOR U1494 ( .A(n1471), .B(e_input[5]), .Z(n1116) );
  OR U1495 ( .A(n1115), .B(n1472), .Z(n1471) );
  XOR U1496 ( .A(n1472), .B(e_input[4]), .Z(n1115) );
  OR U1497 ( .A(n1314), .B(n1473), .Z(n1472) );
  XOR U1498 ( .A(n1473), .B(e_input[3]), .Z(n1314) );
  OR U1499 ( .A(n1313), .B(n1474), .Z(n1473) );
  XOR U1500 ( .A(n1474), .B(e_input[2]), .Z(n1313) );
  NANDN U1501 ( .B(e_input[0]), .A(n1328), .Z(n1474) );
  XNOR U1502 ( .A(e_input[0]), .B(e_input[1]), .Z(n1328) );
  XOR U1503 ( .A(g_input[0]), .B(g_input[1]), .Z(n1457) );
  NANDN U1504 ( .B(n830), .A(n102), .Z(n154) );
  IV U1505 ( .A(rst), .Z(n102) );
  NAND U1506 ( .A(n1475), .B(n1476), .Z(n830) );
  AND U1507 ( .A(n1477), .B(n1478), .Z(n1476) );
  ANDN U1508 ( .A(n1479), .B(\_MxM/n[3] ), .Z(n1478) );
  NOR U1509 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n1479) );
  ANDN U1510 ( .A(n1480), .B(\_MxM/n[13] ), .Z(n1477) );
  NOR U1511 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n1480) );
  AND U1512 ( .A(n1481), .B(n1482), .Z(n1475) );
  ANDN U1513 ( .A(n1483), .B(n1484), .Z(n1482) );
  ANDN U1514 ( .A(\_MxM/N19 ), .B(\_MxM/n[10] ), .Z(n1483) );
  NOR U1515 ( .A(n1485), .B(n1486), .Z(n1481) );
  AND U1516 ( .A(n1487), .B(n1488), .Z(\_MxM/N32 ) );
  XOR U1517 ( .A(\_MxM/n[13] ), .B(\_MxM/add_39/carry[13] ), .Z(n1488) );
  AND U1518 ( .A(\_MxM/N17 ), .B(n1487), .Z(\_MxM/N31 ) );
  AND U1519 ( .A(\_MxM/N16 ), .B(n1487), .Z(\_MxM/N30 ) );
  AND U1520 ( .A(\_MxM/N15 ), .B(n1487), .Z(\_MxM/N29 ) );
  AND U1521 ( .A(\_MxM/N14 ), .B(n1487), .Z(\_MxM/N28 ) );
  AND U1522 ( .A(\_MxM/N13 ), .B(n1487), .Z(\_MxM/N27 ) );
  AND U1523 ( .A(\_MxM/N12 ), .B(n1487), .Z(\_MxM/N26 ) );
  AND U1524 ( .A(\_MxM/N11 ), .B(n1487), .Z(\_MxM/N25 ) );
  AND U1525 ( .A(\_MxM/N10 ), .B(n1487), .Z(\_MxM/N24 ) );
  AND U1526 ( .A(\_MxM/N9 ), .B(n1487), .Z(\_MxM/N23 ) );
  AND U1527 ( .A(\_MxM/N8 ), .B(n1487), .Z(\_MxM/N22 ) );
  AND U1528 ( .A(\_MxM/N7 ), .B(n1487), .Z(\_MxM/N21 ) );
  AND U1529 ( .A(\_MxM/N6 ), .B(n1487), .Z(\_MxM/N20 ) );
  NAND U1530 ( .A(n1489), .B(n1490), .Z(n1487) );
  AND U1531 ( .A(n1491), .B(n1492), .Z(n1490) );
  ANDN U1532 ( .A(n1493), .B(n1486), .Z(n1492) );
  OR U1533 ( .A(\_MxM/n[6] ), .B(\_MxM/n[7] ), .Z(n1486) );
  NOR U1534 ( .A(\_MxM/N19 ), .B(n1484), .Z(n1493) );
  OR U1535 ( .A(\_MxM/n[4] ), .B(\_MxM/n[5] ), .Z(n1484) );
  AND U1536 ( .A(\_MxM/n[13] ), .B(n1494), .Z(n1491) );
  ANDN U1537 ( .A(\_MxM/n[10] ), .B(n1485), .Z(n1494) );
  OR U1538 ( .A(\_MxM/n[12] ), .B(\_MxM/n[11] ), .Z(n1485) );
  AND U1539 ( .A(n1495), .B(n1496), .Z(n1489) );
  AND U1540 ( .A(\_MxM/n[3] ), .B(n1497), .Z(n1496) );
  AND U1541 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n1497) );
  AND U1542 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n1495) );
  IV U1543 ( .A(\_MxM/n[0] ), .Z(\_MxM/N19 ) );
endmodule

