
module MxM_TG_W16_N1000 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MxM/n244 , \_MxM/n243 , \_MxM/n242 , \_MxM/n241 , \_MxM/n240 ,
         \_MxM/n239 , \_MxM/n238 , \_MxM/n237 , \_MxM/n236 , \_MxM/n235 ,
         \_MxM/n234 , \_MxM/n233 , \_MxM/n232 , \_MxM/n231 , \_MxM/n230 ,
         \_MxM/n229 , \_MxM/n228 , \_MxM/n227 , \_MxM/n226 , \_MxM/n225 ,
         \_MxM/n224 , \_MxM/n223 , \_MxM/n222 , \_MxM/n221 , \_MxM/n220 ,
         \_MxM/n219 , \_MxM/n218 , \_MxM/n217 , \_MxM/n216 , \_MxM/n215 ,
         \_MxM/n214 , \_MxM/n213 , \_MxM/n212 , \_MxM/n211 , \_MxM/n210 ,
         \_MxM/n209 , \_MxM/n208 , \_MxM/n207 , \_MxM/n206 , \_MxM/n205 ,
         \_MxM/n204 , \_MxM/n203 , \_MxM/N15 , \_MxM/N14 , \_MxM/N13 ,
         \_MxM/N12 , \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/n[0] ,
         \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] ,
         \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/Y0[0] ,
         \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] , \_MxM/Y0[4] , \_MxM/Y0[5] ,
         \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/Y0[8] , \_MxM/Y0[9] , \_MxM/Y0[10] ,
         \_MxM/Y0[11] , \_MxM/Y0[12] , \_MxM/Y0[13] , \_MxM/Y0[14] ,
         \_MxM/Y0[15] , \_MxM/add_39/carry[9] , \_MxM/add_39/carry[8] ,
         \_MxM/add_39/carry[7] , \_MxM/add_39/carry[6] ,
         \_MxM/add_39/carry[5] , \_MxM/add_39/carry[4] ,
         \_MxM/add_39/carry[3] , \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n203 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n204 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n205 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n206 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n207 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n208 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n209 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n210 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n211 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n212 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n213 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n214 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n215 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n216 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n217 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n218 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/n219 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/n220 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/n221 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/n222 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/n223 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/n224 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/n225 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/n226 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n227 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n228 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n229 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n230 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n231 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n232 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n233 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n234 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/n235 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/n236 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/n237 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n238 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n239 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n240 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n241 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n242 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n243 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n244 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N14 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N15 ) );
  MUX U1 ( .IN0(n1), .IN1(n1317), .SEL(n1318), .F(n1301) );
  IV U2 ( .A(n1319), .Z(n1) );
  MUX U3 ( .IN0(n2), .IN1(n984), .SEL(n985), .F(n961) );
  IV U4 ( .A(n986), .Z(n2) );
  MUX U5 ( .IN0(n1392), .IN1(n1410), .SEL(n1394), .F(n1373) );
  XOR U6 ( .A(n1175), .B(n1165), .Z(n981) );
  XOR U7 ( .A(n987), .B(n969), .Z(n973) );
  MUX U8 ( .IN0(n3), .IN1(n734), .SEL(n735), .F(n664) );
  IV U9 ( .A(n736), .Z(n3) );
  MUX U10 ( .IN0(n4), .IN1(n895), .SEL(n896), .F(n820) );
  IV U11 ( .A(n897), .Z(n4) );
  MUX U12 ( .IN0(n5), .IN1(n961), .SEL(n962), .F(n938) );
  IV U13 ( .A(n963), .Z(n5) );
  MUX U14 ( .IN0(n6), .IN1(n1157), .SEL(n1158), .F(n1147) );
  IV U15 ( .A(n1159), .Z(n6) );
  XOR U16 ( .A(n1160), .B(n1152), .Z(n958) );
  MUX U17 ( .IN0(n1112), .IN1(n1115), .SEL(n1113), .F(n1097) );
  MUX U18 ( .IN0(n7), .IN1(n459), .SEL(n460), .F(n408) );
  IV U19 ( .A(n461), .Z(n7) );
  MUX U20 ( .IN0(n8), .IN1(n811), .SEL(n812), .F(n734) );
  IV U21 ( .A(n813), .Z(n8) );
  XNOR U22 ( .A(n1455), .B(n1456), .Z(n899) );
  XOR U23 ( .A(n962), .B(n963), .Z(n974) );
  MUX U24 ( .IN0(n9), .IN1(n911), .SEL(n912), .F(n849) );
  IV U25 ( .A(n913), .Z(n9) );
  XOR U26 ( .A(n1148), .B(n1149), .Z(n956) );
  MUX U27 ( .IN0(n10), .IN1(n588), .SEL(n589), .F(n523) );
  IV U28 ( .A(n590), .Z(n10) );
  MUX U29 ( .IN0(e_input[8]), .IN1(n1440), .SEL(e_input[15]), .F(n471) );
  MUX U30 ( .IN0(n1153), .IN1(n11), .SEL(n1152), .F(n1144) );
  IV U31 ( .A(n1151), .Z(n11) );
  MUX U32 ( .IN0(e_input[13]), .IN1(n1466), .SEL(e_input[15]), .F(n253) );
  MUX U33 ( .IN0(n1328), .IN1(n1331), .SEL(n1329), .F(n1312) );
  MUX U34 ( .IN0(n12), .IN1(n938), .SEL(n939), .F(n919) );
  IV U35 ( .A(n940), .Z(n12) );
  MUX U36 ( .IN0(n13), .IN1(n1147), .SEL(n1148), .F(n926) );
  IV U37 ( .A(n1149), .Z(n13) );
  XOR U38 ( .A(n964), .B(n946), .Z(n950) );
  MUX U39 ( .IN0(e_input[9]), .IN1(n1441), .SEL(e_input[15]), .F(n417) );
  MUX U40 ( .IN0(n294), .IN1(n14), .SEL(n293), .F(n255) );
  IV U41 ( .A(n292), .Z(n14) );
  MUX U42 ( .IN0(e_input[11]), .IN1(n1421), .SEL(e_input[15]), .F(n323) );
  MUX U43 ( .IN0(n384), .IN1(n382), .SEL(n383), .F(n337) );
  MUX U44 ( .IN0(n15), .IN1(n177), .SEL(n176), .F(n185) );
  IV U45 ( .A(n188), .Z(n15) );
  MUX U46 ( .IN0(n16), .IN1(n1332), .SEL(n1333), .F(n1328) );
  IV U47 ( .A(n1334), .Z(n16) );
  XOR U48 ( .A(n1158), .B(n1159), .Z(n979) );
  MUX U49 ( .IN0(n17), .IN1(n715), .SEL(n716), .F(n646) );
  IV U50 ( .A(n717), .Z(n17) );
  MUX U51 ( .IN0(n18), .IN1(n774), .SEL(n775), .F(n711) );
  IV U52 ( .A(n776), .Z(n18) );
  MUX U53 ( .IN0(e_input[10]), .IN1(n1420), .SEL(e_input[15]), .F(n364) );
  MUX U54 ( .IN0(n474), .IN1(n19), .SEL(n473), .F(n419) );
  IV U55 ( .A(n472), .Z(n19) );
  MUX U56 ( .IN0(n550), .IN1(n548), .SEL(n549), .F(n483) );
  XNOR U57 ( .A(n1442), .B(n896), .Z(n900) );
  XOR U58 ( .A(n186), .B(n207), .Z(n205) );
  MUX U59 ( .IN0(n1373), .IN1(n1391), .SEL(n1375), .F(n1342) );
  MUX U60 ( .IN0(n1261), .IN1(n1283), .SEL(n1263), .F(n1243) );
  MUX U61 ( .IN0(n20), .IN1(n919), .SEL(n920), .F(n857) );
  IV U62 ( .A(n921), .Z(n20) );
  MUX U63 ( .IN0(n21), .IN1(n1164), .SEL(n1165), .F(n1151) );
  IV U64 ( .A(n1166), .Z(n21) );
  MUX U65 ( .IN0(n22), .IN1(n886), .SEL(n887), .F(n811) );
  IV U66 ( .A(n888), .Z(n22) );
  MUX U67 ( .IN0(g_input[11]), .IN1(n1195), .SEL(g_input[15]), .F(n340) );
  MUX U68 ( .IN0(n422), .IN1(n27), .SEL(n421), .F(n371) );
  MUX U69 ( .IN0(n683), .IN1(n681), .SEL(n682), .F(n613) );
  MUX U70 ( .IN0(n713), .IN1(n23), .SEL(n712), .F(n641) );
  IV U71 ( .A(n711), .Z(n23) );
  NAND U72 ( .A(n255), .B(n290), .Z(n289) );
  XOR U73 ( .A(n233), .B(n241), .Z(n239) );
  MUX U74 ( .IN0(n24), .IN1(n1179), .SEL(n1180), .F(n1164) );
  IV U75 ( .A(n1181), .Z(n24) );
  MUX U76 ( .IN0(n25), .IN1(n726), .SEL(n727), .F(n656) );
  IV U77 ( .A(n728), .Z(n25) );
  MUX U78 ( .IN0(n26), .IN1(n782), .SEL(n783), .F(n715) );
  IV U79 ( .A(n784), .Z(n26) );
  MUX U80 ( .IN0(e_input[4]), .IN1(n1126), .SEL(e_input[15]), .F(n710) );
  XOR U81 ( .A(n1422), .B(n1407), .Z(n1347) );
  MUX U82 ( .IN0(n466), .IN1(n468), .SEL(n467), .F(n27) );
  IV U83 ( .A(n27), .Z(n420) );
  MUX U84 ( .IN0(n644), .IN1(n28), .SEL(n643), .F(n571) );
  IV U85 ( .A(n642), .Z(n28) );
  MUX U86 ( .IN0(n751), .IN1(n749), .SEL(n750), .F(n681) );
  MUX U87 ( .IN0(n869), .IN1(n29), .SEL(n868), .F(n792) );
  IV U88 ( .A(n867), .Z(n29) );
  XNOR U89 ( .A(n374), .B(n334), .Z(n338) );
  XOR U90 ( .A(n264), .B(n272), .Z(n270) );
  XOR U91 ( .A(n939), .B(n940), .Z(n951) );
  MUX U92 ( .IN0(n1267), .IN1(n1277), .SEL(n1269), .F(n1253) );
  MUX U93 ( .IN0(n1342), .IN1(n1372), .SEL(n1344), .F(n878) );
  XNOR U94 ( .A(n1119), .B(n1120), .Z(n1103) );
  MUX U95 ( .IN0(g_input[9]), .IN1(n1233), .SEL(g_input[15]), .F(n434) );
  MUX U96 ( .IN0(g_input[12]), .IN1(n1177), .SEL(g_input[15]), .F(n295) );
  XOR U97 ( .A(n343), .B(n386), .Z(n344) );
  MUX U98 ( .IN0(n738), .IN1(n740), .SEL(n739), .F(n670) );
  MUX U99 ( .IN0(n780), .IN1(n778), .SEL(n779), .F(n705) );
  XOR U100 ( .A(n868), .B(n869), .Z(n875) );
  XNOR U101 ( .A(n371), .B(n414), .Z(n372) );
  XNOR U102 ( .A(n475), .B(n428), .Z(n432) );
  MUX U103 ( .IN0(n30), .IN1(n659), .SEL(n660), .F(n591) );
  IV U104 ( .A(n661), .Z(n30) );
  MUX U105 ( .IN0(n518), .IN1(n520), .SEL(n519), .F(n31) );
  IV U106 ( .A(n31), .Z(n454) );
  XOR U107 ( .A(n301), .B(n309), .Z(n307) );
  MUX U108 ( .IN0(n1259), .IN1(n32), .SEL(n1109), .F(n1240) );
  IV U109 ( .A(n1108), .Z(n32) );
  MUX U110 ( .IN0(n1105), .IN1(n1103), .SEL(n1104), .F(n1076) );
  XOR U111 ( .A(n1150), .B(n1144), .Z(n935) );
  MUX U112 ( .IN0(n33), .IN1(n878), .SEL(n879), .F(n803) );
  IV U113 ( .A(n880), .Z(n33) );
  MUX U114 ( .IN0(n34), .IN1(n926), .SEL(n927), .F(n867) );
  IV U115 ( .A(n928), .Z(n34) );
  XOR U116 ( .A(n941), .B(n912), .Z(n916) );
  MUX U117 ( .IN0(n602), .IN1(n604), .SEL(n603), .F(n537) );
  MUX U118 ( .IN0(n828), .IN1(n826), .SEL(n827), .F(n749) );
  XOR U119 ( .A(n1348), .B(n887), .Z(n891) );
  XNOR U120 ( .A(n423), .B(n379), .Z(n383) );
  MUX U121 ( .IN0(n35), .IN1(n462), .SEL(n463), .F(n411) );
  IV U122 ( .A(n464), .Z(n35) );
  MUX U123 ( .IN0(n36), .IN1(n577), .SEL(n578), .F(n517) );
  IV U124 ( .A(n579), .Z(n36) );
  NAND U125 ( .A(n641), .B(n709), .Z(n708) );
  MUX U126 ( .IN0(n583), .IN1(n585), .SEL(n584), .F(n518) );
  MUX U127 ( .IN0(n37), .IN1(n557), .SEL(n558), .F(n492) );
  IV U128 ( .A(\_MxM/Y0[5] ), .Z(n37) );
  XOR U129 ( .A(n346), .B(n354), .Z(n352) );
  MUX U130 ( .IN0(n38), .IN1(n1312), .SEL(n1313), .F(n1295) );
  IV U131 ( .A(n1314), .Z(n38) );
  MUX U132 ( .IN0(g_input[1]), .IN1(n1468), .SEL(g_input[15]), .F(n1122) );
  MUX U133 ( .IN0(n39), .IN1(n523), .SEL(n524), .F(n459) );
  IV U134 ( .A(n525), .Z(n39) );
  MUX U135 ( .IN0(g_input[6]), .IN1(n1364), .SEL(g_input[15]), .F(n616) );
  MUX U136 ( .IN0(g_input[7]), .IN1(n1351), .SEL(g_input[15]), .F(n551) );
  MUX U137 ( .IN0(g_input[5]), .IN1(n1384), .SEL(g_input[15]), .F(n684) );
  MUX U138 ( .IN0(n40), .IN1(n857), .SEL(n858), .F(n782) );
  IV U139 ( .A(n859), .Z(n40) );
  XOR U140 ( .A(n927), .B(n928), .Z(n933) );
  MUX U141 ( .IN0(n670), .IN1(n672), .SEL(n671), .F(n602) );
  XNOR U142 ( .A(n909), .B(n850), .Z(n854) );
  XOR U143 ( .A(n261), .B(n296), .Z(n262) );
  MUX U144 ( .IN0(n41), .IN1(n326), .SEL(n327), .F(n279) );
  IV U145 ( .A(n328), .Z(n41) );
  NAND U146 ( .A(n419), .B(n470), .Z(n469) );
  MUX U147 ( .IN0(n573), .IN1(n571), .SEL(n572), .F(n515) );
  XNOR U148 ( .A(n605), .B(n545), .Z(n549) );
  MUX U149 ( .IN0(n42), .IN1(n806), .SEL(n807), .F(n729) );
  IV U150 ( .A(n808), .Z(n42) );
  MUX U151 ( .IN0(n43), .IN1(n653), .SEL(n652), .F(n583) );
  IV U152 ( .A(n651), .Z(n43) );
  MUX U153 ( .IN0(n44), .IN1(n622), .SEL(n623), .F(n557) );
  IV U154 ( .A(\_MxM/Y0[4] ), .Z(n44) );
  XOR U155 ( .A(n391), .B(n399), .Z(n397) );
  MUX U156 ( .IN0(n1076), .IN1(n45), .SEL(n1077), .F(n1049) );
  IV U157 ( .A(n1078), .Z(n45) );
  MUX U158 ( .IN0(n1168), .IN1(n46), .SEL(n981), .F(n1155) );
  IV U159 ( .A(n979), .Z(n46) );
  XNOR U160 ( .A(n1333), .B(n1334), .Z(n1320) );
  MUX U161 ( .IN0(n47), .IN1(n656), .SEL(n657), .F(n588) );
  IV U162 ( .A(n658), .Z(n47) );
  MUX U163 ( .IN0(g_input[3]), .IN1(n1445), .SEL(g_input[15]), .F(n48) );
  IV U164 ( .A(n48), .Z(n829) );
  MUX U165 ( .IN0(g_input[4]), .IN1(n1402), .SEL(g_input[15]), .F(n49) );
  IV U166 ( .A(n49), .Z(n752) );
  MUX U167 ( .IN0(n915), .IN1(n50), .SEL(n916), .F(n853) );
  IV U168 ( .A(n917), .Z(n50) );
  XOR U169 ( .A(n1246), .B(n1247), .Z(n1108) );
  MUX U170 ( .IN0(n339), .IN1(n337), .SEL(n338), .F(n284) );
  MUX U171 ( .IN0(n51), .IN1(n646), .SEL(n647), .F(n577) );
  IV U172 ( .A(n648), .Z(n51) );
  XOR U173 ( .A(n554), .B(n617), .Z(n555) );
  MUX U174 ( .IN0(n815), .IN1(n817), .SEL(n816), .F(n738) );
  MUX U175 ( .IN0(n901), .IN1(n899), .SEL(n900), .F(n826) );
  MUX U176 ( .IN0(n52), .IN1(n368), .SEL(n369), .F(n326) );
  IV U177 ( .A(n370), .Z(n52) );
  XOR U178 ( .A(n529), .B(n473), .Z(n467) );
  XNOR U179 ( .A(n540), .B(n480), .Z(n484) );
  MUX U180 ( .IN0(n53), .IN1(n591), .SEL(n592), .F(n526) );
  IV U181 ( .A(n593), .Z(n53) );
  XOR U182 ( .A(n704), .B(n642), .Z(n643) );
  MUX U183 ( .IN0(n800), .IN1(n54), .SEL(n799), .F(n721) );
  IV U184 ( .A(n798), .Z(n54) );
  MUX U185 ( .IN0(n718), .IN1(n55), .SEL(n719), .F(n651) );
  IV U186 ( .A(n720), .Z(n55) );
  MUX U187 ( .IN0(n56), .IN1(n690), .SEL(n691), .F(n622) );
  IV U188 ( .A(\_MxM/Y0[3] ), .Z(n56) );
  XOR U189 ( .A(n446), .B(n452), .Z(n441) );
  MUX U190 ( .IN0(n57), .IN1(n1106), .SEL(n923), .F(n1079) );
  IV U191 ( .A(n922), .Z(n57) );
  MUX U192 ( .IN0(n1022), .IN1(n58), .SEL(n1023), .F(n995) );
  IV U193 ( .A(n1024), .Z(n58) );
  MUX U194 ( .IN0(e_input[1]), .IN1(n59), .SEL(e_input[15]), .F(n1139) );
  IV U195 ( .A(n1339), .Z(n59) );
  MUX U196 ( .IN0(e_input[6]), .IN1(n1131), .SEL(e_input[15]), .F(n576) );
  MUX U197 ( .IN0(e_input[3]), .IN1(n1325), .SEL(e_input[15]), .F(n795) );
  MUX U198 ( .IN0(n890), .IN1(n892), .SEL(n891), .F(n815) );
  MUX U199 ( .IN0(e_input[14]), .IN1(n1471), .SEL(e_input[15]), .F(n222) );
  NAND U200 ( .A(n320), .B(n363), .Z(n362) );
  XOR U201 ( .A(n594), .B(n534), .Z(n538) );
  XNOR U202 ( .A(n673), .B(n610), .Z(n614) );
  MUX U203 ( .IN0(n60), .IN1(n729), .SEL(n730), .F(n659) );
  IV U204 ( .A(n731), .Z(n60) );
  XNOR U205 ( .A(n772), .B(n712), .Z(n706) );
  MUX U206 ( .IN0(n785), .IN1(n61), .SEL(n786), .F(n718) );
  IV U207 ( .A(n787), .Z(n61) );
  MUX U208 ( .IN0(n62), .IN1(n264), .SEL(n265), .F(n233) );
  IV U209 ( .A(\_MxM/Y0[11] ), .Z(n62) );
  XOR U210 ( .A(n492), .B(n500), .Z(n498) );
  MUX U211 ( .IN0(n1240), .IN1(n63), .SEL(n1085), .F(n1221) );
  IV U212 ( .A(n1083), .Z(n63) );
  MUX U213 ( .IN0(n1295), .IN1(n1311), .SEL(n1297), .F(n1278) );
  MUX U214 ( .IN0(n972), .IN1(n64), .SEL(n973), .F(n949) );
  IV U215 ( .A(n974), .Z(n64) );
  XOR U216 ( .A(n920), .B(n921), .Z(n917) );
  XOR U217 ( .A(n1318), .B(n1319), .Z(n1133) );
  MUX U218 ( .IN0(n65), .IN1(n803), .SEL(n804), .F(n726) );
  IV U219 ( .A(n805), .Z(n65) );
  MUX U220 ( .IN0(g_input[10]), .IN1(n1213), .SEL(g_input[15]), .F(n385) );
  XNOR U221 ( .A(n1110), .B(n1100), .Z(n1104) );
  XOR U222 ( .A(n437), .B(n487), .Z(n438) );
  MUX U223 ( .IN0(n485), .IN1(n483), .SEL(n484), .F(n431) );
  MUX U224 ( .IN0(n707), .IN1(n705), .SEL(n706), .F(n642) );
  MUX U225 ( .IN0(g_input[13]), .IN1(n1163), .SEL(g_input[15]), .F(n258) );
  MUX U226 ( .IN0(n66), .IN1(n526), .SEL(n527), .F(n462) );
  IV U227 ( .A(n528), .Z(n66) );
  XOR U228 ( .A(n662), .B(n599), .Z(n603) );
  XNOR U229 ( .A(n818), .B(n746), .Z(n750) );
  MUX U230 ( .IN0(n67), .IN1(n881), .SEL(n882), .F(n806) );
  IV U231 ( .A(n883), .Z(n67) );
  MUX U232 ( .IN0(n68), .IN1(n870), .SEL(n871), .F(n798) );
  IV U233 ( .A(n872), .Z(n68) );
  MUX U234 ( .IN0(g_input[14]), .IN1(n1140), .SEL(g_input[15]), .F(n223) );
  MUX U235 ( .IN0(n281), .IN1(n69), .SEL(n280), .F(n249) );
  IV U236 ( .A(n279), .Z(n69) );
  XNOR U237 ( .A(n583), .B(n582), .Z(n635) );
  MUX U238 ( .IN0(\_MxM/Y0[13] ), .IN1(n70), .SEL(n187), .F(n179) );
  IV U239 ( .A(n186), .Z(n70) );
  MUX U240 ( .IN0(n71), .IN1(n346), .SEL(n347), .F(n301) );
  IV U241 ( .A(\_MxM/Y0[9] ), .Z(n71) );
  MUX U242 ( .IN0(n72), .IN1(n835), .SEL(n836), .F(n758) );
  IV U243 ( .A(\_MxM/Y0[1] ), .Z(n72) );
  XOR U244 ( .A(n557), .B(n565), .Z(n563) );
  MUX U245 ( .IN0(n1221), .IN1(n73), .SEL(n1058), .F(n1202) );
  IV U246 ( .A(n1056), .Z(n73) );
  MUX U247 ( .IN0(n995), .IN1(n74), .SEL(n996), .F(n972) );
  IV U248 ( .A(n997), .Z(n74) );
  MUX U249 ( .IN0(n1278), .IN1(n1294), .SEL(n1280), .F(n1267) );
  MUX U250 ( .IN0(n1155), .IN1(n75), .SEL(n958), .F(n1145) );
  IV U251 ( .A(n956), .Z(n75) );
  MUX U252 ( .IN0(g_input[8]), .IN1(n1251), .SEL(g_input[15]), .F(n486) );
  MUX U253 ( .IN0(g_input[2]), .IN1(n1458), .SEL(g_input[15]), .F(n902) );
  MUX U254 ( .IN0(n76), .IN1(n849), .SEL(n850), .F(n774) );
  IV U255 ( .A(n851), .Z(n76) );
  MUX U256 ( .IN0(n77), .IN1(n408), .SEL(n409), .F(n365) );
  IV U257 ( .A(n410), .Z(n77) );
  MUX U258 ( .IN0(n537), .IN1(n539), .SEL(n538), .F(n466) );
  MUX U259 ( .IN0(n615), .IN1(n613), .SEL(n614), .F(n548) );
  XOR U260 ( .A(n832), .B(n903), .Z(n833) );
  MUX U261 ( .IN0(n855), .IN1(n853), .SEL(n854), .F(n778) );
  XNOR U262 ( .A(n284), .B(n285), .Z(n283) );
  MUX U263 ( .IN0(n78), .IN1(n411), .SEL(n412), .F(n368) );
  IV U264 ( .A(n413), .Z(n78) );
  XOR U265 ( .A(n578), .B(n579), .Z(n573) );
  XOR U266 ( .A(n809), .B(n735), .Z(n739) );
  XNOR U267 ( .A(n893), .B(n823), .Z(n827) );
  NAND U268 ( .A(n792), .B(n865), .Z(n864) );
  XNOR U269 ( .A(n288), .B(n287), .Z(n281) );
  XNOR U270 ( .A(n683), .B(n682), .Z(n661) );
  MUX U271 ( .IN0(n723), .IN1(n721), .SEL(n722), .F(n79) );
  IV U272 ( .A(n79), .Z(n650) );
  MUX U273 ( .IN0(n860), .IN1(n80), .SEL(n861), .F(n785) );
  IV U274 ( .A(n862), .Z(n80) );
  MUX U275 ( .IN0(n454), .IN1(n81), .SEL(n455), .F(n405) );
  IV U276 ( .A(n456), .Z(n81) );
  MUX U277 ( .IN0(n82), .IN1(n233), .SEL(n234), .F(n186) );
  IV U278 ( .A(\_MxM/Y0[12] ), .Z(n82) );
  MUX U279 ( .IN0(n83), .IN1(n391), .SEL(n392), .F(n346) );
  IV U280 ( .A(\_MxM/Y0[8] ), .Z(n83) );
  XOR U281 ( .A(n622), .B(n630), .Z(n628) );
  MUX U282 ( .IN0(n1202), .IN1(n84), .SEL(n1031), .F(n1183) );
  IV U283 ( .A(n1029), .Z(n84) );
  MUX U284 ( .IN0(n85), .IN1(n1346), .SEL(n1347), .F(n1396) );
  IV U285 ( .A(n1416), .Z(n85) );
  NOR U286 ( .A(g_input[0]), .B(n1468), .Z(n1459) );
  XOR U287 ( .A(n1326), .B(n1313), .Z(n1134) );
  MUX U288 ( .IN0(n1145), .IN1(n86), .SEL(n935), .F(n873) );
  IV U289 ( .A(n933), .Z(n86) );
  MUX U290 ( .IN0(n433), .IN1(n431), .SEL(n432), .F(n382) );
  XOR U291 ( .A(n687), .B(n753), .Z(n688) );
  MUX U292 ( .IN0(n367), .IN1(n87), .SEL(n366), .F(n320) );
  IV U293 ( .A(n365), .Z(n87) );
  MUX U294 ( .IN0(e_input[7]), .IN1(n1132), .SEL(e_input[15]), .F(n509) );
  XNOR U295 ( .A(n741), .B(n678), .Z(n682) );
  XOR U296 ( .A(n732), .B(n667), .Z(n671) );
  XNOR U297 ( .A(n847), .B(n775), .Z(n779) );
  XNOR U298 ( .A(n901), .B(n900), .Z(n883) );
  MUX U299 ( .IN0(n257), .IN1(n283), .SEL(n256), .F(n228) );
  XNOR U300 ( .A(n339), .B(n338), .Z(n328) );
  XNOR U301 ( .A(n550), .B(n549), .Z(n528) );
  XNOR U302 ( .A(n615), .B(n614), .Z(n593) );
  XNOR U303 ( .A(n721), .B(n788), .Z(n722) );
  XNOR U304 ( .A(n464), .B(n463), .Z(n456) );
  XOR U305 ( .A(n570), .B(n511), .Z(n519) );
  XNOR U306 ( .A(n731), .B(n730), .Z(n720) );
  XNOR U307 ( .A(n808), .B(n807), .Z(n787) );
  XNOR U308 ( .A(n247), .B(n246), .Z(n271) );
  MUX U309 ( .IN0(n88), .IN1(n440), .SEL(n441), .F(n391) );
  IV U310 ( .A(\_MxM/Y0[7] ), .Z(n88) );
  MUX U311 ( .IN0(\_MxM/Y0[14] ), .IN1(n179), .SEL(n180), .F(n169) );
  XOR U312 ( .A(n690), .B(n698), .Z(n696) );
  MUX U313 ( .IN0(n1049), .IN1(n89), .SEL(n1050), .F(n1022) );
  IV U314 ( .A(n1051), .Z(n89) );
  MUX U315 ( .IN0(n90), .IN1(n1133), .SEL(n1134), .F(n1306) );
  IV U316 ( .A(n1320), .Z(n90) );
  MUX U317 ( .IN0(n1183), .IN1(n91), .SEL(n1004), .F(n1168) );
  IV U318 ( .A(n1002), .Z(n91) );
  XOR U319 ( .A(n1444), .B(g_input[3]), .Z(n1445) );
  MUX U320 ( .IN0(n949), .IN1(n92), .SEL(n950), .F(n915) );
  IV U321 ( .A(n951), .Z(n92) );
  XOR U322 ( .A(n1414), .B(n1415), .Z(n1346) );
  XOR U323 ( .A(n1265), .B(n1256), .Z(n1109) );
  MUX U324 ( .IN0(e_input[5]), .IN1(n1127), .SEL(e_input[15]), .F(n639) );
  MUX U325 ( .IN0(e_input[2]), .IN1(n1324), .SEL(e_input[15]), .F(n866) );
  XNOR U326 ( .A(n1105), .B(n1104), .Z(n922) );
  XNOR U327 ( .A(n329), .B(n293), .Z(n287) );
  MUX U328 ( .IN0(n373), .IN1(n371), .SEL(n372), .F(n93) );
  IV U329 ( .A(n93), .Z(n325) );
  XOR U330 ( .A(n647), .B(n648), .Z(n644) );
  XOR U331 ( .A(n884), .B(n812), .Z(n816) );
  MUX U332 ( .IN0(n875), .IN1(n1135), .SEL(n874), .F(n797) );
  XNOR U333 ( .A(n855), .B(n854), .Z(n872) );
  AND U334 ( .A(n217), .B(n194), .Z(n216) );
  XNOR U335 ( .A(n384), .B(n383), .Z(n370) );
  XNOR U336 ( .A(n433), .B(n432), .Z(n413) );
  XNOR U337 ( .A(n485), .B(n484), .Z(n464) );
  XNOR U338 ( .A(n707), .B(n706), .Z(n723) );
  XNOR U339 ( .A(n751), .B(n750), .Z(n731) );
  XNOR U340 ( .A(n828), .B(n827), .Z(n808) );
  XNOR U341 ( .A(n780), .B(n779), .Z(n800) );
  XNOR U342 ( .A(n883), .B(n882), .Z(n862) );
  XNOR U343 ( .A(n248), .B(n249), .Z(n247) );
  XNOR U344 ( .A(n528), .B(n527), .Z(n520) );
  XNOR U345 ( .A(n593), .B(n592), .Z(n585) );
  XNOR U346 ( .A(n661), .B(n660), .Z(n653) );
  MUX U347 ( .IN0(n94), .IN1(n301), .SEL(n302), .F(n264) );
  IV U348 ( .A(\_MxM/Y0[10] ), .Z(n94) );
  MUX U349 ( .IN0(n95), .IN1(n492), .SEL(n493), .F(n440) );
  IV U350 ( .A(\_MxM/Y0[6] ), .Z(n95) );
  MUX U351 ( .IN0(n96), .IN1(n758), .SEL(n759), .F(n690) );
  IV U352 ( .A(\_MxM/Y0[2] ), .Z(n96) );
  MUX U353 ( .IN0(\_MxM/Y0[15] ), .IN1(n169), .SEL(n170), .F(n97) );
  IV U354 ( .A(n97), .Z(n166) );
  XOR U355 ( .A(n836), .B(\_MxM/Y0[1] ), .Z(n111) );
  ANDN U356 ( .A(n98), .B(\_MxM/n[0] ), .Z(\_MxM/n244 ) );
  AND U357 ( .A(\_MxM/N8 ), .B(n98), .Z(\_MxM/n243 ) );
  AND U358 ( .A(\_MxM/N9 ), .B(n98), .Z(\_MxM/n242 ) );
  AND U359 ( .A(\_MxM/N10 ), .B(n98), .Z(\_MxM/n241 ) );
  AND U360 ( .A(\_MxM/N11 ), .B(n98), .Z(\_MxM/n240 ) );
  AND U361 ( .A(\_MxM/N12 ), .B(n98), .Z(\_MxM/n239 ) );
  AND U362 ( .A(\_MxM/N13 ), .B(n98), .Z(\_MxM/n238 ) );
  AND U363 ( .A(\_MxM/N14 ), .B(n98), .Z(\_MxM/n237 ) );
  AND U364 ( .A(\_MxM/N15 ), .B(n98), .Z(\_MxM/n236 ) );
  AND U365 ( .A(n98), .B(n99), .Z(\_MxM/n235 ) );
  XOR U366 ( .A(\_MxM/n[9] ), .B(\_MxM/add_39/carry[9] ), .Z(n99) );
  ANDN U367 ( .A(n100), .B(rst), .Z(n98) );
  NAND U368 ( .A(n101), .B(n102), .Z(n100) );
  AND U369 ( .A(n103), .B(n104), .Z(n102) );
  AND U370 ( .A(\_MxM/n[1] ), .B(n105), .Z(n104) );
  ANDN U371 ( .A(\_MxM/n[0] ), .B(n106), .Z(n105) );
  AND U372 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n103) );
  AND U373 ( .A(n107), .B(n108), .Z(n101) );
  AND U374 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n108) );
  AND U375 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n107) );
  NAND U376 ( .A(n109), .B(n110), .Z(\_MxM/n234 ) );
  OR U377 ( .A(n111), .B(n112), .Z(n110) );
  NANDN U378 ( .B(n113), .A(\_MxM/Y0[0] ), .Z(n109) );
  NAND U379 ( .A(n114), .B(n115), .Z(\_MxM/n233 ) );
  NANDN U380 ( .B(n112), .A(n116), .Z(n115) );
  NANDN U381 ( .B(n117), .A(rst), .Z(n114) );
  NAND U382 ( .A(n118), .B(n119), .Z(\_MxM/n232 ) );
  NANDN U383 ( .B(n112), .A(n120), .Z(n119) );
  NANDN U384 ( .B(n113), .A(\_MxM/Y0[2] ), .Z(n118) );
  NAND U385 ( .A(n121), .B(n122), .Z(\_MxM/n231 ) );
  NANDN U386 ( .B(n112), .A(n123), .Z(n122) );
  NANDN U387 ( .B(n113), .A(\_MxM/Y0[3] ), .Z(n121) );
  NAND U388 ( .A(n124), .B(n125), .Z(\_MxM/n230 ) );
  NANDN U389 ( .B(n112), .A(n126), .Z(n125) );
  NANDN U390 ( .B(n113), .A(\_MxM/Y0[4] ), .Z(n124) );
  NAND U391 ( .A(n127), .B(n128), .Z(\_MxM/n229 ) );
  NANDN U392 ( .B(n112), .A(n129), .Z(n128) );
  NANDN U393 ( .B(n113), .A(\_MxM/Y0[5] ), .Z(n127) );
  NAND U394 ( .A(n130), .B(n131), .Z(\_MxM/n228 ) );
  NANDN U395 ( .B(n112), .A(n132), .Z(n131) );
  NANDN U396 ( .B(n113), .A(\_MxM/Y0[6] ), .Z(n130) );
  NAND U397 ( .A(n133), .B(n134), .Z(\_MxM/n227 ) );
  NANDN U398 ( .B(n112), .A(n135), .Z(n134) );
  NANDN U399 ( .B(n113), .A(\_MxM/Y0[7] ), .Z(n133) );
  NAND U400 ( .A(n136), .B(n137), .Z(\_MxM/n226 ) );
  NANDN U401 ( .B(n112), .A(n138), .Z(n137) );
  NANDN U402 ( .B(n113), .A(\_MxM/Y0[8] ), .Z(n136) );
  NAND U403 ( .A(n139), .B(n140), .Z(\_MxM/n225 ) );
  NANDN U404 ( .B(n112), .A(n141), .Z(n140) );
  NANDN U405 ( .B(n113), .A(\_MxM/Y0[9] ), .Z(n139) );
  NAND U406 ( .A(n142), .B(n143), .Z(\_MxM/n224 ) );
  NANDN U407 ( .B(n112), .A(n144), .Z(n143) );
  NANDN U408 ( .B(n113), .A(\_MxM/Y0[10] ), .Z(n142) );
  NAND U409 ( .A(n145), .B(n146), .Z(\_MxM/n223 ) );
  NANDN U410 ( .B(n112), .A(n147), .Z(n146) );
  NANDN U411 ( .B(n113), .A(\_MxM/Y0[11] ), .Z(n145) );
  NAND U412 ( .A(n148), .B(n149), .Z(\_MxM/n222 ) );
  NANDN U413 ( .B(n112), .A(n150), .Z(n149) );
  NANDN U414 ( .B(n113), .A(\_MxM/Y0[12] ), .Z(n148) );
  NAND U415 ( .A(n151), .B(n152), .Z(\_MxM/n221 ) );
  NANDN U416 ( .B(n112), .A(n153), .Z(n152) );
  NANDN U417 ( .B(n113), .A(\_MxM/Y0[13] ), .Z(n151) );
  NAND U418 ( .A(n154), .B(n155), .Z(\_MxM/n220 ) );
  OR U419 ( .A(n156), .B(n112), .Z(n155) );
  NANDN U420 ( .B(n113), .A(\_MxM/Y0[14] ), .Z(n154) );
  NAND U421 ( .A(n157), .B(n158), .Z(\_MxM/n219 ) );
  OR U422 ( .A(n112), .B(n159), .Z(n158) );
  NANDN U423 ( .B(n160), .A(n113), .Z(n112) );
  NANDN U424 ( .B(n113), .A(\_MxM/Y0[15] ), .Z(n157) );
  NAND U425 ( .A(n161), .B(n162), .Z(\_MxM/n218 ) );
  NANDN U426 ( .B(n113), .A(o[15]), .Z(n162) );
  AND U427 ( .A(n163), .B(n164), .Z(n161) );
  NANDN U428 ( .B(n160), .A(o[15]), .Z(n164) );
  OR U429 ( .A(n159), .B(n165), .Z(n163) );
  XOR U430 ( .A(n166), .B(n167), .Z(n159) );
  XNOR U431 ( .A(\_MxM/Y0[15] ), .B(n168), .Z(n167) );
  NAND U432 ( .A(n171), .B(n172), .Z(\_MxM/n217 ) );
  NANDN U433 ( .B(n113), .A(o[14]), .Z(n172) );
  AND U434 ( .A(n173), .B(n174), .Z(n171) );
  NANDN U435 ( .B(n160), .A(o[14]), .Z(n174) );
  OR U436 ( .A(n156), .B(n165), .Z(n173) );
  XOR U437 ( .A(n170), .B(\_MxM/Y0[15] ), .Z(n156) );
  XOR U438 ( .A(n169), .B(n168), .Z(n170) );
  NAND U439 ( .A(n175), .B(n176), .Z(n168) );
  OR U440 ( .A(n177), .B(n178), .Z(n175) );
  NAND U441 ( .A(n181), .B(n182), .Z(\_MxM/n216 ) );
  NANDN U442 ( .B(n113), .A(o[13]), .Z(n182) );
  AND U443 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U444 ( .B(n160), .A(o[13]), .Z(n184) );
  NANDN U445 ( .B(n165), .A(n153), .Z(n183) );
  XNOR U446 ( .A(n180), .B(\_MxM/Y0[14] ), .Z(n153) );
  XNOR U447 ( .A(n185), .B(n179), .Z(n180) );
  XNOR U448 ( .A(n178), .B(n188), .Z(n177) );
  OR U449 ( .A(n189), .B(n190), .Z(n178) );
  AND U450 ( .A(n191), .B(n192), .Z(n188) );
  OR U451 ( .A(n193), .B(n194), .Z(n192) );
  AND U452 ( .A(n195), .B(n196), .Z(n191) );
  OR U453 ( .A(n197), .B(n198), .Z(n196) );
  OR U454 ( .A(n199), .B(n200), .Z(n195) );
  NAND U455 ( .A(n201), .B(n202), .Z(\_MxM/n215 ) );
  NANDN U456 ( .B(n113), .A(o[12]), .Z(n202) );
  AND U457 ( .A(n203), .B(n204), .Z(n201) );
  NANDN U458 ( .B(n160), .A(o[12]), .Z(n204) );
  NANDN U459 ( .B(n165), .A(n150), .Z(n203) );
  XNOR U460 ( .A(n187), .B(\_MxM/Y0[13] ), .Z(n150) );
  XNOR U461 ( .A(n205), .B(n206), .Z(n187) );
  AND U462 ( .A(n176), .B(n208), .Z(n207) );
  XOR U463 ( .A(n189), .B(n209), .Z(n208) );
  XOR U464 ( .A(n209), .B(n190), .Z(n189) );
  OR U465 ( .A(n210), .B(n211), .Z(n190) );
  IV U466 ( .A(n206), .Z(n209) );
  XNOR U467 ( .A(n200), .B(n199), .Z(n206) );
  OR U468 ( .A(n212), .B(n213), .Z(n199) );
  AND U469 ( .A(n214), .B(n215), .Z(n200) );
  XNOR U470 ( .A(n193), .B(n216), .Z(n215) );
  NAND U471 ( .A(n218), .B(n219), .Z(n194) );
  NANDN U472 ( .B(n220), .A(n221), .Z(n218) );
  NANDN U473 ( .B(n197), .A(n222), .Z(n217) );
  NANDN U474 ( .B(n198), .A(n223), .Z(n193) );
  AND U475 ( .A(n224), .B(n225), .Z(n214) );
  OR U476 ( .A(n226), .B(n227), .Z(n225) );
  XNOR U477 ( .A(n228), .B(n229), .Z(n224) );
  ANDN U478 ( .A(n230), .B(n231), .Z(n229) );
  XOR U479 ( .A(n228), .B(n232), .Z(n230) );
  NAND U480 ( .A(n235), .B(n236), .Z(\_MxM/n214 ) );
  NANDN U481 ( .B(n113), .A(o[11]), .Z(n236) );
  AND U482 ( .A(n237), .B(n238), .Z(n235) );
  NANDN U483 ( .B(n160), .A(o[11]), .Z(n238) );
  NANDN U484 ( .B(n165), .A(n147), .Z(n237) );
  XNOR U485 ( .A(n234), .B(\_MxM/Y0[12] ), .Z(n147) );
  XNOR U486 ( .A(n239), .B(n240), .Z(n234) );
  AND U487 ( .A(n176), .B(n242), .Z(n241) );
  XOR U488 ( .A(n210), .B(n243), .Z(n242) );
  XOR U489 ( .A(n243), .B(n211), .Z(n210) );
  OR U490 ( .A(n244), .B(n245), .Z(n211) );
  IV U491 ( .A(n240), .Z(n243) );
  XNOR U492 ( .A(n213), .B(n212), .Z(n240) );
  OR U493 ( .A(n246), .B(n247), .Z(n212) );
  XNOR U494 ( .A(n227), .B(n226), .Z(n213) );
  OR U495 ( .A(n248), .B(n249), .Z(n226) );
  XOR U496 ( .A(n232), .B(n231), .Z(n227) );
  XOR U497 ( .A(n228), .B(n250), .Z(n231) );
  AND U498 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U499 ( .B(n197), .A(n253), .Z(n252) );
  OR U500 ( .A(n254), .B(n255), .Z(n251) );
  XOR U501 ( .A(n220), .B(n221), .Z(n232) );
  NANDN U502 ( .B(n198), .A(n258), .Z(n221) );
  XNOR U503 ( .A(n219), .B(n259), .Z(n220) );
  AND U504 ( .A(n223), .B(n222), .Z(n259) );
  ANDN U505 ( .A(n260), .B(n261), .Z(n219) );
  NANDN U506 ( .B(n262), .A(n263), .Z(n260) );
  NAND U507 ( .A(n266), .B(n267), .Z(\_MxM/n213 ) );
  NANDN U508 ( .B(n113), .A(o[10]), .Z(n267) );
  AND U509 ( .A(n268), .B(n269), .Z(n266) );
  NANDN U510 ( .B(n160), .A(o[10]), .Z(n269) );
  NANDN U511 ( .B(n165), .A(n144), .Z(n268) );
  XNOR U512 ( .A(n265), .B(\_MxM/Y0[11] ), .Z(n144) );
  XNOR U513 ( .A(n270), .B(n271), .Z(n265) );
  AND U514 ( .A(n176), .B(n273), .Z(n272) );
  XOR U515 ( .A(n244), .B(n274), .Z(n273) );
  XOR U516 ( .A(n274), .B(n245), .Z(n244) );
  OR U517 ( .A(n275), .B(n276), .Z(n245) );
  IV U518 ( .A(n271), .Z(n274) );
  OR U519 ( .A(n277), .B(n278), .Z(n246) );
  XOR U520 ( .A(n257), .B(n256), .Z(n248) );
  XNOR U521 ( .A(n282), .B(n283), .Z(n256) );
  ANDN U522 ( .A(n286), .B(n287), .Z(n285) );
  XOR U523 ( .A(n284), .B(n288), .Z(n286) );
  XNOR U524 ( .A(n289), .B(n254), .Z(n282) );
  NAND U525 ( .A(n253), .B(n223), .Z(n254) );
  NANDN U526 ( .B(n197), .A(n291), .Z(n290) );
  XOR U527 ( .A(n262), .B(n263), .Z(n257) );
  NANDN U528 ( .B(n198), .A(n295), .Z(n263) );
  AND U529 ( .A(n258), .B(n222), .Z(n296) );
  NAND U530 ( .A(n297), .B(n298), .Z(n261) );
  NANDN U531 ( .B(n299), .A(n300), .Z(n297) );
  NAND U532 ( .A(n303), .B(n304), .Z(\_MxM/n212 ) );
  NANDN U533 ( .B(n113), .A(o[9]), .Z(n304) );
  AND U534 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U535 ( .B(n160), .A(o[9]), .Z(n306) );
  NANDN U536 ( .B(n165), .A(n141), .Z(n305) );
  XNOR U537 ( .A(n302), .B(\_MxM/Y0[10] ), .Z(n141) );
  XNOR U538 ( .A(n307), .B(n308), .Z(n302) );
  AND U539 ( .A(n176), .B(n310), .Z(n309) );
  XOR U540 ( .A(n275), .B(n311), .Z(n310) );
  XOR U541 ( .A(n311), .B(n276), .Z(n275) );
  OR U542 ( .A(n312), .B(n313), .Z(n276) );
  IV U543 ( .A(n308), .Z(n311) );
  XNOR U544 ( .A(n278), .B(n277), .Z(n308) );
  OR U545 ( .A(n314), .B(n315), .Z(n277) );
  XNOR U546 ( .A(n281), .B(n280), .Z(n278) );
  XOR U547 ( .A(n279), .B(n316), .Z(n280) );
  AND U548 ( .A(n317), .B(n318), .Z(n316) );
  OR U549 ( .A(n319), .B(n320), .Z(n318) );
  AND U550 ( .A(n321), .B(n322), .Z(n317) );
  NANDN U551 ( .B(n197), .A(n323), .Z(n322) );
  NAND U552 ( .A(n324), .B(n325), .Z(n321) );
  XNOR U553 ( .A(n292), .B(n330), .Z(n293) );
  AND U554 ( .A(n223), .B(n291), .Z(n330) );
  XOR U555 ( .A(n331), .B(n332), .Z(n292) );
  ANDN U556 ( .A(n333), .B(n334), .Z(n332) );
  XNOR U557 ( .A(n335), .B(n331), .Z(n333) );
  XOR U558 ( .A(n336), .B(n294), .Z(n329) );
  NAND U559 ( .A(n253), .B(n258), .Z(n294) );
  IV U560 ( .A(n284), .Z(n336) );
  XNOR U561 ( .A(n299), .B(n300), .Z(n288) );
  NANDN U562 ( .B(n198), .A(n340), .Z(n300) );
  XNOR U563 ( .A(n298), .B(n341), .Z(n299) );
  AND U564 ( .A(n295), .B(n222), .Z(n341) );
  ANDN U565 ( .A(n342), .B(n343), .Z(n298) );
  NANDN U566 ( .B(n344), .A(n345), .Z(n342) );
  NAND U567 ( .A(n348), .B(n349), .Z(\_MxM/n211 ) );
  NANDN U568 ( .B(n113), .A(o[8]), .Z(n349) );
  AND U569 ( .A(n350), .B(n351), .Z(n348) );
  NANDN U570 ( .B(n160), .A(o[8]), .Z(n351) );
  NANDN U571 ( .B(n165), .A(n138), .Z(n350) );
  XNOR U572 ( .A(n347), .B(\_MxM/Y0[9] ), .Z(n138) );
  XNOR U573 ( .A(n352), .B(n353), .Z(n347) );
  AND U574 ( .A(n176), .B(n355), .Z(n354) );
  XOR U575 ( .A(n312), .B(n356), .Z(n355) );
  XOR U576 ( .A(n356), .B(n313), .Z(n312) );
  OR U577 ( .A(n357), .B(n358), .Z(n313) );
  IV U578 ( .A(n353), .Z(n356) );
  XNOR U579 ( .A(n315), .B(n314), .Z(n353) );
  OR U580 ( .A(n359), .B(n360), .Z(n314) );
  XNOR U581 ( .A(n328), .B(n327), .Z(n315) );
  XOR U582 ( .A(n361), .B(n324), .Z(n327) );
  XNOR U583 ( .A(n362), .B(n319), .Z(n324) );
  NAND U584 ( .A(n323), .B(n223), .Z(n319) );
  NANDN U585 ( .B(n197), .A(n364), .Z(n363) );
  XNOR U586 ( .A(n325), .B(n326), .Z(n361) );
  XNOR U587 ( .A(n331), .B(n375), .Z(n334) );
  AND U588 ( .A(n258), .B(n291), .Z(n375) );
  XOR U589 ( .A(n376), .B(n377), .Z(n331) );
  ANDN U590 ( .A(n378), .B(n379), .Z(n377) );
  XNOR U591 ( .A(n380), .B(n376), .Z(n378) );
  XOR U592 ( .A(n381), .B(n335), .Z(n374) );
  NAND U593 ( .A(n253), .B(n295), .Z(n335) );
  IV U594 ( .A(n337), .Z(n381) );
  XNOR U595 ( .A(n344), .B(n345), .Z(n339) );
  NANDN U596 ( .B(n198), .A(n385), .Z(n345) );
  AND U597 ( .A(n340), .B(n222), .Z(n386) );
  NAND U598 ( .A(n387), .B(n388), .Z(n343) );
  NANDN U599 ( .B(n389), .A(n390), .Z(n387) );
  NAND U600 ( .A(n393), .B(n394), .Z(\_MxM/n210 ) );
  NANDN U601 ( .B(n113), .A(o[7]), .Z(n394) );
  AND U602 ( .A(n395), .B(n396), .Z(n393) );
  NANDN U603 ( .B(n160), .A(o[7]), .Z(n396) );
  NANDN U604 ( .B(n165), .A(n135), .Z(n395) );
  XNOR U605 ( .A(n392), .B(\_MxM/Y0[8] ), .Z(n135) );
  XNOR U606 ( .A(n397), .B(n398), .Z(n392) );
  AND U607 ( .A(n176), .B(n400), .Z(n399) );
  XOR U608 ( .A(n357), .B(n401), .Z(n400) );
  XOR U609 ( .A(n401), .B(n358), .Z(n357) );
  OR U610 ( .A(n402), .B(n403), .Z(n358) );
  IV U611 ( .A(n398), .Z(n401) );
  XNOR U612 ( .A(n360), .B(n359), .Z(n398) );
  NANDN U613 ( .B(n404), .A(n405), .Z(n359) );
  XNOR U614 ( .A(n370), .B(n369), .Z(n360) );
  XOR U615 ( .A(n406), .B(n373), .Z(n369) );
  XNOR U616 ( .A(n366), .B(n367), .Z(n373) );
  NAND U617 ( .A(n323), .B(n258), .Z(n367) );
  XNOR U618 ( .A(n365), .B(n407), .Z(n366) );
  AND U619 ( .A(n223), .B(n364), .Z(n407) );
  XNOR U620 ( .A(n372), .B(n368), .Z(n406) );
  AND U621 ( .A(n415), .B(n416), .Z(n414) );
  NANDN U622 ( .B(n197), .A(n417), .Z(n416) );
  OR U623 ( .A(n418), .B(n419), .Z(n415) );
  XNOR U624 ( .A(n376), .B(n424), .Z(n379) );
  AND U625 ( .A(n295), .B(n291), .Z(n424) );
  XOR U626 ( .A(n425), .B(n426), .Z(n376) );
  ANDN U627 ( .A(n427), .B(n428), .Z(n426) );
  XNOR U628 ( .A(n429), .B(n425), .Z(n427) );
  XOR U629 ( .A(n430), .B(n380), .Z(n423) );
  NAND U630 ( .A(n253), .B(n340), .Z(n380) );
  IV U631 ( .A(n382), .Z(n430) );
  XNOR U632 ( .A(n389), .B(n390), .Z(n384) );
  NANDN U633 ( .B(n198), .A(n434), .Z(n390) );
  XNOR U634 ( .A(n388), .B(n435), .Z(n389) );
  AND U635 ( .A(n385), .B(n222), .Z(n435) );
  ANDN U636 ( .A(n436), .B(n437), .Z(n388) );
  NANDN U637 ( .B(n438), .A(n439), .Z(n436) );
  NAND U638 ( .A(n442), .B(n443), .Z(\_MxM/n209 ) );
  NANDN U639 ( .B(n113), .A(o[6]), .Z(n443) );
  AND U640 ( .A(n444), .B(n445), .Z(n442) );
  NANDN U641 ( .B(n160), .A(o[6]), .Z(n445) );
  NANDN U642 ( .B(n165), .A(n132), .Z(n444) );
  XNOR U643 ( .A(n441), .B(\_MxM/Y0[7] ), .Z(n132) );
  XNOR U644 ( .A(n447), .B(n448), .Z(n446) );
  AND U645 ( .A(n176), .B(n449), .Z(n448) );
  XOR U646 ( .A(n402), .B(n452), .Z(n449) );
  XOR U647 ( .A(n452), .B(n403), .Z(n402) );
  OR U648 ( .A(n450), .B(n451), .Z(n403) );
  XNOR U649 ( .A(n404), .B(n405), .Z(n452) );
  XNOR U650 ( .A(n413), .B(n412), .Z(n404) );
  XOR U651 ( .A(n457), .B(n422), .Z(n412) );
  XNOR U652 ( .A(n409), .B(n410), .Z(n422) );
  NAND U653 ( .A(n323), .B(n295), .Z(n410) );
  XNOR U654 ( .A(n408), .B(n458), .Z(n409) );
  AND U655 ( .A(n258), .B(n364), .Z(n458) );
  XNOR U656 ( .A(n421), .B(n411), .Z(n457) );
  XNOR U657 ( .A(n465), .B(n420), .Z(n421) );
  XNOR U658 ( .A(n469), .B(n418), .Z(n465) );
  NAND U659 ( .A(n417), .B(n223), .Z(n418) );
  NANDN U660 ( .B(n197), .A(n471), .Z(n470) );
  XNOR U661 ( .A(n425), .B(n476), .Z(n428) );
  AND U662 ( .A(n340), .B(n291), .Z(n476) );
  XOR U663 ( .A(n477), .B(n478), .Z(n425) );
  ANDN U664 ( .A(n479), .B(n480), .Z(n478) );
  XNOR U665 ( .A(n481), .B(n477), .Z(n479) );
  XOR U666 ( .A(n482), .B(n429), .Z(n475) );
  NAND U667 ( .A(n253), .B(n385), .Z(n429) );
  IV U668 ( .A(n431), .Z(n482) );
  XNOR U669 ( .A(n438), .B(n439), .Z(n433) );
  NANDN U670 ( .B(n198), .A(n486), .Z(n439) );
  AND U671 ( .A(n434), .B(n222), .Z(n487) );
  NAND U672 ( .A(n488), .B(n489), .Z(n437) );
  NANDN U673 ( .B(n490), .A(n491), .Z(n488) );
  IV U674 ( .A(n440), .Z(n447) );
  NAND U675 ( .A(n494), .B(n495), .Z(\_MxM/n208 ) );
  NANDN U676 ( .B(n113), .A(o[5]), .Z(n495) );
  AND U677 ( .A(n496), .B(n497), .Z(n494) );
  NANDN U678 ( .B(n160), .A(o[5]), .Z(n497) );
  NANDN U679 ( .B(n165), .A(n129), .Z(n496) );
  XNOR U680 ( .A(n493), .B(\_MxM/Y0[6] ), .Z(n129) );
  XNOR U681 ( .A(n498), .B(n499), .Z(n493) );
  AND U682 ( .A(n176), .B(n501), .Z(n500) );
  XOR U683 ( .A(n450), .B(n502), .Z(n501) );
  XOR U684 ( .A(n502), .B(n451), .Z(n450) );
  OR U685 ( .A(n503), .B(n504), .Z(n451) );
  IV U686 ( .A(n499), .Z(n502) );
  XOR U687 ( .A(n456), .B(n455), .Z(n499) );
  XNOR U688 ( .A(n454), .B(n505), .Z(n455) );
  AND U689 ( .A(n453), .B(n506), .Z(n505) );
  AND U690 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U691 ( .B(n197), .A(n509), .Z(n508) );
  OR U692 ( .A(n510), .B(n511), .Z(n507) );
  AND U693 ( .A(n512), .B(n513), .Z(n453) );
  NANDN U694 ( .B(n514), .A(n515), .Z(n513) );
  NANDN U695 ( .B(n516), .A(n517), .Z(n512) );
  XNOR U696 ( .A(n521), .B(n468), .Z(n463) );
  XNOR U697 ( .A(n460), .B(n461), .Z(n468) );
  NAND U698 ( .A(n323), .B(n340), .Z(n461) );
  XNOR U699 ( .A(n459), .B(n522), .Z(n460) );
  AND U700 ( .A(n295), .B(n364), .Z(n522) );
  XNOR U701 ( .A(n467), .B(n462), .Z(n521) );
  XNOR U702 ( .A(n472), .B(n530), .Z(n473) );
  AND U703 ( .A(n223), .B(n471), .Z(n530) );
  XOR U704 ( .A(n531), .B(n532), .Z(n472) );
  ANDN U705 ( .A(n533), .B(n534), .Z(n532) );
  XNOR U706 ( .A(n535), .B(n531), .Z(n533) );
  XOR U707 ( .A(n536), .B(n474), .Z(n529) );
  NAND U708 ( .A(n417), .B(n258), .Z(n474) );
  IV U709 ( .A(n466), .Z(n536) );
  XNOR U710 ( .A(n477), .B(n541), .Z(n480) );
  AND U711 ( .A(n385), .B(n291), .Z(n541) );
  XOR U712 ( .A(n542), .B(n543), .Z(n477) );
  ANDN U713 ( .A(n544), .B(n545), .Z(n543) );
  XNOR U714 ( .A(n546), .B(n542), .Z(n544) );
  XOR U715 ( .A(n547), .B(n481), .Z(n540) );
  NAND U716 ( .A(n253), .B(n434), .Z(n481) );
  IV U717 ( .A(n483), .Z(n547) );
  XNOR U718 ( .A(n490), .B(n491), .Z(n485) );
  NANDN U719 ( .B(n198), .A(n551), .Z(n491) );
  XNOR U720 ( .A(n489), .B(n552), .Z(n490) );
  AND U721 ( .A(n486), .B(n222), .Z(n552) );
  ANDN U722 ( .A(n553), .B(n554), .Z(n489) );
  NANDN U723 ( .B(n555), .A(n556), .Z(n553) );
  NAND U724 ( .A(n559), .B(n560), .Z(\_MxM/n207 ) );
  NANDN U725 ( .B(n113), .A(o[4]), .Z(n560) );
  AND U726 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U727 ( .B(n160), .A(o[4]), .Z(n562) );
  NANDN U728 ( .B(n165), .A(n126), .Z(n561) );
  XNOR U729 ( .A(n558), .B(\_MxM/Y0[5] ), .Z(n126) );
  XNOR U730 ( .A(n563), .B(n564), .Z(n558) );
  AND U731 ( .A(n176), .B(n566), .Z(n565) );
  XOR U732 ( .A(n503), .B(n567), .Z(n566) );
  XOR U733 ( .A(n567), .B(n504), .Z(n503) );
  OR U734 ( .A(n568), .B(n569), .Z(n504) );
  IV U735 ( .A(n564), .Z(n567) );
  XOR U736 ( .A(n520), .B(n519), .Z(n564) );
  XOR U737 ( .A(n514), .B(n515), .Z(n511) );
  XOR U738 ( .A(n574), .B(n516), .Z(n514) );
  NAND U739 ( .A(n223), .B(n509), .Z(n516) );
  NANDN U740 ( .B(n517), .A(n575), .Z(n574) );
  NANDN U741 ( .B(n197), .A(n576), .Z(n575) );
  XOR U742 ( .A(n580), .B(n510), .Z(n570) );
  OR U743 ( .A(n581), .B(n582), .Z(n510) );
  IV U744 ( .A(n518), .Z(n580) );
  XNOR U745 ( .A(n586), .B(n539), .Z(n527) );
  XNOR U746 ( .A(n524), .B(n525), .Z(n539) );
  NAND U747 ( .A(n323), .B(n385), .Z(n525) );
  XNOR U748 ( .A(n523), .B(n587), .Z(n524) );
  AND U749 ( .A(n340), .B(n364), .Z(n587) );
  XNOR U750 ( .A(n538), .B(n526), .Z(n586) );
  XNOR U751 ( .A(n531), .B(n595), .Z(n534) );
  AND U752 ( .A(n258), .B(n471), .Z(n595) );
  XOR U753 ( .A(n596), .B(n597), .Z(n531) );
  ANDN U754 ( .A(n598), .B(n599), .Z(n597) );
  XNOR U755 ( .A(n600), .B(n596), .Z(n598) );
  XOR U756 ( .A(n601), .B(n535), .Z(n594) );
  NAND U757 ( .A(n417), .B(n295), .Z(n535) );
  IV U758 ( .A(n537), .Z(n601) );
  XNOR U759 ( .A(n542), .B(n606), .Z(n545) );
  AND U760 ( .A(n434), .B(n291), .Z(n606) );
  XOR U761 ( .A(n607), .B(n608), .Z(n542) );
  ANDN U762 ( .A(n609), .B(n610), .Z(n608) );
  XNOR U763 ( .A(n611), .B(n607), .Z(n609) );
  XOR U764 ( .A(n612), .B(n546), .Z(n605) );
  NAND U765 ( .A(n253), .B(n486), .Z(n546) );
  IV U766 ( .A(n548), .Z(n612) );
  XNOR U767 ( .A(n555), .B(n556), .Z(n550) );
  NANDN U768 ( .B(n198), .A(n616), .Z(n556) );
  AND U769 ( .A(n551), .B(n222), .Z(n617) );
  NAND U770 ( .A(n618), .B(n619), .Z(n554) );
  NANDN U771 ( .B(n620), .A(n621), .Z(n618) );
  NAND U772 ( .A(n624), .B(n625), .Z(\_MxM/n206 ) );
  NANDN U773 ( .B(n113), .A(o[3]), .Z(n625) );
  AND U774 ( .A(n626), .B(n627), .Z(n624) );
  NANDN U775 ( .B(n160), .A(o[3]), .Z(n627) );
  NANDN U776 ( .B(n165), .A(n123), .Z(n626) );
  XNOR U777 ( .A(n623), .B(\_MxM/Y0[4] ), .Z(n123) );
  XNOR U778 ( .A(n628), .B(n629), .Z(n623) );
  AND U779 ( .A(n176), .B(n631), .Z(n630) );
  XOR U780 ( .A(n568), .B(n632), .Z(n631) );
  XOR U781 ( .A(n632), .B(n569), .Z(n568) );
  OR U782 ( .A(n633), .B(n634), .Z(n569) );
  IV U783 ( .A(n629), .Z(n632) );
  XOR U784 ( .A(n585), .B(n584), .Z(n629) );
  XOR U785 ( .A(n635), .B(n581), .Z(n584) );
  XOR U786 ( .A(n573), .B(n572), .Z(n581) );
  XOR U787 ( .A(n571), .B(n636), .Z(n572) );
  AND U788 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U789 ( .B(n197), .A(n639), .Z(n638) );
  OR U790 ( .A(n640), .B(n641), .Z(n637) );
  NAND U791 ( .A(n258), .B(n509), .Z(n579) );
  XNOR U792 ( .A(n577), .B(n645), .Z(n578) );
  AND U793 ( .A(n576), .B(n223), .Z(n645) );
  NANDN U794 ( .B(n649), .A(n650), .Z(n582) );
  XNOR U795 ( .A(n654), .B(n604), .Z(n592) );
  XNOR U796 ( .A(n589), .B(n590), .Z(n604) );
  NAND U797 ( .A(n323), .B(n434), .Z(n590) );
  XNOR U798 ( .A(n588), .B(n655), .Z(n589) );
  AND U799 ( .A(n385), .B(n364), .Z(n655) );
  XNOR U800 ( .A(n603), .B(n591), .Z(n654) );
  XNOR U801 ( .A(n596), .B(n663), .Z(n599) );
  AND U802 ( .A(n295), .B(n471), .Z(n663) );
  XOR U803 ( .A(n664), .B(n665), .Z(n596) );
  ANDN U804 ( .A(n666), .B(n667), .Z(n665) );
  XNOR U805 ( .A(n668), .B(n664), .Z(n666) );
  XOR U806 ( .A(n669), .B(n600), .Z(n662) );
  NAND U807 ( .A(n417), .B(n340), .Z(n600) );
  IV U808 ( .A(n602), .Z(n669) );
  XNOR U809 ( .A(n607), .B(n674), .Z(n610) );
  AND U810 ( .A(n486), .B(n291), .Z(n674) );
  XOR U811 ( .A(n675), .B(n676), .Z(n607) );
  ANDN U812 ( .A(n677), .B(n678), .Z(n676) );
  XNOR U813 ( .A(n679), .B(n675), .Z(n677) );
  XOR U814 ( .A(n680), .B(n611), .Z(n673) );
  NAND U815 ( .A(n253), .B(n551), .Z(n611) );
  IV U816 ( .A(n613), .Z(n680) );
  XNOR U817 ( .A(n620), .B(n621), .Z(n615) );
  NANDN U818 ( .B(n198), .A(n684), .Z(n621) );
  XNOR U819 ( .A(n619), .B(n685), .Z(n620) );
  AND U820 ( .A(n616), .B(n222), .Z(n685) );
  ANDN U821 ( .A(n686), .B(n687), .Z(n619) );
  NANDN U822 ( .B(n688), .A(n689), .Z(n686) );
  NAND U823 ( .A(n692), .B(n693), .Z(\_MxM/n205 ) );
  NANDN U824 ( .B(n113), .A(o[2]), .Z(n693) );
  AND U825 ( .A(n694), .B(n695), .Z(n692) );
  NANDN U826 ( .B(n160), .A(o[2]), .Z(n695) );
  NANDN U827 ( .B(n165), .A(n120), .Z(n694) );
  XNOR U828 ( .A(n691), .B(\_MxM/Y0[3] ), .Z(n120) );
  XNOR U829 ( .A(n696), .B(n697), .Z(n691) );
  AND U830 ( .A(n176), .B(n699), .Z(n698) );
  XOR U831 ( .A(n633), .B(n700), .Z(n699) );
  XOR U832 ( .A(n700), .B(n634), .Z(n633) );
  OR U833 ( .A(n701), .B(n702), .Z(n634) );
  IV U834 ( .A(n697), .Z(n700) );
  XOR U835 ( .A(n653), .B(n652), .Z(n697) );
  XOR U836 ( .A(n703), .B(n649), .Z(n652) );
  XOR U837 ( .A(n644), .B(n643), .Z(n649) );
  XNOR U838 ( .A(n708), .B(n640), .Z(n704) );
  NAND U839 ( .A(n223), .B(n639), .Z(n640) );
  NANDN U840 ( .B(n197), .A(n710), .Z(n709) );
  NAND U841 ( .A(n295), .B(n509), .Z(n648) );
  XNOR U842 ( .A(n646), .B(n714), .Z(n647) );
  AND U843 ( .A(n576), .B(n258), .Z(n714) );
  XNOR U844 ( .A(n650), .B(n651), .Z(n703) );
  XNOR U845 ( .A(n724), .B(n672), .Z(n660) );
  XNOR U846 ( .A(n657), .B(n658), .Z(n672) );
  NAND U847 ( .A(n323), .B(n486), .Z(n658) );
  XNOR U848 ( .A(n656), .B(n725), .Z(n657) );
  AND U849 ( .A(n434), .B(n364), .Z(n725) );
  XNOR U850 ( .A(n671), .B(n659), .Z(n724) );
  XNOR U851 ( .A(n664), .B(n733), .Z(n667) );
  AND U852 ( .A(n340), .B(n471), .Z(n733) );
  XOR U853 ( .A(n737), .B(n668), .Z(n732) );
  NAND U854 ( .A(n417), .B(n385), .Z(n668) );
  IV U855 ( .A(n670), .Z(n737) );
  XNOR U856 ( .A(n675), .B(n742), .Z(n678) );
  AND U857 ( .A(n551), .B(n291), .Z(n742) );
  XOR U858 ( .A(n743), .B(n744), .Z(n675) );
  ANDN U859 ( .A(n745), .B(n746), .Z(n744) );
  XNOR U860 ( .A(n747), .B(n743), .Z(n745) );
  XOR U861 ( .A(n748), .B(n679), .Z(n741) );
  NAND U862 ( .A(n253), .B(n616), .Z(n679) );
  IV U863 ( .A(n681), .Z(n748) );
  XNOR U864 ( .A(n688), .B(n689), .Z(n683) );
  OR U865 ( .A(n752), .B(n198), .Z(n689) );
  AND U866 ( .A(n684), .B(n222), .Z(n753) );
  NAND U867 ( .A(n754), .B(n755), .Z(n687) );
  NANDN U868 ( .B(n756), .A(n757), .Z(n754) );
  NAND U869 ( .A(n760), .B(n761), .Z(\_MxM/n204 ) );
  NANDN U870 ( .B(n113), .A(o[1]), .Z(n761) );
  AND U871 ( .A(n762), .B(n763), .Z(n760) );
  NANDN U872 ( .B(n160), .A(o[1]), .Z(n763) );
  NANDN U873 ( .B(n165), .A(n116), .Z(n762) );
  XNOR U874 ( .A(n759), .B(\_MxM/Y0[2] ), .Z(n116) );
  XNOR U875 ( .A(n764), .B(n765), .Z(n759) );
  XOR U876 ( .A(n758), .B(n766), .Z(n764) );
  AND U877 ( .A(n176), .B(n767), .Z(n766) );
  XOR U878 ( .A(n701), .B(n768), .Z(n767) );
  XOR U879 ( .A(n768), .B(n702), .Z(n701) );
  NANDN U880 ( .B(n769), .A(n770), .Z(n702) );
  IV U881 ( .A(n765), .Z(n768) );
  XOR U882 ( .A(n720), .B(n719), .Z(n765) );
  XNOR U883 ( .A(n771), .B(n723), .Z(n719) );
  XNOR U884 ( .A(n711), .B(n773), .Z(n712) );
  AND U885 ( .A(n710), .B(n223), .Z(n773) );
  XOR U886 ( .A(n777), .B(n713), .Z(n772) );
  NAND U887 ( .A(n258), .B(n639), .Z(n713) );
  IV U888 ( .A(n705), .Z(n777) );
  XNOR U889 ( .A(n716), .B(n717), .Z(n707) );
  NAND U890 ( .A(n340), .B(n509), .Z(n717) );
  XNOR U891 ( .A(n715), .B(n781), .Z(n716) );
  AND U892 ( .A(n576), .B(n295), .Z(n781) );
  XNOR U893 ( .A(n722), .B(n718), .Z(n771) );
  AND U894 ( .A(n789), .B(n790), .Z(n788) );
  OR U895 ( .A(n791), .B(n792), .Z(n790) );
  AND U896 ( .A(n793), .B(n794), .Z(n789) );
  NANDN U897 ( .B(n197), .A(n795), .Z(n794) );
  NANDN U898 ( .B(n796), .A(n797), .Z(n793) );
  XNOR U899 ( .A(n801), .B(n740), .Z(n730) );
  XNOR U900 ( .A(n727), .B(n728), .Z(n740) );
  NAND U901 ( .A(n323), .B(n551), .Z(n728) );
  XNOR U902 ( .A(n726), .B(n802), .Z(n727) );
  AND U903 ( .A(n486), .B(n364), .Z(n802) );
  XNOR U904 ( .A(n739), .B(n729), .Z(n801) );
  XNOR U905 ( .A(n734), .B(n810), .Z(n735) );
  AND U906 ( .A(n385), .B(n471), .Z(n810) );
  XOR U907 ( .A(n814), .B(n736), .Z(n809) );
  NAND U908 ( .A(n417), .B(n434), .Z(n736) );
  IV U909 ( .A(n738), .Z(n814) );
  XNOR U910 ( .A(n743), .B(n819), .Z(n746) );
  AND U911 ( .A(n616), .B(n291), .Z(n819) );
  XOR U912 ( .A(n820), .B(n821), .Z(n743) );
  ANDN U913 ( .A(n822), .B(n823), .Z(n821) );
  XNOR U914 ( .A(n824), .B(n820), .Z(n822) );
  XOR U915 ( .A(n825), .B(n747), .Z(n818) );
  NAND U916 ( .A(n253), .B(n684), .Z(n747) );
  IV U917 ( .A(n749), .Z(n825) );
  XNOR U918 ( .A(n756), .B(n757), .Z(n751) );
  OR U919 ( .A(n829), .B(n198), .Z(n757) );
  XNOR U920 ( .A(n755), .B(n830), .Z(n756) );
  ANDN U921 ( .A(n222), .B(n752), .Z(n830) );
  ANDN U922 ( .A(n831), .B(n832), .Z(n755) );
  NANDN U923 ( .B(n833), .A(n834), .Z(n831) );
  NAND U924 ( .A(n837), .B(n838), .Z(\_MxM/n203 ) );
  NANDN U925 ( .B(n113), .A(o[0]), .Z(n838) );
  AND U926 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U927 ( .B(n160), .A(o[0]), .Z(n840) );
  IV U928 ( .A(n841), .Z(n160) );
  OR U929 ( .A(n165), .B(n111), .Z(n839) );
  IV U930 ( .A(\_MxM/Y0[1] ), .Z(n117) );
  XOR U931 ( .A(n842), .B(n843), .Z(n836) );
  XNOR U932 ( .A(n844), .B(n835), .Z(n842) );
  NAND U933 ( .A(\_MxM/Y0[0] ), .B(n769), .Z(n835) );
  NAND U934 ( .A(n845), .B(n176), .Z(n844) );
  XOR U935 ( .A(e_input[15]), .B(g_input[15]), .Z(n176) );
  XNOR U936 ( .A(n770), .B(n843), .Z(n845) );
  XNOR U937 ( .A(n769), .B(n843), .Z(n770) );
  XNOR U938 ( .A(n787), .B(n786), .Z(n843) );
  XNOR U939 ( .A(n846), .B(n800), .Z(n786) );
  XNOR U940 ( .A(n774), .B(n848), .Z(n775) );
  AND U941 ( .A(n710), .B(n258), .Z(n848) );
  XOR U942 ( .A(n852), .B(n776), .Z(n847) );
  NAND U943 ( .A(n295), .B(n639), .Z(n776) );
  IV U944 ( .A(n778), .Z(n852) );
  XNOR U945 ( .A(n783), .B(n784), .Z(n780) );
  NAND U946 ( .A(n385), .B(n509), .Z(n784) );
  XNOR U947 ( .A(n782), .B(n856), .Z(n783) );
  AND U948 ( .A(n576), .B(n340), .Z(n856) );
  XNOR U949 ( .A(n799), .B(n785), .Z(n846) );
  XNOR U950 ( .A(n863), .B(n796), .Z(n799) );
  XOR U951 ( .A(n864), .B(n791), .Z(n796) );
  NAND U952 ( .A(n223), .B(n795), .Z(n791) );
  NANDN U953 ( .B(n197), .A(n866), .Z(n865) );
  XNOR U954 ( .A(n797), .B(n798), .Z(n863) );
  XNOR U955 ( .A(n876), .B(n817), .Z(n807) );
  XNOR U956 ( .A(n804), .B(n805), .Z(n817) );
  NAND U957 ( .A(n323), .B(n616), .Z(n805) );
  XNOR U958 ( .A(n803), .B(n877), .Z(n804) );
  AND U959 ( .A(n551), .B(n364), .Z(n877) );
  XNOR U960 ( .A(n816), .B(n806), .Z(n876) );
  XNOR U961 ( .A(n811), .B(n885), .Z(n812) );
  AND U962 ( .A(n434), .B(n471), .Z(n885) );
  XOR U963 ( .A(n889), .B(n813), .Z(n884) );
  NAND U964 ( .A(n417), .B(n486), .Z(n813) );
  IV U965 ( .A(n815), .Z(n889) );
  XNOR U966 ( .A(n820), .B(n894), .Z(n823) );
  AND U967 ( .A(n684), .B(n291), .Z(n894) );
  XOR U968 ( .A(n898), .B(n824), .Z(n893) );
  NANDN U969 ( .B(n752), .A(n253), .Z(n824) );
  IV U970 ( .A(n826), .Z(n898) );
  XNOR U971 ( .A(n833), .B(n834), .Z(n828) );
  NANDN U972 ( .B(n198), .A(n902), .Z(n834) );
  ANDN U973 ( .A(n222), .B(n829), .Z(n903) );
  NAND U974 ( .A(n904), .B(n905), .Z(n832) );
  NANDN U975 ( .B(n906), .A(n907), .Z(n904) );
  XNOR U976 ( .A(n862), .B(n861), .Z(n769) );
  XNOR U977 ( .A(n908), .B(n872), .Z(n861) );
  XNOR U978 ( .A(n849), .B(n910), .Z(n850) );
  AND U979 ( .A(n710), .B(n295), .Z(n910) );
  XOR U980 ( .A(n914), .B(n851), .Z(n909) );
  NAND U981 ( .A(n340), .B(n639), .Z(n851) );
  IV U982 ( .A(n853), .Z(n914) );
  XNOR U983 ( .A(n858), .B(n859), .Z(n855) );
  NAND U984 ( .A(n434), .B(n509), .Z(n859) );
  XNOR U985 ( .A(n857), .B(n918), .Z(n858) );
  AND U986 ( .A(n576), .B(n385), .Z(n918) );
  XNOR U987 ( .A(n871), .B(n860), .Z(n908) );
  XOR U988 ( .A(n922), .B(n923), .Z(n860) );
  XNOR U989 ( .A(n924), .B(n875), .Z(n871) );
  NAND U990 ( .A(n258), .B(n795), .Z(n869) );
  XNOR U991 ( .A(n867), .B(n925), .Z(n868) );
  AND U992 ( .A(n866), .B(n223), .Z(n925) );
  XNOR U993 ( .A(n874), .B(n870), .Z(n924) );
  XOR U994 ( .A(n929), .B(n930), .Z(n870) );
  AND U995 ( .A(n931), .B(n932), .Z(n930) );
  XOR U996 ( .A(n933), .B(n934), .Z(n932) );
  XOR U997 ( .A(n929), .B(n935), .Z(n934) );
  XOR U998 ( .A(n916), .B(n936), .Z(n931) );
  XOR U999 ( .A(n929), .B(n917), .Z(n936) );
  NAND U1000 ( .A(n509), .B(n486), .Z(n921) );
  XNOR U1001 ( .A(n919), .B(n937), .Z(n920) );
  AND U1002 ( .A(n576), .B(n434), .Z(n937) );
  XNOR U1003 ( .A(n911), .B(n942), .Z(n912) );
  AND U1004 ( .A(n710), .B(n340), .Z(n942) );
  XOR U1005 ( .A(n943), .B(n944), .Z(n911) );
  ANDN U1006 ( .A(n945), .B(n946), .Z(n944) );
  XNOR U1007 ( .A(n947), .B(n943), .Z(n945) );
  XOR U1008 ( .A(n948), .B(n913), .Z(n941) );
  NAND U1009 ( .A(n385), .B(n639), .Z(n913) );
  IV U1010 ( .A(n915), .Z(n948) );
  XOR U1011 ( .A(n952), .B(n953), .Z(n929) );
  AND U1012 ( .A(n954), .B(n955), .Z(n953) );
  XOR U1013 ( .A(n956), .B(n957), .Z(n955) );
  XOR U1014 ( .A(n952), .B(n958), .Z(n957) );
  XOR U1015 ( .A(n950), .B(n959), .Z(n954) );
  XOR U1016 ( .A(n952), .B(n951), .Z(n959) );
  NAND U1017 ( .A(n509), .B(n551), .Z(n940) );
  XNOR U1018 ( .A(n938), .B(n960), .Z(n939) );
  AND U1019 ( .A(n486), .B(n576), .Z(n960) );
  XNOR U1020 ( .A(n943), .B(n965), .Z(n946) );
  AND U1021 ( .A(n710), .B(n385), .Z(n965) );
  XOR U1022 ( .A(n966), .B(n967), .Z(n943) );
  ANDN U1023 ( .A(n968), .B(n969), .Z(n967) );
  XNOR U1024 ( .A(n970), .B(n966), .Z(n968) );
  XOR U1025 ( .A(n971), .B(n947), .Z(n964) );
  NAND U1026 ( .A(n434), .B(n639), .Z(n947) );
  IV U1027 ( .A(n949), .Z(n971) );
  XOR U1028 ( .A(n975), .B(n976), .Z(n952) );
  AND U1029 ( .A(n977), .B(n978), .Z(n976) );
  XOR U1030 ( .A(n979), .B(n980), .Z(n978) );
  XOR U1031 ( .A(n975), .B(n981), .Z(n980) );
  XOR U1032 ( .A(n973), .B(n982), .Z(n977) );
  XOR U1033 ( .A(n975), .B(n974), .Z(n982) );
  NAND U1034 ( .A(n509), .B(n616), .Z(n963) );
  XNOR U1035 ( .A(n961), .B(n983), .Z(n962) );
  AND U1036 ( .A(n551), .B(n576), .Z(n983) );
  XNOR U1037 ( .A(n966), .B(n988), .Z(n969) );
  AND U1038 ( .A(n710), .B(n434), .Z(n988) );
  XOR U1039 ( .A(n989), .B(n990), .Z(n966) );
  ANDN U1040 ( .A(n991), .B(n992), .Z(n990) );
  XNOR U1041 ( .A(n993), .B(n989), .Z(n991) );
  XOR U1042 ( .A(n994), .B(n970), .Z(n987) );
  NAND U1043 ( .A(n639), .B(n486), .Z(n970) );
  IV U1044 ( .A(n972), .Z(n994) );
  XOR U1045 ( .A(n998), .B(n999), .Z(n975) );
  AND U1046 ( .A(n1000), .B(n1001), .Z(n999) );
  XOR U1047 ( .A(n1002), .B(n1003), .Z(n1001) );
  XOR U1048 ( .A(n998), .B(n1004), .Z(n1003) );
  XOR U1049 ( .A(n996), .B(n1005), .Z(n1000) );
  XOR U1050 ( .A(n998), .B(n997), .Z(n1005) );
  XNOR U1051 ( .A(n1006), .B(n986), .Z(n997) );
  NAND U1052 ( .A(n509), .B(n684), .Z(n986) );
  IV U1053 ( .A(n985), .Z(n1006) );
  XNOR U1054 ( .A(n984), .B(n1007), .Z(n985) );
  AND U1055 ( .A(n616), .B(n576), .Z(n1007) );
  XOR U1056 ( .A(n1008), .B(n1009), .Z(n984) );
  ANDN U1057 ( .A(n1010), .B(n1011), .Z(n1009) );
  XNOR U1058 ( .A(n1012), .B(n1008), .Z(n1010) );
  XNOR U1059 ( .A(n1013), .B(n1014), .Z(n996) );
  IV U1060 ( .A(n992), .Z(n1014) );
  XNOR U1061 ( .A(n989), .B(n1015), .Z(n992) );
  AND U1062 ( .A(n486), .B(n710), .Z(n1015) );
  XOR U1063 ( .A(n1016), .B(n1017), .Z(n989) );
  ANDN U1064 ( .A(n1018), .B(n1019), .Z(n1017) );
  XNOR U1065 ( .A(n1020), .B(n1016), .Z(n1018) );
  XOR U1066 ( .A(n1021), .B(n993), .Z(n1013) );
  NAND U1067 ( .A(n639), .B(n551), .Z(n993) );
  IV U1068 ( .A(n995), .Z(n1021) );
  XOR U1069 ( .A(n1025), .B(n1026), .Z(n998) );
  AND U1070 ( .A(n1027), .B(n1028), .Z(n1026) );
  XOR U1071 ( .A(n1029), .B(n1030), .Z(n1028) );
  XOR U1072 ( .A(n1025), .B(n1031), .Z(n1030) );
  XOR U1073 ( .A(n1023), .B(n1032), .Z(n1027) );
  XOR U1074 ( .A(n1025), .B(n1024), .Z(n1032) );
  XNOR U1075 ( .A(n1033), .B(n1012), .Z(n1024) );
  NANDN U1076 ( .B(n752), .A(n509), .Z(n1012) );
  IV U1077 ( .A(n1011), .Z(n1033) );
  XNOR U1078 ( .A(n1008), .B(n1034), .Z(n1011) );
  AND U1079 ( .A(n684), .B(n576), .Z(n1034) );
  XOR U1080 ( .A(n1035), .B(n1036), .Z(n1008) );
  ANDN U1081 ( .A(n1037), .B(n1038), .Z(n1036) );
  XNOR U1082 ( .A(n1039), .B(n1035), .Z(n1037) );
  XNOR U1083 ( .A(n1040), .B(n1041), .Z(n1023) );
  IV U1084 ( .A(n1019), .Z(n1041) );
  XNOR U1085 ( .A(n1016), .B(n1042), .Z(n1019) );
  AND U1086 ( .A(n551), .B(n710), .Z(n1042) );
  XOR U1087 ( .A(n1043), .B(n1044), .Z(n1016) );
  ANDN U1088 ( .A(n1045), .B(n1046), .Z(n1044) );
  XNOR U1089 ( .A(n1047), .B(n1043), .Z(n1045) );
  XOR U1090 ( .A(n1048), .B(n1020), .Z(n1040) );
  NAND U1091 ( .A(n639), .B(n616), .Z(n1020) );
  IV U1092 ( .A(n1022), .Z(n1048) );
  XOR U1093 ( .A(n1052), .B(n1053), .Z(n1025) );
  AND U1094 ( .A(n1054), .B(n1055), .Z(n1053) );
  XOR U1095 ( .A(n1056), .B(n1057), .Z(n1055) );
  XOR U1096 ( .A(n1052), .B(n1058), .Z(n1057) );
  XOR U1097 ( .A(n1050), .B(n1059), .Z(n1054) );
  XOR U1098 ( .A(n1052), .B(n1051), .Z(n1059) );
  XNOR U1099 ( .A(n1060), .B(n1039), .Z(n1051) );
  NANDN U1100 ( .B(n829), .A(n509), .Z(n1039) );
  IV U1101 ( .A(n1038), .Z(n1060) );
  XNOR U1102 ( .A(n1035), .B(n1061), .Z(n1038) );
  ANDN U1103 ( .A(n576), .B(n752), .Z(n1061) );
  XOR U1104 ( .A(n1062), .B(n1063), .Z(n1035) );
  ANDN U1105 ( .A(n1064), .B(n1065), .Z(n1063) );
  XNOR U1106 ( .A(n1066), .B(n1062), .Z(n1064) );
  XNOR U1107 ( .A(n1067), .B(n1068), .Z(n1050) );
  IV U1108 ( .A(n1046), .Z(n1068) );
  XNOR U1109 ( .A(n1043), .B(n1069), .Z(n1046) );
  AND U1110 ( .A(n616), .B(n710), .Z(n1069) );
  XOR U1111 ( .A(n1070), .B(n1071), .Z(n1043) );
  ANDN U1112 ( .A(n1072), .B(n1073), .Z(n1071) );
  XNOR U1113 ( .A(n1074), .B(n1070), .Z(n1072) );
  XOR U1114 ( .A(n1075), .B(n1047), .Z(n1067) );
  NAND U1115 ( .A(n639), .B(n684), .Z(n1047) );
  IV U1116 ( .A(n1049), .Z(n1075) );
  XOR U1117 ( .A(n1079), .B(n1080), .Z(n1052) );
  AND U1118 ( .A(n1081), .B(n1082), .Z(n1080) );
  XOR U1119 ( .A(n1083), .B(n1084), .Z(n1082) );
  XOR U1120 ( .A(n1079), .B(n1085), .Z(n1084) );
  XOR U1121 ( .A(n1077), .B(n1086), .Z(n1081) );
  XOR U1122 ( .A(n1079), .B(n1078), .Z(n1086) );
  XNOR U1123 ( .A(n1087), .B(n1066), .Z(n1078) );
  NAND U1124 ( .A(n509), .B(n902), .Z(n1066) );
  IV U1125 ( .A(n1065), .Z(n1087) );
  XNOR U1126 ( .A(n1062), .B(n1088), .Z(n1065) );
  ANDN U1127 ( .A(n576), .B(n829), .Z(n1088) );
  XOR U1128 ( .A(n1089), .B(n1090), .Z(n1062) );
  ANDN U1129 ( .A(n1091), .B(n1092), .Z(n1090) );
  XNOR U1130 ( .A(n1093), .B(n1089), .Z(n1091) );
  XNOR U1131 ( .A(n1094), .B(n1095), .Z(n1077) );
  IV U1132 ( .A(n1073), .Z(n1095) );
  XNOR U1133 ( .A(n1070), .B(n1096), .Z(n1073) );
  AND U1134 ( .A(n684), .B(n710), .Z(n1096) );
  XOR U1135 ( .A(n1097), .B(n1098), .Z(n1070) );
  ANDN U1136 ( .A(n1099), .B(n1100), .Z(n1098) );
  XNOR U1137 ( .A(n1101), .B(n1097), .Z(n1099) );
  XOR U1138 ( .A(n1102), .B(n1074), .Z(n1094) );
  NANDN U1139 ( .B(n752), .A(n639), .Z(n1074) );
  IV U1140 ( .A(n1076), .Z(n1102) );
  XOR U1141 ( .A(n1107), .B(n1108), .Z(n923) );
  XNOR U1142 ( .A(n1109), .B(n1106), .Z(n1107) );
  XNOR U1143 ( .A(n1097), .B(n1111), .Z(n1100) );
  ANDN U1144 ( .A(n710), .B(n752), .Z(n1111) );
  XOR U1145 ( .A(n1114), .B(n1112), .Z(n1113) );
  ANDN U1146 ( .A(n710), .B(n829), .Z(n1114) );
  AND U1147 ( .A(n902), .B(n639), .Z(n1115) );
  XOR U1148 ( .A(n1116), .B(n1117), .Z(n1112) );
  ANDN U1149 ( .A(n1118), .B(n1119), .Z(n1117) );
  XNOR U1150 ( .A(n1120), .B(n1116), .Z(n1118) );
  XOR U1151 ( .A(n1121), .B(n1101), .Z(n1110) );
  NANDN U1152 ( .B(n829), .A(n639), .Z(n1101) );
  IV U1153 ( .A(n1103), .Z(n1121) );
  NAND U1154 ( .A(n639), .B(n1122), .Z(n1120) );
  XNOR U1155 ( .A(n1116), .B(n1123), .Z(n1119) );
  AND U1156 ( .A(n902), .B(n710), .Z(n1123) );
  AND U1157 ( .A(n1124), .B(g_input[0]), .Z(n1116) );
  NANDN U1158 ( .B(n639), .A(n1125), .Z(n1124) );
  NAND U1159 ( .A(n1122), .B(n710), .Z(n1125) );
  XNOR U1160 ( .A(n1092), .B(n1093), .Z(n1105) );
  NAND U1161 ( .A(n509), .B(n1122), .Z(n1093) );
  XNOR U1162 ( .A(n1089), .B(n1128), .Z(n1092) );
  AND U1163 ( .A(n902), .B(n576), .Z(n1128) );
  AND U1164 ( .A(n1129), .B(g_input[0]), .Z(n1089) );
  NANDN U1165 ( .B(n509), .A(n1130), .Z(n1129) );
  NAND U1166 ( .A(n1122), .B(n576), .Z(n1130) );
  XOR U1167 ( .A(n1133), .B(n1134), .Z(n1106) );
  XOR U1168 ( .A(n1135), .B(n1136), .Z(n874) );
  AND U1169 ( .A(n1137), .B(n1138), .Z(n1136) );
  NANDN U1170 ( .B(n197), .A(n1139), .Z(n1138) );
  NANDN U1171 ( .B(n1140), .A(n1141), .Z(n197) );
  AND U1172 ( .A(n1142), .B(g_input[15]), .Z(n1141) );
  OR U1173 ( .A(n1143), .B(n1144), .Z(n1137) );
  IV U1174 ( .A(n873), .Z(n1135) );
  NAND U1175 ( .A(n295), .B(n795), .Z(n928) );
  XNOR U1176 ( .A(n926), .B(n1146), .Z(n927) );
  AND U1177 ( .A(n866), .B(n258), .Z(n1146) );
  XOR U1178 ( .A(n1154), .B(n1143), .Z(n1150) );
  NAND U1179 ( .A(n223), .B(n1139), .Z(n1143) );
  IV U1180 ( .A(n1145), .Z(n1154) );
  NAND U1181 ( .A(n340), .B(n795), .Z(n1149) );
  XNOR U1182 ( .A(n1147), .B(n1156), .Z(n1148) );
  AND U1183 ( .A(n866), .B(n295), .Z(n1156) );
  XNOR U1184 ( .A(n1151), .B(n1161), .Z(n1152) );
  AND U1185 ( .A(n223), .B(e_input[0]), .Z(n1161) );
  XNOR U1186 ( .A(n1142), .B(g_input[14]), .Z(n1140) );
  NOR U1187 ( .A(n1162), .B(n1163), .Z(n1142) );
  XOR U1188 ( .A(n1167), .B(n1153), .Z(n1160) );
  NAND U1189 ( .A(n258), .B(n1139), .Z(n1153) );
  IV U1190 ( .A(n1155), .Z(n1167) );
  NAND U1191 ( .A(n385), .B(n795), .Z(n1159) );
  XNOR U1192 ( .A(n1157), .B(n1169), .Z(n1158) );
  AND U1193 ( .A(n866), .B(n340), .Z(n1169) );
  XOR U1194 ( .A(n1170), .B(n1171), .Z(n1157) );
  ANDN U1195 ( .A(n1172), .B(n1173), .Z(n1171) );
  XNOR U1196 ( .A(n1174), .B(n1170), .Z(n1172) );
  XNOR U1197 ( .A(n1164), .B(n1176), .Z(n1165) );
  AND U1198 ( .A(n258), .B(e_input[0]), .Z(n1176) );
  XOR U1199 ( .A(n1162), .B(g_input[13]), .Z(n1163) );
  NANDN U1200 ( .B(n1177), .A(n1178), .Z(n1162) );
  XOR U1201 ( .A(n1182), .B(n1166), .Z(n1175) );
  NAND U1202 ( .A(n295), .B(n1139), .Z(n1166) );
  IV U1203 ( .A(n1168), .Z(n1182) );
  XNOR U1204 ( .A(n1184), .B(n1174), .Z(n1002) );
  NAND U1205 ( .A(n434), .B(n795), .Z(n1174) );
  IV U1206 ( .A(n1173), .Z(n1184) );
  XNOR U1207 ( .A(n1170), .B(n1185), .Z(n1173) );
  AND U1208 ( .A(n866), .B(n385), .Z(n1185) );
  XOR U1209 ( .A(n1186), .B(n1187), .Z(n1170) );
  ANDN U1210 ( .A(n1188), .B(n1189), .Z(n1187) );
  XNOR U1211 ( .A(n1190), .B(n1186), .Z(n1188) );
  XNOR U1212 ( .A(n1191), .B(n1192), .Z(n1004) );
  IV U1213 ( .A(n1180), .Z(n1192) );
  XNOR U1214 ( .A(n1179), .B(n1193), .Z(n1180) );
  AND U1215 ( .A(n295), .B(e_input[0]), .Z(n1193) );
  XNOR U1216 ( .A(n1178), .B(g_input[12]), .Z(n1177) );
  NOR U1217 ( .A(n1194), .B(n1195), .Z(n1178) );
  XOR U1218 ( .A(n1196), .B(n1197), .Z(n1179) );
  ANDN U1219 ( .A(n1198), .B(n1199), .Z(n1197) );
  XNOR U1220 ( .A(n1200), .B(n1196), .Z(n1198) );
  XOR U1221 ( .A(n1201), .B(n1181), .Z(n1191) );
  NAND U1222 ( .A(n340), .B(n1139), .Z(n1181) );
  IV U1223 ( .A(n1183), .Z(n1201) );
  XNOR U1224 ( .A(n1203), .B(n1190), .Z(n1029) );
  NAND U1225 ( .A(n486), .B(n795), .Z(n1190) );
  IV U1226 ( .A(n1189), .Z(n1203) );
  XNOR U1227 ( .A(n1186), .B(n1204), .Z(n1189) );
  AND U1228 ( .A(n866), .B(n434), .Z(n1204) );
  XOR U1229 ( .A(n1205), .B(n1206), .Z(n1186) );
  ANDN U1230 ( .A(n1207), .B(n1208), .Z(n1206) );
  XNOR U1231 ( .A(n1209), .B(n1205), .Z(n1207) );
  XNOR U1232 ( .A(n1210), .B(n1211), .Z(n1031) );
  IV U1233 ( .A(n1199), .Z(n1211) );
  XNOR U1234 ( .A(n1196), .B(n1212), .Z(n1199) );
  AND U1235 ( .A(n340), .B(e_input[0]), .Z(n1212) );
  XOR U1236 ( .A(n1194), .B(g_input[11]), .Z(n1195) );
  NANDN U1237 ( .B(n1213), .A(n1214), .Z(n1194) );
  XOR U1238 ( .A(n1215), .B(n1216), .Z(n1196) );
  ANDN U1239 ( .A(n1217), .B(n1218), .Z(n1216) );
  XNOR U1240 ( .A(n1219), .B(n1215), .Z(n1217) );
  XOR U1241 ( .A(n1220), .B(n1200), .Z(n1210) );
  NAND U1242 ( .A(n385), .B(n1139), .Z(n1200) );
  IV U1243 ( .A(n1202), .Z(n1220) );
  XNOR U1244 ( .A(n1222), .B(n1209), .Z(n1056) );
  NAND U1245 ( .A(n551), .B(n795), .Z(n1209) );
  IV U1246 ( .A(n1208), .Z(n1222) );
  XNOR U1247 ( .A(n1205), .B(n1223), .Z(n1208) );
  AND U1248 ( .A(n866), .B(n486), .Z(n1223) );
  XOR U1249 ( .A(n1224), .B(n1225), .Z(n1205) );
  ANDN U1250 ( .A(n1226), .B(n1227), .Z(n1225) );
  XNOR U1251 ( .A(n1228), .B(n1224), .Z(n1226) );
  XNOR U1252 ( .A(n1229), .B(n1230), .Z(n1058) );
  IV U1253 ( .A(n1218), .Z(n1230) );
  XNOR U1254 ( .A(n1215), .B(n1231), .Z(n1218) );
  AND U1255 ( .A(n385), .B(e_input[0]), .Z(n1231) );
  XNOR U1256 ( .A(n1214), .B(g_input[10]), .Z(n1213) );
  NOR U1257 ( .A(n1232), .B(n1233), .Z(n1214) );
  XOR U1258 ( .A(n1234), .B(n1235), .Z(n1215) );
  ANDN U1259 ( .A(n1236), .B(n1237), .Z(n1235) );
  XNOR U1260 ( .A(n1238), .B(n1234), .Z(n1236) );
  XOR U1261 ( .A(n1239), .B(n1219), .Z(n1229) );
  NAND U1262 ( .A(n434), .B(n1139), .Z(n1219) );
  IV U1263 ( .A(n1221), .Z(n1239) );
  XNOR U1264 ( .A(n1241), .B(n1228), .Z(n1083) );
  NAND U1265 ( .A(n616), .B(n795), .Z(n1228) );
  IV U1266 ( .A(n1227), .Z(n1241) );
  XNOR U1267 ( .A(n1224), .B(n1242), .Z(n1227) );
  AND U1268 ( .A(n866), .B(n551), .Z(n1242) );
  XOR U1269 ( .A(n1243), .B(n1244), .Z(n1224) );
  ANDN U1270 ( .A(n1245), .B(n1246), .Z(n1244) );
  XNOR U1271 ( .A(n1247), .B(n1243), .Z(n1245) );
  XNOR U1272 ( .A(n1248), .B(n1249), .Z(n1085) );
  IV U1273 ( .A(n1237), .Z(n1249) );
  XNOR U1274 ( .A(n1234), .B(n1250), .Z(n1237) );
  AND U1275 ( .A(n434), .B(e_input[0]), .Z(n1250) );
  XOR U1276 ( .A(n1232), .B(g_input[9]), .Z(n1233) );
  NANDN U1277 ( .B(n1251), .A(n1252), .Z(n1232) );
  XOR U1278 ( .A(n1253), .B(n1254), .Z(n1234) );
  ANDN U1279 ( .A(n1255), .B(n1256), .Z(n1254) );
  XNOR U1280 ( .A(n1257), .B(n1253), .Z(n1255) );
  XOR U1281 ( .A(n1258), .B(n1238), .Z(n1248) );
  NAND U1282 ( .A(n486), .B(n1139), .Z(n1238) );
  IV U1283 ( .A(n1240), .Z(n1258) );
  NAND U1284 ( .A(n684), .B(n795), .Z(n1247) );
  XNOR U1285 ( .A(n1243), .B(n1260), .Z(n1246) );
  AND U1286 ( .A(n866), .B(n616), .Z(n1260) );
  XNOR U1287 ( .A(n1264), .B(n1261), .Z(n1263) );
  XNOR U1288 ( .A(n1253), .B(n1266), .Z(n1256) );
  AND U1289 ( .A(n486), .B(e_input[0]), .Z(n1266) );
  XNOR U1290 ( .A(n1270), .B(n1267), .Z(n1269) );
  XOR U1291 ( .A(n1271), .B(n1257), .Z(n1265) );
  NAND U1292 ( .A(n551), .B(n1139), .Z(n1257) );
  IV U1293 ( .A(n1259), .Z(n1271) );
  XNOR U1294 ( .A(n1272), .B(n1273), .Z(n1259) );
  AND U1295 ( .A(n1274), .B(n1275), .Z(n1273) );
  XOR U1296 ( .A(n1268), .B(n1276), .Z(n1275) );
  XNOR U1297 ( .A(n1270), .B(n1272), .Z(n1276) );
  NAND U1298 ( .A(n616), .B(n1139), .Z(n1270) );
  XOR U1299 ( .A(n1267), .B(n1277), .Z(n1268) );
  AND U1300 ( .A(n551), .B(e_input[0]), .Z(n1277) );
  XNOR U1301 ( .A(n1281), .B(n1278), .Z(n1280) );
  XOR U1302 ( .A(n1262), .B(n1282), .Z(n1274) );
  XNOR U1303 ( .A(n1264), .B(n1272), .Z(n1282) );
  NANDN U1304 ( .B(n752), .A(n795), .Z(n1264) );
  XOR U1305 ( .A(n1261), .B(n1283), .Z(n1262) );
  AND U1306 ( .A(n866), .B(n684), .Z(n1283) );
  XOR U1307 ( .A(n1284), .B(n1285), .Z(n1261) );
  AND U1308 ( .A(n1286), .B(n1287), .Z(n1285) );
  XNOR U1309 ( .A(n1288), .B(n1284), .Z(n1287) );
  XOR U1310 ( .A(n1289), .B(n1290), .Z(n1272) );
  AND U1311 ( .A(n1291), .B(n1292), .Z(n1290) );
  XOR U1312 ( .A(n1279), .B(n1293), .Z(n1292) );
  XNOR U1313 ( .A(n1281), .B(n1289), .Z(n1293) );
  NAND U1314 ( .A(n684), .B(n1139), .Z(n1281) );
  XOR U1315 ( .A(n1278), .B(n1294), .Z(n1279) );
  AND U1316 ( .A(n616), .B(e_input[0]), .Z(n1294) );
  XNOR U1317 ( .A(n1298), .B(n1295), .Z(n1297) );
  XOR U1318 ( .A(n1286), .B(n1299), .Z(n1291) );
  XNOR U1319 ( .A(n1288), .B(n1289), .Z(n1299) );
  NANDN U1320 ( .B(n829), .A(n795), .Z(n1288) );
  XOR U1321 ( .A(n1284), .B(n1300), .Z(n1286) );
  ANDN U1322 ( .A(n866), .B(n752), .Z(n1300) );
  XOR U1323 ( .A(n1301), .B(n1302), .Z(n1284) );
  AND U1324 ( .A(n1303), .B(n1304), .Z(n1302) );
  XNOR U1325 ( .A(n1305), .B(n1301), .Z(n1304) );
  XOR U1326 ( .A(n1306), .B(n1307), .Z(n1289) );
  AND U1327 ( .A(n1308), .B(n1309), .Z(n1307) );
  XOR U1328 ( .A(n1296), .B(n1310), .Z(n1309) );
  XNOR U1329 ( .A(n1298), .B(n1306), .Z(n1310) );
  NANDN U1330 ( .B(n752), .A(n1139), .Z(n1298) );
  XOR U1331 ( .A(n1295), .B(n1311), .Z(n1296) );
  AND U1332 ( .A(n684), .B(e_input[0]), .Z(n1311) );
  XOR U1333 ( .A(n1303), .B(n1315), .Z(n1308) );
  XNOR U1334 ( .A(n1305), .B(n1306), .Z(n1315) );
  NAND U1335 ( .A(n795), .B(n902), .Z(n1305) );
  XOR U1336 ( .A(n1301), .B(n1316), .Z(n1303) );
  ANDN U1337 ( .A(n866), .B(n829), .Z(n1316) );
  NAND U1338 ( .A(n795), .B(n1122), .Z(n1319) );
  XNOR U1339 ( .A(n1317), .B(n1321), .Z(n1318) );
  AND U1340 ( .A(n902), .B(n866), .Z(n1321) );
  AND U1341 ( .A(n1322), .B(g_input[0]), .Z(n1317) );
  NANDN U1342 ( .B(n795), .A(n1323), .Z(n1322) );
  NAND U1343 ( .A(n1122), .B(n866), .Z(n1323) );
  XNOR U1344 ( .A(n1312), .B(n1327), .Z(n1313) );
  ANDN U1345 ( .A(e_input[0]), .B(n752), .Z(n1327) );
  XOR U1346 ( .A(n1330), .B(n1328), .Z(n1329) );
  ANDN U1347 ( .A(e_input[0]), .B(n829), .Z(n1330) );
  AND U1348 ( .A(n1139), .B(n902), .Z(n1331) );
  XOR U1349 ( .A(n1335), .B(n1314), .Z(n1326) );
  NANDN U1350 ( .B(n829), .A(n1139), .Z(n1314) );
  IV U1351 ( .A(n1320), .Z(n1335) );
  NAND U1352 ( .A(n1139), .B(n1122), .Z(n1334) );
  XNOR U1353 ( .A(n1332), .B(n1336), .Z(n1333) );
  AND U1354 ( .A(n902), .B(e_input[0]), .Z(n1336) );
  AND U1355 ( .A(n1337), .B(g_input[0]), .Z(n1332) );
  NANDN U1356 ( .B(n1139), .A(n1338), .Z(n1337) );
  NAND U1357 ( .A(n1122), .B(e_input[0]), .Z(n1338) );
  XNOR U1358 ( .A(n1340), .B(n892), .Z(n882) );
  XNOR U1359 ( .A(n879), .B(n880), .Z(n892) );
  NAND U1360 ( .A(n323), .B(n684), .Z(n880) );
  XNOR U1361 ( .A(n878), .B(n1341), .Z(n879) );
  AND U1362 ( .A(n616), .B(n364), .Z(n1341) );
  XNOR U1363 ( .A(n1345), .B(n1342), .Z(n1344) );
  XNOR U1364 ( .A(n891), .B(n881), .Z(n1340) );
  XOR U1365 ( .A(n1346), .B(n1347), .Z(n881) );
  XNOR U1366 ( .A(n886), .B(n1349), .Z(n887) );
  AND U1367 ( .A(n486), .B(n471), .Z(n1349) );
  XNOR U1368 ( .A(n1252), .B(g_input[8]), .Z(n1251) );
  NOR U1369 ( .A(n1350), .B(n1351), .Z(n1252) );
  XOR U1370 ( .A(n1352), .B(n1353), .Z(n886) );
  AND U1371 ( .A(n1354), .B(n1355), .Z(n1353) );
  XNOR U1372 ( .A(n1356), .B(n1352), .Z(n1355) );
  XOR U1373 ( .A(n1357), .B(n888), .Z(n1348) );
  NAND U1374 ( .A(n417), .B(n551), .Z(n888) );
  IV U1375 ( .A(n890), .Z(n1357) );
  XNOR U1376 ( .A(n1358), .B(n1359), .Z(n890) );
  AND U1377 ( .A(n1360), .B(n1361), .Z(n1359) );
  XOR U1378 ( .A(n1354), .B(n1362), .Z(n1361) );
  XNOR U1379 ( .A(n1356), .B(n1358), .Z(n1362) );
  NAND U1380 ( .A(n417), .B(n616), .Z(n1356) );
  XOR U1381 ( .A(n1352), .B(n1363), .Z(n1354) );
  AND U1382 ( .A(n551), .B(n471), .Z(n1363) );
  XOR U1383 ( .A(n1350), .B(g_input[7]), .Z(n1351) );
  NANDN U1384 ( .B(n1364), .A(n1365), .Z(n1350) );
  XOR U1385 ( .A(n1366), .B(n1367), .Z(n1352) );
  AND U1386 ( .A(n1368), .B(n1369), .Z(n1367) );
  XNOR U1387 ( .A(n1370), .B(n1366), .Z(n1369) );
  XOR U1388 ( .A(n1343), .B(n1371), .Z(n1360) );
  XNOR U1389 ( .A(n1345), .B(n1358), .Z(n1371) );
  NANDN U1390 ( .B(n752), .A(n323), .Z(n1345) );
  XOR U1391 ( .A(n1342), .B(n1372), .Z(n1343) );
  AND U1392 ( .A(n684), .B(n364), .Z(n1372) );
  XNOR U1393 ( .A(n1376), .B(n1373), .Z(n1375) );
  XOR U1394 ( .A(n1377), .B(n1378), .Z(n1358) );
  AND U1395 ( .A(n1379), .B(n1380), .Z(n1378) );
  XOR U1396 ( .A(n1368), .B(n1381), .Z(n1380) );
  XNOR U1397 ( .A(n1370), .B(n1377), .Z(n1381) );
  NAND U1398 ( .A(n417), .B(n684), .Z(n1370) );
  XOR U1399 ( .A(n1366), .B(n1382), .Z(n1368) );
  AND U1400 ( .A(n616), .B(n471), .Z(n1382) );
  XNOR U1401 ( .A(n1365), .B(g_input[6]), .Z(n1364) );
  NOR U1402 ( .A(n1383), .B(n1384), .Z(n1365) );
  XOR U1403 ( .A(n1385), .B(n1386), .Z(n1366) );
  AND U1404 ( .A(n1387), .B(n1388), .Z(n1386) );
  XNOR U1405 ( .A(n1389), .B(n1385), .Z(n1388) );
  XOR U1406 ( .A(n1374), .B(n1390), .Z(n1379) );
  XNOR U1407 ( .A(n1376), .B(n1377), .Z(n1390) );
  NANDN U1408 ( .B(n829), .A(n323), .Z(n1376) );
  XOR U1409 ( .A(n1373), .B(n1391), .Z(n1374) );
  ANDN U1410 ( .A(n364), .B(n752), .Z(n1391) );
  XNOR U1411 ( .A(n1395), .B(n1392), .Z(n1394) );
  XOR U1412 ( .A(n1396), .B(n1397), .Z(n1377) );
  AND U1413 ( .A(n1398), .B(n1399), .Z(n1397) );
  XOR U1414 ( .A(n1387), .B(n1400), .Z(n1399) );
  XNOR U1415 ( .A(n1389), .B(n1396), .Z(n1400) );
  NANDN U1416 ( .B(n752), .A(n417), .Z(n1389) );
  XOR U1417 ( .A(n1385), .B(n1401), .Z(n1387) );
  AND U1418 ( .A(n684), .B(n471), .Z(n1401) );
  XOR U1419 ( .A(n1383), .B(g_input[5]), .Z(n1384) );
  NANDN U1420 ( .B(n1402), .A(n1403), .Z(n1383) );
  XOR U1421 ( .A(n1404), .B(n1405), .Z(n1385) );
  ANDN U1422 ( .A(n1406), .B(n1407), .Z(n1405) );
  XNOR U1423 ( .A(n1408), .B(n1404), .Z(n1406) );
  XOR U1424 ( .A(n1393), .B(n1409), .Z(n1398) );
  XNOR U1425 ( .A(n1395), .B(n1396), .Z(n1409) );
  NAND U1426 ( .A(n323), .B(n902), .Z(n1395) );
  XOR U1427 ( .A(n1392), .B(n1410), .Z(n1393) );
  ANDN U1428 ( .A(n364), .B(n829), .Z(n1410) );
  XOR U1429 ( .A(n1411), .B(n1412), .Z(n1392) );
  ANDN U1430 ( .A(n1413), .B(n1414), .Z(n1412) );
  XNOR U1431 ( .A(n1415), .B(n1411), .Z(n1413) );
  NAND U1432 ( .A(n323), .B(n1122), .Z(n1415) );
  XNOR U1433 ( .A(n1411), .B(n1417), .Z(n1414) );
  AND U1434 ( .A(n902), .B(n364), .Z(n1417) );
  AND U1435 ( .A(n1418), .B(g_input[0]), .Z(n1411) );
  NANDN U1436 ( .B(n323), .A(n1419), .Z(n1418) );
  NAND U1437 ( .A(n1122), .B(n364), .Z(n1419) );
  XNOR U1438 ( .A(n1404), .B(n1423), .Z(n1407) );
  ANDN U1439 ( .A(n471), .B(n752), .Z(n1423) );
  XOR U1440 ( .A(n1424), .B(n1425), .Z(n1404) );
  AND U1441 ( .A(n1426), .B(n1427), .Z(n1425) );
  XOR U1442 ( .A(n1428), .B(n1424), .Z(n1427) );
  ANDN U1443 ( .A(n471), .B(n829), .Z(n1428) );
  XOR U1444 ( .A(n1429), .B(n1424), .Z(n1426) );
  AND U1445 ( .A(n902), .B(n417), .Z(n1429) );
  XOR U1446 ( .A(n1430), .B(n1431), .Z(n1424) );
  ANDN U1447 ( .A(n1432), .B(n1433), .Z(n1431) );
  XNOR U1448 ( .A(n1434), .B(n1430), .Z(n1432) );
  XOR U1449 ( .A(n1435), .B(n1408), .Z(n1422) );
  NANDN U1450 ( .B(n829), .A(n417), .Z(n1408) );
  IV U1451 ( .A(n1416), .Z(n1435) );
  XOR U1452 ( .A(n1436), .B(n1434), .Z(n1416) );
  NAND U1453 ( .A(n417), .B(n1122), .Z(n1434) );
  IV U1454 ( .A(n1433), .Z(n1436) );
  XNOR U1455 ( .A(n1430), .B(n1437), .Z(n1433) );
  AND U1456 ( .A(n902), .B(n471), .Z(n1437) );
  AND U1457 ( .A(n1438), .B(g_input[0]), .Z(n1430) );
  NANDN U1458 ( .B(n417), .A(n1439), .Z(n1438) );
  NAND U1459 ( .A(n1122), .B(n471), .Z(n1439) );
  XNOR U1460 ( .A(n895), .B(n1443), .Z(n896) );
  ANDN U1461 ( .A(n291), .B(n752), .Z(n1443) );
  XNOR U1462 ( .A(n1403), .B(g_input[4]), .Z(n1402) );
  NOR U1463 ( .A(n1444), .B(n1445), .Z(n1403) );
  XOR U1464 ( .A(n1446), .B(n1447), .Z(n895) );
  AND U1465 ( .A(n1448), .B(n1449), .Z(n1447) );
  XOR U1466 ( .A(n1450), .B(n1446), .Z(n1449) );
  ANDN U1467 ( .A(n291), .B(n829), .Z(n1450) );
  XOR U1468 ( .A(n1451), .B(n1446), .Z(n1448) );
  AND U1469 ( .A(n902), .B(n253), .Z(n1451) );
  XOR U1470 ( .A(n1452), .B(n1453), .Z(n1446) );
  ANDN U1471 ( .A(n1454), .B(n1455), .Z(n1453) );
  XNOR U1472 ( .A(n1456), .B(n1452), .Z(n1454) );
  XOR U1473 ( .A(n1457), .B(n897), .Z(n1442) );
  NANDN U1474 ( .B(n829), .A(n253), .Z(n897) );
  NANDN U1475 ( .B(n1458), .A(n1459), .Z(n1444) );
  IV U1476 ( .A(n899), .Z(n1457) );
  NAND U1477 ( .A(n253), .B(n1122), .Z(n1456) );
  XNOR U1478 ( .A(n1452), .B(n1460), .Z(n1455) );
  AND U1479 ( .A(n902), .B(n291), .Z(n1460) );
  AND U1480 ( .A(n1461), .B(g_input[0]), .Z(n1452) );
  NANDN U1481 ( .B(n253), .A(n1462), .Z(n1461) );
  NAND U1482 ( .A(n1122), .B(n291), .Z(n1462) );
  XNOR U1483 ( .A(n1463), .B(e_input[12]), .Z(n291) );
  NAND U1484 ( .A(n1464), .B(e_input[15]), .Z(n1463) );
  XOR U1485 ( .A(n1465), .B(e_input[12]), .Z(n1464) );
  XNOR U1486 ( .A(n906), .B(n907), .Z(n901) );
  NANDN U1487 ( .B(n198), .A(n1122), .Z(n907) );
  XNOR U1488 ( .A(n905), .B(n1467), .Z(n906) );
  AND U1489 ( .A(n902), .B(n222), .Z(n1467) );
  XNOR U1490 ( .A(n1459), .B(g_input[2]), .Z(n1458) );
  AND U1491 ( .A(n1469), .B(g_input[0]), .Z(n905) );
  NAND U1492 ( .A(n1470), .B(n198), .Z(n1469) );
  NANDN U1493 ( .B(n1471), .A(n1472), .Z(n198) );
  ANDN U1494 ( .A(e_input[15]), .B(n1473), .Z(n1472) );
  NAND U1495 ( .A(n1122), .B(n222), .Z(n1470) );
  XOR U1496 ( .A(n1473), .B(e_input[14]), .Z(n1471) );
  OR U1497 ( .A(n1466), .B(n1474), .Z(n1473) );
  XOR U1498 ( .A(n1474), .B(e_input[13]), .Z(n1466) );
  OR U1499 ( .A(n1465), .B(n1475), .Z(n1474) );
  XOR U1500 ( .A(n1475), .B(e_input[12]), .Z(n1465) );
  OR U1501 ( .A(n1421), .B(n1476), .Z(n1475) );
  XOR U1502 ( .A(n1476), .B(e_input[11]), .Z(n1421) );
  OR U1503 ( .A(n1420), .B(n1477), .Z(n1476) );
  XOR U1504 ( .A(n1477), .B(e_input[10]), .Z(n1420) );
  OR U1505 ( .A(n1441), .B(n1478), .Z(n1477) );
  XOR U1506 ( .A(n1478), .B(e_input[9]), .Z(n1441) );
  OR U1507 ( .A(n1440), .B(n1479), .Z(n1478) );
  XOR U1508 ( .A(n1479), .B(e_input[8]), .Z(n1440) );
  OR U1509 ( .A(n1132), .B(n1480), .Z(n1479) );
  XOR U1510 ( .A(n1480), .B(e_input[7]), .Z(n1132) );
  OR U1511 ( .A(n1131), .B(n1481), .Z(n1480) );
  XOR U1512 ( .A(n1481), .B(e_input[6]), .Z(n1131) );
  OR U1513 ( .A(n1127), .B(n1482), .Z(n1481) );
  XOR U1514 ( .A(n1482), .B(e_input[5]), .Z(n1127) );
  OR U1515 ( .A(n1126), .B(n1483), .Z(n1482) );
  XOR U1516 ( .A(n1483), .B(e_input[4]), .Z(n1126) );
  OR U1517 ( .A(n1325), .B(n1484), .Z(n1483) );
  XOR U1518 ( .A(n1484), .B(e_input[3]), .Z(n1325) );
  OR U1519 ( .A(n1324), .B(n1485), .Z(n1484) );
  XOR U1520 ( .A(n1485), .B(e_input[2]), .Z(n1324) );
  NANDN U1521 ( .B(e_input[0]), .A(n1339), .Z(n1485) );
  XNOR U1522 ( .A(e_input[0]), .B(e_input[1]), .Z(n1339) );
  XOR U1523 ( .A(g_input[0]), .B(g_input[1]), .Z(n1468) );
  NANDN U1524 ( .B(n841), .A(n113), .Z(n165) );
  IV U1525 ( .A(rst), .Z(n113) );
  NAND U1526 ( .A(n1486), .B(n1487), .Z(n841) );
  AND U1527 ( .A(n1488), .B(n1489), .Z(n1487) );
  ANDN U1528 ( .A(n1490), .B(\_MxM/n[7] ), .Z(n1489) );
  NOR U1529 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n1490) );
  NOR U1530 ( .A(\_MxM/n[5] ), .B(\_MxM/n[6] ), .Z(n1488) );
  AND U1531 ( .A(n1491), .B(n1492), .Z(n1486) );
  NOR U1532 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n1492) );
  NOR U1533 ( .A(\_MxM/n[0] ), .B(n106), .Z(n1491) );
  OR U1534 ( .A(\_MxM/n[3] ), .B(\_MxM/n[4] ), .Z(n106) );
endmodule

