
module MxM_TG_W8_N1000 ( clk, rst, g_input, e_input, o );
  input [7:0] g_input;
  input [7:0] e_input;
  output [7:0] o;
  input clk, rst;
  wire   \_MxM/n148 , \_MxM/n147 , \_MxM/n146 , \_MxM/n145 , \_MxM/n144 ,
         \_MxM/n143 , \_MxM/n142 , \_MxM/n141 , \_MxM/n140 , \_MxM/n139 ,
         \_MxM/n138 , \_MxM/n137 , \_MxM/n136 , \_MxM/n135 , \_MxM/n134 ,
         \_MxM/n133 , \_MxM/n132 , \_MxM/n131 , \_MxM/n130 , \_MxM/n129 ,
         \_MxM/n128 , \_MxM/n127 , \_MxM/n126 , \_MxM/n125 , \_MxM/n124 ,
         \_MxM/n123 , \_MxM/N15 , \_MxM/N14 , \_MxM/N13 , \_MxM/N12 ,
         \_MxM/N11 , \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/n[0] ,
         \_MxM/n[1] , \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] ,
         \_MxM/n[6] , \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/Y0[0] ,
         \_MxM/Y0[1] , \_MxM/Y0[2] , \_MxM/Y0[3] , \_MxM/Y0[4] , \_MxM/Y0[5] ,
         \_MxM/Y0[6] , \_MxM/Y0[7] , \_MxM/add_39/carry[9] ,
         \_MxM/add_39/carry[8] , \_MxM/add_39/carry[7] ,
         \_MxM/add_39/carry[6] , \_MxM/add_39/carry[5] ,
         \_MxM/add_39/carry[4] , \_MxM/add_39/carry[3] ,
         \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n123 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n124 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n125 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n126 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n127 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n128 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n129 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n130 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n131 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n132 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n133 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n134 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n135 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n136 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n137 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n138 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/n139 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/n140 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/n141 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n142 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n143 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n144 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n145 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n146 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n147 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n148 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N14 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N15 ) );
  MUX U1 ( .IN0(n322), .IN1(n338), .SEL(n324), .F(n303) );
  MUX U2 ( .IN0(g_input[3]), .IN1(n387), .SEL(g_input[7]), .F(n1) );
  IV U3 ( .A(n1), .Z(n232) );
  MUX U4 ( .IN0(n272), .IN1(n270), .SEL(n271), .F(n227) );
  NAND U5 ( .A(n145), .B(n179), .Z(n178) );
  MUX U6 ( .IN0(n255), .IN1(n2), .SEL(n254), .F(n210) );
  IV U7 ( .A(n253), .Z(n2) );
  MUX U8 ( .IN0(n3), .IN1(n155), .SEL(n156), .F(n123) );
  IV U9 ( .A(\_MxM/Y0[3] ), .Z(n3) );
  XOR U10 ( .A(n386), .B(g_input[3]), .Z(n387) );
  XNOR U11 ( .A(n374), .B(n375), .Z(n353) );
  MUX U12 ( .IN0(e_input[6]), .IN1(n412), .SEL(e_input[7]), .F(n121) );
  MUX U13 ( .IN0(e_input[3]), .IN1(n362), .SEL(e_input[7]), .F(n213) );
  MUX U14 ( .IN0(n216), .IN1(n4), .SEL(n217), .F(n168) );
  IV U15 ( .A(n218), .Z(n4) );
  XNOR U16 ( .A(n219), .B(n184), .Z(n176) );
  MUX U17 ( .IN0(n5), .IN1(n238), .SEL(n239), .F(n193) );
  IV U18 ( .A(\_MxM/Y0[1] ), .Z(n5) );
  XOR U19 ( .A(n91), .B(n101), .Z(n99) );
  MUX U20 ( .IN0(n6), .IN1(n392), .SEL(n393), .F(n388) );
  IV U21 ( .A(n394), .Z(n6) );
  MUX U22 ( .IN0(g_input[4]), .IN1(n339), .SEL(g_input[7]), .F(n7) );
  IV U23 ( .A(n7), .Z(n186) );
  MUX U24 ( .IN0(g_input[5]), .IN1(n321), .SEL(g_input[7]), .F(n149) );
  XOR U25 ( .A(n235), .B(n274), .Z(n236) );
  MUX U26 ( .IN0(g_input[6]), .IN1(n293), .SEL(g_input[7]), .F(n122) );
  MUX U27 ( .IN0(n256), .IN1(n8), .SEL(n257), .F(n216) );
  IV U28 ( .A(n258), .Z(n8) );
  XNOR U29 ( .A(n138), .B(n139), .Z(n162) );
  XOR U30 ( .A(n123), .B(n133), .Z(n131) );
  NOR U31 ( .A(g_input[0]), .B(n409), .Z(n397) );
  MUX U32 ( .IN0(n9), .IN1(n286), .SEL(n287), .F(n333) );
  IV U33 ( .A(n353), .Z(n9) );
  MUX U34 ( .IN0(n388), .IN1(n391), .SEL(n389), .F(n264) );
  MUX U35 ( .IN0(n303), .IN1(n319), .SEL(n305), .F(n297) );
  MUX U36 ( .IN0(n148), .IN1(n172), .SEL(n147), .F(n110) );
  NAND U37 ( .A(n210), .B(n251), .Z(n250) );
  XNOR U38 ( .A(n272), .B(n271), .Z(n258) );
  XNOR U39 ( .A(n177), .B(n176), .Z(n170) );
  XNOR U40 ( .A(n231), .B(n230), .Z(n218) );
  MUX U41 ( .IN0(\_MxM/Y0[6] ), .IN1(n73), .SEL(n68), .F(n61) );
  XOR U42 ( .A(n155), .B(n163), .Z(n161) );
  MUX U43 ( .IN0(g_input[2]), .IN1(n396), .SEL(g_input[7]), .F(n273) );
  XOR U44 ( .A(n363), .B(n344), .Z(n287) );
  XNOR U45 ( .A(n262), .B(n224), .Z(n230) );
  MUX U46 ( .IN0(n261), .IN1(n259), .SEL(n260), .F(n10) );
  IV U47 ( .A(n10), .Z(n215) );
  AND U48 ( .A(n116), .B(n82), .Z(n115) );
  MUX U49 ( .IN0(n11), .IN1(n170), .SEL(n169), .F(n139) );
  IV U50 ( .A(n168), .Z(n11) );
  MUX U51 ( .IN0(n12), .IN1(n193), .SEL(n194), .F(n155) );
  IV U52 ( .A(\_MxM/Y0[2] ), .Z(n12) );
  MUX U53 ( .IN0(\_MxM/Y0[7] ), .IN1(n61), .SEL(n62), .F(n13) );
  IV U54 ( .A(n13), .Z(n58) );
  XOR U55 ( .A(n239), .B(\_MxM/Y0[1] ), .Z(n27) );
  ANDN U56 ( .A(n14), .B(\_MxM/n[0] ), .Z(\_MxM/n148 ) );
  AND U57 ( .A(\_MxM/N8 ), .B(n14), .Z(\_MxM/n147 ) );
  AND U58 ( .A(\_MxM/N9 ), .B(n14), .Z(\_MxM/n146 ) );
  AND U59 ( .A(\_MxM/N10 ), .B(n14), .Z(\_MxM/n145 ) );
  AND U60 ( .A(\_MxM/N11 ), .B(n14), .Z(\_MxM/n144 ) );
  AND U61 ( .A(\_MxM/N12 ), .B(n14), .Z(\_MxM/n143 ) );
  AND U62 ( .A(\_MxM/N13 ), .B(n14), .Z(\_MxM/n142 ) );
  AND U63 ( .A(\_MxM/N14 ), .B(n14), .Z(\_MxM/n141 ) );
  AND U64 ( .A(\_MxM/N15 ), .B(n14), .Z(\_MxM/n140 ) );
  AND U65 ( .A(n14), .B(n15), .Z(\_MxM/n139 ) );
  XOR U66 ( .A(\_MxM/n[9] ), .B(\_MxM/add_39/carry[9] ), .Z(n15) );
  ANDN U67 ( .A(n16), .B(rst), .Z(n14) );
  NAND U68 ( .A(n17), .B(n18), .Z(n16) );
  AND U69 ( .A(n19), .B(n20), .Z(n18) );
  AND U70 ( .A(\_MxM/n[1] ), .B(n21), .Z(n20) );
  ANDN U71 ( .A(\_MxM/n[0] ), .B(n22), .Z(n21) );
  AND U72 ( .A(\_MxM/n[5] ), .B(\_MxM/n[2] ), .Z(n19) );
  AND U73 ( .A(n23), .B(n24), .Z(n17) );
  AND U74 ( .A(\_MxM/n[7] ), .B(\_MxM/n[6] ), .Z(n24) );
  AND U75 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n23) );
  NAND U76 ( .A(n25), .B(n26), .Z(\_MxM/n138 ) );
  OR U77 ( .A(n27), .B(n28), .Z(n26) );
  NANDN U78 ( .B(n29), .A(\_MxM/Y0[0] ), .Z(n25) );
  NAND U79 ( .A(n30), .B(n31), .Z(\_MxM/n137 ) );
  NANDN U80 ( .B(n28), .A(n32), .Z(n31) );
  NANDN U81 ( .B(n33), .A(rst), .Z(n30) );
  NAND U82 ( .A(n34), .B(n35), .Z(\_MxM/n136 ) );
  NANDN U83 ( .B(n28), .A(n36), .Z(n35) );
  NANDN U84 ( .B(n29), .A(\_MxM/Y0[2] ), .Z(n34) );
  NAND U85 ( .A(n37), .B(n38), .Z(\_MxM/n135 ) );
  NANDN U86 ( .B(n28), .A(n39), .Z(n38) );
  NANDN U87 ( .B(n29), .A(\_MxM/Y0[3] ), .Z(n37) );
  NAND U88 ( .A(n40), .B(n41), .Z(\_MxM/n134 ) );
  NANDN U89 ( .B(n28), .A(n42), .Z(n41) );
  NANDN U90 ( .B(n29), .A(\_MxM/Y0[4] ), .Z(n40) );
  NAND U91 ( .A(n43), .B(n44), .Z(\_MxM/n133 ) );
  NANDN U92 ( .B(n28), .A(n45), .Z(n44) );
  NANDN U93 ( .B(n29), .A(\_MxM/Y0[5] ), .Z(n43) );
  NAND U94 ( .A(n46), .B(n47), .Z(\_MxM/n132 ) );
  OR U95 ( .A(n48), .B(n28), .Z(n47) );
  NANDN U96 ( .B(n29), .A(\_MxM/Y0[6] ), .Z(n46) );
  NAND U97 ( .A(n49), .B(n50), .Z(\_MxM/n131 ) );
  OR U98 ( .A(n28), .B(n51), .Z(n50) );
  NANDN U99 ( .B(n52), .A(n29), .Z(n28) );
  NANDN U100 ( .B(n29), .A(\_MxM/Y0[7] ), .Z(n49) );
  NAND U101 ( .A(n53), .B(n54), .Z(\_MxM/n130 ) );
  NANDN U102 ( .B(n29), .A(o[7]), .Z(n54) );
  AND U103 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U104 ( .B(n52), .A(o[7]), .Z(n56) );
  OR U105 ( .A(n51), .B(n57), .Z(n55) );
  XOR U106 ( .A(n58), .B(n59), .Z(n51) );
  XNOR U107 ( .A(\_MxM/Y0[7] ), .B(n60), .Z(n59) );
  NAND U108 ( .A(n63), .B(n64), .Z(\_MxM/n129 ) );
  NANDN U109 ( .B(n29), .A(o[6]), .Z(n64) );
  AND U110 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U111 ( .B(n52), .A(o[6]), .Z(n66) );
  OR U112 ( .A(n48), .B(n57), .Z(n65) );
  XOR U113 ( .A(n62), .B(\_MxM/Y0[7] ), .Z(n48) );
  XOR U114 ( .A(n61), .B(n60), .Z(n62) );
  NAND U115 ( .A(n69), .B(n70), .Z(\_MxM/n128 ) );
  NANDN U116 ( .B(n29), .A(o[5]), .Z(n70) );
  AND U117 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U118 ( .B(n52), .A(o[5]), .Z(n72) );
  NANDN U119 ( .B(n57), .A(n45), .Z(n71) );
  XNOR U120 ( .A(n68), .B(\_MxM/Y0[6] ), .Z(n45) );
  XOR U121 ( .A(n73), .B(n74), .Z(n68) );
  ANDN U122 ( .A(n60), .B(n75), .Z(n74) );
  NANDN U123 ( .B(n76), .A(n77), .Z(n60) );
  ANDN U124 ( .A(n78), .B(n75), .Z(n76) );
  NAND U125 ( .A(n79), .B(n80), .Z(n75) );
  OR U126 ( .A(n81), .B(n82), .Z(n80) );
  AND U127 ( .A(n83), .B(n84), .Z(n79) );
  OR U128 ( .A(n85), .B(n86), .Z(n84) );
  OR U129 ( .A(n87), .B(n88), .Z(n83) );
  NOR U130 ( .A(n89), .B(n90), .Z(n78) );
  IV U131 ( .A(n67), .Z(n73) );
  XOR U132 ( .A(n91), .B(n92), .Z(n67) );
  ANDN U133 ( .A(n93), .B(n94), .Z(n92) );
  XNOR U134 ( .A(\_MxM/Y0[5] ), .B(n91), .Z(n93) );
  NAND U135 ( .A(n95), .B(n96), .Z(\_MxM/n127 ) );
  NANDN U136 ( .B(n29), .A(o[4]), .Z(n96) );
  AND U137 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U138 ( .B(n52), .A(o[4]), .Z(n98) );
  NANDN U139 ( .B(n57), .A(n42), .Z(n97) );
  XNOR U140 ( .A(n94), .B(\_MxM/Y0[5] ), .Z(n42) );
  XNOR U141 ( .A(n99), .B(n100), .Z(n94) );
  AND U142 ( .A(n77), .B(n102), .Z(n101) );
  XOR U143 ( .A(n89), .B(n103), .Z(n102) );
  XOR U144 ( .A(n103), .B(n90), .Z(n89) );
  OR U145 ( .A(n104), .B(n105), .Z(n90) );
  IV U146 ( .A(n100), .Z(n103) );
  XNOR U147 ( .A(n88), .B(n87), .Z(n100) );
  OR U148 ( .A(n106), .B(n107), .Z(n87) );
  AND U149 ( .A(n108), .B(n109), .Z(n88) );
  XNOR U150 ( .A(n110), .B(n111), .Z(n109) );
  ANDN U151 ( .A(n112), .B(n113), .Z(n111) );
  XOR U152 ( .A(n110), .B(n114), .Z(n112) );
  XNOR U153 ( .A(n81), .B(n115), .Z(n108) );
  NAND U154 ( .A(n117), .B(n118), .Z(n82) );
  NANDN U155 ( .B(n119), .A(n120), .Z(n117) );
  NANDN U156 ( .B(n85), .A(n121), .Z(n116) );
  NANDN U157 ( .B(n86), .A(n122), .Z(n81) );
  XOR U158 ( .A(n123), .B(n124), .Z(n91) );
  ANDN U159 ( .A(n125), .B(n126), .Z(n124) );
  XNOR U160 ( .A(\_MxM/Y0[4] ), .B(n123), .Z(n125) );
  NAND U161 ( .A(n127), .B(n128), .Z(\_MxM/n126 ) );
  NANDN U162 ( .B(n29), .A(o[3]), .Z(n128) );
  AND U163 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U164 ( .B(n52), .A(o[3]), .Z(n130) );
  NANDN U165 ( .B(n57), .A(n39), .Z(n129) );
  XNOR U166 ( .A(n126), .B(\_MxM/Y0[4] ), .Z(n39) );
  XNOR U167 ( .A(n131), .B(n132), .Z(n126) );
  AND U168 ( .A(n77), .B(n134), .Z(n133) );
  XOR U169 ( .A(n104), .B(n135), .Z(n134) );
  XOR U170 ( .A(n135), .B(n105), .Z(n104) );
  OR U171 ( .A(n136), .B(n137), .Z(n105) );
  IV U172 ( .A(n132), .Z(n135) );
  XNOR U173 ( .A(n107), .B(n106), .Z(n132) );
  OR U174 ( .A(n138), .B(n139), .Z(n106) );
  XOR U175 ( .A(n114), .B(n113), .Z(n107) );
  XOR U176 ( .A(n110), .B(n140), .Z(n113) );
  AND U177 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U178 ( .B(n85), .A(n143), .Z(n142) );
  OR U179 ( .A(n144), .B(n145), .Z(n141) );
  XOR U180 ( .A(n119), .B(n120), .Z(n114) );
  NANDN U181 ( .B(n86), .A(n149), .Z(n120) );
  XNOR U182 ( .A(n118), .B(n150), .Z(n119) );
  AND U183 ( .A(n122), .B(n121), .Z(n150) );
  ANDN U184 ( .A(n151), .B(n152), .Z(n118) );
  NANDN U185 ( .B(n153), .A(n154), .Z(n151) );
  NAND U186 ( .A(n157), .B(n158), .Z(\_MxM/n125 ) );
  NANDN U187 ( .B(n29), .A(o[2]), .Z(n158) );
  AND U188 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U189 ( .B(n52), .A(o[2]), .Z(n160) );
  NANDN U190 ( .B(n57), .A(n36), .Z(n159) );
  XNOR U191 ( .A(n156), .B(\_MxM/Y0[3] ), .Z(n36) );
  XNOR U192 ( .A(n161), .B(n162), .Z(n156) );
  AND U193 ( .A(n77), .B(n164), .Z(n163) );
  XOR U194 ( .A(n136), .B(n165), .Z(n164) );
  XOR U195 ( .A(n165), .B(n137), .Z(n136) );
  OR U196 ( .A(n166), .B(n167), .Z(n137) );
  IV U197 ( .A(n162), .Z(n165) );
  XOR U198 ( .A(n148), .B(n147), .Z(n138) );
  XNOR U199 ( .A(n171), .B(n172), .Z(n147) );
  IV U200 ( .A(n146), .Z(n172) );
  XOR U201 ( .A(n173), .B(n174), .Z(n146) );
  ANDN U202 ( .A(n175), .B(n176), .Z(n174) );
  XOR U203 ( .A(n173), .B(n177), .Z(n175) );
  XNOR U204 ( .A(n178), .B(n144), .Z(n171) );
  NAND U205 ( .A(n143), .B(n122), .Z(n144) );
  NANDN U206 ( .B(n85), .A(n180), .Z(n179) );
  XNOR U207 ( .A(n181), .B(n182), .Z(n145) );
  ANDN U208 ( .A(n183), .B(n184), .Z(n182) );
  XNOR U209 ( .A(n185), .B(n181), .Z(n183) );
  XOR U210 ( .A(n153), .B(n154), .Z(n148) );
  OR U211 ( .A(n186), .B(n86), .Z(n154) );
  XNOR U212 ( .A(n187), .B(n188), .Z(n153) );
  AND U213 ( .A(n149), .B(n121), .Z(n188) );
  IV U214 ( .A(n152), .Z(n187) );
  NAND U215 ( .A(n189), .B(n190), .Z(n152) );
  NANDN U216 ( .B(n191), .A(n192), .Z(n189) );
  NAND U217 ( .A(n195), .B(n196), .Z(\_MxM/n124 ) );
  NANDN U218 ( .B(n29), .A(o[1]), .Z(n196) );
  AND U219 ( .A(n197), .B(n198), .Z(n195) );
  NANDN U220 ( .B(n52), .A(o[1]), .Z(n198) );
  NANDN U221 ( .B(n57), .A(n32), .Z(n197) );
  XNOR U222 ( .A(n194), .B(\_MxM/Y0[2] ), .Z(n32) );
  XNOR U223 ( .A(n199), .B(n200), .Z(n194) );
  XOR U224 ( .A(n193), .B(n201), .Z(n199) );
  AND U225 ( .A(n77), .B(n202), .Z(n201) );
  XOR U226 ( .A(n166), .B(n203), .Z(n202) );
  XOR U227 ( .A(n203), .B(n167), .Z(n166) );
  NANDN U228 ( .B(n204), .A(n205), .Z(n167) );
  IV U229 ( .A(n200), .Z(n203) );
  XOR U230 ( .A(n170), .B(n169), .Z(n200) );
  XNOR U231 ( .A(n168), .B(n206), .Z(n169) );
  AND U232 ( .A(n207), .B(n208), .Z(n206) );
  OR U233 ( .A(n209), .B(n210), .Z(n208) );
  AND U234 ( .A(n211), .B(n212), .Z(n207) );
  NANDN U235 ( .B(n85), .A(n213), .Z(n212) );
  NAND U236 ( .A(n214), .B(n215), .Z(n211) );
  XNOR U237 ( .A(n181), .B(n220), .Z(n184) );
  AND U238 ( .A(n122), .B(n180), .Z(n220) );
  XOR U239 ( .A(n221), .B(n222), .Z(n181) );
  ANDN U240 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U241 ( .A(n225), .B(n221), .Z(n223) );
  XOR U242 ( .A(n226), .B(n185), .Z(n219) );
  NAND U243 ( .A(n143), .B(n149), .Z(n185) );
  IV U244 ( .A(n173), .Z(n226) );
  XOR U245 ( .A(n227), .B(n228), .Z(n173) );
  ANDN U246 ( .A(n229), .B(n230), .Z(n228) );
  XOR U247 ( .A(n227), .B(n231), .Z(n229) );
  XNOR U248 ( .A(n191), .B(n192), .Z(n177) );
  OR U249 ( .A(n232), .B(n86), .Z(n192) );
  XNOR U250 ( .A(n190), .B(n233), .Z(n191) );
  ANDN U251 ( .A(n121), .B(n186), .Z(n233) );
  ANDN U252 ( .A(n234), .B(n235), .Z(n190) );
  NANDN U253 ( .B(n236), .A(n237), .Z(n234) );
  NAND U254 ( .A(n240), .B(n241), .Z(\_MxM/n123 ) );
  NANDN U255 ( .B(n29), .A(o[0]), .Z(n241) );
  AND U256 ( .A(n242), .B(n243), .Z(n240) );
  NANDN U257 ( .B(n52), .A(o[0]), .Z(n243) );
  IV U258 ( .A(n244), .Z(n52) );
  OR U259 ( .A(n57), .B(n27), .Z(n242) );
  IV U260 ( .A(\_MxM/Y0[1] ), .Z(n33) );
  XOR U261 ( .A(n245), .B(n246), .Z(n239) );
  XNOR U262 ( .A(n247), .B(n238), .Z(n245) );
  NAND U263 ( .A(\_MxM/Y0[0] ), .B(n204), .Z(n238) );
  NAND U264 ( .A(n248), .B(n77), .Z(n247) );
  XOR U265 ( .A(e_input[7]), .B(g_input[7]), .Z(n77) );
  XNOR U266 ( .A(n205), .B(n246), .Z(n248) );
  XNOR U267 ( .A(n204), .B(n246), .Z(n205) );
  XNOR U268 ( .A(n218), .B(n217), .Z(n246) );
  XNOR U269 ( .A(n249), .B(n214), .Z(n217) );
  XNOR U270 ( .A(n250), .B(n209), .Z(n214) );
  NAND U271 ( .A(n122), .B(n213), .Z(n209) );
  NANDN U272 ( .B(n85), .A(n252), .Z(n251) );
  XNOR U273 ( .A(n215), .B(n216), .Z(n249) );
  XNOR U274 ( .A(n221), .B(n263), .Z(n224) );
  AND U275 ( .A(n149), .B(n180), .Z(n263) );
  XOR U276 ( .A(n264), .B(n265), .Z(n221) );
  ANDN U277 ( .A(n266), .B(n267), .Z(n265) );
  XNOR U278 ( .A(n268), .B(n264), .Z(n266) );
  XOR U279 ( .A(n269), .B(n225), .Z(n262) );
  NANDN U280 ( .B(n186), .A(n143), .Z(n225) );
  IV U281 ( .A(n227), .Z(n269) );
  XNOR U282 ( .A(n236), .B(n237), .Z(n231) );
  NANDN U283 ( .B(n86), .A(n273), .Z(n237) );
  ANDN U284 ( .A(n121), .B(n232), .Z(n274) );
  NAND U285 ( .A(n275), .B(n276), .Z(n235) );
  NANDN U286 ( .B(n277), .A(n278), .Z(n275) );
  XNOR U287 ( .A(n258), .B(n257), .Z(n204) );
  XNOR U288 ( .A(n279), .B(n261), .Z(n257) );
  XNOR U289 ( .A(n254), .B(n255), .Z(n261) );
  NAND U290 ( .A(n149), .B(n213), .Z(n255) );
  XNOR U291 ( .A(n253), .B(n280), .Z(n254) );
  AND U292 ( .A(n252), .B(n122), .Z(n280) );
  XOR U293 ( .A(n281), .B(n282), .Z(n253) );
  AND U294 ( .A(n283), .B(n284), .Z(n282) );
  XNOR U295 ( .A(n285), .B(n281), .Z(n284) );
  XNOR U296 ( .A(n260), .B(n256), .Z(n279) );
  XOR U297 ( .A(n286), .B(n287), .Z(n256) );
  XOR U298 ( .A(n288), .B(n289), .Z(n260) );
  AND U299 ( .A(n290), .B(n291), .Z(n289) );
  NANDN U300 ( .B(n85), .A(n292), .Z(n291) );
  NANDN U301 ( .B(n293), .A(n294), .Z(n85) );
  AND U302 ( .A(n295), .B(g_input[7]), .Z(n294) );
  NANDN U303 ( .B(n296), .A(n297), .Z(n290) );
  IV U304 ( .A(n259), .Z(n288) );
  XNOR U305 ( .A(n298), .B(n299), .Z(n259) );
  AND U306 ( .A(n300), .B(n301), .Z(n299) );
  XOR U307 ( .A(n297), .B(n302), .Z(n301) );
  XNOR U308 ( .A(n296), .B(n298), .Z(n302) );
  NAND U309 ( .A(n122), .B(n292), .Z(n296) );
  XNOR U310 ( .A(n306), .B(n303), .Z(n305) );
  XOR U311 ( .A(n283), .B(n307), .Z(n300) );
  XNOR U312 ( .A(n285), .B(n298), .Z(n307) );
  NANDN U313 ( .B(n186), .A(n213), .Z(n285) );
  XOR U314 ( .A(n281), .B(n308), .Z(n283) );
  AND U315 ( .A(n252), .B(n149), .Z(n308) );
  XOR U316 ( .A(n309), .B(n310), .Z(n281) );
  AND U317 ( .A(n311), .B(n312), .Z(n310) );
  XNOR U318 ( .A(n313), .B(n309), .Z(n312) );
  XOR U319 ( .A(n314), .B(n315), .Z(n298) );
  AND U320 ( .A(n316), .B(n317), .Z(n315) );
  XOR U321 ( .A(n304), .B(n318), .Z(n317) );
  XNOR U322 ( .A(n306), .B(n314), .Z(n318) );
  NAND U323 ( .A(n149), .B(n292), .Z(n306) );
  XOR U324 ( .A(n303), .B(n319), .Z(n304) );
  AND U325 ( .A(n122), .B(e_input[0]), .Z(n319) );
  XNOR U326 ( .A(n295), .B(g_input[6]), .Z(n293) );
  NOR U327 ( .A(n320), .B(n321), .Z(n295) );
  XNOR U328 ( .A(n325), .B(n322), .Z(n324) );
  XOR U329 ( .A(n311), .B(n326), .Z(n316) );
  XNOR U330 ( .A(n313), .B(n314), .Z(n326) );
  NANDN U331 ( .B(n232), .A(n213), .Z(n313) );
  XOR U332 ( .A(n309), .B(n327), .Z(n311) );
  ANDN U333 ( .A(n252), .B(n186), .Z(n327) );
  XOR U334 ( .A(n328), .B(n329), .Z(n309) );
  AND U335 ( .A(n330), .B(n331), .Z(n329) );
  XNOR U336 ( .A(n332), .B(n328), .Z(n331) );
  XOR U337 ( .A(n333), .B(n334), .Z(n314) );
  AND U338 ( .A(n335), .B(n336), .Z(n334) );
  XOR U339 ( .A(n323), .B(n337), .Z(n336) );
  XNOR U340 ( .A(n325), .B(n333), .Z(n337) );
  NANDN U341 ( .B(n186), .A(n292), .Z(n325) );
  XOR U342 ( .A(n322), .B(n338), .Z(n323) );
  AND U343 ( .A(n149), .B(e_input[0]), .Z(n338) );
  XOR U344 ( .A(n320), .B(g_input[5]), .Z(n321) );
  NANDN U345 ( .B(n339), .A(n340), .Z(n320) );
  XOR U346 ( .A(n341), .B(n342), .Z(n322) );
  ANDN U347 ( .A(n343), .B(n344), .Z(n342) );
  XNOR U348 ( .A(n345), .B(n341), .Z(n343) );
  XOR U349 ( .A(n330), .B(n346), .Z(n335) );
  XNOR U350 ( .A(n332), .B(n333), .Z(n346) );
  NAND U351 ( .A(n213), .B(n273), .Z(n332) );
  XOR U352 ( .A(n328), .B(n347), .Z(n330) );
  ANDN U353 ( .A(n252), .B(n232), .Z(n347) );
  XOR U354 ( .A(n348), .B(n349), .Z(n328) );
  ANDN U355 ( .A(n350), .B(n351), .Z(n349) );
  XNOR U356 ( .A(n352), .B(n348), .Z(n350) );
  XNOR U357 ( .A(n354), .B(n352), .Z(n286) );
  NAND U358 ( .A(n213), .B(n355), .Z(n352) );
  IV U359 ( .A(n351), .Z(n354) );
  XNOR U360 ( .A(n348), .B(n356), .Z(n351) );
  AND U361 ( .A(n273), .B(n252), .Z(n356) );
  AND U362 ( .A(n357), .B(g_input[0]), .Z(n348) );
  NANDN U363 ( .B(n213), .A(n358), .Z(n357) );
  NAND U364 ( .A(n355), .B(n252), .Z(n358) );
  XNOR U365 ( .A(n359), .B(e_input[2]), .Z(n252) );
  NAND U366 ( .A(n360), .B(e_input[7]), .Z(n359) );
  XOR U367 ( .A(n361), .B(e_input[2]), .Z(n360) );
  XNOR U368 ( .A(n341), .B(n364), .Z(n344) );
  ANDN U369 ( .A(e_input[0]), .B(n186), .Z(n364) );
  XOR U370 ( .A(n365), .B(n366), .Z(n341) );
  AND U371 ( .A(n367), .B(n368), .Z(n366) );
  XOR U372 ( .A(n369), .B(n365), .Z(n368) );
  ANDN U373 ( .A(e_input[0]), .B(n232), .Z(n369) );
  XOR U374 ( .A(n370), .B(n365), .Z(n367) );
  AND U375 ( .A(n292), .B(n273), .Z(n370) );
  XOR U376 ( .A(n371), .B(n372), .Z(n365) );
  ANDN U377 ( .A(n373), .B(n374), .Z(n372) );
  XNOR U378 ( .A(n375), .B(n371), .Z(n373) );
  XOR U379 ( .A(n376), .B(n345), .Z(n363) );
  NANDN U380 ( .B(n232), .A(n292), .Z(n345) );
  IV U381 ( .A(n353), .Z(n376) );
  NAND U382 ( .A(n292), .B(n355), .Z(n375) );
  XNOR U383 ( .A(n371), .B(n377), .Z(n374) );
  AND U384 ( .A(n273), .B(e_input[0]), .Z(n377) );
  AND U385 ( .A(n378), .B(g_input[0]), .Z(n371) );
  NANDN U386 ( .B(n292), .A(n379), .Z(n378) );
  NAND U387 ( .A(n355), .B(e_input[0]), .Z(n379) );
  XNOR U388 ( .A(n380), .B(e_input[1]), .Z(n292) );
  NAND U389 ( .A(n381), .B(e_input[7]), .Z(n380) );
  XNOR U390 ( .A(e_input[1]), .B(n382), .Z(n381) );
  XOR U391 ( .A(n383), .B(n384), .Z(n271) );
  IV U392 ( .A(n267), .Z(n384) );
  XNOR U393 ( .A(n264), .B(n385), .Z(n267) );
  ANDN U394 ( .A(n180), .B(n186), .Z(n385) );
  XNOR U395 ( .A(n340), .B(g_input[4]), .Z(n339) );
  NOR U396 ( .A(n386), .B(n387), .Z(n340) );
  XOR U397 ( .A(n390), .B(n388), .Z(n389) );
  ANDN U398 ( .A(n180), .B(n232), .Z(n390) );
  AND U399 ( .A(n273), .B(n143), .Z(n391) );
  XOR U400 ( .A(n395), .B(n268), .Z(n383) );
  NANDN U401 ( .B(n232), .A(n143), .Z(n268) );
  NANDN U402 ( .B(n396), .A(n397), .Z(n386) );
  IV U403 ( .A(n270), .Z(n395) );
  XOR U404 ( .A(n398), .B(n394), .Z(n270) );
  NAND U405 ( .A(n143), .B(n355), .Z(n394) );
  IV U406 ( .A(n393), .Z(n398) );
  XNOR U407 ( .A(n392), .B(n399), .Z(n393) );
  AND U408 ( .A(n273), .B(n180), .Z(n399) );
  AND U409 ( .A(n400), .B(g_input[0]), .Z(n392) );
  NANDN U410 ( .B(n143), .A(n401), .Z(n400) );
  NAND U411 ( .A(n355), .B(n180), .Z(n401) );
  XNOR U412 ( .A(n402), .B(e_input[4]), .Z(n180) );
  NAND U413 ( .A(n403), .B(e_input[7]), .Z(n402) );
  XOR U414 ( .A(n404), .B(e_input[4]), .Z(n403) );
  XNOR U415 ( .A(n405), .B(e_input[5]), .Z(n143) );
  NAND U416 ( .A(n406), .B(e_input[7]), .Z(n405) );
  XOR U417 ( .A(n407), .B(e_input[5]), .Z(n406) );
  XNOR U418 ( .A(n277), .B(n278), .Z(n272) );
  NANDN U419 ( .B(n86), .A(n355), .Z(n278) );
  XNOR U420 ( .A(n276), .B(n408), .Z(n277) );
  AND U421 ( .A(n273), .B(n121), .Z(n408) );
  XNOR U422 ( .A(n397), .B(g_input[2]), .Z(n396) );
  AND U423 ( .A(n410), .B(g_input[0]), .Z(n276) );
  NAND U424 ( .A(n411), .B(n86), .Z(n410) );
  NANDN U425 ( .B(n412), .A(n413), .Z(n86) );
  ANDN U426 ( .A(e_input[7]), .B(n414), .Z(n413) );
  NAND U427 ( .A(n355), .B(n121), .Z(n411) );
  XOR U428 ( .A(n414), .B(e_input[6]), .Z(n412) );
  OR U429 ( .A(n407), .B(n415), .Z(n414) );
  XOR U430 ( .A(n415), .B(e_input[5]), .Z(n407) );
  OR U431 ( .A(n404), .B(n416), .Z(n415) );
  XOR U432 ( .A(n416), .B(e_input[4]), .Z(n404) );
  OR U433 ( .A(n362), .B(n417), .Z(n416) );
  XOR U434 ( .A(n417), .B(e_input[3]), .Z(n362) );
  OR U435 ( .A(n361), .B(n418), .Z(n417) );
  XOR U436 ( .A(n418), .B(e_input[2]), .Z(n361) );
  NANDN U437 ( .B(e_input[0]), .A(n382), .Z(n418) );
  XNOR U438 ( .A(e_input[0]), .B(e_input[1]), .Z(n382) );
  XNOR U439 ( .A(n419), .B(g_input[1]), .Z(n355) );
  NAND U440 ( .A(n420), .B(g_input[7]), .Z(n419) );
  XOR U441 ( .A(g_input[1]), .B(n409), .Z(n420) );
  XOR U442 ( .A(g_input[0]), .B(g_input[1]), .Z(n409) );
  NANDN U443 ( .B(n244), .A(n29), .Z(n57) );
  IV U444 ( .A(rst), .Z(n29) );
  NAND U445 ( .A(n421), .B(n422), .Z(n244) );
  AND U446 ( .A(n423), .B(n424), .Z(n422) );
  ANDN U447 ( .A(n425), .B(\_MxM/n[7] ), .Z(n424) );
  NOR U448 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n425) );
  NOR U449 ( .A(\_MxM/n[5] ), .B(\_MxM/n[6] ), .Z(n423) );
  AND U450 ( .A(n426), .B(n427), .Z(n421) );
  NOR U451 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n427) );
  NOR U452 ( .A(\_MxM/n[0] ), .B(n22), .Z(n426) );
  OR U453 ( .A(\_MxM/n[3] ), .B(\_MxM/n[4] ), .Z(n22) );
endmodule

