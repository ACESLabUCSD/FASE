
module MxM_W16_N10000 ( clk, rst, A, X, Y );
  input [15:0] A;
  input [15:0] X;
  output [15:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         \add_25/carry[13] , \add_25/carry[12] , \add_25/carry[11] ,
         \add_25/carry[10] , \add_25/carry[9] , \add_25/carry[8] ,
         \add_25/carry[7] , \add_25/carry[6] , \add_25/carry[5] ,
         \add_25/carry[4] , \add_25/carry[3] , \add_25/carry[2] , n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760;
  wire   [15:0] Y0;
  wire   [13:0] n;

  DFF \n_reg[0]  ( .D(n262), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n261), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n260), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n259), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n258), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n257), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n256), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \n_reg[7]  ( .D(n255), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[7]) );
  DFF \n_reg[8]  ( .D(n254), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[8]) );
  DFF \n_reg[9]  ( .D(n253), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[9]) );
  DFF \n_reg[10]  ( .D(n252), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[10]) );
  DFF \n_reg[11]  ( .D(n251), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[11]) );
  DFF \n_reg[12]  ( .D(n250), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[12]) );
  DFF \n_reg[13]  ( .D(n249), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[13]) );
  DFF \Y0_reg[0]  ( .D(n248), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n247), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n246), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n245), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n244), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n243), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n242), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n241), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y0_reg[8]  ( .D(n240), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[8]) );
  DFF \Y0_reg[9]  ( .D(n239), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[9]) );
  DFF \Y0_reg[10]  ( .D(n238), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[10]) );
  DFF \Y0_reg[11]  ( .D(n237), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[11]) );
  DFF \Y0_reg[12]  ( .D(n236), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[12]) );
  DFF \Y0_reg[13]  ( .D(n235), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[13]) );
  DFF \Y0_reg[14]  ( .D(n234), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[14]) );
  DFF \Y0_reg[15]  ( .D(n233), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[15]) );
  DFF \Y_reg[15]  ( .D(n232), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[15]) );
  DFF \Y_reg[14]  ( .D(n231), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[14]) );
  DFF \Y_reg[13]  ( .D(n230), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[13]) );
  DFF \Y_reg[12]  ( .D(n229), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[12]) );
  DFF \Y_reg[11]  ( .D(n228), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[11]) );
  DFF \Y_reg[10]  ( .D(n227), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[10]) );
  DFF \Y_reg[9]  ( .D(n226), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[9]) );
  DFF \Y_reg[8]  ( .D(n225), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[8]) );
  DFF \Y_reg[7]  ( .D(n224), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n223), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n222), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n221), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n220), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n219), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n218), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n217), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  HADDER \add_25/U1_1_6  ( .IN0(n[6]), .IN1(\add_25/carry[6] ), .COUT(
        \add_25/carry[7] ), .SUM(N13) );
  HADDER \add_25/U1_1_7  ( .IN0(n[7]), .IN1(\add_25/carry[7] ), .COUT(
        \add_25/carry[8] ), .SUM(N14) );
  HADDER \add_25/U1_1_8  ( .IN0(n[8]), .IN1(\add_25/carry[8] ), .COUT(
        \add_25/carry[9] ), .SUM(N15) );
  HADDER \add_25/U1_1_9  ( .IN0(n[9]), .IN1(\add_25/carry[9] ), .COUT(
        \add_25/carry[10] ), .SUM(N16) );
  HADDER \add_25/U1_1_10  ( .IN0(n[10]), .IN1(\add_25/carry[10] ), .COUT(
        \add_25/carry[11] ), .SUM(N17) );
  HADDER \add_25/U1_1_11  ( .IN0(n[11]), .IN1(\add_25/carry[11] ), .COUT(
        \add_25/carry[12] ), .SUM(N18) );
  HADDER \add_25/U1_1_12  ( .IN0(n[12]), .IN1(\add_25/carry[12] ), .COUT(
        \add_25/carry[13] ), .SUM(N19) );
  MUX U265 ( .IN0(n263), .IN1(n1583), .SEL(n1584), .F(n1567) );
  IV U266 ( .A(n1585), .Z(n263) );
  MUX U267 ( .IN0(n264), .IN1(n1250), .SEL(n1251), .F(n1227) );
  IV U268 ( .A(n1252), .Z(n264) );
  MUX U269 ( .IN0(n1658), .IN1(n1676), .SEL(n1660), .F(n1639) );
  XOR U270 ( .A(n1441), .B(n1431), .Z(n1247) );
  XOR U271 ( .A(n1253), .B(n1235), .Z(n1239) );
  MUX U272 ( .IN0(n265), .IN1(n1000), .SEL(n1001), .F(n930) );
  IV U273 ( .A(n1002), .Z(n265) );
  MUX U274 ( .IN0(n266), .IN1(n1161), .SEL(n1162), .F(n1086) );
  IV U275 ( .A(n1163), .Z(n266) );
  MUX U276 ( .IN0(n267), .IN1(n1227), .SEL(n1228), .F(n1204) );
  IV U277 ( .A(n1229), .Z(n267) );
  MUX U278 ( .IN0(n268), .IN1(n1423), .SEL(n1424), .F(n1413) );
  IV U279 ( .A(n1425), .Z(n268) );
  XOR U280 ( .A(n1426), .B(n1418), .Z(n1224) );
  MUX U281 ( .IN0(n1378), .IN1(n1381), .SEL(n1379), .F(n1363) );
  MUX U282 ( .IN0(n269), .IN1(n725), .SEL(n726), .F(n674) );
  IV U283 ( .A(n727), .Z(n269) );
  MUX U284 ( .IN0(n270), .IN1(n1077), .SEL(n1078), .F(n1000) );
  IV U285 ( .A(n1079), .Z(n270) );
  XNOR U286 ( .A(n1721), .B(n1722), .Z(n1165) );
  XOR U287 ( .A(n1228), .B(n1229), .Z(n1240) );
  MUX U288 ( .IN0(n271), .IN1(n1177), .SEL(n1178), .F(n1115) );
  IV U289 ( .A(n1179), .Z(n271) );
  XOR U290 ( .A(n1414), .B(n1415), .Z(n1222) );
  MUX U291 ( .IN0(n272), .IN1(n854), .SEL(n855), .F(n789) );
  IV U292 ( .A(n856), .Z(n272) );
  MUX U293 ( .IN0(X[8]), .IN1(n1706), .SEL(X[15]), .F(n737) );
  MUX U294 ( .IN0(n1419), .IN1(n273), .SEL(n1418), .F(n1410) );
  IV U295 ( .A(n1417), .Z(n273) );
  MUX U296 ( .IN0(X[13]), .IN1(n1732), .SEL(X[15]), .F(n519) );
  MUX U297 ( .IN0(n1594), .IN1(n1597), .SEL(n1595), .F(n1578) );
  MUX U298 ( .IN0(n274), .IN1(n1204), .SEL(n1205), .F(n1185) );
  IV U299 ( .A(n1206), .Z(n274) );
  MUX U300 ( .IN0(n275), .IN1(n1413), .SEL(n1414), .F(n1192) );
  IV U301 ( .A(n1415), .Z(n275) );
  XOR U302 ( .A(n1230), .B(n1212), .Z(n1216) );
  MUX U303 ( .IN0(X[9]), .IN1(n1707), .SEL(X[15]), .F(n683) );
  MUX U304 ( .IN0(n560), .IN1(n276), .SEL(n559), .F(n521) );
  IV U305 ( .A(n558), .Z(n276) );
  MUX U306 ( .IN0(X[11]), .IN1(n1687), .SEL(X[15]), .F(n589) );
  MUX U307 ( .IN0(n650), .IN1(n648), .SEL(n649), .F(n603) );
  MUX U308 ( .IN0(n277), .IN1(n443), .SEL(n442), .F(n451) );
  IV U309 ( .A(n454), .Z(n277) );
  MUX U310 ( .IN0(n278), .IN1(n1598), .SEL(n1599), .F(n1594) );
  IV U311 ( .A(n1600), .Z(n278) );
  XOR U312 ( .A(n1424), .B(n1425), .Z(n1245) );
  MUX U313 ( .IN0(n279), .IN1(n981), .SEL(n982), .F(n912) );
  IV U314 ( .A(n983), .Z(n279) );
  MUX U315 ( .IN0(n280), .IN1(n1040), .SEL(n1041), .F(n977) );
  IV U316 ( .A(n1042), .Z(n280) );
  MUX U317 ( .IN0(X[10]), .IN1(n1686), .SEL(X[15]), .F(n630) );
  MUX U318 ( .IN0(n740), .IN1(n281), .SEL(n739), .F(n685) );
  IV U319 ( .A(n738), .Z(n281) );
  MUX U320 ( .IN0(n816), .IN1(n814), .SEL(n815), .F(n749) );
  XNOR U321 ( .A(n1708), .B(n1162), .Z(n1166) );
  XOR U322 ( .A(n452), .B(n473), .Z(n471) );
  MUX U323 ( .IN0(n1639), .IN1(n1657), .SEL(n1641), .F(n1608) );
  MUX U324 ( .IN0(n1527), .IN1(n1549), .SEL(n1529), .F(n1509) );
  MUX U325 ( .IN0(n282), .IN1(n1185), .SEL(n1186), .F(n1123) );
  IV U326 ( .A(n1187), .Z(n282) );
  MUX U327 ( .IN0(n283), .IN1(n1430), .SEL(n1431), .F(n1417) );
  IV U328 ( .A(n1432), .Z(n283) );
  MUX U329 ( .IN0(n284), .IN1(n1152), .SEL(n1153), .F(n1077) );
  IV U330 ( .A(n1154), .Z(n284) );
  MUX U331 ( .IN0(A[11]), .IN1(n1461), .SEL(A[15]), .F(n606) );
  MUX U332 ( .IN0(n688), .IN1(n289), .SEL(n687), .F(n637) );
  MUX U333 ( .IN0(n949), .IN1(n947), .SEL(n948), .F(n879) );
  MUX U334 ( .IN0(n979), .IN1(n285), .SEL(n978), .F(n907) );
  IV U335 ( .A(n977), .Z(n285) );
  NAND U336 ( .A(n521), .B(n556), .Z(n555) );
  XOR U337 ( .A(n499), .B(n507), .Z(n505) );
  MUX U338 ( .IN0(n286), .IN1(n1445), .SEL(n1446), .F(n1430) );
  IV U339 ( .A(n1447), .Z(n286) );
  MUX U340 ( .IN0(n287), .IN1(n992), .SEL(n993), .F(n922) );
  IV U341 ( .A(n994), .Z(n287) );
  MUX U342 ( .IN0(n288), .IN1(n1048), .SEL(n1049), .F(n981) );
  IV U343 ( .A(n1050), .Z(n288) );
  MUX U344 ( .IN0(X[4]), .IN1(n1392), .SEL(X[15]), .F(n976) );
  XOR U345 ( .A(n1688), .B(n1673), .Z(n1613) );
  MUX U346 ( .IN0(n732), .IN1(n734), .SEL(n733), .F(n289) );
  IV U347 ( .A(n289), .Z(n686) );
  MUX U348 ( .IN0(n910), .IN1(n290), .SEL(n909), .F(n837) );
  IV U349 ( .A(n908), .Z(n290) );
  MUX U350 ( .IN0(n1017), .IN1(n1015), .SEL(n1016), .F(n947) );
  MUX U351 ( .IN0(n1135), .IN1(n291), .SEL(n1134), .F(n1058) );
  IV U352 ( .A(n1133), .Z(n291) );
  XNOR U353 ( .A(n640), .B(n600), .Z(n604) );
  XOR U354 ( .A(n530), .B(n538), .Z(n536) );
  XOR U355 ( .A(n1205), .B(n1206), .Z(n1217) );
  MUX U356 ( .IN0(n1533), .IN1(n1543), .SEL(n1535), .F(n1519) );
  MUX U357 ( .IN0(n1608), .IN1(n1638), .SEL(n1610), .F(n1144) );
  XNOR U358 ( .A(n1385), .B(n1386), .Z(n1369) );
  MUX U359 ( .IN0(A[9]), .IN1(n1499), .SEL(A[15]), .F(n700) );
  MUX U360 ( .IN0(A[12]), .IN1(n1443), .SEL(A[15]), .F(n561) );
  XOR U361 ( .A(n609), .B(n652), .Z(n610) );
  MUX U362 ( .IN0(n1004), .IN1(n1006), .SEL(n1005), .F(n936) );
  MUX U363 ( .IN0(n1046), .IN1(n1044), .SEL(n1045), .F(n971) );
  XOR U364 ( .A(n1134), .B(n1135), .Z(n1141) );
  XNOR U365 ( .A(n637), .B(n680), .Z(n638) );
  XNOR U366 ( .A(n741), .B(n694), .Z(n698) );
  MUX U367 ( .IN0(n292), .IN1(n925), .SEL(n926), .F(n857) );
  IV U368 ( .A(n927), .Z(n292) );
  MUX U369 ( .IN0(n784), .IN1(n786), .SEL(n785), .F(n293) );
  IV U370 ( .A(n293), .Z(n720) );
  XOR U371 ( .A(n567), .B(n575), .Z(n573) );
  MUX U372 ( .IN0(n1525), .IN1(n294), .SEL(n1375), .F(n1506) );
  IV U373 ( .A(n1374), .Z(n294) );
  MUX U374 ( .IN0(n1371), .IN1(n1369), .SEL(n1370), .F(n1342) );
  XOR U375 ( .A(n1416), .B(n1410), .Z(n1201) );
  MUX U376 ( .IN0(n295), .IN1(n1144), .SEL(n1145), .F(n1069) );
  IV U377 ( .A(n1146), .Z(n295) );
  MUX U378 ( .IN0(n296), .IN1(n1192), .SEL(n1193), .F(n1133) );
  IV U379 ( .A(n1194), .Z(n296) );
  XOR U380 ( .A(n1207), .B(n1178), .Z(n1182) );
  MUX U381 ( .IN0(n868), .IN1(n870), .SEL(n869), .F(n803) );
  MUX U382 ( .IN0(n1094), .IN1(n1092), .SEL(n1093), .F(n1015) );
  XOR U383 ( .A(n1614), .B(n1153), .Z(n1157) );
  XNOR U384 ( .A(n689), .B(n645), .Z(n649) );
  MUX U385 ( .IN0(n297), .IN1(n728), .SEL(n729), .F(n677) );
  IV U386 ( .A(n730), .Z(n297) );
  MUX U387 ( .IN0(n298), .IN1(n843), .SEL(n844), .F(n783) );
  IV U388 ( .A(n845), .Z(n298) );
  NAND U389 ( .A(n907), .B(n975), .Z(n974) );
  MUX U390 ( .IN0(n849), .IN1(n851), .SEL(n850), .F(n784) );
  MUX U391 ( .IN0(n299), .IN1(n823), .SEL(n824), .F(n758) );
  IV U392 ( .A(Y0[5]), .Z(n299) );
  XOR U393 ( .A(n612), .B(n620), .Z(n618) );
  MUX U394 ( .IN0(n300), .IN1(n1578), .SEL(n1579), .F(n1561) );
  IV U395 ( .A(n1580), .Z(n300) );
  MUX U396 ( .IN0(A[1]), .IN1(n1734), .SEL(A[15]), .F(n1388) );
  MUX U397 ( .IN0(n301), .IN1(n789), .SEL(n790), .F(n725) );
  IV U398 ( .A(n791), .Z(n301) );
  MUX U399 ( .IN0(A[6]), .IN1(n1630), .SEL(A[15]), .F(n882) );
  MUX U400 ( .IN0(A[7]), .IN1(n1617), .SEL(A[15]), .F(n817) );
  MUX U401 ( .IN0(A[5]), .IN1(n1650), .SEL(A[15]), .F(n950) );
  MUX U402 ( .IN0(n302), .IN1(n1123), .SEL(n1124), .F(n1048) );
  IV U403 ( .A(n1125), .Z(n302) );
  XOR U404 ( .A(n1193), .B(n1194), .Z(n1199) );
  MUX U405 ( .IN0(n936), .IN1(n938), .SEL(n937), .F(n868) );
  XNOR U406 ( .A(n1175), .B(n1116), .Z(n1120) );
  XOR U407 ( .A(n527), .B(n562), .Z(n528) );
  MUX U408 ( .IN0(n303), .IN1(n592), .SEL(n593), .F(n545) );
  IV U409 ( .A(n594), .Z(n303) );
  NAND U410 ( .A(n685), .B(n736), .Z(n735) );
  MUX U411 ( .IN0(n839), .IN1(n837), .SEL(n838), .F(n781) );
  XNOR U412 ( .A(n871), .B(n811), .Z(n815) );
  MUX U413 ( .IN0(n304), .IN1(n1072), .SEL(n1073), .F(n995) );
  IV U414 ( .A(n1074), .Z(n304) );
  MUX U415 ( .IN0(n305), .IN1(n919), .SEL(n918), .F(n849) );
  IV U416 ( .A(n917), .Z(n305) );
  MUX U417 ( .IN0(n306), .IN1(n888), .SEL(n889), .F(n823) );
  IV U418 ( .A(Y0[4]), .Z(n306) );
  XOR U419 ( .A(n657), .B(n665), .Z(n663) );
  MUX U420 ( .IN0(n1342), .IN1(n307), .SEL(n1343), .F(n1315) );
  IV U421 ( .A(n1344), .Z(n307) );
  MUX U422 ( .IN0(n1434), .IN1(n308), .SEL(n1247), .F(n1421) );
  IV U423 ( .A(n1245), .Z(n308) );
  XNOR U424 ( .A(n1599), .B(n1600), .Z(n1586) );
  MUX U425 ( .IN0(n309), .IN1(n922), .SEL(n923), .F(n854) );
  IV U426 ( .A(n924), .Z(n309) );
  MUX U427 ( .IN0(A[3]), .IN1(n1711), .SEL(A[15]), .F(n310) );
  IV U428 ( .A(n310), .Z(n1095) );
  MUX U429 ( .IN0(A[4]), .IN1(n1668), .SEL(A[15]), .F(n311) );
  IV U430 ( .A(n311), .Z(n1018) );
  MUX U431 ( .IN0(n1181), .IN1(n312), .SEL(n1182), .F(n1119) );
  IV U432 ( .A(n1183), .Z(n312) );
  XOR U433 ( .A(n1512), .B(n1513), .Z(n1374) );
  MUX U434 ( .IN0(n605), .IN1(n603), .SEL(n604), .F(n550) );
  MUX U435 ( .IN0(n313), .IN1(n912), .SEL(n913), .F(n843) );
  IV U436 ( .A(n914), .Z(n313) );
  XOR U437 ( .A(n820), .B(n883), .Z(n821) );
  MUX U438 ( .IN0(n1081), .IN1(n1083), .SEL(n1082), .F(n1004) );
  MUX U439 ( .IN0(n1167), .IN1(n1165), .SEL(n1166), .F(n1092) );
  MUX U440 ( .IN0(n314), .IN1(n634), .SEL(n635), .F(n592) );
  IV U441 ( .A(n636), .Z(n314) );
  XOR U442 ( .A(n795), .B(n739), .Z(n733) );
  XNOR U443 ( .A(n806), .B(n746), .Z(n750) );
  MUX U444 ( .IN0(n315), .IN1(n857), .SEL(n858), .F(n792) );
  IV U445 ( .A(n859), .Z(n315) );
  XOR U446 ( .A(n970), .B(n908), .Z(n909) );
  MUX U447 ( .IN0(n1066), .IN1(n316), .SEL(n1065), .F(n987) );
  IV U448 ( .A(n1064), .Z(n316) );
  MUX U449 ( .IN0(n984), .IN1(n317), .SEL(n985), .F(n917) );
  IV U450 ( .A(n986), .Z(n317) );
  MUX U451 ( .IN0(n318), .IN1(n956), .SEL(n957), .F(n888) );
  IV U452 ( .A(Y0[3]), .Z(n318) );
  XOR U453 ( .A(n712), .B(n718), .Z(n707) );
  MUX U454 ( .IN0(n319), .IN1(n1372), .SEL(n1189), .F(n1345) );
  IV U455 ( .A(n1188), .Z(n319) );
  MUX U456 ( .IN0(n1288), .IN1(n320), .SEL(n1289), .F(n1261) );
  IV U457 ( .A(n1290), .Z(n320) );
  MUX U458 ( .IN0(X[1]), .IN1(n321), .SEL(X[15]), .F(n1405) );
  IV U459 ( .A(n1605), .Z(n321) );
  MUX U460 ( .IN0(X[6]), .IN1(n1397), .SEL(X[15]), .F(n842) );
  MUX U461 ( .IN0(X[3]), .IN1(n1591), .SEL(X[15]), .F(n1061) );
  MUX U462 ( .IN0(n1156), .IN1(n1158), .SEL(n1157), .F(n1081) );
  MUX U463 ( .IN0(X[14]), .IN1(n1737), .SEL(X[15]), .F(n488) );
  NAND U464 ( .A(n586), .B(n629), .Z(n628) );
  XOR U465 ( .A(n860), .B(n800), .Z(n804) );
  XNOR U466 ( .A(n939), .B(n876), .Z(n880) );
  MUX U467 ( .IN0(n322), .IN1(n995), .SEL(n996), .F(n925) );
  IV U468 ( .A(n997), .Z(n322) );
  XNOR U469 ( .A(n1038), .B(n978), .Z(n972) );
  MUX U470 ( .IN0(n1051), .IN1(n323), .SEL(n1052), .F(n984) );
  IV U471 ( .A(n1053), .Z(n323) );
  MUX U472 ( .IN0(n324), .IN1(n530), .SEL(n531), .F(n499) );
  IV U473 ( .A(Y0[11]), .Z(n324) );
  XOR U474 ( .A(n758), .B(n766), .Z(n764) );
  MUX U475 ( .IN0(n1506), .IN1(n325), .SEL(n1351), .F(n1487) );
  IV U476 ( .A(n1349), .Z(n325) );
  MUX U477 ( .IN0(n1561), .IN1(n1577), .SEL(n1563), .F(n1544) );
  MUX U478 ( .IN0(n1238), .IN1(n326), .SEL(n1239), .F(n1215) );
  IV U479 ( .A(n1240), .Z(n326) );
  XOR U480 ( .A(n1186), .B(n1187), .Z(n1183) );
  XOR U481 ( .A(n1584), .B(n1585), .Z(n1399) );
  MUX U482 ( .IN0(n327), .IN1(n1069), .SEL(n1070), .F(n992) );
  IV U483 ( .A(n1071), .Z(n327) );
  MUX U484 ( .IN0(A[10]), .IN1(n1479), .SEL(A[15]), .F(n651) );
  XNOR U485 ( .A(n1376), .B(n1366), .Z(n1370) );
  XOR U486 ( .A(n703), .B(n753), .Z(n704) );
  MUX U487 ( .IN0(n751), .IN1(n749), .SEL(n750), .F(n697) );
  MUX U488 ( .IN0(n973), .IN1(n971), .SEL(n972), .F(n908) );
  MUX U489 ( .IN0(A[13]), .IN1(n1429), .SEL(A[15]), .F(n524) );
  MUX U490 ( .IN0(n328), .IN1(n792), .SEL(n793), .F(n728) );
  IV U491 ( .A(n794), .Z(n328) );
  XOR U492 ( .A(n928), .B(n865), .Z(n869) );
  XNOR U493 ( .A(n1084), .B(n1012), .Z(n1016) );
  MUX U494 ( .IN0(n329), .IN1(n1147), .SEL(n1148), .F(n1072) );
  IV U495 ( .A(n1149), .Z(n329) );
  MUX U496 ( .IN0(n330), .IN1(n1136), .SEL(n1137), .F(n1064) );
  IV U497 ( .A(n1138), .Z(n330) );
  MUX U498 ( .IN0(A[14]), .IN1(n1406), .SEL(A[15]), .F(n489) );
  MUX U499 ( .IN0(n547), .IN1(n331), .SEL(n546), .F(n515) );
  IV U500 ( .A(n545), .Z(n331) );
  XNOR U501 ( .A(n849), .B(n848), .Z(n901) );
  MUX U502 ( .IN0(Y0[13]), .IN1(n332), .SEL(n453), .F(n445) );
  IV U503 ( .A(n452), .Z(n332) );
  MUX U504 ( .IN0(n333), .IN1(n612), .SEL(n613), .F(n567) );
  IV U505 ( .A(Y0[9]), .Z(n333) );
  MUX U506 ( .IN0(n334), .IN1(n1101), .SEL(n1102), .F(n1024) );
  IV U507 ( .A(Y0[1]), .Z(n334) );
  XOR U508 ( .A(n823), .B(n831), .Z(n829) );
  MUX U509 ( .IN0(n1487), .IN1(n335), .SEL(n1324), .F(n1468) );
  IV U510 ( .A(n1322), .Z(n335) );
  MUX U511 ( .IN0(n1261), .IN1(n336), .SEL(n1262), .F(n1238) );
  IV U512 ( .A(n1263), .Z(n336) );
  MUX U513 ( .IN0(n1544), .IN1(n1560), .SEL(n1546), .F(n1533) );
  MUX U514 ( .IN0(n1421), .IN1(n337), .SEL(n1224), .F(n1411) );
  IV U515 ( .A(n1222), .Z(n337) );
  MUX U516 ( .IN0(A[8]), .IN1(n1517), .SEL(A[15]), .F(n752) );
  MUX U517 ( .IN0(A[2]), .IN1(n1724), .SEL(A[15]), .F(n1168) );
  MUX U518 ( .IN0(n338), .IN1(n1115), .SEL(n1116), .F(n1040) );
  IV U519 ( .A(n1117), .Z(n338) );
  MUX U520 ( .IN0(n339), .IN1(n674), .SEL(n675), .F(n631) );
  IV U521 ( .A(n676), .Z(n339) );
  MUX U522 ( .IN0(n803), .IN1(n805), .SEL(n804), .F(n732) );
  MUX U523 ( .IN0(n881), .IN1(n879), .SEL(n880), .F(n814) );
  XOR U524 ( .A(n1098), .B(n1169), .Z(n1099) );
  MUX U525 ( .IN0(n1121), .IN1(n1119), .SEL(n1120), .F(n1044) );
  XNOR U526 ( .A(n550), .B(n551), .Z(n549) );
  MUX U527 ( .IN0(n340), .IN1(n677), .SEL(n678), .F(n634) );
  IV U528 ( .A(n679), .Z(n340) );
  XOR U529 ( .A(n844), .B(n845), .Z(n839) );
  XOR U530 ( .A(n1075), .B(n1001), .Z(n1005) );
  XNOR U531 ( .A(n1159), .B(n1089), .Z(n1093) );
  NAND U532 ( .A(n1058), .B(n1131), .Z(n1130) );
  XNOR U533 ( .A(n554), .B(n553), .Z(n547) );
  XNOR U534 ( .A(n949), .B(n948), .Z(n927) );
  MUX U535 ( .IN0(n989), .IN1(n987), .SEL(n988), .F(n341) );
  IV U536 ( .A(n341), .Z(n916) );
  MUX U537 ( .IN0(n1126), .IN1(n342), .SEL(n1127), .F(n1051) );
  IV U538 ( .A(n1128), .Z(n342) );
  MUX U539 ( .IN0(n720), .IN1(n343), .SEL(n721), .F(n671) );
  IV U540 ( .A(n722), .Z(n343) );
  MUX U541 ( .IN0(n344), .IN1(n499), .SEL(n500), .F(n452) );
  IV U542 ( .A(Y0[12]), .Z(n344) );
  MUX U543 ( .IN0(n345), .IN1(n657), .SEL(n658), .F(n612) );
  IV U544 ( .A(Y0[8]), .Z(n345) );
  XOR U545 ( .A(n888), .B(n896), .Z(n894) );
  MUX U546 ( .IN0(n1468), .IN1(n346), .SEL(n1297), .F(n1449) );
  IV U547 ( .A(n1295), .Z(n346) );
  MUX U548 ( .IN0(n347), .IN1(n1612), .SEL(n1613), .F(n1662) );
  IV U549 ( .A(n1682), .Z(n347) );
  NOR U550 ( .A(A[0]), .B(n1734), .Z(n1725) );
  XOR U551 ( .A(n1592), .B(n1579), .Z(n1400) );
  MUX U552 ( .IN0(n1411), .IN1(n348), .SEL(n1201), .F(n1139) );
  IV U553 ( .A(n1199), .Z(n348) );
  MUX U554 ( .IN0(n699), .IN1(n697), .SEL(n698), .F(n648) );
  XOR U555 ( .A(n953), .B(n1019), .Z(n954) );
  MUX U556 ( .IN0(n633), .IN1(n349), .SEL(n632), .F(n586) );
  IV U557 ( .A(n631), .Z(n349) );
  MUX U558 ( .IN0(X[7]), .IN1(n1398), .SEL(X[15]), .F(n775) );
  XNOR U559 ( .A(n1007), .B(n944), .Z(n948) );
  XOR U560 ( .A(n998), .B(n933), .Z(n937) );
  XNOR U561 ( .A(n1113), .B(n1041), .Z(n1045) );
  XNOR U562 ( .A(n1167), .B(n1166), .Z(n1149) );
  MUX U563 ( .IN0(n523), .IN1(n549), .SEL(n522), .F(n494) );
  XNOR U564 ( .A(n605), .B(n604), .Z(n594) );
  XNOR U565 ( .A(n816), .B(n815), .Z(n794) );
  XNOR U566 ( .A(n881), .B(n880), .Z(n859) );
  XNOR U567 ( .A(n987), .B(n1054), .Z(n988) );
  XNOR U568 ( .A(n730), .B(n729), .Z(n722) );
  XOR U569 ( .A(n836), .B(n777), .Z(n785) );
  XNOR U570 ( .A(n997), .B(n996), .Z(n986) );
  XNOR U571 ( .A(n1074), .B(n1073), .Z(n1053) );
  XNOR U572 ( .A(n513), .B(n512), .Z(n537) );
  MUX U573 ( .IN0(n350), .IN1(n706), .SEL(n707), .F(n657) );
  IV U574 ( .A(Y0[7]), .Z(n350) );
  MUX U575 ( .IN0(Y0[14]), .IN1(n445), .SEL(n446), .F(n435) );
  XOR U576 ( .A(n956), .B(n964), .Z(n962) );
  MUX U577 ( .IN0(n1315), .IN1(n351), .SEL(n1316), .F(n1288) );
  IV U578 ( .A(n1317), .Z(n351) );
  MUX U579 ( .IN0(n352), .IN1(n1399), .SEL(n1400), .F(n1572) );
  IV U580 ( .A(n1586), .Z(n352) );
  MUX U581 ( .IN0(n1449), .IN1(n353), .SEL(n1270), .F(n1434) );
  IV U582 ( .A(n1268), .Z(n353) );
  XOR U583 ( .A(n1710), .B(A[3]), .Z(n1711) );
  MUX U584 ( .IN0(n1215), .IN1(n354), .SEL(n1216), .F(n1181) );
  IV U585 ( .A(n1217), .Z(n354) );
  XOR U586 ( .A(n1680), .B(n1681), .Z(n1612) );
  XOR U587 ( .A(n1531), .B(n1522), .Z(n1375) );
  MUX U588 ( .IN0(X[5]), .IN1(n1393), .SEL(X[15]), .F(n905) );
  MUX U589 ( .IN0(X[2]), .IN1(n1590), .SEL(X[15]), .F(n1132) );
  XNOR U590 ( .A(n1371), .B(n1370), .Z(n1188) );
  XNOR U591 ( .A(n595), .B(n559), .Z(n553) );
  MUX U592 ( .IN0(n639), .IN1(n637), .SEL(n638), .F(n355) );
  IV U593 ( .A(n355), .Z(n591) );
  XOR U594 ( .A(n913), .B(n914), .Z(n910) );
  XOR U595 ( .A(n1150), .B(n1078), .Z(n1082) );
  MUX U596 ( .IN0(n1141), .IN1(n1401), .SEL(n1140), .F(n1063) );
  XNOR U597 ( .A(n1121), .B(n1120), .Z(n1138) );
  AND U598 ( .A(n483), .B(n460), .Z(n482) );
  XNOR U599 ( .A(n650), .B(n649), .Z(n636) );
  XNOR U600 ( .A(n699), .B(n698), .Z(n679) );
  XNOR U601 ( .A(n751), .B(n750), .Z(n730) );
  XNOR U602 ( .A(n973), .B(n972), .Z(n989) );
  XNOR U603 ( .A(n1017), .B(n1016), .Z(n997) );
  XNOR U604 ( .A(n1094), .B(n1093), .Z(n1074) );
  XNOR U605 ( .A(n1046), .B(n1045), .Z(n1066) );
  XNOR U606 ( .A(n1149), .B(n1148), .Z(n1128) );
  XNOR U607 ( .A(n514), .B(n515), .Z(n513) );
  XNOR U608 ( .A(n794), .B(n793), .Z(n786) );
  XNOR U609 ( .A(n859), .B(n858), .Z(n851) );
  XNOR U610 ( .A(n927), .B(n926), .Z(n919) );
  MUX U611 ( .IN0(n356), .IN1(n567), .SEL(n568), .F(n530) );
  IV U612 ( .A(Y0[10]), .Z(n356) );
  MUX U613 ( .IN0(n357), .IN1(n758), .SEL(n759), .F(n706) );
  IV U614 ( .A(Y0[6]), .Z(n357) );
  MUX U615 ( .IN0(n358), .IN1(n1024), .SEL(n1025), .F(n956) );
  IV U616 ( .A(Y0[2]), .Z(n358) );
  MUX U617 ( .IN0(Y0[15]), .IN1(n435), .SEL(n436), .F(n359) );
  IV U618 ( .A(n359), .Z(n432) );
  XOR U619 ( .A(n1102), .B(Y0[1]), .Z(n377) );
  ANDN U620 ( .A(n360), .B(n[0]), .Z(n262) );
  AND U621 ( .A(N8), .B(n360), .Z(n261) );
  AND U622 ( .A(N9), .B(n360), .Z(n260) );
  AND U623 ( .A(N10), .B(n360), .Z(n259) );
  AND U624 ( .A(N11), .B(n360), .Z(n258) );
  AND U625 ( .A(N12), .B(n360), .Z(n257) );
  AND U626 ( .A(N13), .B(n360), .Z(n256) );
  AND U627 ( .A(N14), .B(n360), .Z(n255) );
  AND U628 ( .A(N15), .B(n360), .Z(n254) );
  AND U629 ( .A(N16), .B(n360), .Z(n253) );
  AND U630 ( .A(N17), .B(n360), .Z(n252) );
  AND U631 ( .A(N18), .B(n360), .Z(n251) );
  AND U632 ( .A(N19), .B(n360), .Z(n250) );
  AND U633 ( .A(n360), .B(n361), .Z(n249) );
  XOR U634 ( .A(n[13]), .B(\add_25/carry[13] ), .Z(n361) );
  ANDN U635 ( .A(n362), .B(rst), .Z(n360) );
  NAND U636 ( .A(n363), .B(n364), .Z(n362) );
  AND U637 ( .A(n365), .B(n366), .Z(n364) );
  ANDN U638 ( .A(n367), .B(n368), .Z(n366) );
  NOR U639 ( .A(n369), .B(n370), .Z(n367) );
  AND U640 ( .A(n371), .B(n[13]), .Z(n365) );
  AND U641 ( .A(n[10]), .B(n[0]), .Z(n371) );
  AND U642 ( .A(n372), .B(n373), .Z(n363) );
  AND U643 ( .A(n[3]), .B(n374), .Z(n373) );
  AND U644 ( .A(n[2]), .B(n[1]), .Z(n374) );
  AND U645 ( .A(n[9]), .B(n[8]), .Z(n372) );
  NAND U646 ( .A(n375), .B(n376), .Z(n248) );
  OR U647 ( .A(n377), .B(n378), .Z(n376) );
  NANDN U648 ( .B(n379), .A(Y0[0]), .Z(n375) );
  NAND U649 ( .A(n380), .B(n381), .Z(n247) );
  NANDN U650 ( .B(n378), .A(n382), .Z(n381) );
  NANDN U651 ( .B(n383), .A(rst), .Z(n380) );
  NAND U652 ( .A(n384), .B(n385), .Z(n246) );
  NANDN U653 ( .B(n378), .A(n386), .Z(n385) );
  NANDN U654 ( .B(n379), .A(Y0[2]), .Z(n384) );
  NAND U655 ( .A(n387), .B(n388), .Z(n245) );
  NANDN U656 ( .B(n378), .A(n389), .Z(n388) );
  NANDN U657 ( .B(n379), .A(Y0[3]), .Z(n387) );
  NAND U658 ( .A(n390), .B(n391), .Z(n244) );
  NANDN U659 ( .B(n378), .A(n392), .Z(n391) );
  NANDN U660 ( .B(n379), .A(Y0[4]), .Z(n390) );
  NAND U661 ( .A(n393), .B(n394), .Z(n243) );
  NANDN U662 ( .B(n378), .A(n395), .Z(n394) );
  NANDN U663 ( .B(n379), .A(Y0[5]), .Z(n393) );
  NAND U664 ( .A(n396), .B(n397), .Z(n242) );
  NANDN U665 ( .B(n378), .A(n398), .Z(n397) );
  NANDN U666 ( .B(n379), .A(Y0[6]), .Z(n396) );
  NAND U667 ( .A(n399), .B(n400), .Z(n241) );
  NANDN U668 ( .B(n378), .A(n401), .Z(n400) );
  NANDN U669 ( .B(n379), .A(Y0[7]), .Z(n399) );
  NAND U670 ( .A(n402), .B(n403), .Z(n240) );
  NANDN U671 ( .B(n378), .A(n404), .Z(n403) );
  NANDN U672 ( .B(n379), .A(Y0[8]), .Z(n402) );
  NAND U673 ( .A(n405), .B(n406), .Z(n239) );
  NANDN U674 ( .B(n378), .A(n407), .Z(n406) );
  NANDN U675 ( .B(n379), .A(Y0[9]), .Z(n405) );
  NAND U676 ( .A(n408), .B(n409), .Z(n238) );
  NANDN U677 ( .B(n378), .A(n410), .Z(n409) );
  NANDN U678 ( .B(n379), .A(Y0[10]), .Z(n408) );
  NAND U679 ( .A(n411), .B(n412), .Z(n237) );
  NANDN U680 ( .B(n378), .A(n413), .Z(n412) );
  NANDN U681 ( .B(n379), .A(Y0[11]), .Z(n411) );
  NAND U682 ( .A(n414), .B(n415), .Z(n236) );
  NANDN U683 ( .B(n378), .A(n416), .Z(n415) );
  NANDN U684 ( .B(n379), .A(Y0[12]), .Z(n414) );
  NAND U685 ( .A(n417), .B(n418), .Z(n235) );
  NANDN U686 ( .B(n378), .A(n419), .Z(n418) );
  NANDN U687 ( .B(n379), .A(Y0[13]), .Z(n417) );
  NAND U688 ( .A(n420), .B(n421), .Z(n234) );
  OR U689 ( .A(n422), .B(n378), .Z(n421) );
  NANDN U690 ( .B(n379), .A(Y0[14]), .Z(n420) );
  NAND U691 ( .A(n423), .B(n424), .Z(n233) );
  OR U692 ( .A(n378), .B(n425), .Z(n424) );
  NANDN U693 ( .B(n426), .A(n379), .Z(n378) );
  NANDN U694 ( .B(n379), .A(Y0[15]), .Z(n423) );
  NAND U695 ( .A(n427), .B(n428), .Z(n232) );
  NANDN U696 ( .B(n379), .A(Y[15]), .Z(n428) );
  AND U697 ( .A(n429), .B(n430), .Z(n427) );
  NANDN U698 ( .B(n426), .A(Y[15]), .Z(n430) );
  OR U699 ( .A(n425), .B(n431), .Z(n429) );
  XOR U700 ( .A(n432), .B(n433), .Z(n425) );
  XNOR U701 ( .A(Y0[15]), .B(n434), .Z(n433) );
  NAND U702 ( .A(n437), .B(n438), .Z(n231) );
  NANDN U703 ( .B(n379), .A(Y[14]), .Z(n438) );
  AND U704 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U705 ( .B(n426), .A(Y[14]), .Z(n440) );
  OR U706 ( .A(n422), .B(n431), .Z(n439) );
  XOR U707 ( .A(n436), .B(Y0[15]), .Z(n422) );
  XOR U708 ( .A(n435), .B(n434), .Z(n436) );
  NAND U709 ( .A(n441), .B(n442), .Z(n434) );
  OR U710 ( .A(n443), .B(n444), .Z(n441) );
  NAND U711 ( .A(n447), .B(n448), .Z(n230) );
  NANDN U712 ( .B(n379), .A(Y[13]), .Z(n448) );
  AND U713 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U714 ( .B(n426), .A(Y[13]), .Z(n450) );
  NANDN U715 ( .B(n431), .A(n419), .Z(n449) );
  XNOR U716 ( .A(n446), .B(Y0[14]), .Z(n419) );
  XNOR U717 ( .A(n451), .B(n445), .Z(n446) );
  XNOR U718 ( .A(n444), .B(n454), .Z(n443) );
  OR U719 ( .A(n455), .B(n456), .Z(n444) );
  AND U720 ( .A(n457), .B(n458), .Z(n454) );
  OR U721 ( .A(n459), .B(n460), .Z(n458) );
  AND U722 ( .A(n461), .B(n462), .Z(n457) );
  OR U723 ( .A(n463), .B(n464), .Z(n462) );
  OR U724 ( .A(n465), .B(n466), .Z(n461) );
  NAND U725 ( .A(n467), .B(n468), .Z(n229) );
  NANDN U726 ( .B(n379), .A(Y[12]), .Z(n468) );
  AND U727 ( .A(n469), .B(n470), .Z(n467) );
  NANDN U728 ( .B(n426), .A(Y[12]), .Z(n470) );
  NANDN U729 ( .B(n431), .A(n416), .Z(n469) );
  XNOR U730 ( .A(n453), .B(Y0[13]), .Z(n416) );
  XNOR U731 ( .A(n471), .B(n472), .Z(n453) );
  AND U732 ( .A(n442), .B(n474), .Z(n473) );
  XOR U733 ( .A(n455), .B(n475), .Z(n474) );
  XOR U734 ( .A(n475), .B(n456), .Z(n455) );
  OR U735 ( .A(n476), .B(n477), .Z(n456) );
  IV U736 ( .A(n472), .Z(n475) );
  XNOR U737 ( .A(n466), .B(n465), .Z(n472) );
  OR U738 ( .A(n478), .B(n479), .Z(n465) );
  AND U739 ( .A(n480), .B(n481), .Z(n466) );
  XNOR U740 ( .A(n459), .B(n482), .Z(n481) );
  NAND U741 ( .A(n484), .B(n485), .Z(n460) );
  NANDN U742 ( .B(n486), .A(n487), .Z(n484) );
  NANDN U743 ( .B(n463), .A(n488), .Z(n483) );
  NANDN U744 ( .B(n464), .A(n489), .Z(n459) );
  AND U745 ( .A(n490), .B(n491), .Z(n480) );
  OR U746 ( .A(n492), .B(n493), .Z(n491) );
  XNOR U747 ( .A(n494), .B(n495), .Z(n490) );
  ANDN U748 ( .A(n496), .B(n497), .Z(n495) );
  XOR U749 ( .A(n494), .B(n498), .Z(n496) );
  NAND U750 ( .A(n501), .B(n502), .Z(n228) );
  NANDN U751 ( .B(n379), .A(Y[11]), .Z(n502) );
  AND U752 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U753 ( .B(n426), .A(Y[11]), .Z(n504) );
  NANDN U754 ( .B(n431), .A(n413), .Z(n503) );
  XNOR U755 ( .A(n500), .B(Y0[12]), .Z(n413) );
  XNOR U756 ( .A(n505), .B(n506), .Z(n500) );
  AND U757 ( .A(n442), .B(n508), .Z(n507) );
  XOR U758 ( .A(n476), .B(n509), .Z(n508) );
  XOR U759 ( .A(n509), .B(n477), .Z(n476) );
  OR U760 ( .A(n510), .B(n511), .Z(n477) );
  IV U761 ( .A(n506), .Z(n509) );
  XNOR U762 ( .A(n479), .B(n478), .Z(n506) );
  OR U763 ( .A(n512), .B(n513), .Z(n478) );
  XNOR U764 ( .A(n493), .B(n492), .Z(n479) );
  OR U765 ( .A(n514), .B(n515), .Z(n492) );
  XOR U766 ( .A(n498), .B(n497), .Z(n493) );
  XOR U767 ( .A(n494), .B(n516), .Z(n497) );
  AND U768 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U769 ( .B(n463), .A(n519), .Z(n518) );
  OR U770 ( .A(n520), .B(n521), .Z(n517) );
  XOR U771 ( .A(n486), .B(n487), .Z(n498) );
  NANDN U772 ( .B(n464), .A(n524), .Z(n487) );
  XNOR U773 ( .A(n485), .B(n525), .Z(n486) );
  AND U774 ( .A(n489), .B(n488), .Z(n525) );
  ANDN U775 ( .A(n526), .B(n527), .Z(n485) );
  NANDN U776 ( .B(n528), .A(n529), .Z(n526) );
  NAND U777 ( .A(n532), .B(n533), .Z(n227) );
  NANDN U778 ( .B(n379), .A(Y[10]), .Z(n533) );
  AND U779 ( .A(n534), .B(n535), .Z(n532) );
  NANDN U780 ( .B(n426), .A(Y[10]), .Z(n535) );
  NANDN U781 ( .B(n431), .A(n410), .Z(n534) );
  XNOR U782 ( .A(n531), .B(Y0[11]), .Z(n410) );
  XNOR U783 ( .A(n536), .B(n537), .Z(n531) );
  AND U784 ( .A(n442), .B(n539), .Z(n538) );
  XOR U785 ( .A(n510), .B(n540), .Z(n539) );
  XOR U786 ( .A(n540), .B(n511), .Z(n510) );
  OR U787 ( .A(n541), .B(n542), .Z(n511) );
  IV U788 ( .A(n537), .Z(n540) );
  OR U789 ( .A(n543), .B(n544), .Z(n512) );
  XOR U790 ( .A(n523), .B(n522), .Z(n514) );
  XNOR U791 ( .A(n548), .B(n549), .Z(n522) );
  ANDN U792 ( .A(n552), .B(n553), .Z(n551) );
  XOR U793 ( .A(n550), .B(n554), .Z(n552) );
  XNOR U794 ( .A(n555), .B(n520), .Z(n548) );
  NAND U795 ( .A(n519), .B(n489), .Z(n520) );
  NANDN U796 ( .B(n463), .A(n557), .Z(n556) );
  XOR U797 ( .A(n528), .B(n529), .Z(n523) );
  NANDN U798 ( .B(n464), .A(n561), .Z(n529) );
  AND U799 ( .A(n524), .B(n488), .Z(n562) );
  NAND U800 ( .A(n563), .B(n564), .Z(n527) );
  NANDN U801 ( .B(n565), .A(n566), .Z(n563) );
  NAND U802 ( .A(n569), .B(n570), .Z(n226) );
  NANDN U803 ( .B(n379), .A(Y[9]), .Z(n570) );
  AND U804 ( .A(n571), .B(n572), .Z(n569) );
  NANDN U805 ( .B(n426), .A(Y[9]), .Z(n572) );
  NANDN U806 ( .B(n431), .A(n407), .Z(n571) );
  XNOR U807 ( .A(n568), .B(Y0[10]), .Z(n407) );
  XNOR U808 ( .A(n573), .B(n574), .Z(n568) );
  AND U809 ( .A(n442), .B(n576), .Z(n575) );
  XOR U810 ( .A(n541), .B(n577), .Z(n576) );
  XOR U811 ( .A(n577), .B(n542), .Z(n541) );
  OR U812 ( .A(n578), .B(n579), .Z(n542) );
  IV U813 ( .A(n574), .Z(n577) );
  XNOR U814 ( .A(n544), .B(n543), .Z(n574) );
  OR U815 ( .A(n580), .B(n581), .Z(n543) );
  XNOR U816 ( .A(n547), .B(n546), .Z(n544) );
  XOR U817 ( .A(n545), .B(n582), .Z(n546) );
  AND U818 ( .A(n583), .B(n584), .Z(n582) );
  OR U819 ( .A(n585), .B(n586), .Z(n584) );
  AND U820 ( .A(n587), .B(n588), .Z(n583) );
  NANDN U821 ( .B(n463), .A(n589), .Z(n588) );
  NAND U822 ( .A(n590), .B(n591), .Z(n587) );
  XNOR U823 ( .A(n558), .B(n596), .Z(n559) );
  AND U824 ( .A(n489), .B(n557), .Z(n596) );
  XOR U825 ( .A(n597), .B(n598), .Z(n558) );
  ANDN U826 ( .A(n599), .B(n600), .Z(n598) );
  XNOR U827 ( .A(n601), .B(n597), .Z(n599) );
  XOR U828 ( .A(n602), .B(n560), .Z(n595) );
  NAND U829 ( .A(n519), .B(n524), .Z(n560) );
  IV U830 ( .A(n550), .Z(n602) );
  XNOR U831 ( .A(n565), .B(n566), .Z(n554) );
  NANDN U832 ( .B(n464), .A(n606), .Z(n566) );
  XNOR U833 ( .A(n564), .B(n607), .Z(n565) );
  AND U834 ( .A(n561), .B(n488), .Z(n607) );
  ANDN U835 ( .A(n608), .B(n609), .Z(n564) );
  NANDN U836 ( .B(n610), .A(n611), .Z(n608) );
  NAND U837 ( .A(n614), .B(n615), .Z(n225) );
  NANDN U838 ( .B(n379), .A(Y[8]), .Z(n615) );
  AND U839 ( .A(n616), .B(n617), .Z(n614) );
  NANDN U840 ( .B(n426), .A(Y[8]), .Z(n617) );
  NANDN U841 ( .B(n431), .A(n404), .Z(n616) );
  XNOR U842 ( .A(n613), .B(Y0[9]), .Z(n404) );
  XNOR U843 ( .A(n618), .B(n619), .Z(n613) );
  AND U844 ( .A(n442), .B(n621), .Z(n620) );
  XOR U845 ( .A(n578), .B(n622), .Z(n621) );
  XOR U846 ( .A(n622), .B(n579), .Z(n578) );
  OR U847 ( .A(n623), .B(n624), .Z(n579) );
  IV U848 ( .A(n619), .Z(n622) );
  XNOR U849 ( .A(n581), .B(n580), .Z(n619) );
  OR U850 ( .A(n625), .B(n626), .Z(n580) );
  XNOR U851 ( .A(n594), .B(n593), .Z(n581) );
  XOR U852 ( .A(n627), .B(n590), .Z(n593) );
  XNOR U853 ( .A(n628), .B(n585), .Z(n590) );
  NAND U854 ( .A(n589), .B(n489), .Z(n585) );
  NANDN U855 ( .B(n463), .A(n630), .Z(n629) );
  XNOR U856 ( .A(n591), .B(n592), .Z(n627) );
  XNOR U857 ( .A(n597), .B(n641), .Z(n600) );
  AND U858 ( .A(n524), .B(n557), .Z(n641) );
  XOR U859 ( .A(n642), .B(n643), .Z(n597) );
  ANDN U860 ( .A(n644), .B(n645), .Z(n643) );
  XNOR U861 ( .A(n646), .B(n642), .Z(n644) );
  XOR U862 ( .A(n647), .B(n601), .Z(n640) );
  NAND U863 ( .A(n519), .B(n561), .Z(n601) );
  IV U864 ( .A(n603), .Z(n647) );
  XNOR U865 ( .A(n610), .B(n611), .Z(n605) );
  NANDN U866 ( .B(n464), .A(n651), .Z(n611) );
  AND U867 ( .A(n606), .B(n488), .Z(n652) );
  NAND U868 ( .A(n653), .B(n654), .Z(n609) );
  NANDN U869 ( .B(n655), .A(n656), .Z(n653) );
  NAND U870 ( .A(n659), .B(n660), .Z(n224) );
  NANDN U871 ( .B(n379), .A(Y[7]), .Z(n660) );
  AND U872 ( .A(n661), .B(n662), .Z(n659) );
  NANDN U873 ( .B(n426), .A(Y[7]), .Z(n662) );
  NANDN U874 ( .B(n431), .A(n401), .Z(n661) );
  XNOR U875 ( .A(n658), .B(Y0[8]), .Z(n401) );
  XNOR U876 ( .A(n663), .B(n664), .Z(n658) );
  AND U877 ( .A(n442), .B(n666), .Z(n665) );
  XOR U878 ( .A(n623), .B(n667), .Z(n666) );
  XOR U879 ( .A(n667), .B(n624), .Z(n623) );
  OR U880 ( .A(n668), .B(n669), .Z(n624) );
  IV U881 ( .A(n664), .Z(n667) );
  XNOR U882 ( .A(n626), .B(n625), .Z(n664) );
  NANDN U883 ( .B(n670), .A(n671), .Z(n625) );
  XNOR U884 ( .A(n636), .B(n635), .Z(n626) );
  XOR U885 ( .A(n672), .B(n639), .Z(n635) );
  XNOR U886 ( .A(n632), .B(n633), .Z(n639) );
  NAND U887 ( .A(n589), .B(n524), .Z(n633) );
  XNOR U888 ( .A(n631), .B(n673), .Z(n632) );
  AND U889 ( .A(n489), .B(n630), .Z(n673) );
  XNOR U890 ( .A(n638), .B(n634), .Z(n672) );
  AND U891 ( .A(n681), .B(n682), .Z(n680) );
  NANDN U892 ( .B(n463), .A(n683), .Z(n682) );
  OR U893 ( .A(n684), .B(n685), .Z(n681) );
  XNOR U894 ( .A(n642), .B(n690), .Z(n645) );
  AND U895 ( .A(n561), .B(n557), .Z(n690) );
  XOR U896 ( .A(n691), .B(n692), .Z(n642) );
  ANDN U897 ( .A(n693), .B(n694), .Z(n692) );
  XNOR U898 ( .A(n695), .B(n691), .Z(n693) );
  XOR U899 ( .A(n696), .B(n646), .Z(n689) );
  NAND U900 ( .A(n519), .B(n606), .Z(n646) );
  IV U901 ( .A(n648), .Z(n696) );
  XNOR U902 ( .A(n655), .B(n656), .Z(n650) );
  NANDN U903 ( .B(n464), .A(n700), .Z(n656) );
  XNOR U904 ( .A(n654), .B(n701), .Z(n655) );
  AND U905 ( .A(n651), .B(n488), .Z(n701) );
  ANDN U906 ( .A(n702), .B(n703), .Z(n654) );
  NANDN U907 ( .B(n704), .A(n705), .Z(n702) );
  NAND U908 ( .A(n708), .B(n709), .Z(n223) );
  NANDN U909 ( .B(n379), .A(Y[6]), .Z(n709) );
  AND U910 ( .A(n710), .B(n711), .Z(n708) );
  NANDN U911 ( .B(n426), .A(Y[6]), .Z(n711) );
  NANDN U912 ( .B(n431), .A(n398), .Z(n710) );
  XNOR U913 ( .A(n707), .B(Y0[7]), .Z(n398) );
  XNOR U914 ( .A(n713), .B(n714), .Z(n712) );
  AND U915 ( .A(n442), .B(n715), .Z(n714) );
  XOR U916 ( .A(n668), .B(n718), .Z(n715) );
  XOR U917 ( .A(n718), .B(n669), .Z(n668) );
  OR U918 ( .A(n716), .B(n717), .Z(n669) );
  XNOR U919 ( .A(n670), .B(n671), .Z(n718) );
  XNOR U920 ( .A(n679), .B(n678), .Z(n670) );
  XOR U921 ( .A(n723), .B(n688), .Z(n678) );
  XNOR U922 ( .A(n675), .B(n676), .Z(n688) );
  NAND U923 ( .A(n589), .B(n561), .Z(n676) );
  XNOR U924 ( .A(n674), .B(n724), .Z(n675) );
  AND U925 ( .A(n524), .B(n630), .Z(n724) );
  XNOR U926 ( .A(n687), .B(n677), .Z(n723) );
  XNOR U927 ( .A(n731), .B(n686), .Z(n687) );
  XNOR U928 ( .A(n735), .B(n684), .Z(n731) );
  NAND U929 ( .A(n683), .B(n489), .Z(n684) );
  NANDN U930 ( .B(n463), .A(n737), .Z(n736) );
  XNOR U931 ( .A(n691), .B(n742), .Z(n694) );
  AND U932 ( .A(n606), .B(n557), .Z(n742) );
  XOR U933 ( .A(n743), .B(n744), .Z(n691) );
  ANDN U934 ( .A(n745), .B(n746), .Z(n744) );
  XNOR U935 ( .A(n747), .B(n743), .Z(n745) );
  XOR U936 ( .A(n748), .B(n695), .Z(n741) );
  NAND U937 ( .A(n519), .B(n651), .Z(n695) );
  IV U938 ( .A(n697), .Z(n748) );
  XNOR U939 ( .A(n704), .B(n705), .Z(n699) );
  NANDN U940 ( .B(n464), .A(n752), .Z(n705) );
  AND U941 ( .A(n700), .B(n488), .Z(n753) );
  NAND U942 ( .A(n754), .B(n755), .Z(n703) );
  NANDN U943 ( .B(n756), .A(n757), .Z(n754) );
  IV U944 ( .A(n706), .Z(n713) );
  NAND U945 ( .A(n760), .B(n761), .Z(n222) );
  NANDN U946 ( .B(n379), .A(Y[5]), .Z(n761) );
  AND U947 ( .A(n762), .B(n763), .Z(n760) );
  NANDN U948 ( .B(n426), .A(Y[5]), .Z(n763) );
  NANDN U949 ( .B(n431), .A(n395), .Z(n762) );
  XNOR U950 ( .A(n759), .B(Y0[6]), .Z(n395) );
  XNOR U951 ( .A(n764), .B(n765), .Z(n759) );
  AND U952 ( .A(n442), .B(n767), .Z(n766) );
  XOR U953 ( .A(n716), .B(n768), .Z(n767) );
  XOR U954 ( .A(n768), .B(n717), .Z(n716) );
  OR U955 ( .A(n769), .B(n770), .Z(n717) );
  IV U956 ( .A(n765), .Z(n768) );
  XOR U957 ( .A(n722), .B(n721), .Z(n765) );
  XNOR U958 ( .A(n720), .B(n771), .Z(n721) );
  AND U959 ( .A(n719), .B(n772), .Z(n771) );
  AND U960 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U961 ( .B(n463), .A(n775), .Z(n774) );
  OR U962 ( .A(n776), .B(n777), .Z(n773) );
  AND U963 ( .A(n778), .B(n779), .Z(n719) );
  NANDN U964 ( .B(n780), .A(n781), .Z(n779) );
  NANDN U965 ( .B(n782), .A(n783), .Z(n778) );
  XNOR U966 ( .A(n787), .B(n734), .Z(n729) );
  XNOR U967 ( .A(n726), .B(n727), .Z(n734) );
  NAND U968 ( .A(n589), .B(n606), .Z(n727) );
  XNOR U969 ( .A(n725), .B(n788), .Z(n726) );
  AND U970 ( .A(n561), .B(n630), .Z(n788) );
  XNOR U971 ( .A(n733), .B(n728), .Z(n787) );
  XNOR U972 ( .A(n738), .B(n796), .Z(n739) );
  AND U973 ( .A(n489), .B(n737), .Z(n796) );
  XOR U974 ( .A(n797), .B(n798), .Z(n738) );
  ANDN U975 ( .A(n799), .B(n800), .Z(n798) );
  XNOR U976 ( .A(n801), .B(n797), .Z(n799) );
  XOR U977 ( .A(n802), .B(n740), .Z(n795) );
  NAND U978 ( .A(n683), .B(n524), .Z(n740) );
  IV U979 ( .A(n732), .Z(n802) );
  XNOR U980 ( .A(n743), .B(n807), .Z(n746) );
  AND U981 ( .A(n651), .B(n557), .Z(n807) );
  XOR U982 ( .A(n808), .B(n809), .Z(n743) );
  ANDN U983 ( .A(n810), .B(n811), .Z(n809) );
  XNOR U984 ( .A(n812), .B(n808), .Z(n810) );
  XOR U985 ( .A(n813), .B(n747), .Z(n806) );
  NAND U986 ( .A(n519), .B(n700), .Z(n747) );
  IV U987 ( .A(n749), .Z(n813) );
  XNOR U988 ( .A(n756), .B(n757), .Z(n751) );
  NANDN U989 ( .B(n464), .A(n817), .Z(n757) );
  XNOR U990 ( .A(n755), .B(n818), .Z(n756) );
  AND U991 ( .A(n752), .B(n488), .Z(n818) );
  ANDN U992 ( .A(n819), .B(n820), .Z(n755) );
  NANDN U993 ( .B(n821), .A(n822), .Z(n819) );
  NAND U994 ( .A(n825), .B(n826), .Z(n221) );
  NANDN U995 ( .B(n379), .A(Y[4]), .Z(n826) );
  AND U996 ( .A(n827), .B(n828), .Z(n825) );
  NANDN U997 ( .B(n426), .A(Y[4]), .Z(n828) );
  NANDN U998 ( .B(n431), .A(n392), .Z(n827) );
  XNOR U999 ( .A(n824), .B(Y0[5]), .Z(n392) );
  XNOR U1000 ( .A(n829), .B(n830), .Z(n824) );
  AND U1001 ( .A(n442), .B(n832), .Z(n831) );
  XOR U1002 ( .A(n769), .B(n833), .Z(n832) );
  XOR U1003 ( .A(n833), .B(n770), .Z(n769) );
  OR U1004 ( .A(n834), .B(n835), .Z(n770) );
  IV U1005 ( .A(n830), .Z(n833) );
  XOR U1006 ( .A(n786), .B(n785), .Z(n830) );
  XOR U1007 ( .A(n780), .B(n781), .Z(n777) );
  XOR U1008 ( .A(n840), .B(n782), .Z(n780) );
  NAND U1009 ( .A(n489), .B(n775), .Z(n782) );
  NANDN U1010 ( .B(n783), .A(n841), .Z(n840) );
  NANDN U1011 ( .B(n463), .A(n842), .Z(n841) );
  XOR U1012 ( .A(n846), .B(n776), .Z(n836) );
  OR U1013 ( .A(n847), .B(n848), .Z(n776) );
  IV U1014 ( .A(n784), .Z(n846) );
  XNOR U1015 ( .A(n852), .B(n805), .Z(n793) );
  XNOR U1016 ( .A(n790), .B(n791), .Z(n805) );
  NAND U1017 ( .A(n589), .B(n651), .Z(n791) );
  XNOR U1018 ( .A(n789), .B(n853), .Z(n790) );
  AND U1019 ( .A(n606), .B(n630), .Z(n853) );
  XNOR U1020 ( .A(n804), .B(n792), .Z(n852) );
  XNOR U1021 ( .A(n797), .B(n861), .Z(n800) );
  AND U1022 ( .A(n524), .B(n737), .Z(n861) );
  XOR U1023 ( .A(n862), .B(n863), .Z(n797) );
  ANDN U1024 ( .A(n864), .B(n865), .Z(n863) );
  XNOR U1025 ( .A(n866), .B(n862), .Z(n864) );
  XOR U1026 ( .A(n867), .B(n801), .Z(n860) );
  NAND U1027 ( .A(n683), .B(n561), .Z(n801) );
  IV U1028 ( .A(n803), .Z(n867) );
  XNOR U1029 ( .A(n808), .B(n872), .Z(n811) );
  AND U1030 ( .A(n700), .B(n557), .Z(n872) );
  XOR U1031 ( .A(n873), .B(n874), .Z(n808) );
  ANDN U1032 ( .A(n875), .B(n876), .Z(n874) );
  XNOR U1033 ( .A(n877), .B(n873), .Z(n875) );
  XOR U1034 ( .A(n878), .B(n812), .Z(n871) );
  NAND U1035 ( .A(n519), .B(n752), .Z(n812) );
  IV U1036 ( .A(n814), .Z(n878) );
  XNOR U1037 ( .A(n821), .B(n822), .Z(n816) );
  NANDN U1038 ( .B(n464), .A(n882), .Z(n822) );
  AND U1039 ( .A(n817), .B(n488), .Z(n883) );
  NAND U1040 ( .A(n884), .B(n885), .Z(n820) );
  NANDN U1041 ( .B(n886), .A(n887), .Z(n884) );
  NAND U1042 ( .A(n890), .B(n891), .Z(n220) );
  NANDN U1043 ( .B(n379), .A(Y[3]), .Z(n891) );
  AND U1044 ( .A(n892), .B(n893), .Z(n890) );
  NANDN U1045 ( .B(n426), .A(Y[3]), .Z(n893) );
  NANDN U1046 ( .B(n431), .A(n389), .Z(n892) );
  XNOR U1047 ( .A(n889), .B(Y0[4]), .Z(n389) );
  XNOR U1048 ( .A(n894), .B(n895), .Z(n889) );
  AND U1049 ( .A(n442), .B(n897), .Z(n896) );
  XOR U1050 ( .A(n834), .B(n898), .Z(n897) );
  XOR U1051 ( .A(n898), .B(n835), .Z(n834) );
  OR U1052 ( .A(n899), .B(n900), .Z(n835) );
  IV U1053 ( .A(n895), .Z(n898) );
  XOR U1054 ( .A(n851), .B(n850), .Z(n895) );
  XOR U1055 ( .A(n901), .B(n847), .Z(n850) );
  XOR U1056 ( .A(n839), .B(n838), .Z(n847) );
  XOR U1057 ( .A(n837), .B(n902), .Z(n838) );
  AND U1058 ( .A(n903), .B(n904), .Z(n902) );
  NANDN U1059 ( .B(n463), .A(n905), .Z(n904) );
  OR U1060 ( .A(n906), .B(n907), .Z(n903) );
  NAND U1061 ( .A(n524), .B(n775), .Z(n845) );
  XNOR U1062 ( .A(n843), .B(n911), .Z(n844) );
  AND U1063 ( .A(n842), .B(n489), .Z(n911) );
  NANDN U1064 ( .B(n915), .A(n916), .Z(n848) );
  XNOR U1065 ( .A(n920), .B(n870), .Z(n858) );
  XNOR U1066 ( .A(n855), .B(n856), .Z(n870) );
  NAND U1067 ( .A(n589), .B(n700), .Z(n856) );
  XNOR U1068 ( .A(n854), .B(n921), .Z(n855) );
  AND U1069 ( .A(n651), .B(n630), .Z(n921) );
  XNOR U1070 ( .A(n869), .B(n857), .Z(n920) );
  XNOR U1071 ( .A(n862), .B(n929), .Z(n865) );
  AND U1072 ( .A(n561), .B(n737), .Z(n929) );
  XOR U1073 ( .A(n930), .B(n931), .Z(n862) );
  ANDN U1074 ( .A(n932), .B(n933), .Z(n931) );
  XNOR U1075 ( .A(n934), .B(n930), .Z(n932) );
  XOR U1076 ( .A(n935), .B(n866), .Z(n928) );
  NAND U1077 ( .A(n683), .B(n606), .Z(n866) );
  IV U1078 ( .A(n868), .Z(n935) );
  XNOR U1079 ( .A(n873), .B(n940), .Z(n876) );
  AND U1080 ( .A(n752), .B(n557), .Z(n940) );
  XOR U1081 ( .A(n941), .B(n942), .Z(n873) );
  ANDN U1082 ( .A(n943), .B(n944), .Z(n942) );
  XNOR U1083 ( .A(n945), .B(n941), .Z(n943) );
  XOR U1084 ( .A(n946), .B(n877), .Z(n939) );
  NAND U1085 ( .A(n519), .B(n817), .Z(n877) );
  IV U1086 ( .A(n879), .Z(n946) );
  XNOR U1087 ( .A(n886), .B(n887), .Z(n881) );
  NANDN U1088 ( .B(n464), .A(n950), .Z(n887) );
  XNOR U1089 ( .A(n885), .B(n951), .Z(n886) );
  AND U1090 ( .A(n882), .B(n488), .Z(n951) );
  ANDN U1091 ( .A(n952), .B(n953), .Z(n885) );
  NANDN U1092 ( .B(n954), .A(n955), .Z(n952) );
  NAND U1093 ( .A(n958), .B(n959), .Z(n219) );
  NANDN U1094 ( .B(n379), .A(Y[2]), .Z(n959) );
  AND U1095 ( .A(n960), .B(n961), .Z(n958) );
  NANDN U1096 ( .B(n426), .A(Y[2]), .Z(n961) );
  NANDN U1097 ( .B(n431), .A(n386), .Z(n960) );
  XNOR U1098 ( .A(n957), .B(Y0[3]), .Z(n386) );
  XNOR U1099 ( .A(n962), .B(n963), .Z(n957) );
  AND U1100 ( .A(n442), .B(n965), .Z(n964) );
  XOR U1101 ( .A(n899), .B(n966), .Z(n965) );
  XOR U1102 ( .A(n966), .B(n900), .Z(n899) );
  OR U1103 ( .A(n967), .B(n968), .Z(n900) );
  IV U1104 ( .A(n963), .Z(n966) );
  XOR U1105 ( .A(n919), .B(n918), .Z(n963) );
  XOR U1106 ( .A(n969), .B(n915), .Z(n918) );
  XOR U1107 ( .A(n910), .B(n909), .Z(n915) );
  XNOR U1108 ( .A(n974), .B(n906), .Z(n970) );
  NAND U1109 ( .A(n489), .B(n905), .Z(n906) );
  NANDN U1110 ( .B(n463), .A(n976), .Z(n975) );
  NAND U1111 ( .A(n561), .B(n775), .Z(n914) );
  XNOR U1112 ( .A(n912), .B(n980), .Z(n913) );
  AND U1113 ( .A(n842), .B(n524), .Z(n980) );
  XNOR U1114 ( .A(n916), .B(n917), .Z(n969) );
  XNOR U1115 ( .A(n990), .B(n938), .Z(n926) );
  XNOR U1116 ( .A(n923), .B(n924), .Z(n938) );
  NAND U1117 ( .A(n589), .B(n752), .Z(n924) );
  XNOR U1118 ( .A(n922), .B(n991), .Z(n923) );
  AND U1119 ( .A(n700), .B(n630), .Z(n991) );
  XNOR U1120 ( .A(n937), .B(n925), .Z(n990) );
  XNOR U1121 ( .A(n930), .B(n999), .Z(n933) );
  AND U1122 ( .A(n606), .B(n737), .Z(n999) );
  XOR U1123 ( .A(n1003), .B(n934), .Z(n998) );
  NAND U1124 ( .A(n683), .B(n651), .Z(n934) );
  IV U1125 ( .A(n936), .Z(n1003) );
  XNOR U1126 ( .A(n941), .B(n1008), .Z(n944) );
  AND U1127 ( .A(n817), .B(n557), .Z(n1008) );
  XOR U1128 ( .A(n1009), .B(n1010), .Z(n941) );
  ANDN U1129 ( .A(n1011), .B(n1012), .Z(n1010) );
  XNOR U1130 ( .A(n1013), .B(n1009), .Z(n1011) );
  XOR U1131 ( .A(n1014), .B(n945), .Z(n1007) );
  NAND U1132 ( .A(n519), .B(n882), .Z(n945) );
  IV U1133 ( .A(n947), .Z(n1014) );
  XNOR U1134 ( .A(n954), .B(n955), .Z(n949) );
  OR U1135 ( .A(n1018), .B(n464), .Z(n955) );
  AND U1136 ( .A(n950), .B(n488), .Z(n1019) );
  NAND U1137 ( .A(n1020), .B(n1021), .Z(n953) );
  NANDN U1138 ( .B(n1022), .A(n1023), .Z(n1020) );
  NAND U1139 ( .A(n1026), .B(n1027), .Z(n218) );
  NANDN U1140 ( .B(n379), .A(Y[1]), .Z(n1027) );
  AND U1141 ( .A(n1028), .B(n1029), .Z(n1026) );
  NANDN U1142 ( .B(n426), .A(Y[1]), .Z(n1029) );
  NANDN U1143 ( .B(n431), .A(n382), .Z(n1028) );
  XNOR U1144 ( .A(n1025), .B(Y0[2]), .Z(n382) );
  XNOR U1145 ( .A(n1030), .B(n1031), .Z(n1025) );
  XOR U1146 ( .A(n1024), .B(n1032), .Z(n1030) );
  AND U1147 ( .A(n442), .B(n1033), .Z(n1032) );
  XOR U1148 ( .A(n967), .B(n1034), .Z(n1033) );
  XOR U1149 ( .A(n1034), .B(n968), .Z(n967) );
  NANDN U1150 ( .B(n1035), .A(n1036), .Z(n968) );
  IV U1151 ( .A(n1031), .Z(n1034) );
  XOR U1152 ( .A(n986), .B(n985), .Z(n1031) );
  XNOR U1153 ( .A(n1037), .B(n989), .Z(n985) );
  XNOR U1154 ( .A(n977), .B(n1039), .Z(n978) );
  AND U1155 ( .A(n976), .B(n489), .Z(n1039) );
  XOR U1156 ( .A(n1043), .B(n979), .Z(n1038) );
  NAND U1157 ( .A(n524), .B(n905), .Z(n979) );
  IV U1158 ( .A(n971), .Z(n1043) );
  XNOR U1159 ( .A(n982), .B(n983), .Z(n973) );
  NAND U1160 ( .A(n606), .B(n775), .Z(n983) );
  XNOR U1161 ( .A(n981), .B(n1047), .Z(n982) );
  AND U1162 ( .A(n842), .B(n561), .Z(n1047) );
  XNOR U1163 ( .A(n988), .B(n984), .Z(n1037) );
  AND U1164 ( .A(n1055), .B(n1056), .Z(n1054) );
  OR U1165 ( .A(n1057), .B(n1058), .Z(n1056) );
  AND U1166 ( .A(n1059), .B(n1060), .Z(n1055) );
  NANDN U1167 ( .B(n463), .A(n1061), .Z(n1060) );
  NANDN U1168 ( .B(n1062), .A(n1063), .Z(n1059) );
  XNOR U1169 ( .A(n1067), .B(n1006), .Z(n996) );
  XNOR U1170 ( .A(n993), .B(n994), .Z(n1006) );
  NAND U1171 ( .A(n589), .B(n817), .Z(n994) );
  XNOR U1172 ( .A(n992), .B(n1068), .Z(n993) );
  AND U1173 ( .A(n752), .B(n630), .Z(n1068) );
  XNOR U1174 ( .A(n1005), .B(n995), .Z(n1067) );
  XNOR U1175 ( .A(n1000), .B(n1076), .Z(n1001) );
  AND U1176 ( .A(n651), .B(n737), .Z(n1076) );
  XOR U1177 ( .A(n1080), .B(n1002), .Z(n1075) );
  NAND U1178 ( .A(n683), .B(n700), .Z(n1002) );
  IV U1179 ( .A(n1004), .Z(n1080) );
  XNOR U1180 ( .A(n1009), .B(n1085), .Z(n1012) );
  AND U1181 ( .A(n882), .B(n557), .Z(n1085) );
  XOR U1182 ( .A(n1086), .B(n1087), .Z(n1009) );
  ANDN U1183 ( .A(n1088), .B(n1089), .Z(n1087) );
  XNOR U1184 ( .A(n1090), .B(n1086), .Z(n1088) );
  XOR U1185 ( .A(n1091), .B(n1013), .Z(n1084) );
  NAND U1186 ( .A(n519), .B(n950), .Z(n1013) );
  IV U1187 ( .A(n1015), .Z(n1091) );
  XNOR U1188 ( .A(n1022), .B(n1023), .Z(n1017) );
  OR U1189 ( .A(n1095), .B(n464), .Z(n1023) );
  XNOR U1190 ( .A(n1021), .B(n1096), .Z(n1022) );
  ANDN U1191 ( .A(n488), .B(n1018), .Z(n1096) );
  ANDN U1192 ( .A(n1097), .B(n1098), .Z(n1021) );
  NANDN U1193 ( .B(n1099), .A(n1100), .Z(n1097) );
  NAND U1194 ( .A(n1103), .B(n1104), .Z(n217) );
  NANDN U1195 ( .B(n379), .A(Y[0]), .Z(n1104) );
  AND U1196 ( .A(n1105), .B(n1106), .Z(n1103) );
  NANDN U1197 ( .B(n426), .A(Y[0]), .Z(n1106) );
  IV U1198 ( .A(n1107), .Z(n426) );
  OR U1199 ( .A(n431), .B(n377), .Z(n1105) );
  IV U1200 ( .A(Y0[1]), .Z(n383) );
  XOR U1201 ( .A(n1108), .B(n1109), .Z(n1102) );
  XNOR U1202 ( .A(n1110), .B(n1101), .Z(n1108) );
  NAND U1203 ( .A(Y0[0]), .B(n1035), .Z(n1101) );
  NAND U1204 ( .A(n1111), .B(n442), .Z(n1110) );
  XOR U1205 ( .A(A[15]), .B(X[15]), .Z(n442) );
  XNOR U1206 ( .A(n1036), .B(n1109), .Z(n1111) );
  XNOR U1207 ( .A(n1035), .B(n1109), .Z(n1036) );
  XNOR U1208 ( .A(n1053), .B(n1052), .Z(n1109) );
  XNOR U1209 ( .A(n1112), .B(n1066), .Z(n1052) );
  XNOR U1210 ( .A(n1040), .B(n1114), .Z(n1041) );
  AND U1211 ( .A(n976), .B(n524), .Z(n1114) );
  XOR U1212 ( .A(n1118), .B(n1042), .Z(n1113) );
  NAND U1213 ( .A(n561), .B(n905), .Z(n1042) );
  IV U1214 ( .A(n1044), .Z(n1118) );
  XNOR U1215 ( .A(n1049), .B(n1050), .Z(n1046) );
  NAND U1216 ( .A(n651), .B(n775), .Z(n1050) );
  XNOR U1217 ( .A(n1048), .B(n1122), .Z(n1049) );
  AND U1218 ( .A(n842), .B(n606), .Z(n1122) );
  XNOR U1219 ( .A(n1065), .B(n1051), .Z(n1112) );
  XNOR U1220 ( .A(n1129), .B(n1062), .Z(n1065) );
  XOR U1221 ( .A(n1130), .B(n1057), .Z(n1062) );
  NAND U1222 ( .A(n489), .B(n1061), .Z(n1057) );
  NANDN U1223 ( .B(n463), .A(n1132), .Z(n1131) );
  XNOR U1224 ( .A(n1063), .B(n1064), .Z(n1129) );
  XNOR U1225 ( .A(n1142), .B(n1083), .Z(n1073) );
  XNOR U1226 ( .A(n1070), .B(n1071), .Z(n1083) );
  NAND U1227 ( .A(n589), .B(n882), .Z(n1071) );
  XNOR U1228 ( .A(n1069), .B(n1143), .Z(n1070) );
  AND U1229 ( .A(n817), .B(n630), .Z(n1143) );
  XNOR U1230 ( .A(n1082), .B(n1072), .Z(n1142) );
  XNOR U1231 ( .A(n1077), .B(n1151), .Z(n1078) );
  AND U1232 ( .A(n700), .B(n737), .Z(n1151) );
  XOR U1233 ( .A(n1155), .B(n1079), .Z(n1150) );
  NAND U1234 ( .A(n683), .B(n752), .Z(n1079) );
  IV U1235 ( .A(n1081), .Z(n1155) );
  XNOR U1236 ( .A(n1086), .B(n1160), .Z(n1089) );
  AND U1237 ( .A(n950), .B(n557), .Z(n1160) );
  XOR U1238 ( .A(n1164), .B(n1090), .Z(n1159) );
  NANDN U1239 ( .B(n1018), .A(n519), .Z(n1090) );
  IV U1240 ( .A(n1092), .Z(n1164) );
  XNOR U1241 ( .A(n1099), .B(n1100), .Z(n1094) );
  NANDN U1242 ( .B(n464), .A(n1168), .Z(n1100) );
  ANDN U1243 ( .A(n488), .B(n1095), .Z(n1169) );
  NAND U1244 ( .A(n1170), .B(n1171), .Z(n1098) );
  NANDN U1245 ( .B(n1172), .A(n1173), .Z(n1170) );
  XNOR U1246 ( .A(n1128), .B(n1127), .Z(n1035) );
  XNOR U1247 ( .A(n1174), .B(n1138), .Z(n1127) );
  XNOR U1248 ( .A(n1115), .B(n1176), .Z(n1116) );
  AND U1249 ( .A(n976), .B(n561), .Z(n1176) );
  XOR U1250 ( .A(n1180), .B(n1117), .Z(n1175) );
  NAND U1251 ( .A(n606), .B(n905), .Z(n1117) );
  IV U1252 ( .A(n1119), .Z(n1180) );
  XNOR U1253 ( .A(n1124), .B(n1125), .Z(n1121) );
  NAND U1254 ( .A(n700), .B(n775), .Z(n1125) );
  XNOR U1255 ( .A(n1123), .B(n1184), .Z(n1124) );
  AND U1256 ( .A(n842), .B(n651), .Z(n1184) );
  XNOR U1257 ( .A(n1137), .B(n1126), .Z(n1174) );
  XOR U1258 ( .A(n1188), .B(n1189), .Z(n1126) );
  XNOR U1259 ( .A(n1190), .B(n1141), .Z(n1137) );
  NAND U1260 ( .A(n524), .B(n1061), .Z(n1135) );
  XNOR U1261 ( .A(n1133), .B(n1191), .Z(n1134) );
  AND U1262 ( .A(n1132), .B(n489), .Z(n1191) );
  XNOR U1263 ( .A(n1140), .B(n1136), .Z(n1190) );
  XOR U1264 ( .A(n1195), .B(n1196), .Z(n1136) );
  AND U1265 ( .A(n1197), .B(n1198), .Z(n1196) );
  XOR U1266 ( .A(n1199), .B(n1200), .Z(n1198) );
  XOR U1267 ( .A(n1195), .B(n1201), .Z(n1200) );
  XOR U1268 ( .A(n1182), .B(n1202), .Z(n1197) );
  XOR U1269 ( .A(n1195), .B(n1183), .Z(n1202) );
  NAND U1270 ( .A(n775), .B(n752), .Z(n1187) );
  XNOR U1271 ( .A(n1185), .B(n1203), .Z(n1186) );
  AND U1272 ( .A(n842), .B(n700), .Z(n1203) );
  XNOR U1273 ( .A(n1177), .B(n1208), .Z(n1178) );
  AND U1274 ( .A(n976), .B(n606), .Z(n1208) );
  XOR U1275 ( .A(n1209), .B(n1210), .Z(n1177) );
  ANDN U1276 ( .A(n1211), .B(n1212), .Z(n1210) );
  XNOR U1277 ( .A(n1213), .B(n1209), .Z(n1211) );
  XOR U1278 ( .A(n1214), .B(n1179), .Z(n1207) );
  NAND U1279 ( .A(n651), .B(n905), .Z(n1179) );
  IV U1280 ( .A(n1181), .Z(n1214) );
  XOR U1281 ( .A(n1218), .B(n1219), .Z(n1195) );
  AND U1282 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U1283 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U1284 ( .A(n1218), .B(n1224), .Z(n1223) );
  XOR U1285 ( .A(n1216), .B(n1225), .Z(n1220) );
  XOR U1286 ( .A(n1218), .B(n1217), .Z(n1225) );
  NAND U1287 ( .A(n775), .B(n817), .Z(n1206) );
  XNOR U1288 ( .A(n1204), .B(n1226), .Z(n1205) );
  AND U1289 ( .A(n752), .B(n842), .Z(n1226) );
  XNOR U1290 ( .A(n1209), .B(n1231), .Z(n1212) );
  AND U1291 ( .A(n976), .B(n651), .Z(n1231) );
  XOR U1292 ( .A(n1232), .B(n1233), .Z(n1209) );
  ANDN U1293 ( .A(n1234), .B(n1235), .Z(n1233) );
  XNOR U1294 ( .A(n1236), .B(n1232), .Z(n1234) );
  XOR U1295 ( .A(n1237), .B(n1213), .Z(n1230) );
  NAND U1296 ( .A(n700), .B(n905), .Z(n1213) );
  IV U1297 ( .A(n1215), .Z(n1237) );
  XOR U1298 ( .A(n1241), .B(n1242), .Z(n1218) );
  AND U1299 ( .A(n1243), .B(n1244), .Z(n1242) );
  XOR U1300 ( .A(n1245), .B(n1246), .Z(n1244) );
  XOR U1301 ( .A(n1241), .B(n1247), .Z(n1246) );
  XOR U1302 ( .A(n1239), .B(n1248), .Z(n1243) );
  XOR U1303 ( .A(n1241), .B(n1240), .Z(n1248) );
  NAND U1304 ( .A(n775), .B(n882), .Z(n1229) );
  XNOR U1305 ( .A(n1227), .B(n1249), .Z(n1228) );
  AND U1306 ( .A(n817), .B(n842), .Z(n1249) );
  XNOR U1307 ( .A(n1232), .B(n1254), .Z(n1235) );
  AND U1308 ( .A(n976), .B(n700), .Z(n1254) );
  XOR U1309 ( .A(n1255), .B(n1256), .Z(n1232) );
  ANDN U1310 ( .A(n1257), .B(n1258), .Z(n1256) );
  XNOR U1311 ( .A(n1259), .B(n1255), .Z(n1257) );
  XOR U1312 ( .A(n1260), .B(n1236), .Z(n1253) );
  NAND U1313 ( .A(n905), .B(n752), .Z(n1236) );
  IV U1314 ( .A(n1238), .Z(n1260) );
  XOR U1315 ( .A(n1264), .B(n1265), .Z(n1241) );
  AND U1316 ( .A(n1266), .B(n1267), .Z(n1265) );
  XOR U1317 ( .A(n1268), .B(n1269), .Z(n1267) );
  XOR U1318 ( .A(n1264), .B(n1270), .Z(n1269) );
  XOR U1319 ( .A(n1262), .B(n1271), .Z(n1266) );
  XOR U1320 ( .A(n1264), .B(n1263), .Z(n1271) );
  XNOR U1321 ( .A(n1272), .B(n1252), .Z(n1263) );
  NAND U1322 ( .A(n775), .B(n950), .Z(n1252) );
  IV U1323 ( .A(n1251), .Z(n1272) );
  XNOR U1324 ( .A(n1250), .B(n1273), .Z(n1251) );
  AND U1325 ( .A(n882), .B(n842), .Z(n1273) );
  XOR U1326 ( .A(n1274), .B(n1275), .Z(n1250) );
  ANDN U1327 ( .A(n1276), .B(n1277), .Z(n1275) );
  XNOR U1328 ( .A(n1278), .B(n1274), .Z(n1276) );
  XNOR U1329 ( .A(n1279), .B(n1280), .Z(n1262) );
  IV U1330 ( .A(n1258), .Z(n1280) );
  XNOR U1331 ( .A(n1255), .B(n1281), .Z(n1258) );
  AND U1332 ( .A(n752), .B(n976), .Z(n1281) );
  XOR U1333 ( .A(n1282), .B(n1283), .Z(n1255) );
  ANDN U1334 ( .A(n1284), .B(n1285), .Z(n1283) );
  XNOR U1335 ( .A(n1286), .B(n1282), .Z(n1284) );
  XOR U1336 ( .A(n1287), .B(n1259), .Z(n1279) );
  NAND U1337 ( .A(n905), .B(n817), .Z(n1259) );
  IV U1338 ( .A(n1261), .Z(n1287) );
  XOR U1339 ( .A(n1291), .B(n1292), .Z(n1264) );
  AND U1340 ( .A(n1293), .B(n1294), .Z(n1292) );
  XOR U1341 ( .A(n1295), .B(n1296), .Z(n1294) );
  XOR U1342 ( .A(n1291), .B(n1297), .Z(n1296) );
  XOR U1343 ( .A(n1289), .B(n1298), .Z(n1293) );
  XOR U1344 ( .A(n1291), .B(n1290), .Z(n1298) );
  XNOR U1345 ( .A(n1299), .B(n1278), .Z(n1290) );
  NANDN U1346 ( .B(n1018), .A(n775), .Z(n1278) );
  IV U1347 ( .A(n1277), .Z(n1299) );
  XNOR U1348 ( .A(n1274), .B(n1300), .Z(n1277) );
  AND U1349 ( .A(n950), .B(n842), .Z(n1300) );
  XOR U1350 ( .A(n1301), .B(n1302), .Z(n1274) );
  ANDN U1351 ( .A(n1303), .B(n1304), .Z(n1302) );
  XNOR U1352 ( .A(n1305), .B(n1301), .Z(n1303) );
  XNOR U1353 ( .A(n1306), .B(n1307), .Z(n1289) );
  IV U1354 ( .A(n1285), .Z(n1307) );
  XNOR U1355 ( .A(n1282), .B(n1308), .Z(n1285) );
  AND U1356 ( .A(n817), .B(n976), .Z(n1308) );
  XOR U1357 ( .A(n1309), .B(n1310), .Z(n1282) );
  ANDN U1358 ( .A(n1311), .B(n1312), .Z(n1310) );
  XNOR U1359 ( .A(n1313), .B(n1309), .Z(n1311) );
  XOR U1360 ( .A(n1314), .B(n1286), .Z(n1306) );
  NAND U1361 ( .A(n905), .B(n882), .Z(n1286) );
  IV U1362 ( .A(n1288), .Z(n1314) );
  XOR U1363 ( .A(n1318), .B(n1319), .Z(n1291) );
  AND U1364 ( .A(n1320), .B(n1321), .Z(n1319) );
  XOR U1365 ( .A(n1322), .B(n1323), .Z(n1321) );
  XOR U1366 ( .A(n1318), .B(n1324), .Z(n1323) );
  XOR U1367 ( .A(n1316), .B(n1325), .Z(n1320) );
  XOR U1368 ( .A(n1318), .B(n1317), .Z(n1325) );
  XNOR U1369 ( .A(n1326), .B(n1305), .Z(n1317) );
  NANDN U1370 ( .B(n1095), .A(n775), .Z(n1305) );
  IV U1371 ( .A(n1304), .Z(n1326) );
  XNOR U1372 ( .A(n1301), .B(n1327), .Z(n1304) );
  ANDN U1373 ( .A(n842), .B(n1018), .Z(n1327) );
  XOR U1374 ( .A(n1328), .B(n1329), .Z(n1301) );
  ANDN U1375 ( .A(n1330), .B(n1331), .Z(n1329) );
  XNOR U1376 ( .A(n1332), .B(n1328), .Z(n1330) );
  XNOR U1377 ( .A(n1333), .B(n1334), .Z(n1316) );
  IV U1378 ( .A(n1312), .Z(n1334) );
  XNOR U1379 ( .A(n1309), .B(n1335), .Z(n1312) );
  AND U1380 ( .A(n882), .B(n976), .Z(n1335) );
  XOR U1381 ( .A(n1336), .B(n1337), .Z(n1309) );
  ANDN U1382 ( .A(n1338), .B(n1339), .Z(n1337) );
  XNOR U1383 ( .A(n1340), .B(n1336), .Z(n1338) );
  XOR U1384 ( .A(n1341), .B(n1313), .Z(n1333) );
  NAND U1385 ( .A(n905), .B(n950), .Z(n1313) );
  IV U1386 ( .A(n1315), .Z(n1341) );
  XOR U1387 ( .A(n1345), .B(n1346), .Z(n1318) );
  AND U1388 ( .A(n1347), .B(n1348), .Z(n1346) );
  XOR U1389 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U1390 ( .A(n1345), .B(n1351), .Z(n1350) );
  XOR U1391 ( .A(n1343), .B(n1352), .Z(n1347) );
  XOR U1392 ( .A(n1345), .B(n1344), .Z(n1352) );
  XNOR U1393 ( .A(n1353), .B(n1332), .Z(n1344) );
  NAND U1394 ( .A(n775), .B(n1168), .Z(n1332) );
  IV U1395 ( .A(n1331), .Z(n1353) );
  XNOR U1396 ( .A(n1328), .B(n1354), .Z(n1331) );
  ANDN U1397 ( .A(n842), .B(n1095), .Z(n1354) );
  XOR U1398 ( .A(n1355), .B(n1356), .Z(n1328) );
  ANDN U1399 ( .A(n1357), .B(n1358), .Z(n1356) );
  XNOR U1400 ( .A(n1359), .B(n1355), .Z(n1357) );
  XNOR U1401 ( .A(n1360), .B(n1361), .Z(n1343) );
  IV U1402 ( .A(n1339), .Z(n1361) );
  XNOR U1403 ( .A(n1336), .B(n1362), .Z(n1339) );
  AND U1404 ( .A(n950), .B(n976), .Z(n1362) );
  XOR U1405 ( .A(n1363), .B(n1364), .Z(n1336) );
  ANDN U1406 ( .A(n1365), .B(n1366), .Z(n1364) );
  XNOR U1407 ( .A(n1367), .B(n1363), .Z(n1365) );
  XOR U1408 ( .A(n1368), .B(n1340), .Z(n1360) );
  NANDN U1409 ( .B(n1018), .A(n905), .Z(n1340) );
  IV U1410 ( .A(n1342), .Z(n1368) );
  XOR U1411 ( .A(n1373), .B(n1374), .Z(n1189) );
  XNOR U1412 ( .A(n1375), .B(n1372), .Z(n1373) );
  XNOR U1413 ( .A(n1363), .B(n1377), .Z(n1366) );
  ANDN U1414 ( .A(n976), .B(n1018), .Z(n1377) );
  XOR U1415 ( .A(n1380), .B(n1378), .Z(n1379) );
  ANDN U1416 ( .A(n976), .B(n1095), .Z(n1380) );
  AND U1417 ( .A(n1168), .B(n905), .Z(n1381) );
  XOR U1418 ( .A(n1382), .B(n1383), .Z(n1378) );
  ANDN U1419 ( .A(n1384), .B(n1385), .Z(n1383) );
  XNOR U1420 ( .A(n1386), .B(n1382), .Z(n1384) );
  XOR U1421 ( .A(n1387), .B(n1367), .Z(n1376) );
  NANDN U1422 ( .B(n1095), .A(n905), .Z(n1367) );
  IV U1423 ( .A(n1369), .Z(n1387) );
  NAND U1424 ( .A(n905), .B(n1388), .Z(n1386) );
  XNOR U1425 ( .A(n1382), .B(n1389), .Z(n1385) );
  AND U1426 ( .A(n1168), .B(n976), .Z(n1389) );
  AND U1427 ( .A(n1390), .B(A[0]), .Z(n1382) );
  NANDN U1428 ( .B(n905), .A(n1391), .Z(n1390) );
  NAND U1429 ( .A(n1388), .B(n976), .Z(n1391) );
  XNOR U1430 ( .A(n1358), .B(n1359), .Z(n1371) );
  NAND U1431 ( .A(n775), .B(n1388), .Z(n1359) );
  XNOR U1432 ( .A(n1355), .B(n1394), .Z(n1358) );
  AND U1433 ( .A(n1168), .B(n842), .Z(n1394) );
  AND U1434 ( .A(n1395), .B(A[0]), .Z(n1355) );
  NANDN U1435 ( .B(n775), .A(n1396), .Z(n1395) );
  NAND U1436 ( .A(n1388), .B(n842), .Z(n1396) );
  XOR U1437 ( .A(n1399), .B(n1400), .Z(n1372) );
  XOR U1438 ( .A(n1401), .B(n1402), .Z(n1140) );
  AND U1439 ( .A(n1403), .B(n1404), .Z(n1402) );
  NANDN U1440 ( .B(n463), .A(n1405), .Z(n1404) );
  NANDN U1441 ( .B(n1406), .A(n1407), .Z(n463) );
  AND U1442 ( .A(n1408), .B(A[15]), .Z(n1407) );
  OR U1443 ( .A(n1409), .B(n1410), .Z(n1403) );
  IV U1444 ( .A(n1139), .Z(n1401) );
  NAND U1445 ( .A(n561), .B(n1061), .Z(n1194) );
  XNOR U1446 ( .A(n1192), .B(n1412), .Z(n1193) );
  AND U1447 ( .A(n1132), .B(n524), .Z(n1412) );
  XOR U1448 ( .A(n1420), .B(n1409), .Z(n1416) );
  NAND U1449 ( .A(n489), .B(n1405), .Z(n1409) );
  IV U1450 ( .A(n1411), .Z(n1420) );
  NAND U1451 ( .A(n606), .B(n1061), .Z(n1415) );
  XNOR U1452 ( .A(n1413), .B(n1422), .Z(n1414) );
  AND U1453 ( .A(n1132), .B(n561), .Z(n1422) );
  XNOR U1454 ( .A(n1417), .B(n1427), .Z(n1418) );
  AND U1455 ( .A(n489), .B(X[0]), .Z(n1427) );
  XNOR U1456 ( .A(n1408), .B(A[14]), .Z(n1406) );
  NOR U1457 ( .A(n1428), .B(n1429), .Z(n1408) );
  XOR U1458 ( .A(n1433), .B(n1419), .Z(n1426) );
  NAND U1459 ( .A(n524), .B(n1405), .Z(n1419) );
  IV U1460 ( .A(n1421), .Z(n1433) );
  NAND U1461 ( .A(n651), .B(n1061), .Z(n1425) );
  XNOR U1462 ( .A(n1423), .B(n1435), .Z(n1424) );
  AND U1463 ( .A(n1132), .B(n606), .Z(n1435) );
  XOR U1464 ( .A(n1436), .B(n1437), .Z(n1423) );
  ANDN U1465 ( .A(n1438), .B(n1439), .Z(n1437) );
  XNOR U1466 ( .A(n1440), .B(n1436), .Z(n1438) );
  XNOR U1467 ( .A(n1430), .B(n1442), .Z(n1431) );
  AND U1468 ( .A(n524), .B(X[0]), .Z(n1442) );
  XOR U1469 ( .A(n1428), .B(A[13]), .Z(n1429) );
  NANDN U1470 ( .B(n1443), .A(n1444), .Z(n1428) );
  XOR U1471 ( .A(n1448), .B(n1432), .Z(n1441) );
  NAND U1472 ( .A(n561), .B(n1405), .Z(n1432) );
  IV U1473 ( .A(n1434), .Z(n1448) );
  XNOR U1474 ( .A(n1450), .B(n1440), .Z(n1268) );
  NAND U1475 ( .A(n700), .B(n1061), .Z(n1440) );
  IV U1476 ( .A(n1439), .Z(n1450) );
  XNOR U1477 ( .A(n1436), .B(n1451), .Z(n1439) );
  AND U1478 ( .A(n1132), .B(n651), .Z(n1451) );
  XOR U1479 ( .A(n1452), .B(n1453), .Z(n1436) );
  ANDN U1480 ( .A(n1454), .B(n1455), .Z(n1453) );
  XNOR U1481 ( .A(n1456), .B(n1452), .Z(n1454) );
  XNOR U1482 ( .A(n1457), .B(n1458), .Z(n1270) );
  IV U1483 ( .A(n1446), .Z(n1458) );
  XNOR U1484 ( .A(n1445), .B(n1459), .Z(n1446) );
  AND U1485 ( .A(n561), .B(X[0]), .Z(n1459) );
  XNOR U1486 ( .A(n1444), .B(A[12]), .Z(n1443) );
  NOR U1487 ( .A(n1460), .B(n1461), .Z(n1444) );
  XOR U1488 ( .A(n1462), .B(n1463), .Z(n1445) );
  ANDN U1489 ( .A(n1464), .B(n1465), .Z(n1463) );
  XNOR U1490 ( .A(n1466), .B(n1462), .Z(n1464) );
  XOR U1491 ( .A(n1467), .B(n1447), .Z(n1457) );
  NAND U1492 ( .A(n606), .B(n1405), .Z(n1447) );
  IV U1493 ( .A(n1449), .Z(n1467) );
  XNOR U1494 ( .A(n1469), .B(n1456), .Z(n1295) );
  NAND U1495 ( .A(n752), .B(n1061), .Z(n1456) );
  IV U1496 ( .A(n1455), .Z(n1469) );
  XNOR U1497 ( .A(n1452), .B(n1470), .Z(n1455) );
  AND U1498 ( .A(n1132), .B(n700), .Z(n1470) );
  XOR U1499 ( .A(n1471), .B(n1472), .Z(n1452) );
  ANDN U1500 ( .A(n1473), .B(n1474), .Z(n1472) );
  XNOR U1501 ( .A(n1475), .B(n1471), .Z(n1473) );
  XNOR U1502 ( .A(n1476), .B(n1477), .Z(n1297) );
  IV U1503 ( .A(n1465), .Z(n1477) );
  XNOR U1504 ( .A(n1462), .B(n1478), .Z(n1465) );
  AND U1505 ( .A(n606), .B(X[0]), .Z(n1478) );
  XOR U1506 ( .A(n1460), .B(A[11]), .Z(n1461) );
  NANDN U1507 ( .B(n1479), .A(n1480), .Z(n1460) );
  XOR U1508 ( .A(n1481), .B(n1482), .Z(n1462) );
  ANDN U1509 ( .A(n1483), .B(n1484), .Z(n1482) );
  XNOR U1510 ( .A(n1485), .B(n1481), .Z(n1483) );
  XOR U1511 ( .A(n1486), .B(n1466), .Z(n1476) );
  NAND U1512 ( .A(n651), .B(n1405), .Z(n1466) );
  IV U1513 ( .A(n1468), .Z(n1486) );
  XNOR U1514 ( .A(n1488), .B(n1475), .Z(n1322) );
  NAND U1515 ( .A(n817), .B(n1061), .Z(n1475) );
  IV U1516 ( .A(n1474), .Z(n1488) );
  XNOR U1517 ( .A(n1471), .B(n1489), .Z(n1474) );
  AND U1518 ( .A(n1132), .B(n752), .Z(n1489) );
  XOR U1519 ( .A(n1490), .B(n1491), .Z(n1471) );
  ANDN U1520 ( .A(n1492), .B(n1493), .Z(n1491) );
  XNOR U1521 ( .A(n1494), .B(n1490), .Z(n1492) );
  XNOR U1522 ( .A(n1495), .B(n1496), .Z(n1324) );
  IV U1523 ( .A(n1484), .Z(n1496) );
  XNOR U1524 ( .A(n1481), .B(n1497), .Z(n1484) );
  AND U1525 ( .A(n651), .B(X[0]), .Z(n1497) );
  XNOR U1526 ( .A(n1480), .B(A[10]), .Z(n1479) );
  NOR U1527 ( .A(n1498), .B(n1499), .Z(n1480) );
  XOR U1528 ( .A(n1500), .B(n1501), .Z(n1481) );
  ANDN U1529 ( .A(n1502), .B(n1503), .Z(n1501) );
  XNOR U1530 ( .A(n1504), .B(n1500), .Z(n1502) );
  XOR U1531 ( .A(n1505), .B(n1485), .Z(n1495) );
  NAND U1532 ( .A(n700), .B(n1405), .Z(n1485) );
  IV U1533 ( .A(n1487), .Z(n1505) );
  XNOR U1534 ( .A(n1507), .B(n1494), .Z(n1349) );
  NAND U1535 ( .A(n882), .B(n1061), .Z(n1494) );
  IV U1536 ( .A(n1493), .Z(n1507) );
  XNOR U1537 ( .A(n1490), .B(n1508), .Z(n1493) );
  AND U1538 ( .A(n1132), .B(n817), .Z(n1508) );
  XOR U1539 ( .A(n1509), .B(n1510), .Z(n1490) );
  ANDN U1540 ( .A(n1511), .B(n1512), .Z(n1510) );
  XNOR U1541 ( .A(n1513), .B(n1509), .Z(n1511) );
  XNOR U1542 ( .A(n1514), .B(n1515), .Z(n1351) );
  IV U1543 ( .A(n1503), .Z(n1515) );
  XNOR U1544 ( .A(n1500), .B(n1516), .Z(n1503) );
  AND U1545 ( .A(n700), .B(X[0]), .Z(n1516) );
  XOR U1546 ( .A(n1498), .B(A[9]), .Z(n1499) );
  NANDN U1547 ( .B(n1517), .A(n1518), .Z(n1498) );
  XOR U1548 ( .A(n1519), .B(n1520), .Z(n1500) );
  ANDN U1549 ( .A(n1521), .B(n1522), .Z(n1520) );
  XNOR U1550 ( .A(n1523), .B(n1519), .Z(n1521) );
  XOR U1551 ( .A(n1524), .B(n1504), .Z(n1514) );
  NAND U1552 ( .A(n752), .B(n1405), .Z(n1504) );
  IV U1553 ( .A(n1506), .Z(n1524) );
  NAND U1554 ( .A(n950), .B(n1061), .Z(n1513) );
  XNOR U1555 ( .A(n1509), .B(n1526), .Z(n1512) );
  AND U1556 ( .A(n1132), .B(n882), .Z(n1526) );
  XNOR U1557 ( .A(n1530), .B(n1527), .Z(n1529) );
  XNOR U1558 ( .A(n1519), .B(n1532), .Z(n1522) );
  AND U1559 ( .A(n752), .B(X[0]), .Z(n1532) );
  XNOR U1560 ( .A(n1536), .B(n1533), .Z(n1535) );
  XOR U1561 ( .A(n1537), .B(n1523), .Z(n1531) );
  NAND U1562 ( .A(n817), .B(n1405), .Z(n1523) );
  IV U1563 ( .A(n1525), .Z(n1537) );
  XNOR U1564 ( .A(n1538), .B(n1539), .Z(n1525) );
  AND U1565 ( .A(n1540), .B(n1541), .Z(n1539) );
  XOR U1566 ( .A(n1534), .B(n1542), .Z(n1541) );
  XNOR U1567 ( .A(n1536), .B(n1538), .Z(n1542) );
  NAND U1568 ( .A(n882), .B(n1405), .Z(n1536) );
  XOR U1569 ( .A(n1533), .B(n1543), .Z(n1534) );
  AND U1570 ( .A(n817), .B(X[0]), .Z(n1543) );
  XNOR U1571 ( .A(n1547), .B(n1544), .Z(n1546) );
  XOR U1572 ( .A(n1528), .B(n1548), .Z(n1540) );
  XNOR U1573 ( .A(n1530), .B(n1538), .Z(n1548) );
  NANDN U1574 ( .B(n1018), .A(n1061), .Z(n1530) );
  XOR U1575 ( .A(n1527), .B(n1549), .Z(n1528) );
  AND U1576 ( .A(n1132), .B(n950), .Z(n1549) );
  XOR U1577 ( .A(n1550), .B(n1551), .Z(n1527) );
  AND U1578 ( .A(n1552), .B(n1553), .Z(n1551) );
  XNOR U1579 ( .A(n1554), .B(n1550), .Z(n1553) );
  XOR U1580 ( .A(n1555), .B(n1556), .Z(n1538) );
  AND U1581 ( .A(n1557), .B(n1558), .Z(n1556) );
  XOR U1582 ( .A(n1545), .B(n1559), .Z(n1558) );
  XNOR U1583 ( .A(n1547), .B(n1555), .Z(n1559) );
  NAND U1584 ( .A(n950), .B(n1405), .Z(n1547) );
  XOR U1585 ( .A(n1544), .B(n1560), .Z(n1545) );
  AND U1586 ( .A(n882), .B(X[0]), .Z(n1560) );
  XNOR U1587 ( .A(n1564), .B(n1561), .Z(n1563) );
  XOR U1588 ( .A(n1552), .B(n1565), .Z(n1557) );
  XNOR U1589 ( .A(n1554), .B(n1555), .Z(n1565) );
  NANDN U1590 ( .B(n1095), .A(n1061), .Z(n1554) );
  XOR U1591 ( .A(n1550), .B(n1566), .Z(n1552) );
  ANDN U1592 ( .A(n1132), .B(n1018), .Z(n1566) );
  XOR U1593 ( .A(n1567), .B(n1568), .Z(n1550) );
  AND U1594 ( .A(n1569), .B(n1570), .Z(n1568) );
  XNOR U1595 ( .A(n1571), .B(n1567), .Z(n1570) );
  XOR U1596 ( .A(n1572), .B(n1573), .Z(n1555) );
  AND U1597 ( .A(n1574), .B(n1575), .Z(n1573) );
  XOR U1598 ( .A(n1562), .B(n1576), .Z(n1575) );
  XNOR U1599 ( .A(n1564), .B(n1572), .Z(n1576) );
  NANDN U1600 ( .B(n1018), .A(n1405), .Z(n1564) );
  XOR U1601 ( .A(n1561), .B(n1577), .Z(n1562) );
  AND U1602 ( .A(n950), .B(X[0]), .Z(n1577) );
  XOR U1603 ( .A(n1569), .B(n1581), .Z(n1574) );
  XNOR U1604 ( .A(n1571), .B(n1572), .Z(n1581) );
  NAND U1605 ( .A(n1061), .B(n1168), .Z(n1571) );
  XOR U1606 ( .A(n1567), .B(n1582), .Z(n1569) );
  ANDN U1607 ( .A(n1132), .B(n1095), .Z(n1582) );
  NAND U1608 ( .A(n1061), .B(n1388), .Z(n1585) );
  XNOR U1609 ( .A(n1583), .B(n1587), .Z(n1584) );
  AND U1610 ( .A(n1168), .B(n1132), .Z(n1587) );
  AND U1611 ( .A(n1588), .B(A[0]), .Z(n1583) );
  NANDN U1612 ( .B(n1061), .A(n1589), .Z(n1588) );
  NAND U1613 ( .A(n1388), .B(n1132), .Z(n1589) );
  XNOR U1614 ( .A(n1578), .B(n1593), .Z(n1579) );
  ANDN U1615 ( .A(X[0]), .B(n1018), .Z(n1593) );
  XOR U1616 ( .A(n1596), .B(n1594), .Z(n1595) );
  ANDN U1617 ( .A(X[0]), .B(n1095), .Z(n1596) );
  AND U1618 ( .A(n1405), .B(n1168), .Z(n1597) );
  XOR U1619 ( .A(n1601), .B(n1580), .Z(n1592) );
  NANDN U1620 ( .B(n1095), .A(n1405), .Z(n1580) );
  IV U1621 ( .A(n1586), .Z(n1601) );
  NAND U1622 ( .A(n1405), .B(n1388), .Z(n1600) );
  XNOR U1623 ( .A(n1598), .B(n1602), .Z(n1599) );
  AND U1624 ( .A(n1168), .B(X[0]), .Z(n1602) );
  AND U1625 ( .A(n1603), .B(A[0]), .Z(n1598) );
  NANDN U1626 ( .B(n1405), .A(n1604), .Z(n1603) );
  NAND U1627 ( .A(n1388), .B(X[0]), .Z(n1604) );
  XNOR U1628 ( .A(n1606), .B(n1158), .Z(n1148) );
  XNOR U1629 ( .A(n1145), .B(n1146), .Z(n1158) );
  NAND U1630 ( .A(n589), .B(n950), .Z(n1146) );
  XNOR U1631 ( .A(n1144), .B(n1607), .Z(n1145) );
  AND U1632 ( .A(n882), .B(n630), .Z(n1607) );
  XNOR U1633 ( .A(n1611), .B(n1608), .Z(n1610) );
  XNOR U1634 ( .A(n1157), .B(n1147), .Z(n1606) );
  XOR U1635 ( .A(n1612), .B(n1613), .Z(n1147) );
  XNOR U1636 ( .A(n1152), .B(n1615), .Z(n1153) );
  AND U1637 ( .A(n752), .B(n737), .Z(n1615) );
  XNOR U1638 ( .A(n1518), .B(A[8]), .Z(n1517) );
  NOR U1639 ( .A(n1616), .B(n1617), .Z(n1518) );
  XOR U1640 ( .A(n1618), .B(n1619), .Z(n1152) );
  AND U1641 ( .A(n1620), .B(n1621), .Z(n1619) );
  XNOR U1642 ( .A(n1622), .B(n1618), .Z(n1621) );
  XOR U1643 ( .A(n1623), .B(n1154), .Z(n1614) );
  NAND U1644 ( .A(n683), .B(n817), .Z(n1154) );
  IV U1645 ( .A(n1156), .Z(n1623) );
  XNOR U1646 ( .A(n1624), .B(n1625), .Z(n1156) );
  AND U1647 ( .A(n1626), .B(n1627), .Z(n1625) );
  XOR U1648 ( .A(n1620), .B(n1628), .Z(n1627) );
  XNOR U1649 ( .A(n1622), .B(n1624), .Z(n1628) );
  NAND U1650 ( .A(n683), .B(n882), .Z(n1622) );
  XOR U1651 ( .A(n1618), .B(n1629), .Z(n1620) );
  AND U1652 ( .A(n817), .B(n737), .Z(n1629) );
  XOR U1653 ( .A(n1616), .B(A[7]), .Z(n1617) );
  NANDN U1654 ( .B(n1630), .A(n1631), .Z(n1616) );
  XOR U1655 ( .A(n1632), .B(n1633), .Z(n1618) );
  AND U1656 ( .A(n1634), .B(n1635), .Z(n1633) );
  XNOR U1657 ( .A(n1636), .B(n1632), .Z(n1635) );
  XOR U1658 ( .A(n1609), .B(n1637), .Z(n1626) );
  XNOR U1659 ( .A(n1611), .B(n1624), .Z(n1637) );
  NANDN U1660 ( .B(n1018), .A(n589), .Z(n1611) );
  XOR U1661 ( .A(n1608), .B(n1638), .Z(n1609) );
  AND U1662 ( .A(n950), .B(n630), .Z(n1638) );
  XNOR U1663 ( .A(n1642), .B(n1639), .Z(n1641) );
  XOR U1664 ( .A(n1643), .B(n1644), .Z(n1624) );
  AND U1665 ( .A(n1645), .B(n1646), .Z(n1644) );
  XOR U1666 ( .A(n1634), .B(n1647), .Z(n1646) );
  XNOR U1667 ( .A(n1636), .B(n1643), .Z(n1647) );
  NAND U1668 ( .A(n683), .B(n950), .Z(n1636) );
  XOR U1669 ( .A(n1632), .B(n1648), .Z(n1634) );
  AND U1670 ( .A(n882), .B(n737), .Z(n1648) );
  XNOR U1671 ( .A(n1631), .B(A[6]), .Z(n1630) );
  NOR U1672 ( .A(n1649), .B(n1650), .Z(n1631) );
  XOR U1673 ( .A(n1651), .B(n1652), .Z(n1632) );
  AND U1674 ( .A(n1653), .B(n1654), .Z(n1652) );
  XNOR U1675 ( .A(n1655), .B(n1651), .Z(n1654) );
  XOR U1676 ( .A(n1640), .B(n1656), .Z(n1645) );
  XNOR U1677 ( .A(n1642), .B(n1643), .Z(n1656) );
  NANDN U1678 ( .B(n1095), .A(n589), .Z(n1642) );
  XOR U1679 ( .A(n1639), .B(n1657), .Z(n1640) );
  ANDN U1680 ( .A(n630), .B(n1018), .Z(n1657) );
  XNOR U1681 ( .A(n1661), .B(n1658), .Z(n1660) );
  XOR U1682 ( .A(n1662), .B(n1663), .Z(n1643) );
  AND U1683 ( .A(n1664), .B(n1665), .Z(n1663) );
  XOR U1684 ( .A(n1653), .B(n1666), .Z(n1665) );
  XNOR U1685 ( .A(n1655), .B(n1662), .Z(n1666) );
  NANDN U1686 ( .B(n1018), .A(n683), .Z(n1655) );
  XOR U1687 ( .A(n1651), .B(n1667), .Z(n1653) );
  AND U1688 ( .A(n950), .B(n737), .Z(n1667) );
  XOR U1689 ( .A(n1649), .B(A[5]), .Z(n1650) );
  NANDN U1690 ( .B(n1668), .A(n1669), .Z(n1649) );
  XOR U1691 ( .A(n1670), .B(n1671), .Z(n1651) );
  ANDN U1692 ( .A(n1672), .B(n1673), .Z(n1671) );
  XNOR U1693 ( .A(n1674), .B(n1670), .Z(n1672) );
  XOR U1694 ( .A(n1659), .B(n1675), .Z(n1664) );
  XNOR U1695 ( .A(n1661), .B(n1662), .Z(n1675) );
  NAND U1696 ( .A(n589), .B(n1168), .Z(n1661) );
  XOR U1697 ( .A(n1658), .B(n1676), .Z(n1659) );
  ANDN U1698 ( .A(n630), .B(n1095), .Z(n1676) );
  XOR U1699 ( .A(n1677), .B(n1678), .Z(n1658) );
  ANDN U1700 ( .A(n1679), .B(n1680), .Z(n1678) );
  XNOR U1701 ( .A(n1681), .B(n1677), .Z(n1679) );
  NAND U1702 ( .A(n589), .B(n1388), .Z(n1681) );
  XNOR U1703 ( .A(n1677), .B(n1683), .Z(n1680) );
  AND U1704 ( .A(n1168), .B(n630), .Z(n1683) );
  AND U1705 ( .A(n1684), .B(A[0]), .Z(n1677) );
  NANDN U1706 ( .B(n589), .A(n1685), .Z(n1684) );
  NAND U1707 ( .A(n1388), .B(n630), .Z(n1685) );
  XNOR U1708 ( .A(n1670), .B(n1689), .Z(n1673) );
  ANDN U1709 ( .A(n737), .B(n1018), .Z(n1689) );
  XOR U1710 ( .A(n1690), .B(n1691), .Z(n1670) );
  AND U1711 ( .A(n1692), .B(n1693), .Z(n1691) );
  XOR U1712 ( .A(n1694), .B(n1690), .Z(n1693) );
  ANDN U1713 ( .A(n737), .B(n1095), .Z(n1694) );
  XOR U1714 ( .A(n1695), .B(n1690), .Z(n1692) );
  AND U1715 ( .A(n1168), .B(n683), .Z(n1695) );
  XOR U1716 ( .A(n1696), .B(n1697), .Z(n1690) );
  ANDN U1717 ( .A(n1698), .B(n1699), .Z(n1697) );
  XNOR U1718 ( .A(n1700), .B(n1696), .Z(n1698) );
  XOR U1719 ( .A(n1701), .B(n1674), .Z(n1688) );
  NANDN U1720 ( .B(n1095), .A(n683), .Z(n1674) );
  IV U1721 ( .A(n1682), .Z(n1701) );
  XOR U1722 ( .A(n1702), .B(n1700), .Z(n1682) );
  NAND U1723 ( .A(n683), .B(n1388), .Z(n1700) );
  IV U1724 ( .A(n1699), .Z(n1702) );
  XNOR U1725 ( .A(n1696), .B(n1703), .Z(n1699) );
  AND U1726 ( .A(n1168), .B(n737), .Z(n1703) );
  AND U1727 ( .A(n1704), .B(A[0]), .Z(n1696) );
  NANDN U1728 ( .B(n683), .A(n1705), .Z(n1704) );
  NAND U1729 ( .A(n1388), .B(n737), .Z(n1705) );
  XNOR U1730 ( .A(n1161), .B(n1709), .Z(n1162) );
  ANDN U1731 ( .A(n557), .B(n1018), .Z(n1709) );
  XNOR U1732 ( .A(n1669), .B(A[4]), .Z(n1668) );
  NOR U1733 ( .A(n1710), .B(n1711), .Z(n1669) );
  XOR U1734 ( .A(n1712), .B(n1713), .Z(n1161) );
  AND U1735 ( .A(n1714), .B(n1715), .Z(n1713) );
  XOR U1736 ( .A(n1716), .B(n1712), .Z(n1715) );
  ANDN U1737 ( .A(n557), .B(n1095), .Z(n1716) );
  XOR U1738 ( .A(n1717), .B(n1712), .Z(n1714) );
  AND U1739 ( .A(n1168), .B(n519), .Z(n1717) );
  XOR U1740 ( .A(n1718), .B(n1719), .Z(n1712) );
  ANDN U1741 ( .A(n1720), .B(n1721), .Z(n1719) );
  XNOR U1742 ( .A(n1722), .B(n1718), .Z(n1720) );
  XOR U1743 ( .A(n1723), .B(n1163), .Z(n1708) );
  NANDN U1744 ( .B(n1095), .A(n519), .Z(n1163) );
  NANDN U1745 ( .B(n1724), .A(n1725), .Z(n1710) );
  IV U1746 ( .A(n1165), .Z(n1723) );
  NAND U1747 ( .A(n519), .B(n1388), .Z(n1722) );
  XNOR U1748 ( .A(n1718), .B(n1726), .Z(n1721) );
  AND U1749 ( .A(n1168), .B(n557), .Z(n1726) );
  AND U1750 ( .A(n1727), .B(A[0]), .Z(n1718) );
  NANDN U1751 ( .B(n519), .A(n1728), .Z(n1727) );
  NAND U1752 ( .A(n1388), .B(n557), .Z(n1728) );
  XNOR U1753 ( .A(n1729), .B(X[12]), .Z(n557) );
  NAND U1754 ( .A(n1730), .B(X[15]), .Z(n1729) );
  XOR U1755 ( .A(n1731), .B(X[12]), .Z(n1730) );
  XNOR U1756 ( .A(n1172), .B(n1173), .Z(n1167) );
  NANDN U1757 ( .B(n464), .A(n1388), .Z(n1173) );
  XNOR U1758 ( .A(n1171), .B(n1733), .Z(n1172) );
  AND U1759 ( .A(n1168), .B(n488), .Z(n1733) );
  XNOR U1760 ( .A(n1725), .B(A[2]), .Z(n1724) );
  AND U1761 ( .A(n1735), .B(A[0]), .Z(n1171) );
  NAND U1762 ( .A(n1736), .B(n464), .Z(n1735) );
  NANDN U1763 ( .B(n1737), .A(n1738), .Z(n464) );
  ANDN U1764 ( .A(X[15]), .B(n1739), .Z(n1738) );
  NAND U1765 ( .A(n1388), .B(n488), .Z(n1736) );
  XOR U1766 ( .A(n1739), .B(X[14]), .Z(n1737) );
  OR U1767 ( .A(n1732), .B(n1740), .Z(n1739) );
  XOR U1768 ( .A(n1740), .B(X[13]), .Z(n1732) );
  OR U1769 ( .A(n1731), .B(n1741), .Z(n1740) );
  XOR U1770 ( .A(n1741), .B(X[12]), .Z(n1731) );
  OR U1771 ( .A(n1687), .B(n1742), .Z(n1741) );
  XOR U1772 ( .A(n1742), .B(X[11]), .Z(n1687) );
  OR U1773 ( .A(n1686), .B(n1743), .Z(n1742) );
  XOR U1774 ( .A(n1743), .B(X[10]), .Z(n1686) );
  OR U1775 ( .A(n1707), .B(n1744), .Z(n1743) );
  XOR U1776 ( .A(n1744), .B(X[9]), .Z(n1707) );
  OR U1777 ( .A(n1706), .B(n1745), .Z(n1744) );
  XOR U1778 ( .A(n1745), .B(X[8]), .Z(n1706) );
  OR U1779 ( .A(n1398), .B(n1746), .Z(n1745) );
  XOR U1780 ( .A(n1746), .B(X[7]), .Z(n1398) );
  OR U1781 ( .A(n1397), .B(n1747), .Z(n1746) );
  XOR U1782 ( .A(n1747), .B(X[6]), .Z(n1397) );
  OR U1783 ( .A(n1393), .B(n1748), .Z(n1747) );
  XOR U1784 ( .A(n1748), .B(X[5]), .Z(n1393) );
  OR U1785 ( .A(n1392), .B(n1749), .Z(n1748) );
  XOR U1786 ( .A(n1749), .B(X[4]), .Z(n1392) );
  OR U1787 ( .A(n1591), .B(n1750), .Z(n1749) );
  XOR U1788 ( .A(n1750), .B(X[3]), .Z(n1591) );
  OR U1789 ( .A(n1590), .B(n1751), .Z(n1750) );
  XOR U1790 ( .A(n1751), .B(X[2]), .Z(n1590) );
  NANDN U1791 ( .B(X[0]), .A(n1605), .Z(n1751) );
  XNOR U1792 ( .A(X[0]), .B(X[1]), .Z(n1605) );
  XOR U1793 ( .A(A[0]), .B(A[1]), .Z(n1734) );
  NANDN U1794 ( .B(n1107), .A(n379), .Z(n431) );
  IV U1795 ( .A(rst), .Z(n379) );
  NAND U1796 ( .A(n1752), .B(n1753), .Z(n1107) );
  AND U1797 ( .A(n1754), .B(n1755), .Z(n1753) );
  ANDN U1798 ( .A(n1756), .B(n[3]), .Z(n1755) );
  NOR U1799 ( .A(n[8]), .B(n[9]), .Z(n1756) );
  ANDN U1800 ( .A(n1757), .B(n[13]), .Z(n1754) );
  NOR U1801 ( .A(n[1]), .B(n[2]), .Z(n1757) );
  AND U1802 ( .A(n1758), .B(n1759), .Z(n1752) );
  ANDN U1803 ( .A(n1760), .B(n370), .Z(n1759) );
  OR U1804 ( .A(n[6]), .B(n[7]), .Z(n370) );
  NOR U1805 ( .A(n[0]), .B(n[10]), .Z(n1760) );
  NOR U1806 ( .A(n368), .B(n369), .Z(n1758) );
  OR U1807 ( .A(n[4]), .B(n[5]), .Z(n369) );
  OR U1808 ( .A(n[12]), .B(n[11]), .Z(n368) );
endmodule

