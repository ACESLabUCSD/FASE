//TEMP_H.vh

`ifndef _TEMP_H_
`define _TEMP_H_

/*simulation files*/
`define SIM	
parameter CC = 32;
parameter LOC = "/home/siam/git/hostCPU_TG/bin/scd/hw_aclrtr/hamming_32bit_32cc/";
`endif