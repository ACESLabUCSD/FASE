
module MAC_TG_N32 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MAC/AX[31] , \_MAC/AX[30] , \_MAC/AX[29] , \_MAC/AX[28] ,
         \_MAC/AX[27] , \_MAC/AX[26] , \_MAC/AX[25] , \_MAC/AX[24] ,
         \_MAC/AX[23] , \_MAC/AX[22] , \_MAC/AX[21] , \_MAC/AX[20] ,
         \_MAC/AX[19] , \_MAC/AX[18] , \_MAC/AX[17] , \_MAC/AX[16] ,
         \_MAC/AX[15] , \_MAC/AX[14] , \_MAC/AX[13] , \_MAC/AX[12] ,
         \_MAC/AX[11] , \_MAC/AX[10] , \_MAC/AX[9] , \_MAC/AX[8] ,
         \_MAC/AX[7] , \_MAC/AX[6] , \_MAC/AX[5] , \_MAC/AX[4] , \_MAC/AX[3] ,
         \_MAC/AX[2] , \_MAC/AX[1] , \_MAC/AX[0] , \_MAC/_MULT/AX__[31] ,
         \_MAC/_MULT/AX__[30] , \_MAC/_MULT/AX__[29] , \_MAC/_MULT/AX__[28] ,
         \_MAC/_MULT/AX__[27] , \_MAC/_MULT/AX__[26] , \_MAC/_MULT/AX__[25] ,
         \_MAC/_MULT/AX__[24] , \_MAC/_MULT/AX__[23] , \_MAC/_MULT/AX__[22] ,
         \_MAC/_MULT/AX__[21] , \_MAC/_MULT/AX__[20] , \_MAC/_MULT/AX__[19] ,
         \_MAC/_MULT/AX__[18] , \_MAC/_MULT/AX__[17] , \_MAC/_MULT/AX__[16] ,
         \_MAC/_MULT/AX__[15] , \_MAC/_MULT/AX__[14] , \_MAC/_MULT/AX__[13] ,
         \_MAC/_MULT/AX__[12] , \_MAC/_MULT/AX__[11] , \_MAC/_MULT/AX__[10] ,
         \_MAC/_MULT/AX__[9] , \_MAC/_MULT/AX__[8] , \_MAC/_MULT/AX__[7] ,
         \_MAC/_MULT/AX__[6] , \_MAC/_MULT/AX__[5] , \_MAC/_MULT/AX__[4] ,
         \_MAC/_MULT/AX__[3] , \_MAC/_MULT/AX__[2] , \_MAC/_MULT/AX__[1] ,
         \_MAC/_MULT/AX__[0] , \_MAC/_MULT/AX_[0] , \_MAC/_MULT/AX_[1] ,
         \_MAC/_MULT/AX_[2] , \_MAC/_MULT/AX_[3] , \_MAC/_MULT/AX_[4] ,
         \_MAC/_MULT/AX_[5] , \_MAC/_MULT/AX_[6] , \_MAC/_MULT/AX_[7] ,
         \_MAC/_MULT/AX_[8] , \_MAC/_MULT/AX_[9] , \_MAC/_MULT/AX_[10] ,
         \_MAC/_MULT/AX_[11] , \_MAC/_MULT/AX_[12] , \_MAC/_MULT/AX_[13] ,
         \_MAC/_MULT/AX_[14] , \_MAC/_MULT/AX_[15] , \_MAC/_MULT/AX_[16] ,
         \_MAC/_MULT/AX_[17] , \_MAC/_MULT/AX_[18] , \_MAC/_MULT/AX_[19] ,
         \_MAC/_MULT/AX_[20] , \_MAC/_MULT/AX_[21] , \_MAC/_MULT/AX_[22] ,
         \_MAC/_MULT/AX_[23] , \_MAC/_MULT/AX_[24] , \_MAC/_MULT/AX_[25] ,
         \_MAC/_MULT/AX_[26] , \_MAC/_MULT/AX_[27] , \_MAC/_MULT/AX_[28] ,
         \_MAC/_MULT/AX_[29] , \_MAC/_MULT/AX_[30] , \_MAC/_MULT/AX_[31] ,
         \_MAC/_MULT/X_[31] , \_MAC/_MULT/X_[30] , \_MAC/_MULT/X_[29] ,
         \_MAC/_MULT/X_[28] , \_MAC/_MULT/X_[27] , \_MAC/_MULT/X_[26] ,
         \_MAC/_MULT/X_[25] , \_MAC/_MULT/X_[24] , \_MAC/_MULT/X_[23] ,
         \_MAC/_MULT/X_[22] , \_MAC/_MULT/X_[21] , \_MAC/_MULT/X_[20] ,
         \_MAC/_MULT/X_[19] , \_MAC/_MULT/X_[18] , \_MAC/_MULT/X_[17] ,
         \_MAC/_MULT/X_[16] , \_MAC/_MULT/X_[15] , \_MAC/_MULT/X_[14] ,
         \_MAC/_MULT/X_[13] , \_MAC/_MULT/X_[12] , \_MAC/_MULT/X_[11] ,
         \_MAC/_MULT/X_[10] , \_MAC/_MULT/X_[9] , \_MAC/_MULT/X_[8] ,
         \_MAC/_MULT/X_[7] , \_MAC/_MULT/X_[6] , \_MAC/_MULT/X_[5] ,
         \_MAC/_MULT/X_[4] , \_MAC/_MULT/X_[3] , \_MAC/_MULT/X_[2] ,
         \_MAC/_MULT/X_[1] , \_MAC/_MULT/X_[0] , \_MAC/_MULT/A_[31] ,
         \_MAC/_MULT/A_[30] , \_MAC/_MULT/A_[29] , \_MAC/_MULT/A_[28] ,
         \_MAC/_MULT/A_[27] , \_MAC/_MULT/A_[26] , \_MAC/_MULT/A_[25] ,
         \_MAC/_MULT/A_[24] , \_MAC/_MULT/A_[23] , \_MAC/_MULT/A_[22] ,
         \_MAC/_MULT/A_[21] , \_MAC/_MULT/A_[20] , \_MAC/_MULT/A_[19] ,
         \_MAC/_MULT/A_[18] , \_MAC/_MULT/A_[17] , \_MAC/_MULT/A_[16] ,
         \_MAC/_MULT/A_[15] , \_MAC/_MULT/A_[14] , \_MAC/_MULT/A_[13] ,
         \_MAC/_MULT/A_[12] , \_MAC/_MULT/A_[11] , \_MAC/_MULT/A_[10] ,
         \_MAC/_MULT/A_[9] , \_MAC/_MULT/A_[8] , \_MAC/_MULT/A_[7] ,
         \_MAC/_MULT/A_[6] , \_MAC/_MULT/A_[5] , \_MAC/_MULT/A_[4] ,
         \_MAC/_MULT/A_[3] , \_MAC/_MULT/A_[2] , \_MAC/_MULT/A_[1] ,
         \_MAC/_MULT/A_[0] , \_MAC/_MULT/MULT/S[3][1][0] ,
         \_MAC/_MULT/MULT/S[3][1][1] , \_MAC/_MULT/MULT/S[3][1][2] ,
         \_MAC/_MULT/MULT/S[3][1][3] , \_MAC/_MULT/MULT/S[3][1][4] ,
         \_MAC/_MULT/MULT/S[3][1][5] , \_MAC/_MULT/MULT/S[3][1][6] ,
         \_MAC/_MULT/MULT/S[3][1][7] , \_MAC/_MULT/MULT/S[3][1][8] ,
         \_MAC/_MULT/MULT/S[3][1][9] , \_MAC/_MULT/MULT/S[3][1][10] ,
         \_MAC/_MULT/MULT/S[3][1][11] , \_MAC/_MULT/MULT/S[3][1][12] ,
         \_MAC/_MULT/MULT/S[3][1][13] , \_MAC/_MULT/MULT/S[3][1][14] ,
         \_MAC/_MULT/MULT/S[3][1][15] , \_MAC/_MULT/MULT/S[3][1][16] ,
         \_MAC/_MULT/MULT/S[3][1][17] , \_MAC/_MULT/MULT/S[3][1][18] ,
         \_MAC/_MULT/MULT/S[3][1][19] , \_MAC/_MULT/MULT/S[3][1][20] ,
         \_MAC/_MULT/MULT/S[3][1][21] , \_MAC/_MULT/MULT/S[3][1][22] ,
         \_MAC/_MULT/MULT/S[3][1][23] , \_MAC/_MULT/MULT/S[3][1][24] ,
         \_MAC/_MULT/MULT/S[3][1][25] , \_MAC/_MULT/MULT/S[3][1][26] ,
         \_MAC/_MULT/MULT/S[3][1][27] , \_MAC/_MULT/MULT/S[3][1][28] ,
         \_MAC/_MULT/MULT/S[3][1][29] , \_MAC/_MULT/MULT/S[3][1][30] ,
         \_MAC/_MULT/MULT/S[3][1][31] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[31] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[30] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[29] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[28] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[27] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[26] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[25] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[24] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[23] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[22] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[21] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[20] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[19] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[18] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[17] ,
         \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[16] , n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159;
  wire   [31:0] o_reg;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFF \o_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[0])
         );
  DFF \o_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[1])
         );
  DFF \o_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[2])
         );
  DFF \o_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[3])
         );
  DFF \o_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[4])
         );
  DFF \o_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[5])
         );
  DFF \o_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[6])
         );
  DFF \o_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[7])
         );
  DFF \o_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[8])
         );
  DFF \o_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[9])
         );
  DFF \o_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[10]) );
  DFF \o_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[11]) );
  DFF \o_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[12]) );
  DFF \o_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[13]) );
  DFF \o_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[14]) );
  DFF \o_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[15]) );
  DFF \o_reg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[16]) );
  DFF \o_reg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[17]) );
  DFF \o_reg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[18]) );
  DFF \o_reg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[19]) );
  DFF \o_reg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[20]) );
  DFF \o_reg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[21]) );
  DFF \o_reg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[22]) );
  DFF \o_reg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[23]) );
  DFF \o_reg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[24]) );
  DFF \o_reg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[25]) );
  DFF \o_reg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[26]) );
  DFF \o_reg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[27]) );
  DFF \o_reg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[28]) );
  DFF \o_reg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[29]) );
  DFF \o_reg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[30]) );
  DFF \o_reg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[31]) );
  ADD_ \_MAC/_ADD  ( .A({\_MAC/AX[31] , \_MAC/AX[30] , \_MAC/AX[29] , 
        \_MAC/AX[28] , \_MAC/AX[27] , \_MAC/AX[26] , \_MAC/AX[25] , 
        \_MAC/AX[24] , \_MAC/AX[23] , \_MAC/AX[22] , \_MAC/AX[21] , 
        \_MAC/AX[20] , \_MAC/AX[19] , \_MAC/AX[18] , \_MAC/AX[17] , 
        \_MAC/AX[16] , \_MAC/AX[15] , \_MAC/AX[14] , \_MAC/AX[13] , 
        \_MAC/AX[12] , \_MAC/AX[11] , \_MAC/AX[10] , \_MAC/AX[9] , 
        \_MAC/AX[8] , \_MAC/AX[7] , \_MAC/AX[6] , \_MAC/AX[5] , \_MAC/AX[4] , 
        \_MAC/AX[3] , \_MAC/AX[2] , \_MAC/AX[1] , \_MAC/AX[0] }), .B(o_reg), 
        .O({o, SYNOPSYS_UNCONNECTED__0}) );
  TwosComplement \_MAC/_MULT/TwosComplement_O  ( .A({\_MAC/_MULT/AX_[31] , 
        \_MAC/_MULT/AX_[30] , \_MAC/_MULT/AX_[29] , \_MAC/_MULT/AX_[28] , 
        \_MAC/_MULT/AX_[27] , \_MAC/_MULT/AX_[26] , \_MAC/_MULT/AX_[25] , 
        \_MAC/_MULT/AX_[24] , \_MAC/_MULT/AX_[23] , \_MAC/_MULT/AX_[22] , 
        \_MAC/_MULT/AX_[21] , \_MAC/_MULT/AX_[20] , \_MAC/_MULT/AX_[19] , 
        \_MAC/_MULT/AX_[18] , \_MAC/_MULT/AX_[17] , \_MAC/_MULT/AX_[16] , 
        \_MAC/_MULT/AX_[15] , \_MAC/_MULT/AX_[14] , \_MAC/_MULT/AX_[13] , 
        \_MAC/_MULT/AX_[12] , \_MAC/_MULT/AX_[11] , \_MAC/_MULT/AX_[10] , 
        \_MAC/_MULT/AX_[9] , \_MAC/_MULT/AX_[8] , \_MAC/_MULT/AX_[7] , 
        \_MAC/_MULT/AX_[6] , \_MAC/_MULT/AX_[5] , \_MAC/_MULT/AX_[4] , 
        \_MAC/_MULT/AX_[3] , \_MAC/_MULT/AX_[2] , \_MAC/_MULT/AX_[1] , 
        \_MAC/_MULT/AX_[0] }), .O({\_MAC/_MULT/AX__[31] , 
        \_MAC/_MULT/AX__[30] , \_MAC/_MULT/AX__[29] , \_MAC/_MULT/AX__[28] , 
        \_MAC/_MULT/AX__[27] , \_MAC/_MULT/AX__[26] , \_MAC/_MULT/AX__[25] , 
        \_MAC/_MULT/AX__[24] , \_MAC/_MULT/AX__[23] , \_MAC/_MULT/AX__[22] , 
        \_MAC/_MULT/AX__[21] , \_MAC/_MULT/AX__[20] , \_MAC/_MULT/AX__[19] , 
        \_MAC/_MULT/AX__[18] , \_MAC/_MULT/AX__[17] , \_MAC/_MULT/AX__[16] , 
        \_MAC/_MULT/AX__[15] , \_MAC/_MULT/AX__[14] , \_MAC/_MULT/AX__[13] , 
        \_MAC/_MULT/AX__[12] , \_MAC/_MULT/AX__[11] , \_MAC/_MULT/AX__[10] , 
        \_MAC/_MULT/AX__[9] , \_MAC/_MULT/AX__[8] , \_MAC/_MULT/AX__[7] , 
        \_MAC/_MULT/AX__[6] , \_MAC/_MULT/AX__[5] , \_MAC/_MULT/AX__[4] , 
        \_MAC/_MULT/AX__[3] , \_MAC/_MULT/AX__[2] , \_MAC/_MULT/AX__[1] , 
        \_MAC/_MULT/AX__[0] }) );
  TwosComplement \_MAC/_MULT/TwosComplement_B  ( .A(e_input), .O({
        \_MAC/_MULT/X_[31] , \_MAC/_MULT/X_[30] , \_MAC/_MULT/X_[29] , 
        \_MAC/_MULT/X_[28] , \_MAC/_MULT/X_[27] , \_MAC/_MULT/X_[26] , 
        \_MAC/_MULT/X_[25] , \_MAC/_MULT/X_[24] , \_MAC/_MULT/X_[23] , 
        \_MAC/_MULT/X_[22] , \_MAC/_MULT/X_[21] , \_MAC/_MULT/X_[20] , 
        \_MAC/_MULT/X_[19] , \_MAC/_MULT/X_[18] , \_MAC/_MULT/X_[17] , 
        \_MAC/_MULT/X_[16] , \_MAC/_MULT/X_[15] , \_MAC/_MULT/X_[14] , 
        \_MAC/_MULT/X_[13] , \_MAC/_MULT/X_[12] , \_MAC/_MULT/X_[11] , 
        \_MAC/_MULT/X_[10] , \_MAC/_MULT/X_[9] , \_MAC/_MULT/X_[8] , 
        \_MAC/_MULT/X_[7] , \_MAC/_MULT/X_[6] , \_MAC/_MULT/X_[5] , 
        \_MAC/_MULT/X_[4] , \_MAC/_MULT/X_[3] , \_MAC/_MULT/X_[2] , 
        \_MAC/_MULT/X_[1] , \_MAC/_MULT/X_[0] }) );
  TwosComplement \_MAC/_MULT/TwosComplement_A  ( .A(g_input), .O({
        \_MAC/_MULT/A_[31] , \_MAC/_MULT/A_[30] , \_MAC/_MULT/A_[29] , 
        \_MAC/_MULT/A_[28] , \_MAC/_MULT/A_[27] , \_MAC/_MULT/A_[26] , 
        \_MAC/_MULT/A_[25] , \_MAC/_MULT/A_[24] , \_MAC/_MULT/A_[23] , 
        \_MAC/_MULT/A_[22] , \_MAC/_MULT/A_[21] , \_MAC/_MULT/A_[20] , 
        \_MAC/_MULT/A_[19] , \_MAC/_MULT/A_[18] , \_MAC/_MULT/A_[17] , 
        \_MAC/_MULT/A_[16] , \_MAC/_MULT/A_[15] , \_MAC/_MULT/A_[14] , 
        \_MAC/_MULT/A_[13] , \_MAC/_MULT/A_[12] , \_MAC/_MULT/A_[11] , 
        \_MAC/_MULT/A_[10] , \_MAC/_MULT/A_[9] , \_MAC/_MULT/A_[8] , 
        \_MAC/_MULT/A_[7] , \_MAC/_MULT/A_[6] , \_MAC/_MULT/A_[5] , 
        \_MAC/_MULT/A_[4] , \_MAC/_MULT/A_[3] , \_MAC/_MULT/A_[2] , 
        \_MAC/_MULT/A_[1] , \_MAC/_MULT/A_[0] }) );
  XOR \_MAC/_MULT/MUX_O/U94  ( .A(\_MAC/_MULT/AX_[0] ), .B(n5159), .Z(
        \_MAC/AX[0] ) );
  XOR \_MAC/_MULT/MUX_O/U91  ( .A(\_MAC/_MULT/AX_[10] ), .B(n5158), .Z(
        \_MAC/AX[10] ) );
  XOR \_MAC/_MULT/MUX_O/U88  ( .A(\_MAC/_MULT/AX_[11] ), .B(n5157), .Z(
        \_MAC/AX[11] ) );
  XOR \_MAC/_MULT/MUX_O/U85  ( .A(\_MAC/_MULT/AX_[12] ), .B(n5156), .Z(
        \_MAC/AX[12] ) );
  XOR \_MAC/_MULT/MUX_O/U82  ( .A(\_MAC/_MULT/AX_[13] ), .B(n5155), .Z(
        \_MAC/AX[13] ) );
  XOR \_MAC/_MULT/MUX_O/U79  ( .A(\_MAC/_MULT/AX_[14] ), .B(n5154), .Z(
        \_MAC/AX[14] ) );
  XOR \_MAC/_MULT/MUX_O/U76  ( .A(\_MAC/_MULT/AX_[15] ), .B(n5153), .Z(
        \_MAC/AX[15] ) );
  XOR \_MAC/_MULT/MUX_O/U73  ( .A(\_MAC/_MULT/AX_[16] ), .B(n5152), .Z(
        \_MAC/AX[16] ) );
  XOR \_MAC/_MULT/MUX_O/U70  ( .A(\_MAC/_MULT/AX_[17] ), .B(n5151), .Z(
        \_MAC/AX[17] ) );
  XOR \_MAC/_MULT/MUX_O/U67  ( .A(\_MAC/_MULT/AX_[18] ), .B(n5150), .Z(
        \_MAC/AX[18] ) );
  XOR \_MAC/_MULT/MUX_O/U64  ( .A(\_MAC/_MULT/AX_[19] ), .B(n5149), .Z(
        \_MAC/AX[19] ) );
  XOR \_MAC/_MULT/MUX_O/U61  ( .A(\_MAC/_MULT/AX_[1] ), .B(n5148), .Z(
        \_MAC/AX[1] ) );
  XOR \_MAC/_MULT/MUX_O/U58  ( .A(\_MAC/_MULT/AX_[20] ), .B(n5147), .Z(
        \_MAC/AX[20] ) );
  XOR \_MAC/_MULT/MUX_O/U55  ( .A(\_MAC/_MULT/AX_[21] ), .B(n5146), .Z(
        \_MAC/AX[21] ) );
  XOR \_MAC/_MULT/MUX_O/U52  ( .A(\_MAC/_MULT/AX_[22] ), .B(n5145), .Z(
        \_MAC/AX[22] ) );
  XOR \_MAC/_MULT/MUX_O/U49  ( .A(\_MAC/_MULT/AX_[23] ), .B(n5144), .Z(
        \_MAC/AX[23] ) );
  XOR \_MAC/_MULT/MUX_O/U46  ( .A(\_MAC/_MULT/AX_[24] ), .B(n5143), .Z(
        \_MAC/AX[24] ) );
  XOR \_MAC/_MULT/MUX_O/U43  ( .A(\_MAC/_MULT/AX_[25] ), .B(n5142), .Z(
        \_MAC/AX[25] ) );
  XOR \_MAC/_MULT/MUX_O/U40  ( .A(\_MAC/_MULT/AX_[26] ), .B(n5141), .Z(
        \_MAC/AX[26] ) );
  XOR \_MAC/_MULT/MUX_O/U37  ( .A(\_MAC/_MULT/AX_[27] ), .B(n5140), .Z(
        \_MAC/AX[27] ) );
  XOR \_MAC/_MULT/MUX_O/U34  ( .A(\_MAC/_MULT/AX_[28] ), .B(n5139), .Z(
        \_MAC/AX[28] ) );
  XOR \_MAC/_MULT/MUX_O/U31  ( .A(\_MAC/_MULT/AX_[29] ), .B(n5138), .Z(
        \_MAC/AX[29] ) );
  XOR \_MAC/_MULT/MUX_O/U28  ( .A(\_MAC/_MULT/AX_[2] ), .B(n5137), .Z(
        \_MAC/AX[2] ) );
  XOR \_MAC/_MULT/MUX_O/U25  ( .A(\_MAC/_MULT/AX_[30] ), .B(n5136), .Z(
        \_MAC/AX[30] ) );
  XOR \_MAC/_MULT/MUX_O/U22  ( .A(\_MAC/_MULT/AX_[31] ), .B(n5135), .Z(
        \_MAC/AX[31] ) );
  XOR \_MAC/_MULT/MUX_O/U19  ( .A(\_MAC/_MULT/AX_[3] ), .B(n5134), .Z(
        \_MAC/AX[3] ) );
  XOR \_MAC/_MULT/MUX_O/U16  ( .A(\_MAC/_MULT/AX_[4] ), .B(n5133), .Z(
        \_MAC/AX[4] ) );
  XOR \_MAC/_MULT/MUX_O/U13  ( .A(\_MAC/_MULT/AX_[5] ), .B(n5132), .Z(
        \_MAC/AX[5] ) );
  XOR \_MAC/_MULT/MUX_O/U10  ( .A(\_MAC/_MULT/AX_[6] ), .B(n5131), .Z(
        \_MAC/AX[6] ) );
  XOR \_MAC/_MULT/MUX_O/U7  ( .A(\_MAC/_MULT/AX_[7] ), .B(n5130), .Z(
        \_MAC/AX[7] ) );
  XOR \_MAC/_MULT/MUX_O/U4  ( .A(\_MAC/_MULT/AX_[8] ), .B(n5129), .Z(
        \_MAC/AX[8] ) );
  XOR \_MAC/_MULT/MUX_O/U1  ( .A(\_MAC/_MULT/AX_[9] ), .B(n5128), .Z(
        \_MAC/AX[9] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[31].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][31] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[31] ), .Z(
        \_MAC/_MULT/AX_[31] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[30].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][30] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[30] ), .Z(
        \_MAC/_MULT/AX_[30] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[29].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][29] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[29] ), .Z(
        \_MAC/_MULT/AX_[29] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[28].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][28] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[28] ), .Z(
        \_MAC/_MULT/AX_[28] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[27].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][27] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[27] ), .Z(
        \_MAC/_MULT/AX_[27] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[26].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][26] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[26] ), .Z(
        \_MAC/_MULT/AX_[26] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[25].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][25] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[25] ), .Z(
        \_MAC/_MULT/AX_[25] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[24].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][24] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[24] ), .Z(
        \_MAC/_MULT/AX_[24] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[23].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][23] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[23] ), .Z(
        \_MAC/_MULT/AX_[23] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[22].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][22] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[22] ), .Z(
        \_MAC/_MULT/AX_[22] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[21].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][21] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[21] ), .Z(
        \_MAC/_MULT/AX_[21] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[20].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][20] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[20] ), .Z(
        \_MAC/_MULT/AX_[20] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[19].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][19] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[19] ), .Z(
        \_MAC/_MULT/AX_[19] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[18].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][18] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[18] ), .Z(
        \_MAC/_MULT/AX_[18] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[17].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][17] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[17] ), .Z(
        \_MAC/_MULT/AX_[17] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[16].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][16] ), .B(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[16] ), .Z(
        \_MAC/_MULT/AX_[16] ) );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[15].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][15] ), .B(n5127), .Z(\_MAC/_MULT/AX_[15] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[14].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][14] ), .B(n5126), .Z(\_MAC/_MULT/AX_[14] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[13].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][13] ), .B(n5125), .Z(\_MAC/_MULT/AX_[13] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[12].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][12] ), .B(n5124), .Z(\_MAC/_MULT/AX_[12] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[11].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][11] ), .B(n5123), .Z(\_MAC/_MULT/AX_[11] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[10].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][10] ), .B(n5122), .Z(\_MAC/_MULT/AX_[10] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[9].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][9] ), .B(n5121), .Z(\_MAC/_MULT/AX_[9] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[8].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][8] ), .B(n5120), .Z(\_MAC/_MULT/AX_[8] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[7].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][7] ), .B(n5119), .Z(\_MAC/_MULT/AX_[7] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[6].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][6] ), .B(n5118), .Z(\_MAC/_MULT/AX_[6] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[5].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][5] ), .B(n5117), .Z(\_MAC/_MULT/AX_[5] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[4].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][4] ), .B(n5116), .Z(\_MAC/_MULT/AX_[4] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[3].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][3] ), .B(n5115), .Z(\_MAC/_MULT/AX_[3] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[2].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][2] ), .B(n5114), .Z(\_MAC/_MULT/AX_[2] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[1].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][1] ), .B(n5113), .Z(\_MAC/_MULT/AX_[1] )
         );
  XOR \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[0].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[3][1][0] ), .B(n5112), .Z(\_MAC/_MULT/AX_[0] )
         );
  MUX U35 ( .IN0(n2496), .IN1(n33), .SEL(n2497), .F(n2485) );
  IV U36 ( .A(n2498), .Z(n33) );
  MUX U37 ( .IN0(n2002), .IN1(n34), .SEL(n2003), .F(n1961) );
  IV U38 ( .A(n2004), .Z(n34) );
  MUX U39 ( .IN0(n1984), .IN1(n35), .SEL(n1985), .F(n1943) );
  IV U40 ( .A(n1986), .Z(n35) );
  XNOR U41 ( .A(n2284), .B(n2270), .Z(n2274) );
  XNOR U42 ( .A(n1818), .B(n1782), .Z(n1786) );
  XNOR U43 ( .A(n2216), .B(n2202), .Z(n2206) );
  MUX U44 ( .IN0(n2769), .IN1(n36), .SEL(n2770), .F(n2758) );
  IV U45 ( .A(n2771), .Z(n36) );
  MUX U46 ( .IN0(n2643), .IN1(n2645), .SEL(n2644), .F(n2622) );
  MUX U47 ( .IN0(n4869), .IN1(n37), .SEL(n4870), .F(n4856) );
  IV U48 ( .A(n4871), .Z(n37) );
  MUX U49 ( .IN0(n4744), .IN1(n4746), .SEL(n4745), .F(n4723) );
  MUX U50 ( .IN0(n1668), .IN1(n38), .SEL(n1669), .F(n1629) );
  IV U51 ( .A(n1670), .Z(n38) );
  MUX U52 ( .IN0(n1586), .IN1(n39), .SEL(n1587), .F(n1547) );
  IV U53 ( .A(n1588), .Z(n39) );
  MUX U54 ( .IN0(n2751), .IN1(n2608), .SEL(n2610), .F(n2740) );
  MUX U55 ( .IN0(n2576), .IN1(n40), .SEL(n2577), .F(n2555) );
  IV U56 ( .A(n2578), .Z(n40) );
  MUX U57 ( .IN0(n5051), .IN1(n41), .SEL(n5052), .F(n5034) );
  IV U58 ( .A(n5053), .Z(n41) );
  MUX U59 ( .IN0(n4677), .IN1(n42), .SEL(n4678), .F(n4656) );
  IV U60 ( .A(n4679), .Z(n42) );
  MUX U61 ( .IN0(n4847), .IN1(n4688), .SEL(n4690), .F(n4834) );
  XNOR U62 ( .A(n2358), .B(n2350), .Z(n2112) );
  MUX U63 ( .IN0(n2103), .IN1(n43), .SEL(n2104), .F(n2086) );
  IV U64 ( .A(n2105), .Z(n43) );
  MUX U65 ( .IN0(n4167), .IN1(n44), .SEL(n4168), .F(n4150) );
  IV U66 ( .A(n4169), .Z(n44) );
  MUX U67 ( .IN0(n4560), .IN1(n45), .SEL(n4561), .F(n4551) );
  IV U68 ( .A(n4562), .Z(n45) );
  MUX U69 ( .IN0(n1241), .IN1(n46), .SEL(n1242), .F(n1188) );
  IV U70 ( .A(n1243), .Z(n46) );
  MUX U71 ( .IN0(n4227), .IN1(n47), .SEL(n4228), .F(n4214) );
  IV U72 ( .A(n4229), .Z(n47) );
  MUX U73 ( .IN0(n938), .IN1(n48), .SEL(n939), .F(n908) );
  IV U74 ( .A(n940), .Z(n48) );
  MUX U75 ( .IN0(n3915), .IN1(n49), .SEL(n3916), .F(n3849) );
  IV U76 ( .A(n3917), .Z(n49) );
  MUX U77 ( .IN0(n3743), .IN1(n50), .SEL(n3744), .F(n3677) );
  IV U78 ( .A(n3745), .Z(n50) );
  MUX U79 ( .IN0(n3498), .IN1(n51), .SEL(n3499), .F(n3439) );
  IV U80 ( .A(n3500), .Z(n51) );
  MUX U81 ( .IN0(n3363), .IN1(n52), .SEL(n3364), .F(n3313) );
  IV U82 ( .A(n3365), .Z(n52) );
  MUX U83 ( .IN0(n1370), .IN1(n53), .SEL(n1371), .F(n1308) );
  IV U84 ( .A(n1372), .Z(n53) );
  MUX U85 ( .IN0(n4457), .IN1(n54), .SEL(n4358), .F(n4446) );
  IV U86 ( .A(n4357), .Z(n54) );
  MUX U87 ( .IN0(n1236), .IN1(n55), .SEL(n1237), .F(n1183) );
  IV U88 ( .A(n1238), .Z(n55) );
  MUX U89 ( .IN0(n4528), .IN1(n56), .SEL(n4342), .F(n4519) );
  IV U90 ( .A(n4341), .Z(n56) );
  MUX U91 ( .IN0(n4413), .IN1(n57), .SEL(n4334), .F(n4402) );
  IV U92 ( .A(n4333), .Z(n57) );
  MUX U93 ( .IN0(n1207), .IN1(n58), .SEL(n1208), .F(n1154) );
  IV U94 ( .A(n1209), .Z(n58) );
  MUX U95 ( .IN0(n1045), .IN1(n59), .SEL(n1046), .F(n1008) );
  IV U96 ( .A(n1047), .Z(n59) );
  MUX U97 ( .IN0(n4035), .IN1(n60), .SEL(n4036), .F(n3959) );
  IV U98 ( .A(n4037), .Z(n60) );
  MUX U99 ( .IN0(n3936), .IN1(n61), .SEL(n3937), .F(n3870) );
  IV U100 ( .A(n3938), .Z(n61) );
  MUX U101 ( .IN0(n3761), .IN1(n62), .SEL(n3762), .F(n3695) );
  IV U102 ( .A(n3763), .Z(n62) );
  MUX U103 ( .IN0(n881), .IN1(n63), .SEL(n882), .F(n859) );
  IV U104 ( .A(n883), .Z(n63) );
  MUX U105 ( .IN0(n3616), .IN1(n64), .SEL(n3617), .F(n3552) );
  IV U106 ( .A(n3618), .Z(n64) );
  MUX U107 ( .IN0(n3384), .IN1(n65), .SEL(n3385), .F(n3331) );
  IV U108 ( .A(n3386), .Z(n65) );
  MUX U109 ( .IN0(n3086), .IN1(n66), .SEL(n3087), .F(n3056) );
  IV U110 ( .A(n3088), .Z(n66) );
  MUX U111 ( .IN0(n4349), .IN1(n67), .SEL(n4004), .F(n4343) );
  IV U112 ( .A(n4003), .Z(n67) );
  MUX U113 ( .IN0(n1174), .IN1(n68), .SEL(n1175), .F(n1122) );
  IV U114 ( .A(n1176), .Z(n68) );
  MUX U115 ( .IN0(n4319), .IN1(n69), .SEL(n3974), .F(n4313) );
  IV U116 ( .A(n3973), .Z(n69) );
  MUX U117 ( .IN0(n929), .IN1(n70), .SEL(n930), .F(n902) );
  IV U118 ( .A(n931), .Z(n70) );
  MUX U119 ( .IN0(n3206), .IN1(n71), .SEL(n3207), .F(n3160) );
  IV U120 ( .A(n3208), .Z(n71) );
  MUX U121 ( .IN0(n1066), .IN1(n72), .SEL(n1067), .F(n1016) );
  IV U122 ( .A(n1068), .Z(n72) );
  MUX U123 ( .IN0(n2045), .IN1(n73), .SEL(n2046), .F(n2002) );
  IV U124 ( .A(n2047), .Z(n73) );
  XNOR U125 ( .A(n2490), .B(n2482), .Z(n2320) );
  XNOR U126 ( .A(n1976), .B(n1940), .Z(n1944) );
  XNOR U127 ( .A(n2267), .B(n2253), .Z(n2257) );
  XNOR U128 ( .A(n1959), .B(n1923), .Z(n1927) );
  XNOR U129 ( .A(n2457), .B(n2449), .Z(n2265) );
  MUX U130 ( .IN0(n1824), .IN1(n74), .SEL(n1825), .F(n1785) );
  IV U131 ( .A(n1826), .Z(n74) );
  MUX U132 ( .IN0(n1742), .IN1(n75), .SEL(n1743), .F(n1703) );
  IV U133 ( .A(n1744), .Z(n75) );
  XNOR U134 ( .A(n1840), .B(n1804), .Z(n1808) );
  XNOR U135 ( .A(n2778), .B(n2770), .Z(n2652) );
  MUX U136 ( .IN0(n2666), .IN1(n76), .SEL(n2667), .F(n2643) );
  IV U137 ( .A(n2668), .Z(n76) );
  MUX U138 ( .IN0(n4767), .IN1(n77), .SEL(n4768), .F(n4744) );
  IV U139 ( .A(n4769), .Z(n77) );
  XNOR U140 ( .A(n2182), .B(n2168), .Z(n2172) );
  XNOR U141 ( .A(n2402), .B(n2394), .Z(n2180) );
  XNOR U142 ( .A(n4878), .B(n4870), .Z(n4732) );
  XNOR U143 ( .A(n1684), .B(n1648), .Z(n1652) );
  MUX U144 ( .IN0(n4974), .IN1(n78), .SEL(n4975), .F(n4970) );
  IV U145 ( .A(n4976), .Z(n78) );
  MUX U146 ( .IN0(n1590), .IN1(n79), .SEL(n1591), .F(n1551) );
  IV U147 ( .A(n1592), .Z(n79) );
  XNOR U148 ( .A(n2131), .B(n2117), .Z(n2121) );
  MUX U149 ( .IN0(n2740), .IN1(n2587), .SEL(n2589), .F(n2729) );
  MUX U150 ( .IN0(n2580), .IN1(n2582), .SEL(n2581), .F(n2559) );
  MUX U151 ( .IN0(n4681), .IN1(n4683), .SEL(n4682), .F(n4660) );
  XNOR U152 ( .A(n1567), .B(n1531), .Z(n1535) );
  XNOR U153 ( .A(n2347), .B(n2339), .Z(n2095) );
  MUX U154 ( .IN0(n4821), .IN1(n4646), .SEL(n4648), .F(n4808) );
  MUX U155 ( .IN0(n2069), .IN1(n80), .SEL(n2070), .F(n1452) );
  IV U156 ( .A(n2071), .Z(n80) );
  MUX U157 ( .IN0(n1381), .IN1(n81), .SEL(n1382), .F(n1319) );
  IV U158 ( .A(n1383), .Z(n81) );
  MUX U159 ( .IN0(n4150), .IN1(n82), .SEL(n4151), .F(n4133) );
  IV U160 ( .A(n4152), .Z(n82) );
  MUX U161 ( .IN0(n4266), .IN1(n83), .SEL(n4267), .F(n4253) );
  IV U162 ( .A(n4268), .Z(n83) );
  MUX U163 ( .IN0(n1179), .IN1(n84), .SEL(n1180), .F(n1127) );
  IV U164 ( .A(n1181), .Z(n84) );
  MUX U165 ( .IN0(n1136), .IN1(n85), .SEL(n1137), .F(n1090) );
  IV U166 ( .A(n1138), .Z(n85) );
  MUX U167 ( .IN0(n4409), .IN1(n86), .SEL(n4410), .F(n4398) );
  IV U168 ( .A(n4411), .Z(n86) );
  MUX U169 ( .IN0(n4065), .IN1(n87), .SEL(n4066), .F(n4048) );
  IV U170 ( .A(n4067), .Z(n87) );
  MUX U171 ( .IN0(n4504), .IN1(n88), .SEL(n4505), .F(n4493) );
  IV U172 ( .A(n4506), .Z(n88) );
  MUX U173 ( .IN0(n89), .IN1(n947), .SEL(n948), .F(n917) );
  IV U174 ( .A(n949), .Z(n89) );
  MUX U175 ( .IN0(n3875), .IN1(n90), .SEL(n3876), .F(n3809) );
  IV U176 ( .A(n3877), .Z(n90) );
  MUX U177 ( .IN0(n91), .IN1(n3831), .SEL(n3832), .F(n3765) );
  IV U178 ( .A(n3833), .Z(n91) );
  MUX U179 ( .IN0(n3668), .IN1(n92), .SEL(n3669), .F(n3603) );
  IV U180 ( .A(n3670), .Z(n92) );
  MUX U181 ( .IN0(n3651), .IN1(n93), .SEL(n3652), .F(n3585) );
  IV U182 ( .A(n3653), .Z(n93) );
  MUX U183 ( .IN0(n3439), .IN1(n94), .SEL(n3440), .F(n3380) );
  IV U184 ( .A(n3441), .Z(n94) );
  MUX U185 ( .IN0(n3416), .IN1(n95), .SEL(n3417), .F(n3354) );
  IV U186 ( .A(n3418), .Z(n95) );
  MUX U187 ( .IN0(n3313), .IN1(n96), .SEL(n3314), .F(n3264) );
  IV U188 ( .A(n3315), .Z(n96) );
  MUX U189 ( .IN0(n3212), .IN1(n97), .SEL(n3213), .F(n3164) );
  IV U190 ( .A(n3214), .Z(n97) );
  MUX U191 ( .IN0(n4575), .IN1(n98), .SEL(n4576), .F(n4566) );
  IV U192 ( .A(n4577), .Z(n98) );
  MUX U193 ( .IN0(n4171), .IN1(n99), .SEL(n4172), .F(n4154) );
  IV U194 ( .A(n4173), .Z(n99) );
  MUX U195 ( .IN0(n4470), .IN1(n100), .SEL(n4364), .F(n4457) );
  IV U196 ( .A(n4363), .Z(n100) );
  MUX U197 ( .IN0(n1245), .IN1(n101), .SEL(n1246), .F(n1192) );
  IV U198 ( .A(n1247), .Z(n101) );
  MUX U199 ( .IN0(n1261), .IN1(n102), .SEL(n1262), .F(n1207) );
  IV U200 ( .A(n1263), .Z(n102) );
  MUX U201 ( .IN0(n4537), .IN1(n103), .SEL(n4348), .F(n4528) );
  IV U202 ( .A(n4347), .Z(n103) );
  MUX U203 ( .IN0(n4103), .IN1(n104), .SEL(n4104), .F(n4086) );
  IV U204 ( .A(n4105), .Z(n104) );
  MUX U205 ( .IN0(n4244), .IN1(n105), .SEL(n4112), .F(n4231) );
  IV U206 ( .A(n4111), .Z(n105) );
  MUX U207 ( .IN0(n1036), .IN1(n106), .SEL(n1037), .F(n999) );
  IV U208 ( .A(n1038), .Z(n106) );
  MUX U209 ( .IN0(n1008), .IN1(n107), .SEL(n1009), .F(n973) );
  IV U210 ( .A(n1010), .Z(n107) );
  MUX U211 ( .IN0(n4391), .IN1(n108), .SEL(n4322), .F(n4378) );
  IV U212 ( .A(n4321), .Z(n108) );
  MUX U213 ( .IN0(n4490), .IN1(n109), .SEL(n4318), .F(n3945) );
  IV U214 ( .A(n4317), .Z(n109) );
  MUX U215 ( .IN0(n3959), .IN1(n110), .SEL(n3960), .F(n3893) );
  IV U216 ( .A(n3961), .Z(n110) );
  MUX U217 ( .IN0(n4192), .IN1(n111), .SEL(n4044), .F(n3919) );
  IV U218 ( .A(n4043), .Z(n111) );
  MUX U219 ( .IN0(n3804), .IN1(n112), .SEL(n3805), .F(n3738) );
  IV U220 ( .A(n3806), .Z(n112) );
  MUX U221 ( .IN0(n3747), .IN1(n113), .SEL(n3748), .F(n3681) );
  IV U222 ( .A(n3749), .Z(n113) );
  MUX U223 ( .IN0(n3630), .IN1(n114), .SEL(n3631), .F(n3566) );
  IV U224 ( .A(n3632), .Z(n114) );
  MUX U225 ( .IN0(n876), .IN1(n115), .SEL(n877), .F(n857) );
  IV U226 ( .A(n878), .Z(n115) );
  MUX U227 ( .IN0(n3543), .IN1(n116), .SEL(n3544), .F(n3479) );
  IV U228 ( .A(n3545), .Z(n116) );
  MUX U229 ( .IN0(n3488), .IN1(n117), .SEL(n3489), .F(n3429) );
  IV U230 ( .A(n3490), .Z(n117) );
  MUX U231 ( .IN0(n3308), .IN1(n118), .SEL(n3309), .F(n3259) );
  IV U232 ( .A(n3310), .Z(n118) );
  MUX U233 ( .IN0(n3331), .IN1(n119), .SEL(n3332), .F(n3281) );
  IV U234 ( .A(n3333), .Z(n119) );
  MUX U235 ( .IN0(n3225), .IN1(n120), .SEL(n3226), .F(n3178) );
  IV U236 ( .A(n3227), .Z(n120) );
  XNOR U237 ( .A(n1355), .B(n1296), .Z(n1300) );
  MUX U238 ( .IN0(n4355), .IN1(n121), .SEL(n4010), .F(n4349) );
  IV U239 ( .A(n4009), .Z(n121) );
  MUX U240 ( .IN0(n1076), .IN1(n122), .SEL(n1077), .F(n1026) );
  IV U241 ( .A(n1078), .Z(n122) );
  MUX U242 ( .IN0(n4331), .IN1(n123), .SEL(n3986), .F(n4325) );
  IV U243 ( .A(n3985), .Z(n123) );
  MUX U244 ( .IN0(n3861), .IN1(n124), .SEL(n3862), .F(n3795) );
  IV U245 ( .A(n3863), .Z(n124) );
  MUX U246 ( .IN0(n3349), .IN1(n125), .SEL(n3350), .F(n3299) );
  IV U247 ( .A(n3351), .Z(n125) );
  MUX U248 ( .IN0(n3100), .IN1(n126), .SEL(n3101), .F(n3076) );
  IV U249 ( .A(n3102), .Z(n126) );
  MUX U250 ( .IN0(n3056), .IN1(n127), .SEL(n3057), .F(n3037) );
  IV U251 ( .A(n3058), .Z(n127) );
  MUX U252 ( .IN0(n1268), .IN1(n128), .SEL(n1269), .F(n1214) );
  IV U253 ( .A(n1270), .Z(n128) );
  ANDN U254 ( .A(n891), .B(n892), .Z(n870) );
  MUX U255 ( .IN0(n3242), .IN1(n129), .SEL(n3243), .F(n3198) );
  IV U256 ( .A(n3244), .Z(n129) );
  XNOR U257 ( .A(n1016), .B(n1064), .Z(n1053) );
  ANDN U258 ( .A(n3045), .B(\_MAC/_MULT/MULT/S[3][1][28] ), .Z(n3028) );
  MUX U259 ( .IN0(n2485), .IN1(n130), .SEL(n2320), .F(n2474) );
  IV U260 ( .A(n2319), .Z(n130) );
  MUX U261 ( .IN0(n2481), .IN1(n131), .SEL(n2482), .F(n2470) );
  IV U262 ( .A(n2483), .Z(n131) );
  XNOR U263 ( .A(n2043), .B(n2003), .Z(n2007) );
  MUX U264 ( .IN0(n1943), .IN1(n132), .SEL(n1944), .F(n1904) );
  IV U265 ( .A(n1945), .Z(n132) );
  MUX U266 ( .IN0(n1900), .IN1(n133), .SEL(n1901), .F(n1859) );
  IV U267 ( .A(n1902), .Z(n133) );
  XNOR U268 ( .A(n2250), .B(n2236), .Z(n2240) );
  XNOR U269 ( .A(n1920), .B(n1884), .Z(n1888) );
  XNOR U270 ( .A(n2435), .B(n2427), .Z(n2231) );
  MUX U271 ( .IN0(n1746), .IN1(n134), .SEL(n1747), .F(n1707) );
  IV U272 ( .A(n1748), .Z(n134) );
  XNOR U273 ( .A(n2199), .B(n2185), .Z(n2189) );
  XNOR U274 ( .A(n1801), .B(n1765), .Z(n1769) );
  MUX U275 ( .IN0(n2764), .IN1(n135), .SEL(n2765), .F(n2753) );
  IV U276 ( .A(n2766), .Z(n135) );
  MUX U277 ( .IN0(n2758), .IN1(n136), .SEL(n2759), .F(n2747) );
  IV U278 ( .A(n2760), .Z(n136) );
  MUX U279 ( .IN0(n4886), .IN1(n4751), .SEL(n4753), .F(n4873) );
  XNOR U280 ( .A(n4761), .B(n4741), .Z(n4745) );
  XNOR U281 ( .A(n4715), .B(n4716), .Z(n4725) );
  MUX U282 ( .IN0(n2397), .IN1(n137), .SEL(n2180), .F(n2386) );
  IV U283 ( .A(n2179), .Z(n137) );
  XNOR U284 ( .A(n2637), .B(n2619), .Z(n2623) );
  MUX U285 ( .IN0(n4856), .IN1(n138), .SEL(n4857), .F(n4843) );
  IV U286 ( .A(n4858), .Z(n138) );
  XNOR U287 ( .A(n2148), .B(n2134), .Z(n2138) );
  XNOR U288 ( .A(n1645), .B(n1609), .Z(n1613) );
  MUX U289 ( .IN0(n2951), .IN1(n139), .SEL(n2952), .F(n2947) );
  IV U290 ( .A(n2953), .Z(n139) );
  MUX U291 ( .IN0(n1551), .IN1(n140), .SEL(n1552), .F(n1512) );
  IV U292 ( .A(n1553), .Z(n140) );
  MUX U293 ( .IN0(n2729), .IN1(n2566), .SEL(n2568), .F(n2718) );
  MUX U294 ( .IN0(n2559), .IN1(n2561), .SEL(n2560), .F(n2538) );
  MUX U295 ( .IN0(n4834), .IN1(n4667), .SEL(n4669), .F(n4821) );
  MUX U296 ( .IN0(n4660), .IN1(n4662), .SEL(n4661), .F(n4639) );
  MUX U297 ( .IN0(n141), .IN1(n1478), .SEL(n1479), .F(n1442) );
  IV U298 ( .A(n1480), .Z(n141) );
  MUX U299 ( .IN0(n2086), .IN1(n142), .SEL(n2087), .F(n2069) );
  IV U300 ( .A(n2088), .Z(n142) );
  MUX U301 ( .IN0(n4804), .IN1(n143), .SEL(n4805), .F(n4301) );
  IV U302 ( .A(n4806), .Z(n143) );
  MUX U303 ( .IN0(n1433), .IN1(n144), .SEL(n1434), .F(n1366) );
  IV U304 ( .A(n1435), .Z(n144) );
  MUX U305 ( .IN0(n1448), .IN1(n145), .SEL(n1449), .F(n1381) );
  IV U306 ( .A(n1450), .Z(n145) );
  XNOR U307 ( .A(n2335), .B(n2326), .Z(n2078) );
  MUX U308 ( .IN0(n4551), .IN1(n146), .SEL(n4552), .F(n4540) );
  IV U309 ( .A(n4553), .Z(n146) );
  MUX U310 ( .IN0(n4453), .IN1(n147), .SEL(n4454), .F(n4442) );
  IV U311 ( .A(n4455), .Z(n147) );
  MUX U312 ( .IN0(n4133), .IN1(n148), .SEL(n4134), .F(n4116) );
  IV U313 ( .A(n4135), .Z(n148) );
  MUX U314 ( .IN0(n149), .IN1(n1197), .SEL(n1198), .F(n1147) );
  IV U315 ( .A(n1199), .Z(n149) );
  MUX U316 ( .IN0(n1081), .IN1(n150), .SEL(n1082), .F(n1032) );
  IV U317 ( .A(n1083), .Z(n150) );
  MUX U318 ( .IN0(n4398), .IN1(n151), .SEL(n4399), .F(n4387) );
  IV U319 ( .A(n4400), .Z(n151) );
  MUX U320 ( .IN0(n152), .IN1(n4056), .SEL(n4057), .F(n4039) );
  IV U321 ( .A(n4058), .Z(n152) );
  MUX U322 ( .IN0(n4214), .IN1(n153), .SEL(n4215), .F(n4201) );
  IV U323 ( .A(n4216), .Z(n153) );
  MUX U324 ( .IN0(n154), .IN1(n4581), .SEL(n4508), .F(n4579) );
  IV U325 ( .A(n4509), .Z(n154) );
  MUX U326 ( .IN0(n3866), .IN1(n155), .SEL(n3867), .F(n3800) );
  IV U327 ( .A(n3868), .Z(n155) );
  MUX U328 ( .IN0(n156), .IN1(n3817), .SEL(n3818), .F(n3751) );
  IV U329 ( .A(n3819), .Z(n156) );
  MUX U330 ( .IN0(n3757), .IN1(n157), .SEL(n3758), .F(n3691) );
  IV U331 ( .A(n3759), .Z(n157) );
  MUX U332 ( .IN0(n3783), .IN1(n158), .SEL(n3784), .F(n3717) );
  IV U333 ( .A(n3785), .Z(n158) );
  MUX U334 ( .IN0(n159), .IN1(n3447), .SEL(n3448), .F(n3388) );
  IV U335 ( .A(n3449), .Z(n159) );
  MUX U336 ( .IN0(n3264), .IN1(n160), .SEL(n3265), .F(n3221) );
  IV U337 ( .A(n3266), .Z(n160) );
  MUX U338 ( .IN0(n161), .IN1(n3157), .SEL(n3158), .F(n3127) );
  IV U339 ( .A(n3159), .Z(n161) );
  MUX U340 ( .IN0(n3109), .IN1(n162), .SEL(n3110), .F(n3082) );
  IV U341 ( .A(n3111), .Z(n162) );
  XNOR U342 ( .A(n4619), .B(n4620), .Z(n4625) );
  MUX U343 ( .IN0(n1428), .IN1(n163), .SEL(n1429), .F(n1361) );
  IV U344 ( .A(n1430), .Z(n163) );
  MUX U345 ( .IN0(n4566), .IN1(n164), .SEL(n4366), .F(n4557) );
  IV U346 ( .A(n4365), .Z(n164) );
  MUX U347 ( .IN0(n4154), .IN1(n165), .SEL(n4155), .F(n4137) );
  IV U348 ( .A(n4156), .Z(n165) );
  MUX U349 ( .IN0(n1308), .IN1(n166), .SEL(n1309), .F(n1245) );
  IV U350 ( .A(n1310), .Z(n166) );
  MUX U351 ( .IN0(n1323), .IN1(n167), .SEL(n1324), .F(n1261) );
  IV U352 ( .A(n1325), .Z(n167) );
  MUX U353 ( .IN0(n4283), .IN1(n168), .SEL(n4163), .F(n4270) );
  IV U354 ( .A(n4162), .Z(n168) );
  MUX U355 ( .IN0(n1183), .IN1(n169), .SEL(n1184), .F(n1131) );
  IV U356 ( .A(n1185), .Z(n169) );
  MUX U357 ( .IN0(n4435), .IN1(n170), .SEL(n4346), .F(n4424) );
  IV U358 ( .A(n4345), .Z(n170) );
  MUX U359 ( .IN0(n4086), .IN1(n171), .SEL(n4087), .F(n4069) );
  IV U360 ( .A(n4088), .Z(n171) );
  MUX U361 ( .IN0(n1094), .IN1(n172), .SEL(n1095), .F(n1045) );
  IV U362 ( .A(n1096), .Z(n172) );
  MUX U363 ( .IN0(n4519), .IN1(n173), .SEL(n4336), .F(n4510) );
  IV U364 ( .A(n4335), .Z(n173) );
  MUX U365 ( .IN0(n4231), .IN1(n174), .SEL(n4095), .F(n4218) );
  IV U366 ( .A(n4094), .Z(n174) );
  MUX U367 ( .IN0(n1202), .IN1(n175), .SEL(n1203), .F(n1152) );
  IV U368 ( .A(n1204), .Z(n175) );
  MUX U369 ( .IN0(n999), .IN1(n176), .SEL(n1000), .F(n964) );
  IV U370 ( .A(n1001), .Z(n176) );
  MUX U371 ( .IN0(n4378), .IN1(n177), .SEL(n4316), .F(n3936) );
  IV U372 ( .A(n4315), .Z(n177) );
  MUX U373 ( .IN0(n942), .IN1(n178), .SEL(n943), .F(n912) );
  IV U374 ( .A(n944), .Z(n178) );
  MUX U375 ( .IN0(n3945), .IN1(n179), .SEL(n3946), .F(n3879) );
  IV U376 ( .A(n3947), .Z(n179) );
  MUX U377 ( .IN0(n3893), .IN1(n180), .SEL(n3894), .F(n3827) );
  IV U378 ( .A(n3895), .Z(n180) );
  MUX U379 ( .IN0(n3919), .IN1(n181), .SEL(n3920), .F(n3853) );
  IV U380 ( .A(n3921), .Z(n181) );
  MUX U381 ( .IN0(n3738), .IN1(n182), .SEL(n3739), .F(n3672) );
  IV U382 ( .A(n3740), .Z(n182) );
  MUX U383 ( .IN0(n3681), .IN1(n183), .SEL(n3682), .F(n3616) );
  IV U384 ( .A(n3683), .Z(n183) );
  MUX U385 ( .IN0(n3655), .IN1(n184), .SEL(n3656), .F(n3590) );
  IV U386 ( .A(n3657), .Z(n184) );
  MUX U387 ( .IN0(n3566), .IN1(n185), .SEL(n3567), .F(n3502) );
  IV U388 ( .A(n3568), .Z(n185) );
  MUX U389 ( .IN0(n3479), .IN1(n186), .SEL(n3480), .F(n3420) );
  IV U390 ( .A(n3481), .Z(n186) );
  MUX U391 ( .IN0(n3429), .IN1(n187), .SEL(n3430), .F(n3367) );
  IV U392 ( .A(n3431), .Z(n187) );
  MUX U393 ( .IN0(n3259), .IN1(n188), .SEL(n3260), .F(n3216) );
  IV U394 ( .A(n3261), .Z(n188) );
  MUX U395 ( .IN0(n3178), .IN1(n189), .SEL(n3179), .F(n3145) );
  IV U396 ( .A(n3180), .Z(n189) );
  MUX U397 ( .IN0(n1352), .IN1(n190), .SEL(n1353), .F(n1290) );
  IV U398 ( .A(n1354), .Z(n190) );
  MUX U399 ( .IN0(n4337), .IN1(n191), .SEL(n3992), .F(n4331) );
  IV U400 ( .A(n3991), .Z(n191) );
  MUX U401 ( .IN0(n3795), .IN1(n192), .SEL(n3796), .F(n3729) );
  IV U402 ( .A(n3797), .Z(n192) );
  MUX U403 ( .IN0(n3534), .IN1(n193), .SEL(n3535), .F(n3470) );
  IV U404 ( .A(n3536), .Z(n193) );
  XNOR U405 ( .A(n3377), .B(n3327), .Z(n3332) );
  MUX U406 ( .IN0(n3299), .IN1(n194), .SEL(n3300), .F(n3250) );
  IV U407 ( .A(n3301), .Z(n194) );
  MUX U408 ( .IN0(n3103), .IN1(n3133), .SEL(n3105), .F(n3070) );
  MUX U409 ( .IN0(n3037), .IN1(n195), .SEL(n3038), .F(n3021) );
  IV U410 ( .A(n3039), .Z(n195) );
  MUX U411 ( .IN0(n1164), .IN1(n196), .SEL(n1165), .F(n1112) );
  IV U412 ( .A(n1166), .Z(n196) );
  MUX U413 ( .IN0(n3978), .IN1(n197), .SEL(n2991), .F(n3972) );
  IV U414 ( .A(n2990), .Z(n197) );
  XOR U415 ( .A(n844), .B(n843), .Z(n840) );
  MUX U416 ( .IN0(n3637), .IN1(n198), .SEL(n3638), .F(n3573) );
  IV U417 ( .A(n3639), .Z(n198) );
  XNOR U418 ( .A(n3341), .B(n3401), .Z(n3394) );
  MUX U419 ( .IN0(n199), .IN1(n3198), .SEL(n3199), .F(n3152) );
  IV U420 ( .A(n3200), .Z(n199) );
  ANDN U421 ( .A(n981), .B(n982), .Z(n922) );
  ANDN U422 ( .A(n3028), .B(\_MAC/_MULT/MULT/S[3][1][29] ), .Z(n3014) );
  MUX U423 ( .IN0(n200), .IN1(n2487), .SEL(n2488), .F(n2476) );
  IV U424 ( .A(n2489), .Z(n200) );
  XNOR U425 ( .A(n2017), .B(n1981), .Z(n1985) );
  MUX U426 ( .IN0(n2321), .IN1(n201), .SEL(n2322), .F(n2302) );
  IV U427 ( .A(n2323), .Z(n201) );
  XNOR U428 ( .A(n2303), .B(n2287), .Z(n2293) );
  XNOR U429 ( .A(n2479), .B(n2471), .Z(n2301) );
  MUX U430 ( .IN0(n202), .IN1(n2277), .SEL(n2278), .F(n2260) );
  IV U431 ( .A(n2279), .Z(n202) );
  MUX U432 ( .IN0(n2006), .IN1(n203), .SEL(n2007), .F(n1965) );
  IV U433 ( .A(n2008), .Z(n203) );
  MUX U434 ( .IN0(n1961), .IN1(n204), .SEL(n1962), .F(n1922) );
  IV U435 ( .A(n1963), .Z(n204) );
  XNOR U436 ( .A(n1898), .B(n1860), .Z(n1866) );
  XNOR U437 ( .A(n2446), .B(n2438), .Z(n2248) );
  MUX U438 ( .IN0(n2239), .IN1(n205), .SEL(n2240), .F(n2222) );
  IV U439 ( .A(n2241), .Z(n205) );
  XNOR U440 ( .A(n1881), .B(n1843), .Z(n1847) );
  MUX U441 ( .IN0(n206), .IN1(n2209), .SEL(n2210), .F(n2192) );
  IV U442 ( .A(n2211), .Z(n206) );
  MUX U443 ( .IN0(n207), .IN1(n1751), .SEL(n1752), .F(n1712) );
  IV U444 ( .A(n1753), .Z(n207) );
  MUX U445 ( .IN0(n208), .IN1(n1756), .SEL(n1757), .F(n1717) );
  IV U446 ( .A(n1758), .Z(n208) );
  XNOR U447 ( .A(n1779), .B(n1743), .Z(n1747) );
  MUX U448 ( .IN0(n4763), .IN1(n209), .SEL(n4764), .F(n4740) );
  IV U449 ( .A(n4765), .Z(n209) );
  XNOR U450 ( .A(n2413), .B(n2405), .Z(n2197) );
  MUX U451 ( .IN0(n4875), .IN1(n210), .SEL(n4876), .F(n4862) );
  IV U452 ( .A(n4877), .Z(n210) );
  XNOR U453 ( .A(n1762), .B(n1726), .Z(n1730) );
  MUX U454 ( .IN0(n2171), .IN1(n211), .SEL(n2172), .F(n2154) );
  IV U455 ( .A(n2173), .Z(n211) );
  MUX U456 ( .IN0(n2773), .IN1(n2650), .SEL(n2652), .F(n2762) );
  MUX U457 ( .IN0(n212), .IN1(n2669), .SEL(n2514), .F(n2646) );
  IV U458 ( .A(n2513), .Z(n212) );
  MUX U459 ( .IN0(n2753), .IN1(n213), .SEL(n2754), .F(n2742) );
  IV U460 ( .A(n2755), .Z(n213) );
  MUX U461 ( .IN0(n214), .IN1(n2141), .SEL(n2142), .F(n2124) );
  IV U462 ( .A(n2143), .Z(n214) );
  XNOR U463 ( .A(n1662), .B(n1626), .Z(n1630) );
  MUX U464 ( .IN0(n2747), .IN1(n215), .SEL(n2748), .F(n2736) );
  IV U465 ( .A(n2749), .Z(n215) );
  MUX U466 ( .IN0(n2622), .IN1(n2624), .SEL(n2623), .F(n2601) );
  XNOR U467 ( .A(n2380), .B(n2372), .Z(n2146) );
  MUX U468 ( .IN0(n216), .IN1(n1600), .SEL(n1601), .F(n1561) );
  IV U469 ( .A(n1602), .Z(n216) );
  XNOR U470 ( .A(n2572), .B(n2573), .Z(n2582) );
  MUX U471 ( .IN0(n4860), .IN1(n4709), .SEL(n4711), .F(n4847) );
  MUX U472 ( .IN0(n4702), .IN1(n4704), .SEL(n4703), .F(n4681) );
  MUX U473 ( .IN0(n1547), .IN1(n217), .SEL(n1548), .F(n1508) );
  IV U474 ( .A(n1549), .Z(n217) );
  XNOR U475 ( .A(n2551), .B(n2552), .Z(n2561) );
  MUX U476 ( .IN0(n5068), .IN1(n218), .SEL(n5069), .F(n5064) );
  IV U477 ( .A(n5070), .Z(n218) );
  XNOR U478 ( .A(n4652), .B(n4653), .Z(n4662) );
  XNOR U479 ( .A(n2114), .B(n2100), .Z(n2104) );
  XNOR U480 ( .A(n1606), .B(n1570), .Z(n1574) );
  XNOR U481 ( .A(n2723), .B(n2715), .Z(n2547) );
  XNOR U482 ( .A(n2530), .B(n2531), .Z(n2540) );
  MUX U483 ( .IN0(n2534), .IN1(n219), .SEL(n2535), .F(n2502) );
  IV U484 ( .A(n2536), .Z(n219) );
  XNOR U485 ( .A(n4631), .B(n4632), .Z(n4641) );
  MUX U486 ( .IN0(n4635), .IN1(n220), .SEL(n4636), .F(n4603) );
  IV U487 ( .A(n4637), .Z(n220) );
  XNOR U488 ( .A(n4813), .B(n4805), .Z(n4627) );
  XNOR U489 ( .A(n4612), .B(n4613), .Z(n4609) );
  MUX U490 ( .IN0(n1473), .IN1(n221), .SEL(n1474), .F(n1437) );
  IV U491 ( .A(n1475), .Z(n221) );
  MUX U492 ( .IN0(n1366), .IN1(n222), .SEL(n1367), .F(n1304) );
  IV U493 ( .A(n1368), .Z(n222) );
  MUX U494 ( .IN0(n1319), .IN1(n223), .SEL(n1320), .F(n1257) );
  IV U495 ( .A(n1321), .Z(n223) );
  MUX U496 ( .IN0(n4540), .IN1(n224), .SEL(n4541), .F(n4531) );
  IV U497 ( .A(n4542), .Z(n224) );
  MUX U498 ( .IN0(n4442), .IN1(n225), .SEL(n4443), .F(n4431) );
  IV U499 ( .A(n4444), .Z(n225) );
  MUX U500 ( .IN0(n4116), .IN1(n226), .SEL(n4117), .F(n4099) );
  IV U501 ( .A(n4118), .Z(n226) );
  MUX U502 ( .IN0(n227), .IN1(n4107), .SEL(n4108), .F(n4090) );
  IV U503 ( .A(n4109), .Z(n227) );
  MUX U504 ( .IN0(n228), .IN1(n4585), .SEL(n4526), .F(n4583) );
  IV U505 ( .A(n4527), .Z(n228) );
  MUX U506 ( .IN0(n4048), .IN1(n229), .SEL(n4049), .F(n4031) );
  IV U507 ( .A(n4050), .Z(n229) );
  MUX U508 ( .IN0(n230), .IN1(n3949), .SEL(n3950), .F(n3883) );
  IV U509 ( .A(n3951), .Z(n230) );
  MUX U510 ( .IN0(n3941), .IN1(n231), .SEL(n3942), .F(n3875) );
  IV U511 ( .A(n3943), .Z(n231) );
  MUX U512 ( .IN0(n3734), .IN1(n232), .SEL(n3735), .F(n3668) );
  IV U513 ( .A(n3736), .Z(n232) );
  MUX U514 ( .IN0(n3691), .IN1(n233), .SEL(n3692), .F(n3626) );
  IV U515 ( .A(n3693), .Z(n233) );
  MUX U516 ( .IN0(n234), .IN1(n3685), .SEL(n3686), .F(n3620) );
  IV U517 ( .A(n3687), .Z(n234) );
  MUX U518 ( .IN0(n3677), .IN1(n235), .SEL(n3678), .F(n3612) );
  IV U519 ( .A(n3679), .Z(n235) );
  MUX U520 ( .IN0(n3475), .IN1(n236), .SEL(n3476), .F(n3416) );
  IV U521 ( .A(n3477), .Z(n236) );
  MUX U522 ( .IN0(n237), .IN1(n3433), .SEL(n3434), .F(n3371) );
  IV U523 ( .A(n3435), .Z(n237) );
  MUX U524 ( .IN0(n3425), .IN1(n238), .SEL(n3426), .F(n3363) );
  IV U525 ( .A(n3427), .Z(n238) );
  MUX U526 ( .IN0(n3255), .IN1(n239), .SEL(n3256), .F(n3212) );
  IV U527 ( .A(n3257), .Z(n239) );
  MUX U528 ( .IN0(n3174), .IN1(n240), .SEL(n3175), .F(n3141) );
  IV U529 ( .A(n3176), .Z(n240) );
  XNOR U530 ( .A(n5088), .B(n5089), .Z(n4575) );
  MUX U531 ( .IN0(n1452), .IN1(n241), .SEL(n1453), .F(n1385) );
  IV U532 ( .A(n1454), .Z(n241) );
  MUX U533 ( .IN0(n2330), .IN1(n242), .SEL(n2078), .F(n1409) );
  IV U534 ( .A(n2077), .Z(n242) );
  XNOR U535 ( .A(n1489), .B(n1425), .Z(n1429) );
  MUX U536 ( .IN0(n4481), .IN1(n243), .SEL(n4482), .F(n4470) );
  IV U537 ( .A(n4483), .Z(n243) );
  MUX U538 ( .IN0(n4137), .IN1(n244), .SEL(n4138), .F(n4120) );
  IV U539 ( .A(n4139), .Z(n244) );
  MUX U540 ( .IN0(n1192), .IN1(n245), .SEL(n1193), .F(n1140) );
  IV U541 ( .A(n1194), .Z(n245) );
  MUX U542 ( .IN0(n1131), .IN1(n246), .SEL(n1132), .F(n1085) );
  IV U543 ( .A(n1133), .Z(n246) );
  MUX U544 ( .IN0(n4424), .IN1(n247), .SEL(n4340), .F(n4413) );
  IV U545 ( .A(n4339), .Z(n247) );
  MUX U546 ( .IN0(n4069), .IN1(n248), .SEL(n4070), .F(n4052) );
  IV U547 ( .A(n4071), .Z(n248) );
  MUX U548 ( .IN0(n994), .IN1(n249), .SEL(n995), .F(n962) );
  IV U549 ( .A(n996), .Z(n249) );
  MUX U550 ( .IN0(n912), .IN1(n250), .SEL(n913), .F(n881) );
  IV U551 ( .A(n914), .Z(n250) );
  MUX U552 ( .IN0(n3827), .IN1(n251), .SEL(n3828), .F(n3761) );
  IV U553 ( .A(n3829), .Z(n251) );
  MUX U554 ( .IN0(n3853), .IN1(n252), .SEL(n3854), .F(n3787) );
  IV U555 ( .A(n3855), .Z(n252) );
  MUX U556 ( .IN0(n3813), .IN1(n253), .SEL(n3814), .F(n3747) );
  IV U557 ( .A(n3815), .Z(n253) );
  MUX U558 ( .IN0(n3607), .IN1(n254), .SEL(n3608), .F(n3543) );
  IV U559 ( .A(n3609), .Z(n254) );
  MUX U560 ( .IN0(n3590), .IN1(n255), .SEL(n3591), .F(n3526) );
  IV U561 ( .A(n3592), .Z(n255) );
  MUX U562 ( .IN0(n3552), .IN1(n256), .SEL(n3553), .F(n3488) );
  IV U563 ( .A(n3554), .Z(n256) );
  MUX U564 ( .IN0(n3443), .IN1(n257), .SEL(n3444), .F(n3384) );
  IV U565 ( .A(n3445), .Z(n257) );
  MUX U566 ( .IN0(n3358), .IN1(n258), .SEL(n3359), .F(n3308) );
  IV U567 ( .A(n3360), .Z(n258) );
  MUX U568 ( .IN0(n3317), .IN1(n259), .SEL(n3318), .F(n3268) );
  IV U569 ( .A(n3319), .Z(n259) );
  MUX U570 ( .IN0(n3169), .IN1(n260), .SEL(n3170), .F(n3136) );
  IV U571 ( .A(n3171), .Z(n260) );
  MUX U572 ( .IN0(n4181), .IN1(n261), .SEL(n4182), .F(n4164) );
  IV U573 ( .A(n4183), .Z(n261) );
  MUX U574 ( .IN0(n4361), .IN1(n262), .SEL(n4016), .F(n4355) );
  IV U575 ( .A(n4015), .Z(n262) );
  XNOR U576 ( .A(n4288), .B(n4280), .Z(n4163) );
  MUX U577 ( .IN0(n1338), .IN1(n263), .SEL(n1339), .F(n1280) );
  IV U578 ( .A(n1340), .Z(n263) );
  MUX U579 ( .IN0(n1227), .IN1(n264), .SEL(n1228), .F(n1174) );
  IV U580 ( .A(n1229), .Z(n264) );
  MUX U581 ( .IN0(n4113), .IN1(n265), .SEL(n4001), .F(n4096) );
  IV U582 ( .A(n4000), .Z(n265) );
  XNOR U583 ( .A(n4520), .B(n4514), .Z(n4336) );
  MUX U584 ( .IN0(n1154), .IN1(n266), .SEL(n1155), .F(n1103) );
  IV U585 ( .A(n1156), .Z(n266) );
  XNOR U586 ( .A(n1039), .B(n1005), .Z(n1009) );
  MUX U587 ( .IN0(n1026), .IN1(n267), .SEL(n1027), .F(n990) );
  IV U588 ( .A(n1028), .Z(n267) );
  MUX U589 ( .IN0(n4325), .IN1(n268), .SEL(n3980), .F(n4319) );
  IV U590 ( .A(n3979), .Z(n268) );
  XNOR U591 ( .A(n4210), .B(n4202), .Z(n4061) );
  XNOR U592 ( .A(n4383), .B(n4375), .Z(n4316) );
  MUX U593 ( .IN0(n3710), .IN1(n269), .SEL(n3711), .F(n3645) );
  IV U594 ( .A(n3712), .Z(n269) );
  MUX U595 ( .IN0(n3663), .IN1(n270), .SEL(n3664), .F(n3598) );
  IV U596 ( .A(n3665), .Z(n270) );
  MUX U597 ( .IN0(n3411), .IN1(n271), .SEL(n3412), .F(n3349) );
  IV U598 ( .A(n3413), .Z(n271) );
  MUX U599 ( .IN0(n3130), .IN1(n272), .SEL(n3131), .F(n3100) );
  IV U600 ( .A(n3132), .Z(n272) );
  XNOR U601 ( .A(n3107), .B(n3083), .Z(n3087) );
  MUX U602 ( .IN0(n1394), .IN1(n273), .SEL(n1395), .F(n1330) );
  IV U603 ( .A(n1396), .Z(n273) );
  MUX U604 ( .IN0(n4002), .IN1(n274), .SEL(n2999), .F(n3996) );
  IV U605 ( .A(n2998), .Z(n274) );
  MUX U606 ( .IN0(n1112), .IN1(n275), .SEL(n1113), .F(n1066) );
  IV U607 ( .A(n1114), .Z(n275) );
  MUX U608 ( .IN0(n3900), .IN1(n276), .SEL(n3901), .F(n3834) );
  IV U609 ( .A(n3902), .Z(n276) );
  XNOR U610 ( .A(n827), .B(n828), .Z(n833) );
  MUX U611 ( .IN0(n3511), .IN1(n277), .SEL(n3512), .F(n3450) );
  IV U612 ( .A(n3513), .Z(n277) );
  MUX U613 ( .IN0(n3291), .IN1(n278), .SEL(n3292), .F(n3242) );
  IV U614 ( .A(n3293), .Z(n278) );
  MUX U615 ( .IN0(n3233), .IN1(n279), .SEL(n3234), .F(n3187) );
  IV U616 ( .A(n3235), .Z(n279) );
  MUX U617 ( .IN0(n3021), .IN1(n280), .SEL(n3022), .F(n3011) );
  IV U618 ( .A(n3023), .Z(n280) );
  MUX U619 ( .IN0(n1069), .IN1(\_MAC/_MULT/MULT/S[3][1][6] ), .SEL(n5118), .F(
        n1019) );
  XOR U620 ( .A(n931), .B(n930), .Z(n923) );
  XOR U621 ( .A(n854), .B(n855), .Z(n853) );
  XOR U622 ( .A(n3208), .B(n3207), .Z(n3200) );
  XOR U623 ( .A(n3032), .B(n3033), .Z(n3046) );
  MUX U624 ( .IN0(n2305), .IN1(n281), .SEL(n2306), .F(n2286) );
  IV U625 ( .A(n2307), .Z(n281) );
  MUX U626 ( .IN0(n2492), .IN1(n282), .SEL(n2493), .F(n2481) );
  IV U627 ( .A(n2494), .Z(n282) );
  MUX U628 ( .IN0(n283), .IN1(n2296), .SEL(n2297), .F(n2277) );
  IV U629 ( .A(n2298), .Z(n283) );
  MUX U630 ( .IN0(n2040), .IN1(n284), .SEL(n2041), .F(n1997) );
  IV U631 ( .A(n2042), .Z(n284) );
  MUX U632 ( .IN0(n285), .IN1(n2465), .SEL(n2466), .F(n2454) );
  IV U633 ( .A(n2467), .Z(n285) );
  MUX U634 ( .IN0(n286), .IN1(n1909), .SEL(n1910), .F(n1870) );
  IV U635 ( .A(n1911), .Z(n286) );
  MUX U636 ( .IN0(n2302), .IN1(n287), .SEL(n2015), .F(n2283) );
  IV U637 ( .A(n2013), .Z(n287) );
  XNOR U638 ( .A(n2000), .B(n1962), .Z(n1966) );
  XNOR U639 ( .A(n2468), .B(n2460), .Z(n2282) );
  MUX U640 ( .IN0(n288), .IN1(n1914), .SEL(n1915), .F(n1875) );
  IV U641 ( .A(n1916), .Z(n288) );
  XNOR U642 ( .A(n1937), .B(n1901), .Z(n1905) );
  MUX U643 ( .IN0(n2256), .IN1(n289), .SEL(n2257), .F(n2239) );
  IV U644 ( .A(n2258), .Z(n289) );
  MUX U645 ( .IN0(n290), .IN1(n2226), .SEL(n2227), .F(n2209) );
  IV U646 ( .A(n2228), .Z(n290) );
  MUX U647 ( .IN0(n2218), .IN1(n291), .SEL(n2219), .F(n2201) );
  IV U648 ( .A(n2220), .Z(n291) );
  MUX U649 ( .IN0(n1878), .IN1(n292), .SEL(n1879), .F(n1837) );
  IV U650 ( .A(n1880), .Z(n292) );
  MUX U651 ( .IN0(n293), .IN1(n2421), .SEL(n2422), .F(n2410) );
  IV U652 ( .A(n2423), .Z(n293) );
  MUX U653 ( .IN0(n1785), .IN1(n294), .SEL(n1786), .F(n1746) );
  IV U654 ( .A(n1787), .Z(n294) );
  MUX U655 ( .IN0(n2232), .IN1(n295), .SEL(n1855), .F(n2215) );
  IV U656 ( .A(n1853), .Z(n295) );
  XNOR U657 ( .A(n2424), .B(n2416), .Z(n2214) );
  MUX U658 ( .IN0(n2780), .IN1(n296), .SEL(n2781), .F(n2769) );
  IV U659 ( .A(n2782), .Z(n296) );
  MUX U660 ( .IN0(n4895), .IN1(n297), .SEL(n4896), .F(n4882) );
  IV U661 ( .A(n4897), .Z(n297) );
  MUX U662 ( .IN0(n4888), .IN1(n298), .SEL(n4889), .F(n4875) );
  IV U663 ( .A(n4890), .Z(n298) );
  MUX U664 ( .IN0(n299), .IN1(n1712), .SEL(n1713), .F(n1673) );
  IV U665 ( .A(n1714), .Z(n299) );
  MUX U666 ( .IN0(n1703), .IN1(n300), .SEL(n1704), .F(n1664) );
  IV U667 ( .A(n1705), .Z(n300) );
  MUX U668 ( .IN0(n2188), .IN1(n301), .SEL(n2189), .F(n2171) );
  IV U669 ( .A(n2190), .Z(n301) );
  MUX U670 ( .IN0(n1768), .IN1(n302), .SEL(n1769), .F(n1729) );
  IV U671 ( .A(n1770), .Z(n302) );
  MUX U672 ( .IN0(n1725), .IN1(n303), .SEL(n1726), .F(n1686) );
  IV U673 ( .A(n1727), .Z(n303) );
  MUX U674 ( .IN0(n304), .IN1(n2158), .SEL(n2159), .F(n2141) );
  IV U675 ( .A(n2160), .Z(n304) );
  MUX U676 ( .IN0(n2150), .IN1(n305), .SEL(n2151), .F(n2133) );
  IV U677 ( .A(n2152), .Z(n305) );
  MUX U678 ( .IN0(n306), .IN1(n1678), .SEL(n1679), .F(n1639) );
  IV U679 ( .A(n1680), .Z(n306) );
  XNOR U680 ( .A(n2660), .B(n2640), .Z(n2644) );
  XNOR U681 ( .A(n2614), .B(n2615), .Z(n2624) );
  MUX U682 ( .IN0(n307), .IN1(n4770), .SEL(n4615), .F(n4747) );
  IV U683 ( .A(n4614), .Z(n307) );
  MUX U684 ( .IN0(n1720), .IN1(n308), .SEL(n1721), .F(n1681) );
  IV U685 ( .A(n1722), .Z(n308) );
  XNOR U686 ( .A(n2756), .B(n2748), .Z(n2610) );
  XNOR U687 ( .A(n2593), .B(n2594), .Z(n2603) );
  MUX U688 ( .IN0(n2597), .IN1(n309), .SEL(n2598), .F(n2576) );
  IV U689 ( .A(n2599), .Z(n309) );
  MUX U690 ( .IN0(n2837), .IN1(n310), .SEL(n2838), .F(n2821) );
  IV U691 ( .A(n2839), .Z(n310) );
  MUX U692 ( .IN0(n4873), .IN1(n4730), .SEL(n4732), .F(n4860) );
  XNOR U693 ( .A(n4738), .B(n4720), .Z(n4724) );
  XNOR U694 ( .A(n4694), .B(n4695), .Z(n4704) );
  MUX U695 ( .IN0(n4950), .IN1(n311), .SEL(n4951), .F(n4934) );
  IV U696 ( .A(n4952), .Z(n311) );
  MUX U697 ( .IN0(n1629), .IN1(n312), .SEL(n1630), .F(n1590) );
  IV U698 ( .A(n1631), .Z(n312) );
  MUX U699 ( .IN0(n2382), .IN1(n313), .SEL(n2383), .F(n2371) );
  IV U700 ( .A(n2384), .Z(n313) );
  MUX U701 ( .IN0(n2164), .IN1(n314), .SEL(n1699), .F(n2147) );
  IV U702 ( .A(n1697), .Z(n314) );
  MUX U703 ( .IN0(n2927), .IN1(n315), .SEL(n2928), .F(n2911) );
  IV U704 ( .A(n2929), .Z(n315) );
  MUX U705 ( .IN0(n2731), .IN1(n316), .SEL(n2732), .F(n2720) );
  IV U706 ( .A(n2733), .Z(n316) );
  MUX U707 ( .IN0(n4843), .IN1(n317), .SEL(n4844), .F(n4830) );
  IV U708 ( .A(n4845), .Z(n317) );
  MUX U709 ( .IN0(n4836), .IN1(n318), .SEL(n4837), .F(n4823) );
  IV U710 ( .A(n4838), .Z(n318) );
  XNOR U711 ( .A(n4673), .B(n4674), .Z(n4683) );
  MUX U712 ( .IN0(n319), .IN1(n1556), .SEL(n1557), .F(n1517) );
  IV U713 ( .A(n1558), .Z(n319) );
  MUX U714 ( .IN0(n2375), .IN1(n320), .SEL(n2146), .F(n2364) );
  IV U715 ( .A(n2145), .Z(n320) );
  MUX U716 ( .IN0(n2120), .IN1(n321), .SEL(n2121), .F(n2103) );
  IV U717 ( .A(n2122), .Z(n321) );
  MUX U718 ( .IN0(n1612), .IN1(n322), .SEL(n1613), .F(n1573) );
  IV U719 ( .A(n1614), .Z(n322) );
  MUX U720 ( .IN0(n2679), .IN1(n323), .SEL(n2680), .F(n2675) );
  IV U721 ( .A(n2681), .Z(n323) );
  MUX U722 ( .IN0(n5028), .IN1(n5043), .SEL(n5030), .F(n5010) );
  MUX U723 ( .IN0(n4656), .IN1(n324), .SEL(n4657), .F(n4635) );
  IV U724 ( .A(n4658), .Z(n324) );
  MUX U725 ( .IN0(n1508), .IN1(n325), .SEL(n1509), .F(n1469) );
  IV U726 ( .A(n1510), .Z(n325) );
  MUX U727 ( .IN0(n326), .IN1(n2090), .SEL(n2091), .F(n2073) );
  IV U728 ( .A(n2092), .Z(n326) );
  MUX U729 ( .IN0(n2082), .IN1(n327), .SEL(n2083), .F(n2065) );
  IV U730 ( .A(n2084), .Z(n327) );
  MUX U731 ( .IN0(n328), .IN1(n1522), .SEL(n1523), .F(n1483) );
  IV U732 ( .A(n1524), .Z(n328) );
  MUX U733 ( .IN0(n1491), .IN1(n329), .SEL(n1492), .F(n1424) );
  IV U734 ( .A(n1493), .Z(n329) );
  MUX U735 ( .IN0(n1564), .IN1(n330), .SEL(n1565), .F(n1525) );
  IV U736 ( .A(n1566), .Z(n330) );
  MUX U737 ( .IN0(n2718), .IN1(n2545), .SEL(n2547), .F(n2707) );
  XNOR U738 ( .A(n2553), .B(n2535), .Z(n2539) );
  XNOR U739 ( .A(n2511), .B(n2512), .Z(n2508) );
  MUX U740 ( .IN0(n2096), .IN1(n331), .SEL(n1543), .F(n2079) );
  IV U741 ( .A(n1541), .Z(n331) );
  MUX U742 ( .IN0(n4569), .IN1(n332), .SEL(n4570), .F(n4560) );
  IV U743 ( .A(n4571), .Z(n332) );
  MUX U744 ( .IN0(n333), .IN1(n4175), .SEL(n4176), .F(n4158) );
  IV U745 ( .A(n4177), .Z(n333) );
  MUX U746 ( .IN0(n334), .IN1(n4296), .SEL(n4297), .F(n4285) );
  IV U747 ( .A(n4298), .Z(n334) );
  MUX U748 ( .IN0(n4301), .IN1(n335), .SEL(n4302), .F(n4290) );
  IV U749 ( .A(n4303), .Z(n335) );
  MUX U750 ( .IN0(n1304), .IN1(n336), .SEL(n1305), .F(n1241) );
  IV U751 ( .A(n1306), .Z(n336) );
  MUX U752 ( .IN0(n337), .IN1(n1327), .SEL(n1328), .F(n1265) );
  IV U753 ( .A(n1329), .Z(n337) );
  MUX U754 ( .IN0(n4531), .IN1(n338), .SEL(n4532), .F(n4522) );
  IV U755 ( .A(n4533), .Z(n338) );
  MUX U756 ( .IN0(n4431), .IN1(n339), .SEL(n4432), .F(n4420) );
  IV U757 ( .A(n4433), .Z(n339) );
  MUX U758 ( .IN0(n4099), .IN1(n340), .SEL(n4100), .F(n4082) );
  IV U759 ( .A(n4101), .Z(n340) );
  MUX U760 ( .IN0(n4253), .IN1(n341), .SEL(n4254), .F(n4240) );
  IV U761 ( .A(n4255), .Z(n341) );
  MUX U762 ( .IN0(n342), .IN1(n1099), .SEL(n1100), .F(n1050) );
  IV U763 ( .A(n1101), .Z(n342) );
  MUX U764 ( .IN0(n1041), .IN1(n343), .SEL(n1042), .F(n1004) );
  IV U765 ( .A(n1043), .Z(n343) );
  MUX U766 ( .IN0(n4493), .IN1(n344), .SEL(n4494), .F(n4486) );
  IV U767 ( .A(n4495), .Z(n344) );
  MUX U768 ( .IN0(n4031), .IN1(n345), .SEL(n4032), .F(n3955) );
  IV U769 ( .A(n4033), .Z(n345) );
  MUX U770 ( .IN0(n3849), .IN1(n346), .SEL(n3850), .F(n3783) );
  IV U771 ( .A(n3851), .Z(n346) );
  MUX U772 ( .IN0(n3809), .IN1(n347), .SEL(n3810), .F(n3743) );
  IV U773 ( .A(n3811), .Z(n347) );
  MUX U774 ( .IN0(n3800), .IN1(n348), .SEL(n3801), .F(n3734) );
  IV U775 ( .A(n3802), .Z(n348) );
  MUX U776 ( .IN0(n349), .IN1(n3699), .SEL(n3700), .F(n3634) );
  IV U777 ( .A(n3701), .Z(n349) );
  MUX U778 ( .IN0(n350), .IN1(n3620), .SEL(n3621), .F(n3556) );
  IV U779 ( .A(n3622), .Z(n350) );
  MUX U780 ( .IN0(n351), .IN1(n3595), .SEL(n3596), .F(n3531) );
  IV U781 ( .A(n3597), .Z(n351) );
  MUX U782 ( .IN0(n3484), .IN1(n352), .SEL(n3485), .F(n3425) );
  IV U783 ( .A(n3486), .Z(n352) );
  MUX U784 ( .IN0(n3354), .IN1(n353), .SEL(n3355), .F(n3304) );
  IV U785 ( .A(n3356), .Z(n353) );
  MUX U786 ( .IN0(n354), .IN1(n3274), .SEL(n3275), .F(n3229) );
  IV U787 ( .A(n3276), .Z(n354) );
  MUX U788 ( .IN0(n355), .IN1(n3388), .SEL(n3389), .F(n3335) );
  IV U789 ( .A(n3390), .Z(n355) );
  MUX U790 ( .IN0(n3221), .IN1(n356), .SEL(n3222), .F(n3174) );
  IV U791 ( .A(n3223), .Z(n356) );
  MUX U792 ( .IN0(n4607), .IN1(n4609), .SEL(n4608), .F(n4171) );
  MUX U793 ( .IN0(n4808), .IN1(n4625), .SEL(n4627), .F(n4305) );
  MUX U794 ( .IN0(n1437), .IN1(n357), .SEL(n1438), .F(n1370) );
  IV U795 ( .A(n1439), .Z(n357) );
  MUX U796 ( .IN0(n1361), .IN1(n358), .SEL(n1362), .F(n1299) );
  IV U797 ( .A(n1363), .Z(n358) );
  MUX U798 ( .IN0(n4557), .IN1(n359), .SEL(n4360), .F(n4546) );
  IV U799 ( .A(n4359), .Z(n359) );
  MUX U800 ( .IN0(n1409), .IN1(n360), .SEL(n1410), .F(n1341) );
  IV U801 ( .A(n1411), .Z(n360) );
  MUX U802 ( .IN0(n4446), .IN1(n361), .SEL(n4352), .F(n4435) );
  IV U803 ( .A(n4351), .Z(n361) );
  MUX U804 ( .IN0(n4120), .IN1(n362), .SEL(n4121), .F(n4103) );
  IV U805 ( .A(n4122), .Z(n362) );
  MUX U806 ( .IN0(n4270), .IN1(n363), .SEL(n4146), .F(n4257) );
  IV U807 ( .A(n4145), .Z(n363) );
  MUX U808 ( .IN0(n4510), .IN1(n364), .SEL(n4330), .F(n4499) );
  IV U809 ( .A(n4329), .Z(n364) );
  MUX U810 ( .IN0(n4402), .IN1(n365), .SEL(n4328), .F(n4391) );
  IV U811 ( .A(n4327), .Z(n365) );
  MUX U812 ( .IN0(n4052), .IN1(n366), .SEL(n4053), .F(n4035) );
  IV U813 ( .A(n4054), .Z(n366) );
  MUX U814 ( .IN0(n4218), .IN1(n367), .SEL(n4078), .F(n4205) );
  IV U815 ( .A(n4077), .Z(n367) );
  MUX U816 ( .IN0(n973), .IN1(n368), .SEL(n974), .F(n942) );
  IV U817 ( .A(n975), .Z(n368) );
  MUX U818 ( .IN0(n964), .IN1(n369), .SEL(n965), .F(n932) );
  IV U819 ( .A(n966), .Z(n369) );
  MUX U820 ( .IN0(n3879), .IN1(n370), .SEL(n3880), .F(n3813) );
  IV U821 ( .A(n3881), .Z(n370) );
  MUX U822 ( .IN0(n3870), .IN1(n371), .SEL(n3871), .F(n3804) );
  IV U823 ( .A(n3872), .Z(n371) );
  MUX U824 ( .IN0(n3721), .IN1(n372), .SEL(n3722), .F(n3655) );
  IV U825 ( .A(n3723), .Z(n372) );
  MUX U826 ( .IN0(n3585), .IN1(n373), .SEL(n3586), .F(n3524) );
  IV U827 ( .A(n3587), .Z(n373) );
  MUX U828 ( .IN0(n3420), .IN1(n374), .SEL(n3421), .F(n3358) );
  IV U829 ( .A(n3422), .Z(n374) );
  MUX U830 ( .IN0(n3367), .IN1(n375), .SEL(n3368), .F(n3317) );
  IV U831 ( .A(n3369), .Z(n375) );
  MUX U832 ( .IN0(n3326), .IN1(n376), .SEL(n3327), .F(n3279) );
  IV U833 ( .A(n3328), .Z(n376) );
  MUX U834 ( .IN0(n3216), .IN1(n377), .SEL(n3217), .F(n3169) );
  IV U835 ( .A(n3218), .Z(n377) );
  MUX U836 ( .IN0(n3145), .IN1(n378), .SEL(n3146), .F(n3113) );
  IV U837 ( .A(n3147), .Z(n378) );
  MUX U838 ( .IN0(n3164), .IN1(n379), .SEL(n3165), .F(n3134) );
  IV U839 ( .A(n3166), .Z(n379) );
  MUX U840 ( .IN0(n3082), .IN1(n380), .SEL(n3083), .F(n3051) );
  IV U841 ( .A(n3084), .Z(n380) );
  XNOR U842 ( .A(n1446), .B(n1382), .Z(n1388) );
  MUX U843 ( .IN0(n4367), .IN1(n381), .SEL(n4368), .F(n4361) );
  IV U844 ( .A(n4369), .Z(n381) );
  MUX U845 ( .IN0(n4164), .IN1(n382), .SEL(n4019), .F(n4147) );
  IV U846 ( .A(n4018), .Z(n382) );
  MUX U847 ( .IN0(n1290), .IN1(n383), .SEL(n1291), .F(n1227) );
  IV U848 ( .A(n1292), .Z(n383) );
  XNOR U849 ( .A(n1186), .B(n1137), .Z(n1143) );
  XNOR U850 ( .A(n1177), .B(n1128), .Z(n1132) );
  MUX U851 ( .IN0(n384), .IN1(n1280), .SEL(n1281), .F(n1217) );
  IV U852 ( .A(n1282), .Z(n384) );
  MUX U853 ( .IN0(n4343), .IN1(n385), .SEL(n3998), .F(n4337) );
  IV U854 ( .A(n3997), .Z(n385) );
  MUX U855 ( .IN0(n4096), .IN1(n386), .SEL(n3995), .F(n4079) );
  IV U856 ( .A(n3994), .Z(n386) );
  MUX U857 ( .IN0(n990), .IN1(n387), .SEL(n991), .F(n958) );
  IV U858 ( .A(n992), .Z(n387) );
  MUX U859 ( .IN0(n4313), .IN1(n388), .SEL(n3968), .F(n3927) );
  IV U860 ( .A(n3967), .Z(n388) );
  MUX U861 ( .IN0(n4028), .IN1(n389), .SEL(n3971), .F(n3908) );
  IV U862 ( .A(n3970), .Z(n389) );
  XNOR U863 ( .A(n3887), .B(n3824), .Z(n3828) );
  XNOR U864 ( .A(n875), .B(n857), .Z(n860) );
  MUX U865 ( .IN0(n3729), .IN1(n390), .SEL(n3730), .F(n3663) );
  IV U866 ( .A(n3731), .Z(n390) );
  XNOR U867 ( .A(n3675), .B(n3613), .Z(n3617) );
  XNOR U868 ( .A(n3666), .B(n3604), .Z(n3608) );
  XNOR U869 ( .A(n3624), .B(n3563), .Z(n3567) );
  MUX U870 ( .IN0(n3645), .IN1(n391), .SEL(n3646), .F(n3581) );
  IV U871 ( .A(n3647), .Z(n391) );
  MUX U872 ( .IN0(n3470), .IN1(n392), .SEL(n3471), .F(n3411) );
  IV U873 ( .A(n3472), .Z(n392) );
  MUX U874 ( .IN0(n393), .IN1(n3403), .SEL(n3404), .F(n3341) );
  IV U875 ( .A(n3405), .Z(n393) );
  MUX U876 ( .IN0(n3250), .IN1(n394), .SEL(n3251), .F(n3206) );
  IV U877 ( .A(n3252), .Z(n394) );
  MUX U878 ( .IN0(n4008), .IN1(n395), .SEL(n3030), .F(n4002) );
  IV U879 ( .A(n3029), .Z(n395) );
  MUX U880 ( .IN0(n396), .IN1(n1214), .SEL(n1215), .F(n1164) );
  IV U881 ( .A(n1216), .Z(n396) );
  MUX U882 ( .IN0(n3984), .IN1(n397), .SEL(n2993), .F(n3978) );
  IV U883 ( .A(n2992), .Z(n397) );
  MUX U884 ( .IN0(n1103), .IN1(n398), .SEL(n1104), .F(n1055) );
  IV U885 ( .A(n1105), .Z(n398) );
  MUX U886 ( .IN0(n399), .IN1(n872), .SEL(n873), .F(n855) );
  IV U887 ( .A(n874), .Z(n399) );
  MUX U888 ( .IN0(n3768), .IN1(n400), .SEL(n3769), .F(n3702) );
  IV U889 ( .A(n3770), .Z(n400) );
  MUX U890 ( .IN0(n401), .IN1(n847), .SEL(n848), .F(n826) );
  IV U891 ( .A(n849), .Z(n401) );
  MUX U892 ( .IN0(n3338), .IN1(n402), .SEL(n3339), .F(n3291) );
  IV U893 ( .A(n3340), .Z(n402) );
  MUX U894 ( .IN0(n3076), .IN1(n403), .SEL(n3077), .F(n3047) );
  IV U895 ( .A(n3078), .Z(n403) );
  MUX U896 ( .IN0(n404), .IN1(n3060), .SEL(n3061), .F(n3042) );
  IV U897 ( .A(n3062), .Z(n404) );
  XOR U898 ( .A(n1078), .B(n1077), .Z(n1114) );
  MUX U899 ( .IN0(n983), .IN1(\_MAC/_MULT/MULT/S[3][1][8] ), .SEL(n5120), .F(
        n950) );
  ANDN U900 ( .A(n870), .B(n871), .Z(n852) );
  MUX U901 ( .IN0(n836), .IN1(\_MAC/_MULT/MULT/S[3][1][14] ), .SEL(n5126), .F(
        n816) );
  MUX U902 ( .IN0(n3152), .IN1(n405), .SEL(n3153), .F(n3123) );
  IV U903 ( .A(n3154), .Z(n405) );
  AND U904 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[27] ), .B(
        \_MAC/_MULT/MULT/S[3][1][27] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[28] ) );
  XOR U905 ( .A(n3015), .B(n3004), .Z(n3018) );
  MUX U906 ( .IN0(n2019), .IN1(n406), .SEL(n2020), .F(n1978) );
  IV U907 ( .A(n2021), .Z(n406) );
  MUX U908 ( .IN0(n407), .IN1(n2315), .SEL(n2316), .F(n2296) );
  IV U909 ( .A(n2317), .Z(n407) );
  MUX U910 ( .IN0(n408), .IN1(n2037), .SEL(n2038), .F(n1994) );
  IV U911 ( .A(n2039), .Z(n408) );
  MUX U912 ( .IN0(n2054), .IN1(n409), .SEL(n2055), .F(n2009) );
  IV U913 ( .A(n2056), .Z(n409) );
  MUX U914 ( .IN0(n2273), .IN1(n410), .SEL(n2274), .F(n2256) );
  IV U915 ( .A(n2275), .Z(n410) );
  MUX U916 ( .IN0(n1965), .IN1(n411), .SEL(n1966), .F(n1926) );
  IV U917 ( .A(n1967), .Z(n411) );
  MUX U918 ( .IN0(n2470), .IN1(n412), .SEL(n2471), .F(n2459) );
  IV U919 ( .A(n2472), .Z(n412) );
  MUX U920 ( .IN0(n413), .IN1(n2454), .SEL(n2455), .F(n2443) );
  IV U921 ( .A(n2456), .Z(n413) );
  MUX U922 ( .IN0(n414), .IN1(n1870), .SEL(n1871), .F(n1829) );
  IV U923 ( .A(n1872), .Z(n414) );
  MUX U924 ( .IN0(n1859), .IN1(n415), .SEL(n1860), .F(n1820) );
  IV U925 ( .A(n1861), .Z(n415) );
  MUX U926 ( .IN0(n2235), .IN1(n416), .SEL(n2236), .F(n2218) );
  IV U927 ( .A(n2237), .Z(n416) );
  MUX U928 ( .IN0(n417), .IN1(n1875), .SEL(n1876), .F(n1834) );
  IV U929 ( .A(n1877), .Z(n417) );
  MUX U930 ( .IN0(n1883), .IN1(n418), .SEL(n1884), .F(n1842) );
  IV U931 ( .A(n1885), .Z(n418) );
  MUX U932 ( .IN0(n1917), .IN1(n419), .SEL(n1918), .F(n1878) );
  IV U933 ( .A(n1919), .Z(n419) );
  MUX U934 ( .IN0(n2441), .IN1(n420), .SEL(n2248), .F(n2430) );
  IV U935 ( .A(n2247), .Z(n420) );
  MUX U936 ( .IN0(n2249), .IN1(n421), .SEL(n1896), .F(n2232) );
  IV U937 ( .A(n1894), .Z(n421) );
  MUX U938 ( .IN0(n2205), .IN1(n422), .SEL(n2206), .F(n2188) );
  IV U939 ( .A(n2207), .Z(n422) );
  MUX U940 ( .IN0(n1807), .IN1(n423), .SEL(n1808), .F(n1768) );
  IV U941 ( .A(n1809), .Z(n423) );
  MUX U942 ( .IN0(n424), .IN1(n2775), .SEL(n2776), .F(n2764) );
  IV U943 ( .A(n2777), .Z(n424) );
  MUX U944 ( .IN0(n2662), .IN1(n425), .SEL(n2663), .F(n2639) );
  IV U945 ( .A(n2664), .Z(n425) );
  MUX U946 ( .IN0(n2426), .IN1(n426), .SEL(n2427), .F(n2415) );
  IV U947 ( .A(n2428), .Z(n426) );
  MUX U948 ( .IN0(n427), .IN1(n2410), .SEL(n2411), .F(n2399) );
  IV U949 ( .A(n2412), .Z(n427) );
  MUX U950 ( .IN0(n2167), .IN1(n428), .SEL(n2168), .F(n2150) );
  IV U951 ( .A(n2169), .Z(n428) );
  MUX U952 ( .IN0(n4899), .IN1(n4772), .SEL(n4773), .F(n4886) );
  MUX U953 ( .IN0(n4882), .IN1(n429), .SEL(n4883), .F(n4869) );
  IV U954 ( .A(n4884), .Z(n429) );
  MUX U955 ( .IN0(n1707), .IN1(n430), .SEL(n1708), .F(n1668) );
  IV U956 ( .A(n1709), .Z(n430) );
  MUX U957 ( .IN0(n1664), .IN1(n431), .SEL(n1665), .F(n1625) );
  IV U958 ( .A(n1666), .Z(n431) );
  MUX U959 ( .IN0(n1759), .IN1(n432), .SEL(n1760), .F(n1720) );
  IV U960 ( .A(n1761), .Z(n432) );
  MUX U961 ( .IN0(n2181), .IN1(n433), .SEL(n1738), .F(n2164) );
  IV U962 ( .A(n1736), .Z(n433) );
  XNOR U963 ( .A(n2391), .B(n2383), .Z(n2163) );
  MUX U964 ( .IN0(n1647), .IN1(n434), .SEL(n1648), .F(n1608) );
  IV U965 ( .A(n1649), .Z(n434) );
  MUX U966 ( .IN0(n2762), .IN1(n2629), .SEL(n2631), .F(n2751) );
  XNOR U967 ( .A(n4863), .B(n4864), .Z(n4730) );
  MUX U968 ( .IN0(n4723), .IN1(n4725), .SEL(n4724), .F(n4702) );
  MUX U969 ( .IN0(n4698), .IN1(n435), .SEL(n4699), .F(n4677) );
  IV U970 ( .A(n4700), .Z(n435) );
  MUX U971 ( .IN0(n436), .IN1(n1595), .SEL(n1596), .F(n1556) );
  IV U972 ( .A(n1597), .Z(n436) );
  MUX U973 ( .IN0(n2137), .IN1(n437), .SEL(n2138), .F(n2120) );
  IV U974 ( .A(n2139), .Z(n437) );
  MUX U975 ( .IN0(n1651), .IN1(n438), .SEL(n1652), .F(n1612) );
  IV U976 ( .A(n1653), .Z(n438) );
  MUX U977 ( .IN0(n2571), .IN1(n439), .SEL(n2572), .F(n2550) );
  IV U978 ( .A(n2573), .Z(n439) );
  MUX U979 ( .IN0(n2736), .IN1(n440), .SEL(n2737), .F(n2725) );
  IV U980 ( .A(n2738), .Z(n440) );
  XNOR U981 ( .A(n2616), .B(n2598), .Z(n2602) );
  MUX U982 ( .IN0(n2847), .IN1(n2699), .SEL(n2700), .F(n2831) );
  MUX U983 ( .IN0(n2821), .IN1(n2836), .SEL(n2823), .F(n2805) );
  MUX U984 ( .IN0(n441), .IN1(n2366), .SEL(n2367), .F(n2355) );
  IV U985 ( .A(n2368), .Z(n441) );
  MUX U986 ( .IN0(n4672), .IN1(n442), .SEL(n4673), .F(n4651) );
  IV U987 ( .A(n4674), .Z(n442) );
  XNOR U988 ( .A(n4850), .B(n4851), .Z(n4709) );
  MUX U989 ( .IN0(n4960), .IN1(n4798), .SEL(n4799), .F(n4944) );
  MUX U990 ( .IN0(n4940), .IN1(n4954), .SEL(n4942), .F(n4924) );
  MUX U991 ( .IN0(n4934), .IN1(n4949), .SEL(n4936), .F(n4918) );
  MUX U992 ( .IN0(n2099), .IN1(n443), .SEL(n2100), .F(n2082) );
  IV U993 ( .A(n2101), .Z(n443) );
  XNOR U994 ( .A(n1584), .B(n1548), .Z(n1552) );
  MUX U995 ( .IN0(n2937), .IN1(n2880), .SEL(n2881), .F(n2921) );
  MUX U996 ( .IN0(n2911), .IN1(n2926), .SEL(n2913), .F(n2895) );
  XNOR U997 ( .A(n2732), .B(n2733), .Z(n2587) );
  MUX U998 ( .IN0(n5054), .IN1(n4991), .SEL(n4992), .F(n5038) );
  MUX U999 ( .IN0(n4830), .IN1(n444), .SEL(n4831), .F(n4817) );
  IV U1000 ( .A(n4832), .Z(n444) );
  XNOR U1001 ( .A(n4837), .B(n4838), .Z(n4688) );
  MUX U1002 ( .IN0(n4780), .IN1(n445), .SEL(n4781), .F(n4776) );
  IV U1003 ( .A(n4782), .Z(n445) );
  MUX U1004 ( .IN0(n1603), .IN1(n446), .SEL(n1604), .F(n1564) );
  IV U1005 ( .A(n1605), .Z(n446) );
  MUX U1006 ( .IN0(n2709), .IN1(n447), .SEL(n2710), .F(n2517) );
  IV U1007 ( .A(n2711), .Z(n447) );
  MUX U1008 ( .IN0(n4810), .IN1(n448), .SEL(n4811), .F(n4618) );
  IV U1009 ( .A(n4812), .Z(n448) );
  MUX U1010 ( .IN0(n2353), .IN1(n449), .SEL(n2112), .F(n2342) );
  IV U1011 ( .A(n2111), .Z(n449) );
  MUX U1012 ( .IN0(n2113), .IN1(n450), .SEL(n1582), .F(n2096) );
  IV U1013 ( .A(n1580), .Z(n450) );
  MUX U1014 ( .IN0(n451), .IN1(n2073), .SEL(n2074), .F(n1456) );
  IV U1015 ( .A(n2075), .Z(n451) );
  XOR U1016 ( .A(n1514), .B(n1513), .Z(n1527) );
  MUX U1017 ( .IN0(n2502), .IN1(n452), .SEL(n2503), .F(n2305) );
  IV U1018 ( .A(n2504), .Z(n452) );
  XNOR U1019 ( .A(n2712), .B(n2704), .Z(n2526) );
  MUX U1020 ( .IN0(n2538), .IN1(n2540), .SEL(n2539), .F(n2506) );
  MUX U1021 ( .IN0(n2349), .IN1(n453), .SEL(n2350), .F(n2338) );
  IV U1022 ( .A(n2351), .Z(n453) );
  MUX U1023 ( .IN0(n5083), .IN1(n5086), .SEL(n5084), .F(n4569) );
  MUX U1024 ( .IN0(n4987), .IN1(n5015), .SEL(n4989), .F(n4472) );
  MUX U1025 ( .IN0(n4997), .IN1(n5007), .SEL(n4999), .F(n4477) );
  MUX U1026 ( .IN0(n4603), .IN1(n454), .SEL(n4604), .F(n4167) );
  IV U1027 ( .A(n4605), .Z(n454) );
  MUX U1028 ( .IN0(n4639), .IN1(n4641), .SEL(n4640), .F(n4607) );
  MUX U1029 ( .IN0(n455), .IN1(n1416), .SEL(n1417), .F(n1349) );
  IV U1030 ( .A(n1418), .Z(n455) );
  XNOR U1031 ( .A(n1528), .B(n1492), .Z(n1496) );
  XNOR U1032 ( .A(n1467), .B(n1434), .Z(n1438) );
  XOR U1033 ( .A(n1475), .B(n1474), .Z(n1488) );
  XNOR U1034 ( .A(n2969), .B(n2970), .Z(n2023) );
  MUX U1035 ( .IN0(n456), .IN1(n4158), .SEL(n4159), .F(n4141) );
  IV U1036 ( .A(n4160), .Z(n456) );
  MUX U1037 ( .IN0(n4290), .IN1(n457), .SEL(n4291), .F(n4279) );
  IV U1038 ( .A(n4292), .Z(n457) );
  MUX U1039 ( .IN0(n458), .IN1(n1313), .SEL(n1314), .F(n1250) );
  IV U1040 ( .A(n1315), .Z(n458) );
  MUX U1041 ( .IN0(n1295), .IN1(n459), .SEL(n1296), .F(n1232) );
  IV U1042 ( .A(n1297), .Z(n459) );
  MUX U1043 ( .IN0(n460), .IN1(n4272), .SEL(n4273), .F(n4259) );
  IV U1044 ( .A(n4274), .Z(n460) );
  MUX U1045 ( .IN0(n461), .IN1(n2059), .SEL(n2060), .F(n1400) );
  IV U1046 ( .A(n2061), .Z(n461) );
  MUX U1047 ( .IN0(n462), .IN1(n4591), .SEL(n4555), .F(n4589) );
  IV U1048 ( .A(n4556), .Z(n462) );
  MUX U1049 ( .IN0(n463), .IN1(n4437), .SEL(n4438), .F(n4426) );
  IV U1050 ( .A(n4439), .Z(n463) );
  MUX U1051 ( .IN0(n464), .IN1(n1171), .SEL(n1172), .F(n1119) );
  IV U1052 ( .A(n1173), .Z(n464) );
  MUX U1053 ( .IN0(n465), .IN1(n4090), .SEL(n4091), .F(n4073) );
  IV U1054 ( .A(n4092), .Z(n465) );
  MUX U1055 ( .IN0(n4240), .IN1(n466), .SEL(n4241), .F(n4227) );
  IV U1056 ( .A(n4242), .Z(n466) );
  MUX U1057 ( .IN0(n467), .IN1(n4220), .SEL(n4221), .F(n4207) );
  IV U1058 ( .A(n4222), .Z(n467) );
  MUX U1059 ( .IN0(n468), .IN1(n1265), .SEL(n1266), .F(n1211) );
  IV U1060 ( .A(n1267), .Z(n468) );
  MUX U1061 ( .IN0(n469), .IN1(n1050), .SEL(n1051), .F(n1013) );
  IV U1062 ( .A(n1052), .Z(n469) );
  MUX U1063 ( .IN0(n470), .IN1(n4393), .SEL(n4394), .F(n4380) );
  IV U1064 ( .A(n4395), .Z(n470) );
  MUX U1065 ( .IN0(n1004), .IN1(n471), .SEL(n1005), .F(n969) );
  IV U1066 ( .A(n1006), .Z(n471) );
  MUX U1067 ( .IN0(n4387), .IN1(n472), .SEL(n4388), .F(n4374) );
  IV U1068 ( .A(n4389), .Z(n472) );
  MUX U1069 ( .IN0(n1032), .IN1(n473), .SEL(n1033), .F(n994) );
  IV U1070 ( .A(n1034), .Z(n473) );
  MUX U1071 ( .IN0(n474), .IN1(n3963), .SEL(n3964), .F(n3897) );
  IV U1072 ( .A(n3965), .Z(n474) );
  MUX U1073 ( .IN0(n4188), .IN1(n475), .SEL(n4189), .F(n3915) );
  IV U1074 ( .A(n4190), .Z(n475) );
  MUX U1075 ( .IN0(n476), .IN1(n3905), .SEL(n3906), .F(n3839) );
  IV U1076 ( .A(n3907), .Z(n476) );
  MUX U1077 ( .IN0(n477), .IN1(n987), .SEL(n988), .F(n955) );
  IV U1078 ( .A(n989), .Z(n477) );
  MUX U1079 ( .IN0(n478), .IN1(n3858), .SEL(n3859), .F(n3792) );
  IV U1080 ( .A(n3860), .Z(n478) );
  MUX U1081 ( .IN0(n3823), .IN1(n479), .SEL(n3824), .F(n3757) );
  IV U1082 ( .A(n3825), .Z(n479) );
  MUX U1083 ( .IN0(n3717), .IN1(n480), .SEL(n3718), .F(n3651) );
  IV U1084 ( .A(n3719), .Z(n480) );
  MUX U1085 ( .IN0(n481), .IN1(n3634), .SEL(n3635), .F(n3570) );
  IV U1086 ( .A(n3636), .Z(n481) );
  MUX U1087 ( .IN0(n482), .IN1(n3642), .SEL(n3643), .F(n3578) );
  IV U1088 ( .A(n3644), .Z(n482) );
  MUX U1089 ( .IN0(n3603), .IN1(n483), .SEL(n3604), .F(n3539) );
  IV U1090 ( .A(n3605), .Z(n483) );
  MUX U1091 ( .IN0(n3562), .IN1(n484), .SEL(n3563), .F(n3498) );
  IV U1092 ( .A(n3564), .Z(n484) );
  MUX U1093 ( .IN0(n485), .IN1(n3556), .SEL(n3557), .F(n3492) );
  IV U1094 ( .A(n3558), .Z(n485) );
  MUX U1095 ( .IN0(n3548), .IN1(n486), .SEL(n3549), .F(n3484) );
  IV U1096 ( .A(n3550), .Z(n486) );
  MUX U1097 ( .IN0(n487), .IN1(n3346), .SEL(n3347), .F(n3296) );
  IV U1098 ( .A(n3348), .Z(n487) );
  MUX U1099 ( .IN0(n3304), .IN1(n488), .SEL(n3305), .F(n3255) );
  IV U1100 ( .A(n3306), .Z(n488) );
  MUX U1101 ( .IN0(n489), .IN1(n3182), .SEL(n3183), .F(n3149) );
  IV U1102 ( .A(n3184), .Z(n489) );
  XNOR U1103 ( .A(n2063), .B(n1449), .Z(n1453) );
  MUX U1104 ( .IN0(n4305), .IN1(n490), .SEL(n4306), .F(n4294) );
  IV U1105 ( .A(n4307), .Z(n490) );
  MUX U1106 ( .IN0(n1299), .IN1(n491), .SEL(n1300), .F(n1236) );
  IV U1107 ( .A(n1301), .Z(n491) );
  MUX U1108 ( .IN0(n4257), .IN1(n492), .SEL(n4129), .F(n4244) );
  IV U1109 ( .A(n4128), .Z(n492) );
  MUX U1110 ( .IN0(n1085), .IN1(n493), .SEL(n1086), .F(n1036) );
  IV U1111 ( .A(n1087), .Z(n493) );
  MUX U1112 ( .IN0(n4205), .IN1(n494), .SEL(n4061), .F(n4192) );
  IV U1113 ( .A(n4060), .Z(n494) );
  MUX U1114 ( .IN0(n3787), .IN1(n495), .SEL(n3788), .F(n3721) );
  IV U1115 ( .A(n3789), .Z(n495) );
  MUX U1116 ( .IN0(n3695), .IN1(n496), .SEL(n3696), .F(n3630) );
  IV U1117 ( .A(n3697), .Z(n496) );
  MUX U1118 ( .IN0(n3672), .IN1(n497), .SEL(n3673), .F(n3607) );
  IV U1119 ( .A(n3674), .Z(n497) );
  MUX U1120 ( .IN0(n3526), .IN1(n498), .SEL(n3527), .F(n3461) );
  IV U1121 ( .A(n3528), .Z(n498) );
  MUX U1122 ( .IN0(n499), .IN1(n3335), .SEL(n3336), .F(n3286) );
  IV U1123 ( .A(n3337), .Z(n499) );
  MUX U1124 ( .IN0(n1403), .IN1(n500), .SEL(n1404), .F(n1338) );
  IV U1125 ( .A(n1405), .Z(n500) );
  XNOR U1126 ( .A(n4558), .B(n4552), .Z(n4360) );
  XNOR U1127 ( .A(n4462), .B(n4454), .Z(n4358) );
  XNOR U1128 ( .A(n4148), .B(n4134), .Z(n4138) );
  XNOR U1129 ( .A(n1302), .B(n1242), .Z(n1246) );
  MUX U1130 ( .IN0(n1341), .IN1(n1406), .SEL(n1343), .F(n1274) );
  XNOR U1131 ( .A(n1254), .B(n1203), .Z(n1208) );
  MUX U1132 ( .IN0(n4130), .IN1(n501), .SEL(n4007), .F(n4113) );
  IV U1133 ( .A(n4006), .Z(n501) );
  MUX U1134 ( .IN0(n1122), .IN1(n502), .SEL(n1123), .F(n1076) );
  IV U1135 ( .A(n1124), .Z(n502) );
  XNOR U1136 ( .A(n4418), .B(n4410), .Z(n4334) );
  XNOR U1137 ( .A(n4080), .B(n4066), .Z(n4070) );
  XNOR U1138 ( .A(n4511), .B(n4505), .Z(n4330) );
  MUX U1139 ( .IN0(n4062), .IN1(n503), .SEL(n3983), .F(n4045) );
  IV U1140 ( .A(n3982), .Z(n503) );
  XNOR U1141 ( .A(n4029), .B(n3956), .Z(n3960) );
  XNOR U1142 ( .A(n4484), .B(n3942), .Z(n3946) );
  XNOR U1143 ( .A(n936), .B(n909), .Z(n913) );
  XNOR U1144 ( .A(n3930), .B(n3867), .Z(n3871) );
  MUX U1145 ( .IN0(n932), .IN1(n961), .SEL(n934), .F(n896) );
  MUX U1146 ( .IN0(n3842), .IN1(n504), .SEL(n3843), .F(n3776) );
  IV U1147 ( .A(n3844), .Z(n504) );
  XNOR U1148 ( .A(n3741), .B(n3678), .Z(n3682) );
  MUX U1149 ( .IN0(n505), .IN1(n865), .SEL(n866), .F(n847) );
  IV U1150 ( .A(n867), .Z(n505) );
  MUX U1151 ( .IN0(n3598), .IN1(n506), .SEL(n3599), .F(n3534) );
  IV U1152 ( .A(n3600), .Z(n506) );
  MUX U1153 ( .IN0(n3581), .IN1(n507), .SEL(n3582), .F(n3520) );
  IV U1154 ( .A(n3583), .Z(n507) );
  XNOR U1155 ( .A(n3473), .B(n3417), .Z(n3421) );
  XNOR U1156 ( .A(n3437), .B(n3381), .Z(n3385) );
  XNOR U1157 ( .A(n3423), .B(n3364), .Z(n3368) );
  XNOR U1158 ( .A(n3219), .B(n3175), .Z(n3179) );
  XNOR U1159 ( .A(n3209), .B(n3165), .Z(n3170) );
  MUX U1160 ( .IN0(n508), .IN1(n3097), .SEL(n3098), .F(n3074) );
  IV U1161 ( .A(n3099), .Z(n508) );
  XOR U1162 ( .A(n4365), .B(n4366), .Z(n4015) );
  MUX U1163 ( .IN0(n4020), .IN1(n509), .SEL(n4021), .F(n4014) );
  IV U1164 ( .A(n4022), .Z(n509) );
  MUX U1165 ( .IN0(n1330), .IN1(n510), .SEL(n1331), .F(n1268) );
  IV U1166 ( .A(n1332), .Z(n510) );
  XOR U1167 ( .A(n4341), .B(n4342), .Z(n3991) );
  MUX U1168 ( .IN0(n3996), .IN1(n511), .SEL(n2997), .F(n3990) );
  IV U1169 ( .A(n2996), .Z(n511) );
  XOR U1170 ( .A(n4317), .B(n4318), .Z(n3967) );
  MUX U1171 ( .IN0(n3972), .IN1(n512), .SEL(n2989), .F(n3966) );
  IV U1172 ( .A(n2988), .Z(n512) );
  XOR U1173 ( .A(n944), .B(n943), .Z(n931) );
  XOR U1174 ( .A(n3881), .B(n3880), .Z(n3863) );
  MUX U1175 ( .IN0(n3702), .IN1(n513), .SEL(n3703), .F(n3637) );
  IV U1176 ( .A(n3704), .Z(n513) );
  XOR U1177 ( .A(n3431), .B(n3430), .Z(n3413) );
  MUX U1178 ( .IN0(n3450), .IN1(n514), .SEL(n3451), .F(n3391) );
  IV U1179 ( .A(n3452), .Z(n514) );
  MUX U1180 ( .IN0(n515), .IN1(n3341), .SEL(n3342), .F(n3290) );
  IV U1181 ( .A(n3343), .Z(n515) );
  XOR U1182 ( .A(n3235), .B(n3234), .Z(n3241) );
  XOR U1183 ( .A(n3117), .B(n3116), .Z(n3102) );
  XOR U1184 ( .A(n3088), .B(n3087), .Z(n3078) );
  XOR U1185 ( .A(n3058), .B(n3057), .Z(n3049) );
  MUX U1186 ( .IN0(n1283), .IN1(\_MAC/_MULT/MULT/S[3][1][2] ), .SEL(n5114), 
        .F(n1220) );
  XOR U1187 ( .A(n1112), .B(n1110), .Z(n1150) );
  XOR U1188 ( .A(n1028), .B(n1027), .Z(n1068) );
  XOR U1189 ( .A(n992), .B(n991), .Z(n1018) );
  XOR U1190 ( .A(n960), .B(n959), .Z(n982) );
  MUX U1191 ( .IN0(n920), .IN1(\_MAC/_MULT/MULT/S[3][1][10] ), .SEL(n5122), 
        .F(n516) );
  IV U1192 ( .A(n516), .Z(n889) );
  ANDN U1193 ( .A(n852), .B(n853), .Z(n838) );
  XOR U1194 ( .A(n833), .B(n822), .Z(n832) );
  XOR U1195 ( .A(n3252), .B(n3251), .Z(n3244) );
  MUX U1196 ( .IN0(n816), .IN1(\_MAC/_MULT/MULT/S[3][1][15] ), .SEL(n5127), 
        .F(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[16] ) );
  AND U1197 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[19] ), .B(
        \_MAC/_MULT/MULT/S[3][1][19] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[20] ) );
  AND U1198 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[23] ), .B(
        \_MAC/_MULT/MULT/S[3][1][23] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[24] ) );
  AND U1199 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[28] ), .B(
        \_MAC/_MULT/MULT/S[3][1][28] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[29] ) );
  MUX U1200 ( .IN0(n517), .IN1(n3025), .SEL(n3026), .F(n3009) );
  IV U1201 ( .A(n3027), .Z(n517) );
  MUX U1202 ( .IN0(n518), .IN1(n1989), .SEL(n1990), .F(n1948) );
  IV U1203 ( .A(n1991), .Z(n518) );
  MUX U1204 ( .IN0(n2286), .IN1(n519), .SEL(n2287), .F(n2269) );
  IV U1205 ( .A(n2288), .Z(n519) );
  MUX U1206 ( .IN0(n520), .IN1(n1994), .SEL(n1995), .F(n1953) );
  IV U1207 ( .A(n1996), .Z(n520) );
  MUX U1208 ( .IN0(n521), .IN1(n2476), .SEL(n2477), .F(n2465) );
  IV U1209 ( .A(n2478), .Z(n521) );
  MUX U1210 ( .IN0(n1997), .IN1(n522), .SEL(n1998), .F(n1956) );
  IV U1211 ( .A(n1999), .Z(n522) );
  MUX U1212 ( .IN0(n1904), .IN1(n523), .SEL(n1905), .F(n1863) );
  IV U1213 ( .A(n1906), .Z(n523) );
  MUX U1214 ( .IN0(n2463), .IN1(n524), .SEL(n2282), .F(n2452) );
  IV U1215 ( .A(n2281), .Z(n524) );
  MUX U1216 ( .IN0(n2283), .IN1(n525), .SEL(n1974), .F(n2266) );
  IV U1217 ( .A(n1972), .Z(n525) );
  MUX U1218 ( .IN0(n526), .IN1(n2243), .SEL(n2244), .F(n2226) );
  IV U1219 ( .A(n2245), .Z(n526) );
  MUX U1220 ( .IN0(n1926), .IN1(n527), .SEL(n1927), .F(n1887) );
  IV U1221 ( .A(n1928), .Z(n527) );
  MUX U1222 ( .IN0(n528), .IN1(n1829), .SEL(n1830), .F(n1790) );
  IV U1223 ( .A(n1831), .Z(n528) );
  MUX U1224 ( .IN0(n1820), .IN1(n529), .SEL(n1821), .F(n1781) );
  IV U1225 ( .A(n1822), .Z(n529) );
  MUX U1226 ( .IN0(n530), .IN1(n1834), .SEL(n1835), .F(n1795) );
  IV U1227 ( .A(n1836), .Z(n530) );
  MUX U1228 ( .IN0(n1842), .IN1(n531), .SEL(n1843), .F(n1803) );
  IV U1229 ( .A(n1844), .Z(n531) );
  XNOR U1230 ( .A(n2233), .B(n2219), .Z(n2223) );
  MUX U1231 ( .IN0(n2437), .IN1(n532), .SEL(n2438), .F(n2426) );
  IV U1232 ( .A(n2439), .Z(n532) );
  MUX U1233 ( .IN0(n1837), .IN1(n533), .SEL(n1838), .F(n1798) );
  IV U1234 ( .A(n1839), .Z(n533) );
  MUX U1235 ( .IN0(n2419), .IN1(n534), .SEL(n2214), .F(n2408) );
  IV U1236 ( .A(n2213), .Z(n534) );
  MUX U1237 ( .IN0(n2215), .IN1(n535), .SEL(n1816), .F(n2198) );
  IV U1238 ( .A(n1814), .Z(n535) );
  MUX U1239 ( .IN0(n536), .IN1(n2175), .SEL(n2176), .F(n2158) );
  IV U1240 ( .A(n2177), .Z(n536) );
  XNOR U1241 ( .A(n1740), .B(n1704), .Z(n1708) );
  MUX U1242 ( .IN0(n2634), .IN1(n537), .SEL(n2635), .F(n2613) );
  IV U1243 ( .A(n2636), .Z(n537) );
  MUX U1244 ( .IN0(n2639), .IN1(n538), .SEL(n2640), .F(n2618) );
  IV U1245 ( .A(n2641), .Z(n538) );
  MUX U1246 ( .IN0(n4735), .IN1(n539), .SEL(n4736), .F(n4714) );
  IV U1247 ( .A(n4737), .Z(n539) );
  XNOR U1248 ( .A(n4891), .B(n4883), .Z(n4753) );
  MUX U1249 ( .IN0(n4740), .IN1(n540), .SEL(n4741), .F(n4719) );
  IV U1250 ( .A(n4742), .Z(n540) );
  MUX U1251 ( .IN0(n541), .IN1(n1673), .SEL(n1674), .F(n1634) );
  IV U1252 ( .A(n1675), .Z(n541) );
  MUX U1253 ( .IN0(n1729), .IN1(n542), .SEL(n1730), .F(n1690) );
  IV U1254 ( .A(n1731), .Z(n542) );
  MUX U1255 ( .IN0(n1686), .IN1(n543), .SEL(n1687), .F(n1647) );
  IV U1256 ( .A(n1688), .Z(n543) );
  XNOR U1257 ( .A(n2765), .B(n2766), .Z(n2650) );
  MUX U1258 ( .IN0(n4862), .IN1(n544), .SEL(n4863), .F(n4849) );
  IV U1259 ( .A(n4864), .Z(n544) );
  XNOR U1260 ( .A(n2165), .B(n2151), .Z(n2155) );
  MUX U1261 ( .IN0(n2393), .IN1(n545), .SEL(n2394), .F(n2382) );
  IV U1262 ( .A(n2395), .Z(n545) );
  MUX U1263 ( .IN0(n546), .IN1(n2377), .SEL(n2378), .F(n2366) );
  IV U1264 ( .A(n2379), .Z(n546) );
  MUX U1265 ( .IN0(n1681), .IN1(n547), .SEL(n1682), .F(n1642) );
  IV U1266 ( .A(n1683), .Z(n547) );
  XNOR U1267 ( .A(n1623), .B(n1587), .Z(n1591) );
  XNOR U1268 ( .A(n2745), .B(n2737), .Z(n2589) );
  MUX U1269 ( .IN0(n2601), .IN1(n2603), .SEL(n2602), .F(n2580) );
  MUX U1270 ( .IN0(n2827), .IN1(n2841), .SEL(n2829), .F(n2811) );
  MUX U1271 ( .IN0(n5046), .IN1(n548), .SEL(n5047), .F(n5028) );
  IV U1272 ( .A(n5048), .Z(n548) );
  XNOR U1273 ( .A(n4852), .B(n4844), .Z(n4690) );
  MUX U1274 ( .IN0(n2147), .IN1(n549), .SEL(n1660), .F(n2130) );
  IV U1275 ( .A(n1658), .Z(n549) );
  XNOR U1276 ( .A(n2369), .B(n2361), .Z(n2129) );
  MUX U1277 ( .IN0(n550), .IN1(n2107), .SEL(n2108), .F(n2090) );
  IV U1278 ( .A(n2109), .Z(n550) );
  MUX U1279 ( .IN0(n2917), .IN1(n2931), .SEL(n2919), .F(n2901) );
  MUX U1280 ( .IN0(n2550), .IN1(n551), .SEL(n2551), .F(n2529) );
  IV U1281 ( .A(n2552), .Z(n551) );
  MUX U1282 ( .IN0(n2720), .IN1(n552), .SEL(n2721), .F(n2709) );
  IV U1283 ( .A(n2722), .Z(n552) );
  MUX U1284 ( .IN0(n2555), .IN1(n553), .SEL(n2556), .F(n2534) );
  IV U1285 ( .A(n2557), .Z(n553) );
  MUX U1286 ( .IN0(n2805), .IN1(n2820), .SEL(n2807), .F(n2794) );
  MUX U1287 ( .IN0(n5034), .IN1(n5050), .SEL(n5036), .F(n5016) );
  MUX U1288 ( .IN0(n4651), .IN1(n554), .SEL(n4652), .F(n4630) );
  IV U1289 ( .A(n4653), .Z(n554) );
  XNOR U1290 ( .A(n4696), .B(n4678), .Z(n4682) );
  MUX U1291 ( .IN0(n4924), .IN1(n4939), .SEL(n4926), .F(n4901) );
  MUX U1292 ( .IN0(n4918), .IN1(n4933), .SEL(n4920), .F(n4907) );
  MUX U1293 ( .IN0(n555), .IN1(n1517), .SEL(n1518), .F(n1478) );
  IV U1294 ( .A(n1519), .Z(n555) );
  MUX U1295 ( .IN0(n1573), .IN1(n556), .SEL(n1574), .F(n1534) );
  IV U1296 ( .A(n1575), .Z(n556) );
  MUX U1297 ( .IN0(n1530), .IN1(n557), .SEL(n1531), .F(n1491) );
  IV U1298 ( .A(n1532), .Z(n557) );
  MUX U1299 ( .IN0(n2895), .IN1(n2910), .SEL(n2897), .F(n2884) );
  MUX U1300 ( .IN0(n2968), .IN1(n558), .SEL(n2969), .F(n2964) );
  IV U1301 ( .A(n2970), .Z(n558) );
  MUX U1302 ( .IN0(n2714), .IN1(n559), .SEL(n2715), .F(n2703) );
  IV U1303 ( .A(n2716), .Z(n559) );
  XNOR U1304 ( .A(n2864), .B(n2865), .Z(n2847) );
  MUX U1305 ( .IN0(n4817), .IN1(n560), .SEL(n4818), .F(n4804) );
  IV U1306 ( .A(n4819), .Z(n560) );
  XNOR U1307 ( .A(n4824), .B(n4825), .Z(n4667) );
  XNOR U1308 ( .A(n4975), .B(n4976), .Z(n4960) );
  XNOR U1309 ( .A(n2097), .B(n2083), .Z(n2087) );
  XNOR U1310 ( .A(n1506), .B(n1470), .Z(n1474) );
  XNOR U1311 ( .A(n2952), .B(n2953), .Z(n2937) );
  XNOR U1312 ( .A(n2680), .B(n2681), .Z(n2666) );
  MUX U1313 ( .IN0(n561), .IN1(n2332), .SEL(n2333), .F(n2059) );
  IV U1314 ( .A(n2334), .Z(n561) );
  XNOR U1315 ( .A(n5069), .B(n5070), .Z(n5054) );
  XNOR U1316 ( .A(n4811), .B(n4812), .Z(n4646) );
  XNOR U1317 ( .A(n4781), .B(n4782), .Z(n4767) );
  MUX U1318 ( .IN0(n1525), .IN1(n562), .SEL(n1526), .F(n1486) );
  IV U1319 ( .A(n1527), .Z(n562) );
  MUX U1320 ( .IN0(n2506), .IN1(n2508), .SEL(n2507), .F(n2309) );
  MUX U1321 ( .IN0(n2707), .IN1(n2524), .SEL(n2526), .F(n2496) );
  MUX U1322 ( .IN0(n4477), .IN1(n563), .SEL(n4478), .F(n4464) );
  IV U1323 ( .A(n4479), .Z(n563) );
  MUX U1324 ( .IN0(n564), .IN1(n1349), .SEL(n1350), .F(n1287) );
  IV U1325 ( .A(n1351), .Z(n564) );
  MUX U1326 ( .IN0(n565), .IN1(n1391), .SEL(n1392), .F(n1327) );
  IV U1327 ( .A(n1393), .Z(n565) );
  MUX U1328 ( .IN0(n2338), .IN1(n566), .SEL(n2339), .F(n2325) );
  IV U1329 ( .A(n2340), .Z(n566) );
  MUX U1330 ( .IN0(n567), .IN1(n4459), .SEL(n4460), .F(n4448) );
  IV U1331 ( .A(n4461), .Z(n567) );
  MUX U1332 ( .IN0(n568), .IN1(n4593), .SEL(n4564), .F(n4591) );
  IV U1333 ( .A(n4565), .Z(n568) );
  MUX U1334 ( .IN0(n569), .IN1(n4141), .SEL(n4142), .F(n4124) );
  IV U1335 ( .A(n4143), .Z(n569) );
  MUX U1336 ( .IN0(n4279), .IN1(n570), .SEL(n4280), .F(n4266) );
  IV U1337 ( .A(n4281), .Z(n570) );
  MUX U1338 ( .IN0(n571), .IN1(n1250), .SEL(n1251), .F(n1197) );
  IV U1339 ( .A(n1252), .Z(n571) );
  MUX U1340 ( .IN0(n1232), .IN1(n572), .SEL(n1233), .F(n1179) );
  IV U1341 ( .A(n1234), .Z(n572) );
  MUX U1342 ( .IN0(n573), .IN1(n4246), .SEL(n4247), .F(n4233) );
  IV U1343 ( .A(n4248), .Z(n573) );
  MUX U1344 ( .IN0(n574), .IN1(n1119), .SEL(n1120), .F(n1073) );
  IV U1345 ( .A(n1121), .Z(n574) );
  MUX U1346 ( .IN0(n4522), .IN1(n575), .SEL(n4523), .F(n4513) );
  IV U1347 ( .A(n4524), .Z(n575) );
  MUX U1348 ( .IN0(n576), .IN1(n4415), .SEL(n4416), .F(n4404) );
  IV U1349 ( .A(n4417), .Z(n576) );
  MUX U1350 ( .IN0(n4420), .IN1(n577), .SEL(n4421), .F(n4409) );
  IV U1351 ( .A(n4422), .Z(n577) );
  MUX U1352 ( .IN0(n4082), .IN1(n578), .SEL(n4083), .F(n4065) );
  IV U1353 ( .A(n4084), .Z(n578) );
  MUX U1354 ( .IN0(n1090), .IN1(n579), .SEL(n1091), .F(n1041) );
  IV U1355 ( .A(n1092), .Z(n579) );
  MUX U1356 ( .IN0(n580), .IN1(n4073), .SEL(n4074), .F(n4056) );
  IV U1357 ( .A(n4075), .Z(n580) );
  MUX U1358 ( .IN0(n581), .IN1(n4583), .SEL(n4517), .F(n4581) );
  IV U1359 ( .A(n4518), .Z(n581) );
  MUX U1360 ( .IN0(n582), .IN1(n1013), .SEL(n1014), .F(n978) );
  IV U1361 ( .A(n1015), .Z(n582) );
  MUX U1362 ( .IN0(n583), .IN1(n4194), .SEL(n4195), .F(n4025) );
  IV U1363 ( .A(n4196), .Z(n583) );
  MUX U1364 ( .IN0(n584), .IN1(n4310), .SEL(n4311), .F(n3924) );
  IV U1365 ( .A(n4312), .Z(n584) );
  MUX U1366 ( .IN0(n3932), .IN1(n585), .SEL(n3933), .F(n3866) );
  IV U1367 ( .A(n3934), .Z(n585) );
  MUX U1368 ( .IN0(n586), .IN1(n3897), .SEL(n3898), .F(n3831) );
  IV U1369 ( .A(n3899), .Z(n586) );
  MUX U1370 ( .IN0(n3889), .IN1(n587), .SEL(n3890), .F(n3823) );
  IV U1371 ( .A(n3891), .Z(n587) );
  MUX U1372 ( .IN0(n588), .IN1(n3883), .SEL(n3884), .F(n3817) );
  IV U1373 ( .A(n3885), .Z(n588) );
  MUX U1374 ( .IN0(n589), .IN1(n3773), .SEL(n3774), .F(n3707) );
  IV U1375 ( .A(n3775), .Z(n589) );
  MUX U1376 ( .IN0(n590), .IN1(n3726), .SEL(n3727), .F(n3660) );
  IV U1377 ( .A(n3728), .Z(n590) );
  MUX U1378 ( .IN0(n908), .IN1(n591), .SEL(n909), .F(n876) );
  IV U1379 ( .A(n910), .Z(n591) );
  MUX U1380 ( .IN0(n592), .IN1(n3570), .SEL(n3571), .F(n3508) );
  IV U1381 ( .A(n3572), .Z(n592) );
  MUX U1382 ( .IN0(n593), .IN1(n3467), .SEL(n3468), .F(n3408) );
  IV U1383 ( .A(n3469), .Z(n593) );
  MUX U1384 ( .IN0(n594), .IN1(n3371), .SEL(n3372), .F(n3321) );
  IV U1385 ( .A(n3373), .Z(n594) );
  MUX U1386 ( .IN0(n595), .IN1(n3247), .SEL(n3248), .F(n3203) );
  IV U1387 ( .A(n3249), .Z(n595) );
  MUX U1388 ( .IN0(n596), .IN1(n3149), .SEL(n3150), .F(n3119) );
  IV U1389 ( .A(n3151), .Z(n596) );
  XNOR U1390 ( .A(n4633), .B(n4604), .Z(n4608) );
  MUX U1391 ( .IN0(n2079), .IN1(n597), .SEL(n1504), .F(n2062) );
  IV U1392 ( .A(n1502), .Z(n597) );
  XOR U1393 ( .A(n1439), .B(n1438), .Z(n1421) );
  MUX U1394 ( .IN0(n4294), .IN1(n598), .SEL(n4180), .F(n4283) );
  IV U1395 ( .A(n4179), .Z(n598) );
  MUX U1396 ( .IN0(n599), .IN1(n955), .SEL(n956), .F(n926) );
  IV U1397 ( .A(n957), .Z(n599) );
  MUX U1398 ( .IN0(n600), .IN1(n886), .SEL(n887), .F(n865) );
  IV U1399 ( .A(n888), .Z(n600) );
  MUX U1400 ( .IN0(n601), .IN1(n3517), .SEL(n3518), .F(n3455) );
  IV U1401 ( .A(n3519), .Z(n601) );
  MUX U1402 ( .IN0(n3136), .IN1(n602), .SEL(n3137), .F(n3103) );
  IV U1403 ( .A(n3138), .Z(n602) );
  XNOR U1404 ( .A(n1422), .B(n1358), .Z(n1362) );
  XNOR U1405 ( .A(n1379), .B(n1320), .Z(n1324) );
  XNOR U1406 ( .A(n4549), .B(n4541), .Z(n4354) );
  XNOR U1407 ( .A(n4451), .B(n4443), .Z(n4352) );
  XNOR U1408 ( .A(n4131), .B(n4117), .Z(n4121) );
  MUX U1409 ( .IN0(n4147), .IN1(n603), .SEL(n4013), .F(n4130) );
  IV U1410 ( .A(n4012), .Z(n603) );
  XNOR U1411 ( .A(n1239), .B(n1189), .Z(n1193) );
  XNOR U1412 ( .A(n1201), .B(n1152), .Z(n1155) );
  XNOR U1413 ( .A(n4249), .B(n4241), .Z(n4112) );
  XNOR U1414 ( .A(n1125), .B(n1082), .Z(n1086) );
  MUX U1415 ( .IN0(n4079), .IN1(n604), .SEL(n3989), .F(n4062) );
  IV U1416 ( .A(n3988), .Z(n604) );
  MUX U1417 ( .IN0(n605), .IN1(n1159), .SEL(n1160), .F(n1107) );
  IV U1418 ( .A(n1161), .Z(n605) );
  XNOR U1419 ( .A(n4502), .B(n4494), .Z(n4324) );
  XNOR U1420 ( .A(n4396), .B(n4388), .Z(n4322) );
  XNOR U1421 ( .A(n4046), .B(n4032), .Z(n4036) );
  XNOR U1422 ( .A(n1002), .B(n970), .Z(n974) );
  XNOR U1423 ( .A(n993), .B(n962), .Z(n965) );
  XNOR U1424 ( .A(n4197), .B(n4189), .Z(n4044) );
  XNOR U1425 ( .A(n3939), .B(n3876), .Z(n3880) );
  MUX U1426 ( .IN0(n3927), .IN1(n606), .SEL(n3928), .F(n3861) );
  IV U1427 ( .A(n3929), .Z(n606) );
  MUX U1428 ( .IN0(n3908), .IN1(n607), .SEL(n3909), .F(n3842) );
  IV U1429 ( .A(n3910), .Z(n607) );
  XNOR U1430 ( .A(n3845), .B(n3784), .Z(n3788) );
  MUX U1431 ( .IN0(n902), .IN1(n608), .SEL(n903), .F(n872) );
  IV U1432 ( .A(n904), .Z(n608) );
  XNOR U1433 ( .A(n3798), .B(n3735), .Z(n3739) );
  XNOR U1434 ( .A(n3755), .B(n3692), .Z(n3696) );
  XNOR U1435 ( .A(n3648), .B(n3586), .Z(n3591) );
  XNOR U1436 ( .A(n3610), .B(n3549), .Z(n3553) );
  XNOR U1437 ( .A(n3601), .B(n3540), .Z(n3544) );
  XNOR U1438 ( .A(n3560), .B(n3499), .Z(n3505) );
  MUX U1439 ( .IN0(n3458), .IN1(n609), .SEL(n3459), .F(n3403) );
  IV U1440 ( .A(n3460), .Z(n609) );
  XNOR U1441 ( .A(n3361), .B(n3314), .Z(n3318) );
  XNOR U1442 ( .A(n3352), .B(n3305), .Z(n3309) );
  XNOR U1443 ( .A(n3325), .B(n3279), .Z(n3282) );
  MUX U1444 ( .IN0(n610), .IN1(n3286), .SEL(n3287), .F(n3237) );
  IV U1445 ( .A(n3288), .Z(n610) );
  XNOR U1446 ( .A(n3172), .B(n3142), .Z(n3146) );
  MUX U1447 ( .IN0(n3160), .IN1(n611), .SEL(n3161), .F(n3130) );
  IV U1448 ( .A(n3162), .Z(n611) );
  MUX U1449 ( .IN0(n3051), .IN1(n612), .SEL(n3052), .F(n3035) );
  IV U1450 ( .A(n3053), .Z(n612) );
  XOR U1451 ( .A(n4577), .B(n4576), .Z(n4369) );
  XOR U1452 ( .A(n1372), .B(n1371), .Z(n1354) );
  XOR U1453 ( .A(n2042), .B(n2041), .Z(n2056) );
  MUX U1454 ( .IN0(n4014), .IN1(n613), .SEL(n3375), .F(n4008) );
  IV U1455 ( .A(n3374), .Z(n613) );
  XNOR U1456 ( .A(n1217), .B(n1278), .Z(n1271) );
  XOR U1457 ( .A(n4347), .B(n4348), .Z(n3997) );
  XOR U1458 ( .A(n1144), .B(n1143), .Z(n1124) );
  MUX U1459 ( .IN0(n3990), .IN1(n614), .SEL(n2995), .F(n3984) );
  IV U1460 ( .A(n2994), .Z(n614) );
  MUX U1461 ( .IN0(n3966), .IN1(n615), .SEL(n2987), .F(n3900) );
  IV U1462 ( .A(n2986), .Z(n615) );
  XOR U1463 ( .A(n3763), .B(n3762), .Z(n3778) );
  XOR U1464 ( .A(n3749), .B(n3748), .Z(n3731) );
  XOR U1465 ( .A(n3618), .B(n3617), .Z(n3600) );
  MUX U1466 ( .IN0(n842), .IN1(n616), .SEL(n843), .F(n828) );
  IV U1467 ( .A(n844), .Z(n616) );
  XOR U1468 ( .A(n3490), .B(n3489), .Z(n3472) );
  MUX U1469 ( .IN0(n3391), .IN1(n617), .SEL(n3392), .F(n3338) );
  IV U1470 ( .A(n3393), .Z(n617) );
  XOR U1471 ( .A(n1292), .B(n1291), .Z(n1332) );
  MUX U1472 ( .IN0(n1220), .IN1(\_MAC/_MULT/MULT/S[3][1][3] ), .SEL(n5115), 
        .F(n1167) );
  XOR U1473 ( .A(n1066), .B(n1059), .Z(n1102) );
  MUX U1474 ( .IN0(n1019), .IN1(\_MAC/_MULT/MULT/S[3][1][7] ), .SEL(n5119), 
        .F(n983) );
  ANDN U1475 ( .A(n922), .B(n923), .Z(n891) );
  XOR U1476 ( .A(n3797), .B(n3796), .Z(n3770) );
  MUX U1477 ( .IN0(n618), .IN1(\_MAC/_MULT/MULT/S[3][1][11] ), .SEL(n5123), 
        .F(n868) );
  IV U1478 ( .A(n889), .Z(n618) );
  AND U1479 ( .A(n838), .B(n839), .Z(n831) );
  XOR U1480 ( .A(n3198), .B(n3191), .Z(n3232) );
  XOR U1481 ( .A(n3102), .B(n3101), .Z(n3093) );
  XOR U1482 ( .A(n3078), .B(n3077), .Z(n3066) );
  MUX U1483 ( .IN0(n3047), .IN1(n619), .SEL(n3048), .F(n3033) );
  IV U1484 ( .A(n3049), .Z(n619) );
  MUX U1485 ( .IN0(n620), .IN1(n3042), .SEL(n3043), .F(n3025) );
  IV U1486 ( .A(n3044), .Z(n620) );
  AND U1487 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[16] ), .B(
        \_MAC/_MULT/MULT/S[3][1][16] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[17] ) );
  AND U1488 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[20] ), .B(
        \_MAC/_MULT/MULT/S[3][1][20] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[21] ) );
  AND U1489 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[24] ), .B(
        \_MAC/_MULT/MULT/S[3][1][24] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[25] ) );
  AND U1490 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[29] ), .B(
        \_MAC/_MULT/MULT/S[3][1][29] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[30] ) );
  MUX U1491 ( .IN0(n621), .IN1(n1948), .SEL(n1949), .F(n1909) );
  IV U1492 ( .A(n1950), .Z(n621) );
  MUX U1493 ( .IN0(n1939), .IN1(n622), .SEL(n1940), .F(n1900) );
  IV U1494 ( .A(n1941), .Z(n622) );
  MUX U1495 ( .IN0(n623), .IN1(n1953), .SEL(n1954), .F(n1914) );
  IV U1496 ( .A(n1955), .Z(n623) );
  MUX U1497 ( .IN0(n2474), .IN1(n624), .SEL(n2301), .F(n2463) );
  IV U1498 ( .A(n2300), .Z(n624) );
  MUX U1499 ( .IN0(n625), .IN1(n2260), .SEL(n2261), .F(n2243) );
  IV U1500 ( .A(n2262), .Z(n625) );
  MUX U1501 ( .IN0(n2252), .IN1(n626), .SEL(n2253), .F(n2235) );
  IV U1502 ( .A(n2254), .Z(n626) );
  MUX U1503 ( .IN0(n1956), .IN1(n627), .SEL(n1957), .F(n1917) );
  IV U1504 ( .A(n1958), .Z(n627) );
  MUX U1505 ( .IN0(n2459), .IN1(n628), .SEL(n2460), .F(n2448) );
  IV U1506 ( .A(n2461), .Z(n628) );
  MUX U1507 ( .IN0(n629), .IN1(n2443), .SEL(n2444), .F(n2432) );
  IV U1508 ( .A(n2445), .Z(n629) );
  MUX U1509 ( .IN0(n2266), .IN1(n630), .SEL(n1935), .F(n2249) );
  IV U1510 ( .A(n1933), .Z(n630) );
  MUX U1511 ( .IN0(n1887), .IN1(n631), .SEL(n1888), .F(n1846) );
  IV U1512 ( .A(n1889), .Z(n631) );
  XNOR U1513 ( .A(n1857), .B(n1821), .Z(n1825) );
  MUX U1514 ( .IN0(n632), .IN1(n1790), .SEL(n1791), .F(n1751) );
  IV U1515 ( .A(n1792), .Z(n632) );
  MUX U1516 ( .IN0(n2222), .IN1(n633), .SEL(n2223), .F(n2205) );
  IV U1517 ( .A(n2224), .Z(n633) );
  MUX U1518 ( .IN0(n1803), .IN1(n634), .SEL(n1804), .F(n1764) );
  IV U1519 ( .A(n1805), .Z(n634) );
  MUX U1520 ( .IN0(n2430), .IN1(n635), .SEL(n2231), .F(n2419) );
  IV U1521 ( .A(n2230), .Z(n635) );
  MUX U1522 ( .IN0(n636), .IN1(n2192), .SEL(n2193), .F(n2175) );
  IV U1523 ( .A(n2194), .Z(n636) );
  MUX U1524 ( .IN0(n2184), .IN1(n637), .SEL(n2185), .F(n2167) );
  IV U1525 ( .A(n2186), .Z(n637) );
  MUX U1526 ( .IN0(n638), .IN1(n1717), .SEL(n1718), .F(n1678) );
  IV U1527 ( .A(n1719), .Z(n638) );
  MUX U1528 ( .IN0(n1798), .IN1(n639), .SEL(n1799), .F(n1759) );
  IV U1529 ( .A(n1800), .Z(n639) );
  XNOR U1530 ( .A(n2635), .B(n2636), .Z(n2645) );
  MUX U1531 ( .IN0(n2415), .IN1(n640), .SEL(n2416), .F(n2404) );
  IV U1532 ( .A(n2417), .Z(n640) );
  MUX U1533 ( .IN0(n641), .IN1(n2399), .SEL(n2400), .F(n2388) );
  IV U1534 ( .A(n2401), .Z(n641) );
  XNOR U1535 ( .A(n4736), .B(n4737), .Z(n4746) );
  MUX U1536 ( .IN0(n2198), .IN1(n642), .SEL(n1777), .F(n2181) );
  IV U1537 ( .A(n1775), .Z(n642) );
  XNOR U1538 ( .A(n1701), .B(n1665), .Z(n1669) );
  XNOR U1539 ( .A(n2767), .B(n2759), .Z(n2631) );
  MUX U1540 ( .IN0(n2618), .IN1(n643), .SEL(n2619), .F(n2597) );
  IV U1541 ( .A(n2620), .Z(n643) );
  XNOR U1542 ( .A(n4876), .B(n4877), .Z(n4751) );
  MUX U1543 ( .IN0(n4719), .IN1(n644), .SEL(n4720), .F(n4698) );
  IV U1544 ( .A(n4721), .Z(n644) );
  MUX U1545 ( .IN0(n645), .IN1(n1634), .SEL(n1635), .F(n1595) );
  IV U1546 ( .A(n1636), .Z(n645) );
  XNOR U1547 ( .A(n1723), .B(n1687), .Z(n1691) );
  MUX U1548 ( .IN0(n2154), .IN1(n646), .SEL(n2155), .F(n2137) );
  IV U1549 ( .A(n2156), .Z(n646) );
  MUX U1550 ( .IN0(n2592), .IN1(n647), .SEL(n2593), .F(n2571) );
  IV U1551 ( .A(n2594), .Z(n647) );
  MUX U1552 ( .IN0(n2742), .IN1(n648), .SEL(n2743), .F(n2731) );
  IV U1553 ( .A(n2744), .Z(n648) );
  MUX U1554 ( .IN0(n4693), .IN1(n649), .SEL(n4694), .F(n4672) );
  IV U1555 ( .A(n4695), .Z(n649) );
  MUX U1556 ( .IN0(n4849), .IN1(n650), .SEL(n4850), .F(n4836) );
  IV U1557 ( .A(n4851), .Z(n650) );
  MUX U1558 ( .IN0(n2386), .IN1(n651), .SEL(n2163), .F(n2375) );
  IV U1559 ( .A(n2162), .Z(n651) );
  MUX U1560 ( .IN0(n652), .IN1(n2124), .SEL(n2125), .F(n2107) );
  IV U1561 ( .A(n2126), .Z(n652) );
  MUX U1562 ( .IN0(n2116), .IN1(n653), .SEL(n2117), .F(n2099) );
  IV U1563 ( .A(n2118), .Z(n653) );
  MUX U1564 ( .IN0(n654), .IN1(n1561), .SEL(n1562), .F(n1522) );
  IV U1565 ( .A(n1563), .Z(n654) );
  MUX U1566 ( .IN0(n1569), .IN1(n655), .SEL(n1570), .F(n1530) );
  IV U1567 ( .A(n1571), .Z(n655) );
  MUX U1568 ( .IN0(n1642), .IN1(n656), .SEL(n1643), .F(n1603) );
  IV U1569 ( .A(n1644), .Z(n656) );
  XNOR U1570 ( .A(n2734), .B(n2726), .Z(n2568) );
  MUX U1571 ( .IN0(n2811), .IN1(n2826), .SEL(n2813), .F(n2788) );
  MUX U1572 ( .IN0(n2857), .IN1(n2860), .SEL(n2858), .F(n2837) );
  MUX U1573 ( .IN0(n2371), .IN1(n657), .SEL(n2372), .F(n2360) );
  IV U1574 ( .A(n2373), .Z(n657) );
  MUX U1575 ( .IN0(n658), .IN1(n2355), .SEL(n2356), .F(n2344) );
  IV U1576 ( .A(n2357), .Z(n658) );
  XNOR U1577 ( .A(n4839), .B(n4831), .Z(n4669) );
  MUX U1578 ( .IN0(n4970), .IN1(n4973), .SEL(n4971), .F(n4950) );
  MUX U1579 ( .IN0(n2130), .IN1(n659), .SEL(n1621), .F(n2113) );
  IV U1580 ( .A(n1619), .Z(n659) );
  XOR U1581 ( .A(n1553), .B(n1552), .Z(n1566) );
  XNOR U1582 ( .A(n1545), .B(n1509), .Z(n1513) );
  MUX U1583 ( .IN0(n2901), .IN1(n2916), .SEL(n2903), .F(n2876) );
  MUX U1584 ( .IN0(n2947), .IN1(n2950), .SEL(n2948), .F(n2927) );
  XNOR U1585 ( .A(n2574), .B(n2556), .Z(n2560) );
  MUX U1586 ( .IN0(n2794), .IN1(n2804), .SEL(n2796), .F(n2780) );
  MUX U1587 ( .IN0(n5064), .IN1(n5067), .SEL(n5065), .F(n5046) );
  XNOR U1588 ( .A(n4675), .B(n4657), .Z(n4661) );
  MUX U1589 ( .IN0(n4907), .IN1(n4917), .SEL(n4909), .F(n4895) );
  MUX U1590 ( .IN0(n2884), .IN1(n2894), .SEL(n2886), .F(n2045) );
  MUX U1591 ( .IN0(n2510), .IN1(n660), .SEL(n2511), .F(n2315) );
  IV U1592 ( .A(n2512), .Z(n660) );
  MUX U1593 ( .IN0(n2703), .IN1(n661), .SEL(n2704), .F(n2492) );
  IV U1594 ( .A(n2705), .Z(n661) );
  XNOR U1595 ( .A(n2710), .B(n2711), .Z(n2545) );
  XNOR U1596 ( .A(n2845), .B(n2846), .Z(n2699) );
  MUX U1597 ( .IN0(n4611), .IN1(n662), .SEL(n4612), .F(n4175) );
  IV U1598 ( .A(n4613), .Z(n662) );
  MUX U1599 ( .IN0(n4618), .IN1(n663), .SEL(n4619), .F(n4296) );
  IV U1600 ( .A(n4620), .Z(n663) );
  XNOR U1601 ( .A(n4958), .B(n4959), .Z(n4798) );
  MUX U1602 ( .IN0(n664), .IN1(n1442), .SEL(n1443), .F(n1375) );
  IV U1603 ( .A(n1444), .Z(n664) );
  MUX U1604 ( .IN0(n665), .IN1(n1456), .SEL(n1457), .F(n1391) );
  IV U1605 ( .A(n1458), .Z(n665) );
  MUX U1606 ( .IN0(n2342), .IN1(n666), .SEL(n2095), .F(n2330) );
  IV U1607 ( .A(n2094), .Z(n666) );
  XNOR U1608 ( .A(n2080), .B(n2066), .Z(n2070) );
  MUX U1609 ( .IN0(n1495), .IN1(n667), .SEL(n1496), .F(n1428) );
  IV U1610 ( .A(n1497), .Z(n667) );
  XNOR U1611 ( .A(n2935), .B(n2936), .Z(n2880) );
  XNOR U1612 ( .A(n2518), .B(n2519), .Z(n2524) );
  XNOR U1613 ( .A(n2673), .B(n2663), .Z(n2667) );
  MUX U1614 ( .IN0(n668), .IN1(n4597), .SEL(n4598), .F(n4595) );
  IV U1615 ( .A(n4599), .Z(n668) );
  MUX U1616 ( .IN0(n669), .IN1(n4472), .SEL(n4473), .F(n4459) );
  IV U1617 ( .A(n4474), .Z(n669) );
  MUX U1618 ( .IN0(n1357), .IN1(n670), .SEL(n1358), .F(n1295) );
  IV U1619 ( .A(n1359), .Z(n670) );
  MUX U1620 ( .IN0(n671), .IN1(n1287), .SEL(n1288), .F(n1224) );
  IV U1621 ( .A(n1289), .Z(n671) );
  MUX U1622 ( .IN0(n672), .IN1(n4124), .SEL(n4125), .F(n4107) );
  IV U1623 ( .A(n4126), .Z(n672) );
  MUX U1624 ( .IN0(n673), .IN1(n4259), .SEL(n4260), .F(n4246) );
  IV U1625 ( .A(n4261), .Z(n673) );
  MUX U1626 ( .IN0(n1188), .IN1(n674), .SEL(n1189), .F(n1136) );
  IV U1627 ( .A(n1190), .Z(n674) );
  MUX U1628 ( .IN0(n675), .IN1(n4589), .SEL(n4544), .F(n4587) );
  IV U1629 ( .A(n4545), .Z(n675) );
  MUX U1630 ( .IN0(n676), .IN1(n4426), .SEL(n4427), .F(n4415) );
  IV U1631 ( .A(n4428), .Z(n676) );
  MUX U1632 ( .IN0(n677), .IN1(n1073), .SEL(n1074), .F(n1023) );
  IV U1633 ( .A(n1075), .Z(n677) );
  MUX U1634 ( .IN0(n4513), .IN1(n678), .SEL(n4514), .F(n4504) );
  IV U1635 ( .A(n4515), .Z(n678) );
  MUX U1636 ( .IN0(n679), .IN1(n4207), .SEL(n4208), .F(n4194) );
  IV U1637 ( .A(n4209), .Z(n679) );
  MUX U1638 ( .IN0(n680), .IN1(n4380), .SEL(n4381), .F(n4310) );
  IV U1639 ( .A(n4382), .Z(n680) );
  MUX U1640 ( .IN0(n681), .IN1(n4039), .SEL(n4040), .F(n3963) );
  IV U1641 ( .A(n4041), .Z(n681) );
  MUX U1642 ( .IN0(n4201), .IN1(n682), .SEL(n4202), .F(n4188) );
  IV U1643 ( .A(n4203), .Z(n682) );
  MUX U1644 ( .IN0(n683), .IN1(n978), .SEL(n979), .F(n947) );
  IV U1645 ( .A(n980), .Z(n683) );
  MUX U1646 ( .IN0(n684), .IN1(n3839), .SEL(n3840), .F(n3773) );
  IV U1647 ( .A(n3841), .Z(n684) );
  MUX U1648 ( .IN0(n685), .IN1(n3792), .SEL(n3793), .F(n3726) );
  IV U1649 ( .A(n3794), .Z(n685) );
  MUX U1650 ( .IN0(n686), .IN1(n3765), .SEL(n3766), .F(n3699) );
  IV U1651 ( .A(n3767), .Z(n686) );
  MUX U1652 ( .IN0(n687), .IN1(n3531), .SEL(n3532), .F(n3467) );
  IV U1653 ( .A(n3533), .Z(n687) );
  MUX U1654 ( .IN0(n688), .IN1(n3508), .SEL(n3509), .F(n3447) );
  IV U1655 ( .A(n3510), .Z(n688) );
  MUX U1656 ( .IN0(n689), .IN1(n3578), .SEL(n3579), .F(n3517) );
  IV U1657 ( .A(n3580), .Z(n689) );
  MUX U1658 ( .IN0(n690), .IN1(n3321), .SEL(n3322), .F(n3274) );
  IV U1659 ( .A(n3323), .Z(n690) );
  MUX U1660 ( .IN0(n691), .IN1(n3296), .SEL(n3297), .F(n3247) );
  IV U1661 ( .A(n3298), .Z(n691) );
  XNOR U1662 ( .A(n5052), .B(n5053), .Z(n4991) );
  XNOR U1663 ( .A(n4774), .B(n4764), .Z(n4768) );
  XNOR U1664 ( .A(n4889), .B(n4890), .Z(n4772) );
  XNOR U1665 ( .A(n2962), .B(n2020), .Z(n2026) );
  XNOR U1666 ( .A(n2500), .B(n2306), .Z(n2312) );
  MUX U1667 ( .IN0(n2325), .IN1(n692), .SEL(n2326), .F(n1407) );
  IV U1668 ( .A(n2327), .Z(n692) );
  MUX U1669 ( .IN0(n693), .IN1(n1400), .SEL(n1401), .F(n1335) );
  IV U1670 ( .A(n1402), .Z(n693) );
  MUX U1671 ( .IN0(n694), .IN1(n1211), .SEL(n1212), .F(n1159) );
  IV U1672 ( .A(n1213), .Z(n694) );
  MUX U1673 ( .IN0(n695), .IN1(n3127), .SEL(n3128), .F(n3097) );
  IV U1674 ( .A(n3129), .Z(n695) );
  MUX U1675 ( .IN0(n696), .IN1(n3119), .SEL(n3120), .F(n3090) );
  IV U1676 ( .A(n3121), .Z(n696) );
  XNOR U1677 ( .A(n5079), .B(n4570), .Z(n4576) );
  XNOR U1678 ( .A(n4993), .B(n4478), .Z(n4482) );
  XNOR U1679 ( .A(n4601), .B(n4168), .Z(n4172) );
  XNOR U1680 ( .A(n4800), .B(n4302), .Z(n4306) );
  XNOR U1681 ( .A(n1431), .B(n1367), .Z(n1371) );
  MUX U1682 ( .IN0(n1419), .IN1(n697), .SEL(n1420), .F(n1352) );
  IV U1683 ( .A(n1421), .Z(n697) );
  MUX U1684 ( .IN0(n2062), .IN1(n698), .SEL(n1465), .F(n1403) );
  IV U1685 ( .A(n1463), .Z(n698) );
  XNOR U1686 ( .A(n1317), .B(n1258), .Z(n1262) );
  XNOR U1687 ( .A(n4275), .B(n4267), .Z(n4146) );
  XNOR U1688 ( .A(n1230), .B(n1180), .Z(n1184) );
  XNOR U1689 ( .A(n4538), .B(n4532), .Z(n4348) );
  XNOR U1690 ( .A(n4440), .B(n4432), .Z(n4346) );
  XNOR U1691 ( .A(n4114), .B(n4100), .Z(n4104) );
  XNOR U1692 ( .A(n4236), .B(n4228), .Z(n4095) );
  XNOR U1693 ( .A(n1088), .B(n1042), .Z(n1046) );
  XNOR U1694 ( .A(n1079), .B(n1033), .Z(n1037) );
  XNOR U1695 ( .A(n4407), .B(n4399), .Z(n4328) );
  XNOR U1696 ( .A(n4063), .B(n4049), .Z(n4053) );
  XNOR U1697 ( .A(n4491), .B(n4487), .Z(n4318) );
  MUX U1698 ( .IN0(n4045), .IN1(n699), .SEL(n3977), .F(n4028) );
  IV U1699 ( .A(n3976), .Z(n699) );
  XNOR U1700 ( .A(n967), .B(n939), .Z(n943) );
  MUX U1701 ( .IN0(n958), .IN1(n700), .SEL(n959), .F(n929) );
  IV U1702 ( .A(n960), .Z(n700) );
  XNOR U1703 ( .A(n4370), .B(n3933), .Z(n3937) );
  XNOR U1704 ( .A(n3953), .B(n3890), .Z(n3894) );
  XNOR U1705 ( .A(n3911), .B(n3850), .Z(n3854) );
  MUX U1706 ( .IN0(n701), .IN1(n926), .SEL(n927), .F(n900) );
  IV U1707 ( .A(n928), .Z(n701) );
  XNOR U1708 ( .A(n3807), .B(n3744), .Z(n3748) );
  MUX U1709 ( .IN0(n3776), .IN1(n702), .SEL(n3777), .F(n3710) );
  IV U1710 ( .A(n3778), .Z(n702) );
  XNOR U1711 ( .A(n3732), .B(n3669), .Z(n3673) );
  XNOR U1712 ( .A(n3689), .B(n3627), .Z(n3631) );
  XNOR U1713 ( .A(n3713), .B(n3652), .Z(n3656) );
  MUX U1714 ( .IN0(n859), .IN1(n703), .SEL(n860), .F(n842) );
  IV U1715 ( .A(n861), .Z(n703) );
  XNOR U1716 ( .A(n3546), .B(n3485), .Z(n3489) );
  XNOR U1717 ( .A(n3537), .B(n3476), .Z(n3480) );
  XNOR U1718 ( .A(n3496), .B(n3440), .Z(n3444) );
  MUX U1719 ( .IN0(n3520), .IN1(n704), .SEL(n3521), .F(n3458) );
  IV U1720 ( .A(n3522), .Z(n704) );
  MUX U1721 ( .IN0(n3461), .IN1(n3523), .SEL(n3463), .F(n3397) );
  XNOR U1722 ( .A(n3311), .B(n3265), .Z(n3271) );
  XNOR U1723 ( .A(n3302), .B(n3256), .Z(n3260) );
  XNOR U1724 ( .A(n3163), .B(n3134), .Z(n3137) );
  XNOR U1725 ( .A(n3139), .B(n3110), .Z(n3116) );
  XOR U1726 ( .A(n4156), .B(n4155), .Z(n4018) );
  XOR U1727 ( .A(n1310), .B(n1309), .Z(n1292) );
  XOR U1728 ( .A(n4359), .B(n4360), .Z(n4009) );
  XOR U1729 ( .A(n4353), .B(n4354), .Z(n4003) );
  XOR U1730 ( .A(n1194), .B(n1193), .Z(n1176) );
  MUX U1731 ( .IN0(n705), .IN1(n1217), .SEL(n1218), .F(n1163) );
  IV U1732 ( .A(n1219), .Z(n705) );
  XOR U1733 ( .A(n4088), .B(n4087), .Z(n3994) );
  XOR U1734 ( .A(n1096), .B(n1095), .Z(n1078) );
  XOR U1735 ( .A(n1105), .B(n1104), .Z(n1111) );
  XOR U1736 ( .A(n4335), .B(n4336), .Z(n3985) );
  XOR U1737 ( .A(n4329), .B(n4330), .Z(n3979) );
  XOR U1738 ( .A(n4323), .B(n4324), .Z(n3973) );
  XOR U1739 ( .A(n3947), .B(n3946), .Z(n3929) );
  XOR U1740 ( .A(n914), .B(n913), .Z(n904) );
  XOR U1741 ( .A(n883), .B(n882), .Z(n874) );
  XOR U1742 ( .A(n3815), .B(n3814), .Z(n3797) );
  MUX U1743 ( .IN0(n3834), .IN1(n706), .SEL(n3835), .F(n3768) );
  IV U1744 ( .A(n3836), .Z(n706) );
  XOR U1745 ( .A(n3683), .B(n3682), .Z(n3665) );
  XOR U1746 ( .A(n3554), .B(n3553), .Z(n3536) );
  MUX U1747 ( .IN0(n3573), .IN1(n707), .SEL(n3574), .F(n3511) );
  IV U1748 ( .A(n3575), .Z(n707) );
  XOR U1749 ( .A(n3386), .B(n3385), .Z(n3405) );
  XOR U1750 ( .A(n3333), .B(n3332), .Z(n3343) );
  XOR U1751 ( .A(n3283), .B(n3282), .Z(n3289) );
  XOR U1752 ( .A(n3227), .B(n3226), .Z(n3208) );
  XOR U1753 ( .A(n3180), .B(n3179), .Z(n3162) );
  XOR U1754 ( .A(n3147), .B(n3146), .Z(n3132) );
  XNOR U1755 ( .A(n3050), .B(n3035), .Z(n3038) );
  XOR U1756 ( .A(n4015), .B(n4016), .Z(n3374) );
  MUX U1757 ( .IN0(n1412), .IN1(\_MAC/_MULT/MULT/S[3][1][0] ), .SEL(n5112), 
        .F(n1345) );
  XOR U1758 ( .A(n1229), .B(n1228), .Z(n1270) );
  XOR U1759 ( .A(n3991), .B(n3992), .Z(n2994) );
  MUX U1760 ( .IN0(n1167), .IN1(\_MAC/_MULT/MULT/S[3][1][4] ), .SEL(n5116), 
        .F(n1115) );
  MUX U1761 ( .IN0(n708), .IN1(n1016), .SEL(n1017), .F(n981) );
  IV U1762 ( .A(n1018), .Z(n708) );
  MUX U1763 ( .IN0(n950), .IN1(\_MAC/_MULT/MULT/S[3][1][9] ), .SEL(n5121), .F(
        n920) );
  MUX U1764 ( .IN0(n850), .IN1(\_MAC/_MULT/MULT/S[3][1][13] ), .SEL(n5125), 
        .F(n836) );
  ANDN U1765 ( .A(n831), .B(n832), .Z(n830) );
  XOR U1766 ( .A(n3413), .B(n3412), .Z(n3393) );
  XOR U1767 ( .A(n3351), .B(n3350), .Z(n3340) );
  XOR U1768 ( .A(n3301), .B(n3300), .Z(n3293) );
  XNOR U1769 ( .A(n3152), .B(n3196), .Z(n3185) );
  ANDN U1770 ( .A(n3064), .B(n3063), .Z(n3045) );
  AND U1771 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[17] ), .B(
        \_MAC/_MULT/MULT/S[3][1][17] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[18] ) );
  AND U1772 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[21] ), .B(
        \_MAC/_MULT/MULT/S[3][1][21] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[22] ) );
  AND U1773 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[25] ), .B(
        \_MAC/_MULT/MULT/S[3][1][25] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[26] ) );
  AND U1774 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[30] ), .B(
        \_MAC/_MULT/MULT/S[3][1][30] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[31] ) );
  MUX U1775 ( .IN0(n2269), .IN1(n709), .SEL(n2270), .F(n2252) );
  IV U1776 ( .A(n2271), .Z(n709) );
  XOR U1777 ( .A(n1986), .B(n1985), .Z(n1999) );
  XOR U1778 ( .A(n2294), .B(n2293), .Z(n2013) );
  MUX U1779 ( .IN0(n1922), .IN1(n710), .SEL(n1923), .F(n1883) );
  IV U1780 ( .A(n1924), .Z(n710) );
  XOR U1781 ( .A(n1945), .B(n1944), .Z(n1958) );
  XOR U1782 ( .A(n2275), .B(n2274), .Z(n1972) );
  XOR U1783 ( .A(n1906), .B(n1905), .Z(n1919) );
  MUX U1784 ( .IN0(n2452), .IN1(n711), .SEL(n2265), .F(n2441) );
  IV U1785 ( .A(n2264), .Z(n711) );
  XOR U1786 ( .A(n2258), .B(n2257), .Z(n1933) );
  XOR U1787 ( .A(n1867), .B(n1866), .Z(n1880) );
  MUX U1788 ( .IN0(n2448), .IN1(n712), .SEL(n2449), .F(n2437) );
  IV U1789 ( .A(n2450), .Z(n712) );
  MUX U1790 ( .IN0(n713), .IN1(n2432), .SEL(n2433), .F(n2421) );
  IV U1791 ( .A(n2434), .Z(n713) );
  MUX U1792 ( .IN0(n1781), .IN1(n714), .SEL(n1782), .F(n1742) );
  IV U1793 ( .A(n1783), .Z(n714) );
  XOR U1794 ( .A(n2241), .B(n2240), .Z(n1894) );
  MUX U1795 ( .IN0(n2201), .IN1(n715), .SEL(n2202), .F(n2184) );
  IV U1796 ( .A(n2203), .Z(n715) );
  MUX U1797 ( .IN0(n716), .IN1(n1795), .SEL(n1796), .F(n1756) );
  IV U1798 ( .A(n1797), .Z(n716) );
  MUX U1799 ( .IN0(n1846), .IN1(n717), .SEL(n1847), .F(n1807) );
  IV U1800 ( .A(n1848), .Z(n717) );
  XOR U1801 ( .A(n1826), .B(n1825), .Z(n1839) );
  XOR U1802 ( .A(n2224), .B(n2223), .Z(n1853) );
  MUX U1803 ( .IN0(n1764), .IN1(n718), .SEL(n1765), .F(n1725) );
  IV U1804 ( .A(n1766), .Z(n718) );
  XOR U1805 ( .A(n1787), .B(n1786), .Z(n1800) );
  XOR U1806 ( .A(n2207), .B(n2206), .Z(n1814) );
  XOR U1807 ( .A(n1748), .B(n1747), .Z(n1761) );
  MUX U1808 ( .IN0(n2408), .IN1(n719), .SEL(n2197), .F(n2397) );
  IV U1809 ( .A(n2196), .Z(n719) );
  XOR U1810 ( .A(n2190), .B(n2189), .Z(n1775) );
  XOR U1811 ( .A(n1709), .B(n1708), .Z(n1722) );
  MUX U1812 ( .IN0(n2613), .IN1(n720), .SEL(n2614), .F(n2592) );
  IV U1813 ( .A(n2615), .Z(n720) );
  MUX U1814 ( .IN0(n2404), .IN1(n721), .SEL(n2405), .F(n2393) );
  IV U1815 ( .A(n2406), .Z(n721) );
  MUX U1816 ( .IN0(n722), .IN1(n2388), .SEL(n2389), .F(n2377) );
  IV U1817 ( .A(n2390), .Z(n722) );
  MUX U1818 ( .IN0(n4714), .IN1(n723), .SEL(n4715), .F(n4693) );
  IV U1819 ( .A(n4716), .Z(n723) );
  MUX U1820 ( .IN0(n1625), .IN1(n724), .SEL(n1626), .F(n1586) );
  IV U1821 ( .A(n1627), .Z(n724) );
  XOR U1822 ( .A(n2173), .B(n2172), .Z(n1736) );
  MUX U1823 ( .IN0(n2133), .IN1(n725), .SEL(n2134), .F(n2116) );
  IV U1824 ( .A(n2135), .Z(n725) );
  MUX U1825 ( .IN0(n726), .IN1(n1639), .SEL(n1640), .F(n1600) );
  IV U1826 ( .A(n1641), .Z(n726) );
  MUX U1827 ( .IN0(n1690), .IN1(n727), .SEL(n1691), .F(n1651) );
  IV U1828 ( .A(n1692), .Z(n727) );
  XOR U1829 ( .A(n1670), .B(n1669), .Z(n1683) );
  XNOR U1830 ( .A(n2754), .B(n2755), .Z(n2629) );
  XNOR U1831 ( .A(n4865), .B(n4857), .Z(n4711) );
  XOR U1832 ( .A(n2156), .B(n2155), .Z(n1697) );
  MUX U1833 ( .IN0(n1608), .IN1(n728), .SEL(n1609), .F(n1569) );
  IV U1834 ( .A(n1610), .Z(n728) );
  XOR U1835 ( .A(n1631), .B(n1630), .Z(n1644) );
  XNOR U1836 ( .A(n2743), .B(n2744), .Z(n2608) );
  XNOR U1837 ( .A(n4717), .B(n4699), .Z(n4703) );
  XOR U1838 ( .A(n2139), .B(n2138), .Z(n1658) );
  XOR U1839 ( .A(n1592), .B(n1591), .Z(n1605) );
  MUX U1840 ( .IN0(n2725), .IN1(n729), .SEL(n2726), .F(n2714) );
  IV U1841 ( .A(n2727), .Z(n729) );
  XNOR U1842 ( .A(n2595), .B(n2577), .Z(n2581) );
  MUX U1843 ( .IN0(n4823), .IN1(n730), .SEL(n4824), .F(n4810) );
  IV U1844 ( .A(n4825), .Z(n730) );
  MUX U1845 ( .IN0(n2364), .IN1(n731), .SEL(n2129), .F(n2353) );
  IV U1846 ( .A(n2128), .Z(n731) );
  XOR U1847 ( .A(n2122), .B(n2121), .Z(n1619) );
  MUX U1848 ( .IN0(n2529), .IN1(n732), .SEL(n2530), .F(n2510) );
  IV U1849 ( .A(n2531), .Z(n732) );
  XNOR U1850 ( .A(n2721), .B(n2722), .Z(n2566) );
  MUX U1851 ( .IN0(n2675), .IN1(n2678), .SEL(n2676), .F(n2662) );
  MUX U1852 ( .IN0(n2788), .IN1(n2810), .SEL(n2790), .F(n2775) );
  MUX U1853 ( .IN0(n2360), .IN1(n733), .SEL(n2361), .F(n2349) );
  IV U1854 ( .A(n2362), .Z(n733) );
  MUX U1855 ( .IN0(n734), .IN1(n2344), .SEL(n2345), .F(n2332) );
  IV U1856 ( .A(n2346), .Z(n734) );
  MUX U1857 ( .IN0(n5087), .IN1(n735), .SEL(n5088), .F(n5083) );
  IV U1858 ( .A(n5089), .Z(n735) );
  MUX U1859 ( .IN0(n5016), .IN1(n5033), .SEL(n5018), .F(n4987) );
  MUX U1860 ( .IN0(n5010), .IN1(n5025), .SEL(n5012), .F(n4997) );
  MUX U1861 ( .IN0(n4630), .IN1(n736), .SEL(n4631), .F(n4611) );
  IV U1862 ( .A(n4632), .Z(n736) );
  XNOR U1863 ( .A(n4826), .B(n4818), .Z(n4648) );
  MUX U1864 ( .IN0(n4776), .IN1(n4779), .SEL(n4777), .F(n4763) );
  MUX U1865 ( .IN0(n4901), .IN1(n4923), .SEL(n4903), .F(n4888) );
  MUX U1866 ( .IN0(n1512), .IN1(n737), .SEL(n1513), .F(n1473) );
  IV U1867 ( .A(n1514), .Z(n737) );
  MUX U1868 ( .IN0(n1469), .IN1(n738), .SEL(n1470), .F(n1433) );
  IV U1869 ( .A(n1471), .Z(n738) );
  XOR U1870 ( .A(n2105), .B(n2104), .Z(n1580) );
  MUX U1871 ( .IN0(n2065), .IN1(n739), .SEL(n2066), .F(n1448) );
  IV U1872 ( .A(n2067), .Z(n739) );
  MUX U1873 ( .IN0(n740), .IN1(n1483), .SEL(n1484), .F(n1416) );
  IV U1874 ( .A(n1485), .Z(n740) );
  MUX U1875 ( .IN0(n1534), .IN1(n741), .SEL(n1535), .F(n1495) );
  IV U1876 ( .A(n1536), .Z(n741) );
  MUX U1877 ( .IN0(n2876), .IN1(n2900), .SEL(n2878), .F(n2037) );
  MUX U1878 ( .IN0(n2964), .IN1(n2967), .SEL(n2965), .F(n2019) );
  MUX U1879 ( .IN0(n2517), .IN1(n742), .SEL(n2518), .F(n2487) );
  IV U1880 ( .A(n2519), .Z(n742) );
  XNOR U1881 ( .A(n2855), .B(n2838), .Z(n2700) );
  XNOR U1882 ( .A(n4654), .B(n4636), .Z(n4640) );
  XNOR U1883 ( .A(n4968), .B(n4951), .Z(n4799) );
  MUX U1884 ( .IN0(n1424), .IN1(n743), .SEL(n1425), .F(n1357) );
  IV U1885 ( .A(n1426), .Z(n743) );
  XOR U1886 ( .A(n2088), .B(n2087), .Z(n1541) );
  XNOR U1887 ( .A(n2945), .B(n2928), .Z(n2881) );
  XNOR U1888 ( .A(n2532), .B(n2503), .Z(n2507) );
  XNOR U1889 ( .A(n2792), .B(n2781), .Z(n2672) );
  MUX U1890 ( .IN0(n744), .IN1(n1375), .SEL(n1376), .F(n1313) );
  IV U1891 ( .A(n1377), .Z(n744) );
  MUX U1892 ( .IN0(n745), .IN1(n4595), .SEL(n4573), .F(n4593) );
  IV U1893 ( .A(n4574), .Z(n745) );
  MUX U1894 ( .IN0(n746), .IN1(n4285), .SEL(n4286), .F(n4272) );
  IV U1895 ( .A(n4287), .Z(n746) );
  MUX U1896 ( .IN0(n747), .IN1(n4448), .SEL(n4449), .F(n4437) );
  IV U1897 ( .A(n4450), .Z(n747) );
  MUX U1898 ( .IN0(n748), .IN1(n1224), .SEL(n1225), .F(n1171) );
  IV U1899 ( .A(n1226), .Z(n748) );
  MUX U1900 ( .IN0(n1127), .IN1(n749), .SEL(n1128), .F(n1081) );
  IV U1901 ( .A(n1129), .Z(n749) );
  MUX U1902 ( .IN0(n750), .IN1(n1147), .SEL(n1148), .F(n1099) );
  IV U1903 ( .A(n1149), .Z(n750) );
  MUX U1904 ( .IN0(n751), .IN1(n4587), .SEL(n4535), .F(n4585) );
  IV U1905 ( .A(n4536), .Z(n751) );
  MUX U1906 ( .IN0(n752), .IN1(n4233), .SEL(n4234), .F(n4220) );
  IV U1907 ( .A(n4235), .Z(n752) );
  MUX U1908 ( .IN0(n753), .IN1(n4404), .SEL(n4405), .F(n4393) );
  IV U1909 ( .A(n4406), .Z(n753) );
  MUX U1910 ( .IN0(n1257), .IN1(n754), .SEL(n1258), .F(n1202) );
  IV U1911 ( .A(n1259), .Z(n754) );
  MUX U1912 ( .IN0(n755), .IN1(n1023), .SEL(n1024), .F(n987) );
  IV U1913 ( .A(n1025), .Z(n755) );
  MUX U1914 ( .IN0(n969), .IN1(n756), .SEL(n970), .F(n938) );
  IV U1915 ( .A(n971), .Z(n756) );
  MUX U1916 ( .IN0(n757), .IN1(n4579), .SEL(n4497), .F(n3949) );
  IV U1917 ( .A(n4498), .Z(n757) );
  MUX U1918 ( .IN0(n4486), .IN1(n758), .SEL(n4487), .F(n3941) );
  IV U1919 ( .A(n4488), .Z(n758) );
  MUX U1920 ( .IN0(n4374), .IN1(n759), .SEL(n4375), .F(n3932) );
  IV U1921 ( .A(n4376), .Z(n759) );
  MUX U1922 ( .IN0(n3955), .IN1(n760), .SEL(n3956), .F(n3889) );
  IV U1923 ( .A(n3957), .Z(n760) );
  MUX U1924 ( .IN0(n761), .IN1(n4025), .SEL(n4026), .F(n3905) );
  IV U1925 ( .A(n4027), .Z(n761) );
  MUX U1926 ( .IN0(n762), .IN1(n3924), .SEL(n3925), .F(n3858) );
  IV U1927 ( .A(n3926), .Z(n762) );
  MUX U1928 ( .IN0(n763), .IN1(n3751), .SEL(n3752), .F(n3685) );
  IV U1929 ( .A(n3753), .Z(n763) );
  MUX U1930 ( .IN0(n764), .IN1(n3707), .SEL(n3708), .F(n3642) );
  IV U1931 ( .A(n3709), .Z(n764) );
  MUX U1932 ( .IN0(n765), .IN1(n3660), .SEL(n3661), .F(n3595) );
  IV U1933 ( .A(n3662), .Z(n765) );
  MUX U1934 ( .IN0(n3626), .IN1(n766), .SEL(n3627), .F(n3562) );
  IV U1935 ( .A(n3628), .Z(n766) );
  MUX U1936 ( .IN0(n767), .IN1(n917), .SEL(n918), .F(n886) );
  IV U1937 ( .A(n919), .Z(n767) );
  MUX U1938 ( .IN0(n3612), .IN1(n768), .SEL(n3613), .F(n3548) );
  IV U1939 ( .A(n3614), .Z(n768) );
  MUX U1940 ( .IN0(n3539), .IN1(n769), .SEL(n3540), .F(n3475) );
  IV U1941 ( .A(n3541), .Z(n769) );
  MUX U1942 ( .IN0(n770), .IN1(n3492), .SEL(n3493), .F(n3433) );
  IV U1943 ( .A(n3494), .Z(n770) );
  MUX U1944 ( .IN0(n771), .IN1(n3408), .SEL(n3409), .F(n3346) );
  IV U1945 ( .A(n3410), .Z(n771) );
  MUX U1946 ( .IN0(n3380), .IN1(n772), .SEL(n3381), .F(n3326) );
  IV U1947 ( .A(n3382), .Z(n772) );
  MUX U1948 ( .IN0(n773), .IN1(n3229), .SEL(n3230), .F(n3182) );
  IV U1949 ( .A(n3231), .Z(n773) );
  MUX U1950 ( .IN0(n774), .IN1(n3203), .SEL(n3204), .F(n3157) );
  IV U1951 ( .A(n3205), .Z(n774) );
  MUX U1952 ( .IN0(n3141), .IN1(n775), .SEL(n3142), .F(n3109) );
  IV U1953 ( .A(n3143), .Z(n775) );
  XNOR U1954 ( .A(n5062), .B(n5047), .Z(n4992) );
  XNOR U1955 ( .A(n4905), .B(n4896), .Z(n4773) );
  XOR U1956 ( .A(n2071), .B(n2070), .Z(n1502) );
  MUX U1957 ( .IN0(n1486), .IN1(n776), .SEL(n1487), .F(n1419) );
  IV U1958 ( .A(n1488), .Z(n776) );
  XNOR U1959 ( .A(n2882), .B(n2046), .Z(n2051) );
  XNOR U1960 ( .A(n2701), .B(n2493), .Z(n2497) );
  XOR U1961 ( .A(n2668), .B(n2667), .Z(n2513) );
  XOR U1962 ( .A(n4769), .B(n4768), .Z(n4614) );
  XNOR U1963 ( .A(n2324), .B(n1407), .Z(n1410) );
  XOR U1964 ( .A(n1454), .B(n1453), .Z(n1463) );
  XOR U1965 ( .A(n2027), .B(n2026), .Z(n2042) );
  XOR U1966 ( .A(n2313), .B(n2312), .Z(n2323) );
  XNOR U1967 ( .A(n4567), .B(n4561), .Z(n4366) );
  XNOR U1968 ( .A(n4475), .B(n4467), .Z(n4364) );
  XNOR U1969 ( .A(n4165), .B(n4151), .Z(n4155) );
  XNOR U1970 ( .A(n4299), .B(n4291), .Z(n4180) );
  XNOR U1971 ( .A(n1364), .B(n1305), .Z(n1309) );
  XNOR U1972 ( .A(n1293), .B(n1233), .Z(n1237) );
  MUX U1973 ( .IN0(n777), .IN1(n1335), .SEL(n1336), .F(n1278) );
  IV U1974 ( .A(n1337), .Z(n777) );
  XNOR U1975 ( .A(n4262), .B(n4254), .Z(n4129) );
  XNOR U1976 ( .A(n4529), .B(n4523), .Z(n4342) );
  XNOR U1977 ( .A(n4429), .B(n4421), .Z(n4340) );
  XNOR U1978 ( .A(n4097), .B(n4083), .Z(n4087) );
  XNOR U1979 ( .A(n1134), .B(n1091), .Z(n1095) );
  XNOR U1980 ( .A(n4223), .B(n4215), .Z(n4078) );
  XNOR U1981 ( .A(n1029), .B(n995), .Z(n1000) );
  XNOR U1982 ( .A(n4184), .B(n3916), .Z(n3920) );
  XNOR U1983 ( .A(n905), .B(n877), .Z(n882) );
  XNOR U1984 ( .A(n3873), .B(n3810), .Z(n3814) );
  XNOR U1985 ( .A(n3864), .B(n3801), .Z(n3805) );
  XNOR U1986 ( .A(n3821), .B(n3758), .Z(n3762) );
  XNOR U1987 ( .A(n3779), .B(n3718), .Z(n3722) );
  XNOR U1988 ( .A(n3584), .B(n3524), .Z(n3527) );
  XNOR U1989 ( .A(n3482), .B(n3426), .Z(n3430) );
  XNOR U1990 ( .A(n3414), .B(n3355), .Z(n3359) );
  MUX U1991 ( .IN0(n778), .IN1(n3455), .SEL(n3456), .F(n3401) );
  IV U1992 ( .A(n3457), .Z(n778) );
  XNOR U1993 ( .A(n3262), .B(n3222), .Z(n3226) );
  XNOR U1994 ( .A(n3253), .B(n3213), .Z(n3217) );
  MUX U1995 ( .IN0(n3281), .IN1(n779), .SEL(n3282), .F(n3233) );
  IV U1996 ( .A(n3283), .Z(n779) );
  XNOR U1997 ( .A(n3079), .B(n3052), .Z(n3057) );
  MUX U1998 ( .IN0(n780), .IN1(n3090), .SEL(n3091), .F(n3060) );
  IV U1999 ( .A(n3092), .Z(n780) );
  XOR U2000 ( .A(n4173), .B(n4172), .Z(n4183) );
  XOR U2001 ( .A(n1389), .B(n1388), .Z(n1405) );
  XOR U2002 ( .A(n1325), .B(n1324), .Z(n1340) );
  XOR U2003 ( .A(n4139), .B(n4138), .Z(n4012) );
  XOR U2004 ( .A(n1247), .B(n1246), .Z(n1229) );
  XOR U2005 ( .A(n1263), .B(n1262), .Z(n1282) );
  XOR U2006 ( .A(n4122), .B(n4121), .Z(n4006) );
  XOR U2007 ( .A(n1209), .B(n1208), .Z(n1219) );
  XOR U2008 ( .A(n4105), .B(n4104), .Z(n4000) );
  XOR U2009 ( .A(n1156), .B(n1155), .Z(n1162) );
  XOR U2010 ( .A(n4071), .B(n4070), .Z(n3988) );
  XOR U2011 ( .A(n1047), .B(n1046), .Z(n1028) );
  XOR U2012 ( .A(n4054), .B(n4053), .Z(n3982) );
  MUX U2013 ( .IN0(n781), .IN1(n1107), .SEL(n1108), .F(n1064) );
  IV U2014 ( .A(n1109), .Z(n781) );
  XOR U2015 ( .A(n1010), .B(n1009), .Z(n992) );
  XOR U2016 ( .A(n4037), .B(n4036), .Z(n3976) );
  XOR U2017 ( .A(n975), .B(n974), .Z(n960) );
  XOR U2018 ( .A(n3961), .B(n3960), .Z(n3970) );
  XOR U2019 ( .A(n3895), .B(n3894), .Z(n3910) );
  XOR U2020 ( .A(n3829), .B(n3828), .Z(n3844) );
  XNOR U2021 ( .A(n872), .B(n900), .Z(n893) );
  XOR U2022 ( .A(n861), .B(n860), .Z(n854) );
  XOR U2023 ( .A(n3697), .B(n3696), .Z(n3712) );
  XOR U2024 ( .A(n3632), .B(n3631), .Z(n3647) );
  XOR U2025 ( .A(n3568), .B(n3567), .Z(n3583) );
  XOR U2026 ( .A(n3506), .B(n3505), .Z(n3522) );
  XOR U2027 ( .A(n3445), .B(n3444), .Z(n3460) );
  XOR U2028 ( .A(n3369), .B(n3368), .Z(n3351) );
  XOR U2029 ( .A(n3319), .B(n3318), .Z(n3301) );
  XOR U2030 ( .A(n3272), .B(n3271), .Z(n3252) );
  MUX U2031 ( .IN0(n782), .IN1(n3237), .SEL(n3238), .F(n3196) );
  IV U2032 ( .A(n3239), .Z(n782) );
  XNOR U2033 ( .A(n3047), .B(n3074), .Z(n3067) );
  XOR U2034 ( .A(n4369), .B(n4368), .Z(n4022) );
  XOR U2035 ( .A(n1354), .B(n1353), .Z(n1396) );
  XOR U2036 ( .A(n4009), .B(n4010), .Z(n3029) );
  MUX U2037 ( .IN0(n1345), .IN1(\_MAC/_MULT/MULT/S[3][1][1] ), .SEL(n5113), 
        .F(n1283) );
  XOR U2038 ( .A(n4003), .B(n4004), .Z(n2998) );
  XOR U2039 ( .A(n1176), .B(n1175), .Z(n1216) );
  XOR U2040 ( .A(n3997), .B(n3998), .Z(n2996) );
  XOR U2041 ( .A(n1124), .B(n1123), .Z(n1166) );
  XOR U2042 ( .A(n3985), .B(n3986), .Z(n2992) );
  MUX U2043 ( .IN0(n1115), .IN1(\_MAC/_MULT/MULT/S[3][1][5] ), .SEL(n5117), 
        .F(n1069) );
  XOR U2044 ( .A(n3979), .B(n3980), .Z(n2990) );
  XOR U2045 ( .A(n3973), .B(n3974), .Z(n2988) );
  XOR U2046 ( .A(n3967), .B(n3968), .Z(n2986) );
  XOR U2047 ( .A(n3929), .B(n3928), .Z(n3902) );
  XOR U2048 ( .A(n904), .B(n903), .Z(n892) );
  XOR U2049 ( .A(n3863), .B(n3862), .Z(n3836) );
  XOR U2050 ( .A(n3731), .B(n3730), .Z(n3704) );
  MUX U2051 ( .IN0(n868), .IN1(\_MAC/_MULT/MULT/S[3][1][12] ), .SEL(n5124), 
        .F(n850) );
  XOR U2052 ( .A(n3665), .B(n3664), .Z(n3639) );
  XOR U2053 ( .A(n3600), .B(n3599), .Z(n3575) );
  XOR U2054 ( .A(n3536), .B(n3535), .Z(n3513) );
  XOR U2055 ( .A(n3472), .B(n3471), .Z(n3452) );
  XOR U2056 ( .A(n3242), .B(n3240), .Z(n3277) );
  XOR U2057 ( .A(n3162), .B(n3161), .Z(n3154) );
  XOR U2058 ( .A(n3132), .B(n3131), .Z(n3122) );
  XOR U2059 ( .A(n3039), .B(n3038), .Z(n3032) );
  XOR U2060 ( .A(n3023), .B(n3022), .Z(n3019) );
  XNOR U2061 ( .A(n922), .B(n950), .Z(n951) );
  XNOR U2062 ( .A(n816), .B(n831), .Z(n834) );
  AND U2063 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[18] ), .B(
        \_MAC/_MULT/MULT/S[3][1][18] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[19] ) );
  AND U2064 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[22] ), .B(
        \_MAC/_MULT/MULT/S[3][1][22] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[23] ) );
  AND U2065 ( .A(\_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[26] ), .B(
        \_MAC/_MULT/MULT/S[3][1][26] ), .Z(
        \_MAC/_MULT/MULT/col[3].row[0]._SHIFT_ADD/_ADD/C[27] ) );
  AND U2066 ( .A(n783), .B(n784), .Z(n5132) );
  XOR U2067 ( .A(\_MAC/_MULT/AX__[5] ), .B(\_MAC/_MULT/AX_[5] ), .Z(n784) );
  AND U2068 ( .A(n783), .B(n785), .Z(n5131) );
  XOR U2069 ( .A(\_MAC/_MULT/AX__[6] ), .B(\_MAC/_MULT/AX_[6] ), .Z(n785) );
  AND U2070 ( .A(n783), .B(n786), .Z(n5159) );
  XOR U2071 ( .A(\_MAC/_MULT/AX__[0] ), .B(\_MAC/_MULT/AX_[0] ), .Z(n786) );
  AND U2072 ( .A(n783), .B(n787), .Z(n5158) );
  XOR U2073 ( .A(\_MAC/_MULT/AX__[10] ), .B(\_MAC/_MULT/AX_[10] ), .Z(n787) );
  AND U2074 ( .A(n783), .B(n788), .Z(n5157) );
  XOR U2075 ( .A(\_MAC/_MULT/AX__[11] ), .B(\_MAC/_MULT/AX_[11] ), .Z(n788) );
  AND U2076 ( .A(n783), .B(n789), .Z(n5156) );
  XOR U2077 ( .A(\_MAC/_MULT/AX__[12] ), .B(\_MAC/_MULT/AX_[12] ), .Z(n789) );
  AND U2078 ( .A(n783), .B(n790), .Z(n5155) );
  XOR U2079 ( .A(\_MAC/_MULT/AX__[13] ), .B(\_MAC/_MULT/AX_[13] ), .Z(n790) );
  AND U2080 ( .A(n783), .B(n791), .Z(n5154) );
  XOR U2081 ( .A(\_MAC/_MULT/AX__[14] ), .B(\_MAC/_MULT/AX_[14] ), .Z(n791) );
  AND U2082 ( .A(n783), .B(n792), .Z(n5153) );
  XOR U2083 ( .A(\_MAC/_MULT/AX__[15] ), .B(\_MAC/_MULT/AX_[15] ), .Z(n792) );
  AND U2084 ( .A(n783), .B(n793), .Z(n5130) );
  XOR U2085 ( .A(\_MAC/_MULT/AX__[7] ), .B(\_MAC/_MULT/AX_[7] ), .Z(n793) );
  AND U2086 ( .A(n783), .B(n794), .Z(n5152) );
  XOR U2087 ( .A(\_MAC/_MULT/AX__[16] ), .B(\_MAC/_MULT/AX_[16] ), .Z(n794) );
  AND U2088 ( .A(n783), .B(n795), .Z(n5151) );
  XOR U2089 ( .A(\_MAC/_MULT/AX__[17] ), .B(\_MAC/_MULT/AX_[17] ), .Z(n795) );
  AND U2090 ( .A(n783), .B(n796), .Z(n5150) );
  XOR U2091 ( .A(\_MAC/_MULT/AX__[18] ), .B(\_MAC/_MULT/AX_[18] ), .Z(n796) );
  AND U2092 ( .A(n783), .B(n797), .Z(n5149) );
  XOR U2093 ( .A(\_MAC/_MULT/AX__[19] ), .B(\_MAC/_MULT/AX_[19] ), .Z(n797) );
  AND U2094 ( .A(n783), .B(n798), .Z(n5148) );
  XOR U2095 ( .A(\_MAC/_MULT/AX__[1] ), .B(\_MAC/_MULT/AX_[1] ), .Z(n798) );
  AND U2096 ( .A(n783), .B(n799), .Z(n5147) );
  XOR U2097 ( .A(\_MAC/_MULT/AX__[20] ), .B(\_MAC/_MULT/AX_[20] ), .Z(n799) );
  AND U2098 ( .A(n783), .B(n800), .Z(n5146) );
  XOR U2099 ( .A(\_MAC/_MULT/AX__[21] ), .B(\_MAC/_MULT/AX_[21] ), .Z(n800) );
  AND U2100 ( .A(n783), .B(n801), .Z(n5145) );
  XOR U2101 ( .A(\_MAC/_MULT/AX__[22] ), .B(\_MAC/_MULT/AX_[22] ), .Z(n801) );
  AND U2102 ( .A(n783), .B(n802), .Z(n5144) );
  XOR U2103 ( .A(\_MAC/_MULT/AX__[23] ), .B(\_MAC/_MULT/AX_[23] ), .Z(n802) );
  AND U2104 ( .A(n783), .B(n803), .Z(n5143) );
  XOR U2105 ( .A(\_MAC/_MULT/AX__[24] ), .B(\_MAC/_MULT/AX_[24] ), .Z(n803) );
  AND U2106 ( .A(n783), .B(n804), .Z(n5129) );
  XOR U2107 ( .A(\_MAC/_MULT/AX__[8] ), .B(\_MAC/_MULT/AX_[8] ), .Z(n804) );
  AND U2108 ( .A(n783), .B(n805), .Z(n5142) );
  XOR U2109 ( .A(\_MAC/_MULT/AX__[25] ), .B(\_MAC/_MULT/AX_[25] ), .Z(n805) );
  AND U2110 ( .A(n783), .B(n806), .Z(n5141) );
  XOR U2111 ( .A(\_MAC/_MULT/AX__[26] ), .B(\_MAC/_MULT/AX_[26] ), .Z(n806) );
  AND U2112 ( .A(n783), .B(n807), .Z(n5140) );
  XOR U2113 ( .A(\_MAC/_MULT/AX__[27] ), .B(\_MAC/_MULT/AX_[27] ), .Z(n807) );
  AND U2114 ( .A(n783), .B(n808), .Z(n5139) );
  XOR U2115 ( .A(\_MAC/_MULT/AX__[28] ), .B(\_MAC/_MULT/AX_[28] ), .Z(n808) );
  AND U2116 ( .A(n783), .B(n809), .Z(n5138) );
  XOR U2117 ( .A(\_MAC/_MULT/AX__[29] ), .B(\_MAC/_MULT/AX_[29] ), .Z(n809) );
  AND U2118 ( .A(n783), .B(n810), .Z(n5137) );
  XOR U2119 ( .A(\_MAC/_MULT/AX__[2] ), .B(\_MAC/_MULT/AX_[2] ), .Z(n810) );
  AND U2120 ( .A(n783), .B(n811), .Z(n5136) );
  XOR U2121 ( .A(\_MAC/_MULT/AX__[30] ), .B(\_MAC/_MULT/AX_[30] ), .Z(n811) );
  AND U2122 ( .A(n783), .B(n812), .Z(n5135) );
  XOR U2123 ( .A(\_MAC/_MULT/AX__[31] ), .B(\_MAC/_MULT/AX_[31] ), .Z(n812) );
  AND U2124 ( .A(n783), .B(n813), .Z(n5134) );
  XOR U2125 ( .A(\_MAC/_MULT/AX__[3] ), .B(\_MAC/_MULT/AX_[3] ), .Z(n813) );
  AND U2126 ( .A(n783), .B(n814), .Z(n5133) );
  XOR U2127 ( .A(\_MAC/_MULT/AX__[4] ), .B(\_MAC/_MULT/AX_[4] ), .Z(n814) );
  AND U2128 ( .A(n783), .B(n815), .Z(n5128) );
  XOR U2129 ( .A(\_MAC/_MULT/AX__[9] ), .B(\_MAC/_MULT/AX_[9] ), .Z(n815) );
  XOR U2130 ( .A(e_input[31]), .B(g_input[31]), .Z(n783) );
  XOR U2131 ( .A(n817), .B(n818), .Z(n5127) );
  XOR U2132 ( .A(n819), .B(n820), .Z(n818) );
  XNOR U2133 ( .A(n821), .B(n822), .Z(n820) );
  AND U2134 ( .A(n823), .B(n824), .Z(n821) );
  NAND U2135 ( .A(n825), .B(n826), .Z(n824) );
  NANDN U2136 ( .B(n827), .A(n828), .Z(n823) );
  XOR U2137 ( .A(n829), .B(n830), .Z(n819) );
  ANDN U2138 ( .A(n833), .B(n822), .Z(n829) );
  XOR U2139 ( .A(n834), .B(n835), .Z(n817) );
  XOR U2140 ( .A(n826), .B(n828), .Z(n835) );
  XNOR U2141 ( .A(n837), .B(n836), .Z(n5126) );
  XNOR U2142 ( .A(n832), .B(n831), .Z(n837) );
  OR U2143 ( .A(n840), .B(n841), .Z(n822) );
  XNOR U2144 ( .A(n826), .B(n825), .Z(n827) );
  NANDN U2145 ( .B(n845), .A(n846), .Z(n825) );
  XNOR U2146 ( .A(n851), .B(n850), .Z(n5125) );
  XNOR U2147 ( .A(n839), .B(n838), .Z(n851) );
  XOR U2148 ( .A(n840), .B(n841), .Z(n839) );
  NANDN U2149 ( .B(n854), .A(n855), .Z(n841) );
  XOR U2150 ( .A(n842), .B(n856), .Z(n843) );
  ANDN U2151 ( .A(n857), .B(n858), .Z(n856) );
  XNOR U2152 ( .A(n848), .B(n849), .Z(n844) );
  NAND U2153 ( .A(n862), .B(n846), .Z(n849) );
  XNOR U2154 ( .A(n847), .B(n863), .Z(n848) );
  ANDN U2155 ( .A(n864), .B(n845), .Z(n863) );
  XNOR U2156 ( .A(n869), .B(n868), .Z(n5124) );
  XOR U2157 ( .A(n853), .B(n852), .Z(n869) );
  XNOR U2158 ( .A(n879), .B(n858), .Z(n875) );
  NANDN U2159 ( .B(n845), .A(n880), .Z(n858) );
  IV U2160 ( .A(n859), .Z(n879) );
  XNOR U2161 ( .A(n866), .B(n867), .Z(n861) );
  NAND U2162 ( .A(n884), .B(n846), .Z(n867) );
  XNOR U2163 ( .A(n865), .B(n885), .Z(n866) );
  AND U2164 ( .A(n864), .B(n862), .Z(n885) );
  XNOR U2165 ( .A(n871), .B(n889), .Z(n5123) );
  XNOR U2166 ( .A(n890), .B(n870), .Z(n871) );
  XNOR U2167 ( .A(n874), .B(n873), .Z(n890) );
  XNOR U2168 ( .A(n893), .B(n894), .Z(n873) );
  XOR U2169 ( .A(n895), .B(n896), .Z(n894) );
  AND U2170 ( .A(n897), .B(n898), .Z(n895) );
  NAND U2171 ( .A(n899), .B(n900), .Z(n898) );
  NANDN U2172 ( .B(n901), .A(n896), .Z(n897) );
  XOR U2173 ( .A(n876), .B(n906), .Z(n877) );
  ANDN U2174 ( .A(n907), .B(n845), .Z(n906) );
  XNOR U2175 ( .A(n911), .B(n878), .Z(n905) );
  NAND U2176 ( .A(n862), .B(n880), .Z(n878) );
  IV U2177 ( .A(n881), .Z(n911) );
  XNOR U2178 ( .A(n887), .B(n888), .Z(n883) );
  NAND U2179 ( .A(n915), .B(n846), .Z(n888) );
  XNOR U2180 ( .A(n886), .B(n916), .Z(n887) );
  AND U2181 ( .A(n864), .B(n884), .Z(n916) );
  XNOR U2182 ( .A(n921), .B(n920), .Z(n5122) );
  XOR U2183 ( .A(n892), .B(n891), .Z(n921) );
  XNOR U2184 ( .A(n924), .B(n901), .Z(n903) );
  XNOR U2185 ( .A(n900), .B(n899), .Z(n901) );
  NANDN U2186 ( .B(n845), .A(n925), .Z(n899) );
  XNOR U2187 ( .A(n896), .B(n902), .Z(n924) );
  XNOR U2188 ( .A(n932), .B(n935), .Z(n934) );
  XOR U2189 ( .A(n908), .B(n937), .Z(n909) );
  AND U2190 ( .A(n907), .B(n862), .Z(n937) );
  XNOR U2191 ( .A(n941), .B(n910), .Z(n936) );
  NAND U2192 ( .A(n884), .B(n880), .Z(n910) );
  IV U2193 ( .A(n912), .Z(n941) );
  XNOR U2194 ( .A(n918), .B(n919), .Z(n914) );
  NAND U2195 ( .A(n945), .B(n846), .Z(n919) );
  XNOR U2196 ( .A(n917), .B(n946), .Z(n918) );
  AND U2197 ( .A(n864), .B(n915), .Z(n946) );
  XOR U2198 ( .A(n951), .B(n923), .Z(n5121) );
  XOR U2199 ( .A(n952), .B(n935), .Z(n930) );
  XNOR U2200 ( .A(n927), .B(n928), .Z(n935) );
  NAND U2201 ( .A(n862), .B(n925), .Z(n928) );
  XNOR U2202 ( .A(n926), .B(n953), .Z(n927) );
  ANDN U2203 ( .A(n954), .B(n845), .Z(n953) );
  XNOR U2204 ( .A(n933), .B(n929), .Z(n952) );
  XOR U2205 ( .A(n932), .B(n961), .Z(n933) );
  ANDN U2206 ( .A(n962), .B(n963), .Z(n961) );
  XOR U2207 ( .A(n938), .B(n968), .Z(n939) );
  AND U2208 ( .A(n907), .B(n884), .Z(n968) );
  XNOR U2209 ( .A(n972), .B(n940), .Z(n967) );
  NAND U2210 ( .A(n915), .B(n880), .Z(n940) );
  IV U2211 ( .A(n942), .Z(n972) );
  XNOR U2212 ( .A(n948), .B(n949), .Z(n944) );
  NAND U2213 ( .A(n976), .B(n846), .Z(n949) );
  XNOR U2214 ( .A(n947), .B(n977), .Z(n948) );
  AND U2215 ( .A(n864), .B(n945), .Z(n977) );
  XOR U2216 ( .A(n984), .B(n982), .Z(n5120) );
  XOR U2217 ( .A(n985), .B(n966), .Z(n959) );
  XNOR U2218 ( .A(n956), .B(n957), .Z(n966) );
  NAND U2219 ( .A(n884), .B(n925), .Z(n957) );
  XNOR U2220 ( .A(n955), .B(n986), .Z(n956) );
  AND U2221 ( .A(n954), .B(n862), .Z(n986) );
  XNOR U2222 ( .A(n965), .B(n958), .Z(n985) );
  XNOR U2223 ( .A(n997), .B(n963), .Z(n993) );
  NANDN U2224 ( .B(n845), .A(n998), .Z(n963) );
  IV U2225 ( .A(n964), .Z(n997) );
  XOR U2226 ( .A(n969), .B(n1003), .Z(n970) );
  AND U2227 ( .A(n907), .B(n915), .Z(n1003) );
  XNOR U2228 ( .A(n1007), .B(n971), .Z(n1002) );
  NAND U2229 ( .A(n945), .B(n880), .Z(n971) );
  IV U2230 ( .A(n973), .Z(n1007) );
  XNOR U2231 ( .A(n979), .B(n980), .Z(n975) );
  NAND U2232 ( .A(n1011), .B(n846), .Z(n980) );
  XNOR U2233 ( .A(n978), .B(n1012), .Z(n979) );
  AND U2234 ( .A(n864), .B(n976), .Z(n1012) );
  XNOR U2235 ( .A(n981), .B(n983), .Z(n984) );
  XNOR U2236 ( .A(n1020), .B(n1018), .Z(n5119) );
  XOR U2237 ( .A(n1021), .B(n1001), .Z(n991) );
  XNOR U2238 ( .A(n988), .B(n989), .Z(n1001) );
  NAND U2239 ( .A(n915), .B(n925), .Z(n989) );
  XNOR U2240 ( .A(n987), .B(n1022), .Z(n988) );
  AND U2241 ( .A(n954), .B(n884), .Z(n1022) );
  XNOR U2242 ( .A(n1000), .B(n990), .Z(n1021) );
  XOR U2243 ( .A(n994), .B(n1030), .Z(n995) );
  ANDN U2244 ( .A(n1031), .B(n845), .Z(n1030) );
  XNOR U2245 ( .A(n1035), .B(n996), .Z(n1029) );
  NAND U2246 ( .A(n862), .B(n998), .Z(n996) );
  IV U2247 ( .A(n999), .Z(n1035) );
  XOR U2248 ( .A(n1004), .B(n1040), .Z(n1005) );
  AND U2249 ( .A(n907), .B(n945), .Z(n1040) );
  XNOR U2250 ( .A(n1044), .B(n1006), .Z(n1039) );
  NAND U2251 ( .A(n976), .B(n880), .Z(n1006) );
  IV U2252 ( .A(n1008), .Z(n1044) );
  XNOR U2253 ( .A(n1014), .B(n1015), .Z(n1010) );
  NAND U2254 ( .A(n1048), .B(n846), .Z(n1015) );
  XNOR U2255 ( .A(n1013), .B(n1049), .Z(n1014) );
  AND U2256 ( .A(n864), .B(n1011), .Z(n1049) );
  XNOR U2257 ( .A(n1017), .B(n1019), .Z(n1020) );
  XNOR U2258 ( .A(n1053), .B(n1054), .Z(n1017) );
  XOR U2259 ( .A(n1055), .B(n1056), .Z(n1054) );
  XOR U2260 ( .A(n1057), .B(n1058), .Z(n1056) );
  NOR U2261 ( .A(n1059), .B(n1060), .Z(n1058) );
  AND U2262 ( .A(n1061), .B(n1062), .Z(n1057) );
  NAND U2263 ( .A(n1063), .B(n1064), .Z(n1062) );
  NANDN U2264 ( .B(n1065), .A(n1055), .Z(n1061) );
  XOR U2265 ( .A(n1070), .B(n1068), .Z(n5118) );
  XOR U2266 ( .A(n1071), .B(n1038), .Z(n1027) );
  XNOR U2267 ( .A(n1024), .B(n1025), .Z(n1038) );
  NAND U2268 ( .A(n945), .B(n925), .Z(n1025) );
  XNOR U2269 ( .A(n1023), .B(n1072), .Z(n1024) );
  AND U2270 ( .A(n954), .B(n915), .Z(n1072) );
  XNOR U2271 ( .A(n1037), .B(n1026), .Z(n1071) );
  XOR U2272 ( .A(n1032), .B(n1080), .Z(n1033) );
  AND U2273 ( .A(n1031), .B(n862), .Z(n1080) );
  XNOR U2274 ( .A(n1084), .B(n1034), .Z(n1079) );
  NAND U2275 ( .A(n884), .B(n998), .Z(n1034) );
  IV U2276 ( .A(n1036), .Z(n1084) );
  XOR U2277 ( .A(n1041), .B(n1089), .Z(n1042) );
  AND U2278 ( .A(n907), .B(n976), .Z(n1089) );
  XNOR U2279 ( .A(n1093), .B(n1043), .Z(n1088) );
  NAND U2280 ( .A(n1011), .B(n880), .Z(n1043) );
  IV U2281 ( .A(n1045), .Z(n1093) );
  XNOR U2282 ( .A(n1051), .B(n1052), .Z(n1047) );
  NAND U2283 ( .A(n1097), .B(n846), .Z(n1052) );
  XNOR U2284 ( .A(n1050), .B(n1098), .Z(n1051) );
  AND U2285 ( .A(n864), .B(n1048), .Z(n1098) );
  XNOR U2286 ( .A(n1067), .B(n1069), .Z(n1070) );
  XOR U2287 ( .A(n1102), .B(n1060), .Z(n1067) );
  XNOR U2288 ( .A(n1065), .B(n1055), .Z(n1060) );
  XNOR U2289 ( .A(n1064), .B(n1063), .Z(n1065) );
  NANDN U2290 ( .B(n845), .A(n1106), .Z(n1063) );
  OR U2291 ( .A(n1110), .B(n1111), .Z(n1059) );
  XOR U2292 ( .A(n1116), .B(n1114), .Z(n5117) );
  XOR U2293 ( .A(n1117), .B(n1087), .Z(n1077) );
  XNOR U2294 ( .A(n1074), .B(n1075), .Z(n1087) );
  NAND U2295 ( .A(n976), .B(n925), .Z(n1075) );
  XNOR U2296 ( .A(n1073), .B(n1118), .Z(n1074) );
  AND U2297 ( .A(n954), .B(n945), .Z(n1118) );
  XNOR U2298 ( .A(n1086), .B(n1076), .Z(n1117) );
  XOR U2299 ( .A(n1081), .B(n1126), .Z(n1082) );
  AND U2300 ( .A(n1031), .B(n884), .Z(n1126) );
  XNOR U2301 ( .A(n1130), .B(n1083), .Z(n1125) );
  NAND U2302 ( .A(n915), .B(n998), .Z(n1083) );
  IV U2303 ( .A(n1085), .Z(n1130) );
  XOR U2304 ( .A(n1090), .B(n1135), .Z(n1091) );
  AND U2305 ( .A(n907), .B(n1011), .Z(n1135) );
  XNOR U2306 ( .A(n1139), .B(n1092), .Z(n1134) );
  NAND U2307 ( .A(n1048), .B(n880), .Z(n1092) );
  IV U2308 ( .A(n1094), .Z(n1139) );
  XOR U2309 ( .A(n1140), .B(n1141), .Z(n1094) );
  AND U2310 ( .A(n1142), .B(n1143), .Z(n1141) );
  XNOR U2311 ( .A(n1140), .B(n1144), .Z(n1142) );
  XNOR U2312 ( .A(n1100), .B(n1101), .Z(n1096) );
  NAND U2313 ( .A(n1145), .B(n846), .Z(n1101) );
  XNOR U2314 ( .A(n1099), .B(n1146), .Z(n1100) );
  AND U2315 ( .A(n864), .B(n1097), .Z(n1146) );
  XNOR U2316 ( .A(n1113), .B(n1115), .Z(n1116) );
  XOR U2317 ( .A(n1150), .B(n1111), .Z(n1113) );
  XOR U2318 ( .A(n1103), .B(n1151), .Z(n1104) );
  ANDN U2319 ( .A(n1152), .B(n1153), .Z(n1151) );
  XNOR U2320 ( .A(n1108), .B(n1109), .Z(n1105) );
  NAND U2321 ( .A(n862), .B(n1106), .Z(n1109) );
  XNOR U2322 ( .A(n1107), .B(n1157), .Z(n1108) );
  ANDN U2323 ( .A(n1158), .B(n845), .Z(n1157) );
  NANDN U2324 ( .B(n1162), .A(n1163), .Z(n1110) );
  XOR U2325 ( .A(n1168), .B(n1166), .Z(n5116) );
  XOR U2326 ( .A(n1169), .B(n1133), .Z(n1123) );
  XNOR U2327 ( .A(n1120), .B(n1121), .Z(n1133) );
  NAND U2328 ( .A(n1011), .B(n925), .Z(n1121) );
  XNOR U2329 ( .A(n1119), .B(n1170), .Z(n1120) );
  AND U2330 ( .A(n954), .B(n976), .Z(n1170) );
  XNOR U2331 ( .A(n1132), .B(n1122), .Z(n1169) );
  XOR U2332 ( .A(n1127), .B(n1178), .Z(n1128) );
  AND U2333 ( .A(n1031), .B(n915), .Z(n1178) );
  XNOR U2334 ( .A(n1182), .B(n1129), .Z(n1177) );
  NAND U2335 ( .A(n945), .B(n998), .Z(n1129) );
  IV U2336 ( .A(n1131), .Z(n1182) );
  XOR U2337 ( .A(n1136), .B(n1187), .Z(n1137) );
  AND U2338 ( .A(n907), .B(n1048), .Z(n1187) );
  XNOR U2339 ( .A(n1191), .B(n1138), .Z(n1186) );
  NAND U2340 ( .A(n1097), .B(n880), .Z(n1138) );
  IV U2341 ( .A(n1140), .Z(n1191) );
  XNOR U2342 ( .A(n1148), .B(n1149), .Z(n1144) );
  NAND U2343 ( .A(n1195), .B(n846), .Z(n1149) );
  XNOR U2344 ( .A(n1147), .B(n1196), .Z(n1148) );
  AND U2345 ( .A(n864), .B(n1145), .Z(n1196) );
  XNOR U2346 ( .A(n1165), .B(n1167), .Z(n1168) );
  XOR U2347 ( .A(n1200), .B(n1162), .Z(n1165) );
  XNOR U2348 ( .A(n1205), .B(n1153), .Z(n1201) );
  NANDN U2349 ( .B(n845), .A(n1206), .Z(n1153) );
  IV U2350 ( .A(n1154), .Z(n1205) );
  XNOR U2351 ( .A(n1160), .B(n1161), .Z(n1156) );
  NAND U2352 ( .A(n884), .B(n1106), .Z(n1161) );
  XNOR U2353 ( .A(n1159), .B(n1210), .Z(n1160) );
  AND U2354 ( .A(n1158), .B(n862), .Z(n1210) );
  XNOR U2355 ( .A(n1163), .B(n1164), .Z(n1200) );
  XNOR U2356 ( .A(n1221), .B(n1216), .Z(n5115) );
  XOR U2357 ( .A(n1222), .B(n1185), .Z(n1175) );
  XNOR U2358 ( .A(n1172), .B(n1173), .Z(n1185) );
  NAND U2359 ( .A(n1048), .B(n925), .Z(n1173) );
  XNOR U2360 ( .A(n1171), .B(n1223), .Z(n1172) );
  AND U2361 ( .A(n954), .B(n1011), .Z(n1223) );
  XNOR U2362 ( .A(n1184), .B(n1174), .Z(n1222) );
  XOR U2363 ( .A(n1179), .B(n1231), .Z(n1180) );
  AND U2364 ( .A(n1031), .B(n945), .Z(n1231) );
  XNOR U2365 ( .A(n1235), .B(n1181), .Z(n1230) );
  NAND U2366 ( .A(n976), .B(n998), .Z(n1181) );
  IV U2367 ( .A(n1183), .Z(n1235) );
  XOR U2368 ( .A(n1188), .B(n1240), .Z(n1189) );
  AND U2369 ( .A(n907), .B(n1097), .Z(n1240) );
  XNOR U2370 ( .A(n1244), .B(n1190), .Z(n1239) );
  NAND U2371 ( .A(n1145), .B(n880), .Z(n1190) );
  IV U2372 ( .A(n1192), .Z(n1244) );
  XNOR U2373 ( .A(n1198), .B(n1199), .Z(n1194) );
  NAND U2374 ( .A(n1248), .B(n846), .Z(n1199) );
  XNOR U2375 ( .A(n1197), .B(n1249), .Z(n1198) );
  AND U2376 ( .A(n864), .B(n1195), .Z(n1249) );
  XNOR U2377 ( .A(n1215), .B(n1220), .Z(n1221) );
  XOR U2378 ( .A(n1253), .B(n1219), .Z(n1215) );
  XOR U2379 ( .A(n1202), .B(n1255), .Z(n1203) );
  ANDN U2380 ( .A(n1256), .B(n845), .Z(n1255) );
  XNOR U2381 ( .A(n1260), .B(n1204), .Z(n1254) );
  NAND U2382 ( .A(n862), .B(n1206), .Z(n1204) );
  IV U2383 ( .A(n1207), .Z(n1260) );
  XNOR U2384 ( .A(n1212), .B(n1213), .Z(n1209) );
  NAND U2385 ( .A(n915), .B(n1106), .Z(n1213) );
  XNOR U2386 ( .A(n1211), .B(n1264), .Z(n1212) );
  AND U2387 ( .A(n1158), .B(n884), .Z(n1264) );
  XNOR U2388 ( .A(n1218), .B(n1214), .Z(n1253) );
  XNOR U2389 ( .A(n1271), .B(n1272), .Z(n1218) );
  XOR U2390 ( .A(n1273), .B(n1274), .Z(n1272) );
  AND U2391 ( .A(n1275), .B(n1276), .Z(n1273) );
  NAND U2392 ( .A(n1277), .B(n1278), .Z(n1276) );
  NANDN U2393 ( .B(n1279), .A(n1274), .Z(n1275) );
  XOR U2394 ( .A(n1284), .B(n1270), .Z(n5114) );
  XOR U2395 ( .A(n1285), .B(n1238), .Z(n1228) );
  XNOR U2396 ( .A(n1225), .B(n1226), .Z(n1238) );
  NAND U2397 ( .A(n1097), .B(n925), .Z(n1226) );
  XNOR U2398 ( .A(n1224), .B(n1286), .Z(n1225) );
  AND U2399 ( .A(n954), .B(n1048), .Z(n1286) );
  XNOR U2400 ( .A(n1237), .B(n1227), .Z(n1285) );
  XOR U2401 ( .A(n1232), .B(n1294), .Z(n1233) );
  AND U2402 ( .A(n1031), .B(n976), .Z(n1294) );
  XNOR U2403 ( .A(n1298), .B(n1234), .Z(n1293) );
  NAND U2404 ( .A(n1011), .B(n998), .Z(n1234) );
  IV U2405 ( .A(n1236), .Z(n1298) );
  XOR U2406 ( .A(n1241), .B(n1303), .Z(n1242) );
  AND U2407 ( .A(n907), .B(n1145), .Z(n1303) );
  XNOR U2408 ( .A(n1307), .B(n1243), .Z(n1302) );
  NAND U2409 ( .A(n1195), .B(n880), .Z(n1243) );
  IV U2410 ( .A(n1245), .Z(n1307) );
  XNOR U2411 ( .A(n1251), .B(n1252), .Z(n1247) );
  NAND U2412 ( .A(n1311), .B(n846), .Z(n1252) );
  XNOR U2413 ( .A(n1250), .B(n1312), .Z(n1251) );
  AND U2414 ( .A(n864), .B(n1248), .Z(n1312) );
  XNOR U2415 ( .A(n1269), .B(n1283), .Z(n1284) );
  XOR U2416 ( .A(n1316), .B(n1282), .Z(n1269) );
  XOR U2417 ( .A(n1257), .B(n1318), .Z(n1258) );
  AND U2418 ( .A(n1256), .B(n862), .Z(n1318) );
  XNOR U2419 ( .A(n1322), .B(n1259), .Z(n1317) );
  NAND U2420 ( .A(n884), .B(n1206), .Z(n1259) );
  IV U2421 ( .A(n1261), .Z(n1322) );
  XNOR U2422 ( .A(n1266), .B(n1267), .Z(n1263) );
  NAND U2423 ( .A(n945), .B(n1106), .Z(n1267) );
  XNOR U2424 ( .A(n1265), .B(n1326), .Z(n1266) );
  AND U2425 ( .A(n1158), .B(n915), .Z(n1326) );
  XOR U2426 ( .A(n1281), .B(n1268), .Z(n1316) );
  XOR U2427 ( .A(n1333), .B(n1279), .Z(n1281) );
  XNOR U2428 ( .A(n1278), .B(n1277), .Z(n1279) );
  NANDN U2429 ( .B(n845), .A(n1334), .Z(n1277) );
  XNOR U2430 ( .A(n1274), .B(n1280), .Z(n1333) );
  XNOR U2431 ( .A(n1341), .B(n1344), .Z(n1343) );
  XOR U2432 ( .A(n1346), .B(n1332), .Z(n5113) );
  XOR U2433 ( .A(n1347), .B(n1301), .Z(n1291) );
  XNOR U2434 ( .A(n1288), .B(n1289), .Z(n1301) );
  NAND U2435 ( .A(n1145), .B(n925), .Z(n1289) );
  XNOR U2436 ( .A(n1287), .B(n1348), .Z(n1288) );
  AND U2437 ( .A(n954), .B(n1097), .Z(n1348) );
  XNOR U2438 ( .A(n1300), .B(n1290), .Z(n1347) );
  XOR U2439 ( .A(n1295), .B(n1356), .Z(n1296) );
  AND U2440 ( .A(n1031), .B(n1011), .Z(n1356) );
  XNOR U2441 ( .A(n1360), .B(n1297), .Z(n1355) );
  NAND U2442 ( .A(n1048), .B(n998), .Z(n1297) );
  IV U2443 ( .A(n1299), .Z(n1360) );
  XOR U2444 ( .A(n1304), .B(n1365), .Z(n1305) );
  AND U2445 ( .A(n907), .B(n1195), .Z(n1365) );
  XNOR U2446 ( .A(n1369), .B(n1306), .Z(n1364) );
  NAND U2447 ( .A(n1248), .B(n880), .Z(n1306) );
  IV U2448 ( .A(n1308), .Z(n1369) );
  XNOR U2449 ( .A(n1314), .B(n1315), .Z(n1310) );
  NAND U2450 ( .A(n1373), .B(n846), .Z(n1315) );
  XNOR U2451 ( .A(n1313), .B(n1374), .Z(n1314) );
  AND U2452 ( .A(n864), .B(n1311), .Z(n1374) );
  XNOR U2453 ( .A(n1331), .B(n1345), .Z(n1346) );
  XOR U2454 ( .A(n1378), .B(n1340), .Z(n1331) );
  XOR U2455 ( .A(n1319), .B(n1380), .Z(n1320) );
  AND U2456 ( .A(n1256), .B(n884), .Z(n1380) );
  XNOR U2457 ( .A(n1384), .B(n1321), .Z(n1379) );
  NAND U2458 ( .A(n915), .B(n1206), .Z(n1321) );
  IV U2459 ( .A(n1323), .Z(n1384) );
  XOR U2460 ( .A(n1385), .B(n1386), .Z(n1323) );
  AND U2461 ( .A(n1387), .B(n1388), .Z(n1386) );
  XNOR U2462 ( .A(n1385), .B(n1389), .Z(n1387) );
  XNOR U2463 ( .A(n1328), .B(n1329), .Z(n1325) );
  NAND U2464 ( .A(n976), .B(n1106), .Z(n1329) );
  XNOR U2465 ( .A(n1327), .B(n1390), .Z(n1328) );
  AND U2466 ( .A(n1158), .B(n945), .Z(n1390) );
  XNOR U2467 ( .A(n1339), .B(n1330), .Z(n1378) );
  XOR U2468 ( .A(n1397), .B(n1344), .Z(n1339) );
  XNOR U2469 ( .A(n1336), .B(n1337), .Z(n1344) );
  NAND U2470 ( .A(n862), .B(n1334), .Z(n1337) );
  XNOR U2471 ( .A(n1335), .B(n1398), .Z(n1336) );
  ANDN U2472 ( .A(n1399), .B(n845), .Z(n1398) );
  XNOR U2473 ( .A(n1342), .B(n1338), .Z(n1397) );
  XOR U2474 ( .A(n1341), .B(n1406), .Z(n1342) );
  ANDN U2475 ( .A(n1407), .B(n1408), .Z(n1406) );
  XOR U2476 ( .A(n1413), .B(n1396), .Z(n5112) );
  XOR U2477 ( .A(n1414), .B(n1363), .Z(n1353) );
  XNOR U2478 ( .A(n1350), .B(n1351), .Z(n1363) );
  NAND U2479 ( .A(n1195), .B(n925), .Z(n1351) );
  XNOR U2480 ( .A(n1349), .B(n1415), .Z(n1350) );
  AND U2481 ( .A(n954), .B(n1145), .Z(n1415) );
  XNOR U2482 ( .A(n1362), .B(n1352), .Z(n1414) );
  XOR U2483 ( .A(n1357), .B(n1423), .Z(n1358) );
  AND U2484 ( .A(n1031), .B(n1048), .Z(n1423) );
  XNOR U2485 ( .A(n1427), .B(n1359), .Z(n1422) );
  NAND U2486 ( .A(n1097), .B(n998), .Z(n1359) );
  IV U2487 ( .A(n1361), .Z(n1427) );
  XOR U2488 ( .A(n1366), .B(n1432), .Z(n1367) );
  AND U2489 ( .A(n907), .B(n1248), .Z(n1432) );
  XNOR U2490 ( .A(n1436), .B(n1368), .Z(n1431) );
  NAND U2491 ( .A(n1311), .B(n880), .Z(n1368) );
  IV U2492 ( .A(n1370), .Z(n1436) );
  XNOR U2493 ( .A(n1376), .B(n1377), .Z(n1372) );
  NAND U2494 ( .A(n1440), .B(n846), .Z(n1377) );
  XNOR U2495 ( .A(n1375), .B(n1441), .Z(n1376) );
  AND U2496 ( .A(n864), .B(n1373), .Z(n1441) );
  XNOR U2497 ( .A(n1395), .B(n1412), .Z(n1413) );
  XOR U2498 ( .A(n1445), .B(n1405), .Z(n1395) );
  XOR U2499 ( .A(n1381), .B(n1447), .Z(n1382) );
  AND U2500 ( .A(n1256), .B(n915), .Z(n1447) );
  XNOR U2501 ( .A(n1451), .B(n1383), .Z(n1446) );
  NAND U2502 ( .A(n945), .B(n1206), .Z(n1383) );
  IV U2503 ( .A(n1385), .Z(n1451) );
  XNOR U2504 ( .A(n1392), .B(n1393), .Z(n1389) );
  NAND U2505 ( .A(n1011), .B(n1106), .Z(n1393) );
  XNOR U2506 ( .A(n1391), .B(n1455), .Z(n1392) );
  AND U2507 ( .A(n1158), .B(n976), .Z(n1455) );
  XNOR U2508 ( .A(n1404), .B(n1394), .Z(n1445) );
  XOR U2509 ( .A(n1459), .B(n1460), .Z(n1394) );
  AND U2510 ( .A(n1461), .B(n1462), .Z(n1460) );
  XNOR U2511 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U2512 ( .A(n1459), .B(n1465), .Z(n1464) );
  XOR U2513 ( .A(n1420), .B(n1466), .Z(n1461) );
  XNOR U2514 ( .A(n1459), .B(n1421), .Z(n1466) );
  XOR U2515 ( .A(n1433), .B(n1468), .Z(n1434) );
  AND U2516 ( .A(n907), .B(n1311), .Z(n1468) );
  XNOR U2517 ( .A(n1472), .B(n1435), .Z(n1467) );
  NAND U2518 ( .A(n1373), .B(n880), .Z(n1435) );
  IV U2519 ( .A(n1437), .Z(n1472) );
  XNOR U2520 ( .A(n1443), .B(n1444), .Z(n1439) );
  NAND U2521 ( .A(n846), .B(n1476), .Z(n1444) );
  XNOR U2522 ( .A(n1442), .B(n1477), .Z(n1443) );
  AND U2523 ( .A(n864), .B(n1440), .Z(n1477) );
  XOR U2524 ( .A(n1481), .B(n1430), .Z(n1420) );
  XNOR U2525 ( .A(n1417), .B(n1418), .Z(n1430) );
  NAND U2526 ( .A(n1248), .B(n925), .Z(n1418) );
  XNOR U2527 ( .A(n1416), .B(n1482), .Z(n1417) );
  AND U2528 ( .A(n954), .B(n1195), .Z(n1482) );
  XNOR U2529 ( .A(n1429), .B(n1419), .Z(n1481) );
  XOR U2530 ( .A(n1424), .B(n1490), .Z(n1425) );
  AND U2531 ( .A(n1031), .B(n1097), .Z(n1490) );
  XNOR U2532 ( .A(n1494), .B(n1426), .Z(n1489) );
  NAND U2533 ( .A(n1145), .B(n998), .Z(n1426) );
  IV U2534 ( .A(n1428), .Z(n1494) );
  XOR U2535 ( .A(n1498), .B(n1499), .Z(n1459) );
  AND U2536 ( .A(n1500), .B(n1501), .Z(n1499) );
  XNOR U2537 ( .A(n1502), .B(n1503), .Z(n1501) );
  XOR U2538 ( .A(n1498), .B(n1504), .Z(n1503) );
  XOR U2539 ( .A(n1487), .B(n1505), .Z(n1500) );
  XNOR U2540 ( .A(n1498), .B(n1488), .Z(n1505) );
  XOR U2541 ( .A(n1469), .B(n1507), .Z(n1470) );
  AND U2542 ( .A(n907), .B(n1373), .Z(n1507) );
  XNOR U2543 ( .A(n1511), .B(n1471), .Z(n1506) );
  NAND U2544 ( .A(n1440), .B(n880), .Z(n1471) );
  IV U2545 ( .A(n1473), .Z(n1511) );
  XNOR U2546 ( .A(n1479), .B(n1480), .Z(n1475) );
  NAND U2547 ( .A(n846), .B(n1515), .Z(n1480) );
  XNOR U2548 ( .A(n1478), .B(n1516), .Z(n1479) );
  AND U2549 ( .A(n1476), .B(n864), .Z(n1516) );
  XOR U2550 ( .A(n1520), .B(n1497), .Z(n1487) );
  XNOR U2551 ( .A(n1484), .B(n1485), .Z(n1497) );
  NAND U2552 ( .A(n1311), .B(n925), .Z(n1485) );
  XNOR U2553 ( .A(n1483), .B(n1521), .Z(n1484) );
  AND U2554 ( .A(n954), .B(n1248), .Z(n1521) );
  XNOR U2555 ( .A(n1496), .B(n1486), .Z(n1520) );
  XOR U2556 ( .A(n1491), .B(n1529), .Z(n1492) );
  AND U2557 ( .A(n1031), .B(n1145), .Z(n1529) );
  XNOR U2558 ( .A(n1533), .B(n1493), .Z(n1528) );
  NAND U2559 ( .A(n1195), .B(n998), .Z(n1493) );
  IV U2560 ( .A(n1495), .Z(n1533) );
  XOR U2561 ( .A(n1537), .B(n1538), .Z(n1498) );
  AND U2562 ( .A(n1539), .B(n1540), .Z(n1538) );
  XNOR U2563 ( .A(n1541), .B(n1542), .Z(n1540) );
  XOR U2564 ( .A(n1537), .B(n1543), .Z(n1542) );
  XOR U2565 ( .A(n1526), .B(n1544), .Z(n1539) );
  XNOR U2566 ( .A(n1537), .B(n1527), .Z(n1544) );
  XOR U2567 ( .A(n1508), .B(n1546), .Z(n1509) );
  AND U2568 ( .A(n907), .B(n1440), .Z(n1546) );
  XNOR U2569 ( .A(n1550), .B(n1510), .Z(n1545) );
  NAND U2570 ( .A(n880), .B(n1476), .Z(n1510) );
  IV U2571 ( .A(n1512), .Z(n1550) );
  XNOR U2572 ( .A(n1518), .B(n1519), .Z(n1514) );
  NAND U2573 ( .A(n846), .B(n1554), .Z(n1519) );
  XNOR U2574 ( .A(n1517), .B(n1555), .Z(n1518) );
  AND U2575 ( .A(n1515), .B(n864), .Z(n1555) );
  XOR U2576 ( .A(n1559), .B(n1536), .Z(n1526) );
  XNOR U2577 ( .A(n1523), .B(n1524), .Z(n1536) );
  NAND U2578 ( .A(n1373), .B(n925), .Z(n1524) );
  XNOR U2579 ( .A(n1522), .B(n1560), .Z(n1523) );
  AND U2580 ( .A(n954), .B(n1311), .Z(n1560) );
  XNOR U2581 ( .A(n1535), .B(n1525), .Z(n1559) );
  XOR U2582 ( .A(n1530), .B(n1568), .Z(n1531) );
  AND U2583 ( .A(n1031), .B(n1195), .Z(n1568) );
  XNOR U2584 ( .A(n1572), .B(n1532), .Z(n1567) );
  NAND U2585 ( .A(n1248), .B(n998), .Z(n1532) );
  IV U2586 ( .A(n1534), .Z(n1572) );
  XOR U2587 ( .A(n1576), .B(n1577), .Z(n1537) );
  AND U2588 ( .A(n1578), .B(n1579), .Z(n1577) );
  XNOR U2589 ( .A(n1580), .B(n1581), .Z(n1579) );
  XOR U2590 ( .A(n1576), .B(n1582), .Z(n1581) );
  XOR U2591 ( .A(n1565), .B(n1583), .Z(n1578) );
  XNOR U2592 ( .A(n1576), .B(n1566), .Z(n1583) );
  XOR U2593 ( .A(n1547), .B(n1585), .Z(n1548) );
  AND U2594 ( .A(n1476), .B(n907), .Z(n1585) );
  XNOR U2595 ( .A(n1589), .B(n1549), .Z(n1584) );
  NAND U2596 ( .A(n880), .B(n1515), .Z(n1549) );
  IV U2597 ( .A(n1551), .Z(n1589) );
  XNOR U2598 ( .A(n1557), .B(n1558), .Z(n1553) );
  NAND U2599 ( .A(n846), .B(n1593), .Z(n1558) );
  XNOR U2600 ( .A(n1556), .B(n1594), .Z(n1557) );
  AND U2601 ( .A(n1554), .B(n864), .Z(n1594) );
  XOR U2602 ( .A(n1598), .B(n1575), .Z(n1565) );
  XNOR U2603 ( .A(n1562), .B(n1563), .Z(n1575) );
  NAND U2604 ( .A(n1440), .B(n925), .Z(n1563) );
  XNOR U2605 ( .A(n1561), .B(n1599), .Z(n1562) );
  AND U2606 ( .A(n954), .B(n1373), .Z(n1599) );
  XNOR U2607 ( .A(n1574), .B(n1564), .Z(n1598) );
  XOR U2608 ( .A(n1569), .B(n1607), .Z(n1570) );
  AND U2609 ( .A(n1031), .B(n1248), .Z(n1607) );
  XNOR U2610 ( .A(n1611), .B(n1571), .Z(n1606) );
  NAND U2611 ( .A(n1311), .B(n998), .Z(n1571) );
  IV U2612 ( .A(n1573), .Z(n1611) );
  XOR U2613 ( .A(n1615), .B(n1616), .Z(n1576) );
  AND U2614 ( .A(n1617), .B(n1618), .Z(n1616) );
  XNOR U2615 ( .A(n1619), .B(n1620), .Z(n1618) );
  XOR U2616 ( .A(n1615), .B(n1621), .Z(n1620) );
  XOR U2617 ( .A(n1604), .B(n1622), .Z(n1617) );
  XNOR U2618 ( .A(n1615), .B(n1605), .Z(n1622) );
  XOR U2619 ( .A(n1586), .B(n1624), .Z(n1587) );
  AND U2620 ( .A(n1515), .B(n907), .Z(n1624) );
  XNOR U2621 ( .A(n1628), .B(n1588), .Z(n1623) );
  NAND U2622 ( .A(n880), .B(n1554), .Z(n1588) );
  IV U2623 ( .A(n1590), .Z(n1628) );
  XNOR U2624 ( .A(n1596), .B(n1597), .Z(n1592) );
  NAND U2625 ( .A(n846), .B(n1632), .Z(n1597) );
  XNOR U2626 ( .A(n1595), .B(n1633), .Z(n1596) );
  AND U2627 ( .A(n1593), .B(n864), .Z(n1633) );
  XOR U2628 ( .A(n1637), .B(n1614), .Z(n1604) );
  XNOR U2629 ( .A(n1601), .B(n1602), .Z(n1614) );
  NAND U2630 ( .A(n925), .B(n1476), .Z(n1602) );
  XNOR U2631 ( .A(n1600), .B(n1638), .Z(n1601) );
  AND U2632 ( .A(n954), .B(n1440), .Z(n1638) );
  XNOR U2633 ( .A(n1613), .B(n1603), .Z(n1637) );
  XOR U2634 ( .A(n1608), .B(n1646), .Z(n1609) );
  AND U2635 ( .A(n1031), .B(n1311), .Z(n1646) );
  XNOR U2636 ( .A(n1650), .B(n1610), .Z(n1645) );
  NAND U2637 ( .A(n1373), .B(n998), .Z(n1610) );
  IV U2638 ( .A(n1612), .Z(n1650) );
  XOR U2639 ( .A(n1654), .B(n1655), .Z(n1615) );
  AND U2640 ( .A(n1656), .B(n1657), .Z(n1655) );
  XNOR U2641 ( .A(n1658), .B(n1659), .Z(n1657) );
  XOR U2642 ( .A(n1654), .B(n1660), .Z(n1659) );
  XOR U2643 ( .A(n1643), .B(n1661), .Z(n1656) );
  XNOR U2644 ( .A(n1654), .B(n1644), .Z(n1661) );
  XOR U2645 ( .A(n1625), .B(n1663), .Z(n1626) );
  AND U2646 ( .A(n1554), .B(n907), .Z(n1663) );
  XNOR U2647 ( .A(n1667), .B(n1627), .Z(n1662) );
  NAND U2648 ( .A(n880), .B(n1593), .Z(n1627) );
  IV U2649 ( .A(n1629), .Z(n1667) );
  XNOR U2650 ( .A(n1635), .B(n1636), .Z(n1631) );
  NAND U2651 ( .A(n846), .B(n1671), .Z(n1636) );
  XNOR U2652 ( .A(n1634), .B(n1672), .Z(n1635) );
  AND U2653 ( .A(n1632), .B(n864), .Z(n1672) );
  XOR U2654 ( .A(n1676), .B(n1653), .Z(n1643) );
  XNOR U2655 ( .A(n1640), .B(n1641), .Z(n1653) );
  NAND U2656 ( .A(n925), .B(n1515), .Z(n1641) );
  XNOR U2657 ( .A(n1639), .B(n1677), .Z(n1640) );
  AND U2658 ( .A(n1476), .B(n954), .Z(n1677) );
  XNOR U2659 ( .A(n1652), .B(n1642), .Z(n1676) );
  XOR U2660 ( .A(n1647), .B(n1685), .Z(n1648) );
  AND U2661 ( .A(n1031), .B(n1373), .Z(n1685) );
  XNOR U2662 ( .A(n1689), .B(n1649), .Z(n1684) );
  NAND U2663 ( .A(n1440), .B(n998), .Z(n1649) );
  IV U2664 ( .A(n1651), .Z(n1689) );
  XOR U2665 ( .A(n1693), .B(n1694), .Z(n1654) );
  AND U2666 ( .A(n1695), .B(n1696), .Z(n1694) );
  XNOR U2667 ( .A(n1697), .B(n1698), .Z(n1696) );
  XOR U2668 ( .A(n1693), .B(n1699), .Z(n1698) );
  XOR U2669 ( .A(n1682), .B(n1700), .Z(n1695) );
  XNOR U2670 ( .A(n1693), .B(n1683), .Z(n1700) );
  XOR U2671 ( .A(n1664), .B(n1702), .Z(n1665) );
  AND U2672 ( .A(n1593), .B(n907), .Z(n1702) );
  XNOR U2673 ( .A(n1706), .B(n1666), .Z(n1701) );
  NAND U2674 ( .A(n880), .B(n1632), .Z(n1666) );
  IV U2675 ( .A(n1668), .Z(n1706) );
  XNOR U2676 ( .A(n1674), .B(n1675), .Z(n1670) );
  NAND U2677 ( .A(n846), .B(n1710), .Z(n1675) );
  XNOR U2678 ( .A(n1673), .B(n1711), .Z(n1674) );
  AND U2679 ( .A(n1671), .B(n864), .Z(n1711) );
  XOR U2680 ( .A(n1715), .B(n1692), .Z(n1682) );
  XNOR U2681 ( .A(n1679), .B(n1680), .Z(n1692) );
  NAND U2682 ( .A(n925), .B(n1554), .Z(n1680) );
  XNOR U2683 ( .A(n1678), .B(n1716), .Z(n1679) );
  AND U2684 ( .A(n1515), .B(n954), .Z(n1716) );
  XNOR U2685 ( .A(n1691), .B(n1681), .Z(n1715) );
  XOR U2686 ( .A(n1686), .B(n1724), .Z(n1687) );
  AND U2687 ( .A(n1031), .B(n1440), .Z(n1724) );
  XNOR U2688 ( .A(n1728), .B(n1688), .Z(n1723) );
  NAND U2689 ( .A(n998), .B(n1476), .Z(n1688) );
  IV U2690 ( .A(n1690), .Z(n1728) );
  XOR U2691 ( .A(n1732), .B(n1733), .Z(n1693) );
  AND U2692 ( .A(n1734), .B(n1735), .Z(n1733) );
  XNOR U2693 ( .A(n1736), .B(n1737), .Z(n1735) );
  XOR U2694 ( .A(n1732), .B(n1738), .Z(n1737) );
  XOR U2695 ( .A(n1721), .B(n1739), .Z(n1734) );
  XNOR U2696 ( .A(n1732), .B(n1722), .Z(n1739) );
  XOR U2697 ( .A(n1703), .B(n1741), .Z(n1704) );
  AND U2698 ( .A(n1632), .B(n907), .Z(n1741) );
  XNOR U2699 ( .A(n1745), .B(n1705), .Z(n1740) );
  NAND U2700 ( .A(n880), .B(n1671), .Z(n1705) );
  IV U2701 ( .A(n1707), .Z(n1745) );
  XNOR U2702 ( .A(n1713), .B(n1714), .Z(n1709) );
  NAND U2703 ( .A(n846), .B(n1749), .Z(n1714) );
  XNOR U2704 ( .A(n1712), .B(n1750), .Z(n1713) );
  AND U2705 ( .A(n1710), .B(n864), .Z(n1750) );
  XOR U2706 ( .A(n1754), .B(n1731), .Z(n1721) );
  XNOR U2707 ( .A(n1718), .B(n1719), .Z(n1731) );
  NAND U2708 ( .A(n925), .B(n1593), .Z(n1719) );
  XNOR U2709 ( .A(n1717), .B(n1755), .Z(n1718) );
  AND U2710 ( .A(n1554), .B(n954), .Z(n1755) );
  XNOR U2711 ( .A(n1730), .B(n1720), .Z(n1754) );
  XOR U2712 ( .A(n1725), .B(n1763), .Z(n1726) );
  AND U2713 ( .A(n1476), .B(n1031), .Z(n1763) );
  XNOR U2714 ( .A(n1767), .B(n1727), .Z(n1762) );
  NAND U2715 ( .A(n998), .B(n1515), .Z(n1727) );
  IV U2716 ( .A(n1729), .Z(n1767) );
  XOR U2717 ( .A(n1771), .B(n1772), .Z(n1732) );
  AND U2718 ( .A(n1773), .B(n1774), .Z(n1772) );
  XNOR U2719 ( .A(n1775), .B(n1776), .Z(n1774) );
  XOR U2720 ( .A(n1771), .B(n1777), .Z(n1776) );
  XOR U2721 ( .A(n1760), .B(n1778), .Z(n1773) );
  XNOR U2722 ( .A(n1771), .B(n1761), .Z(n1778) );
  XOR U2723 ( .A(n1742), .B(n1780), .Z(n1743) );
  AND U2724 ( .A(n1671), .B(n907), .Z(n1780) );
  XNOR U2725 ( .A(n1784), .B(n1744), .Z(n1779) );
  NAND U2726 ( .A(n880), .B(n1710), .Z(n1744) );
  IV U2727 ( .A(n1746), .Z(n1784) );
  XNOR U2728 ( .A(n1752), .B(n1753), .Z(n1748) );
  NAND U2729 ( .A(n846), .B(n1788), .Z(n1753) );
  XNOR U2730 ( .A(n1751), .B(n1789), .Z(n1752) );
  AND U2731 ( .A(n1749), .B(n864), .Z(n1789) );
  XOR U2732 ( .A(n1793), .B(n1770), .Z(n1760) );
  XNOR U2733 ( .A(n1757), .B(n1758), .Z(n1770) );
  NAND U2734 ( .A(n925), .B(n1632), .Z(n1758) );
  XNOR U2735 ( .A(n1756), .B(n1794), .Z(n1757) );
  AND U2736 ( .A(n1593), .B(n954), .Z(n1794) );
  XNOR U2737 ( .A(n1769), .B(n1759), .Z(n1793) );
  XOR U2738 ( .A(n1764), .B(n1802), .Z(n1765) );
  AND U2739 ( .A(n1515), .B(n1031), .Z(n1802) );
  XNOR U2740 ( .A(n1806), .B(n1766), .Z(n1801) );
  NAND U2741 ( .A(n998), .B(n1554), .Z(n1766) );
  IV U2742 ( .A(n1768), .Z(n1806) );
  XOR U2743 ( .A(n1810), .B(n1811), .Z(n1771) );
  AND U2744 ( .A(n1812), .B(n1813), .Z(n1811) );
  XNOR U2745 ( .A(n1814), .B(n1815), .Z(n1813) );
  XOR U2746 ( .A(n1810), .B(n1816), .Z(n1815) );
  XOR U2747 ( .A(n1799), .B(n1817), .Z(n1812) );
  XNOR U2748 ( .A(n1810), .B(n1800), .Z(n1817) );
  XOR U2749 ( .A(n1781), .B(n1819), .Z(n1782) );
  AND U2750 ( .A(n1710), .B(n907), .Z(n1819) );
  XNOR U2751 ( .A(n1823), .B(n1783), .Z(n1818) );
  NAND U2752 ( .A(n880), .B(n1749), .Z(n1783) );
  IV U2753 ( .A(n1785), .Z(n1823) );
  XNOR U2754 ( .A(n1791), .B(n1792), .Z(n1787) );
  NAND U2755 ( .A(n846), .B(n1827), .Z(n1792) );
  XNOR U2756 ( .A(n1790), .B(n1828), .Z(n1791) );
  AND U2757 ( .A(n1788), .B(n864), .Z(n1828) );
  XOR U2758 ( .A(n1832), .B(n1809), .Z(n1799) );
  XNOR U2759 ( .A(n1796), .B(n1797), .Z(n1809) );
  NAND U2760 ( .A(n925), .B(n1671), .Z(n1797) );
  XNOR U2761 ( .A(n1795), .B(n1833), .Z(n1796) );
  AND U2762 ( .A(n1632), .B(n954), .Z(n1833) );
  XNOR U2763 ( .A(n1808), .B(n1798), .Z(n1832) );
  XOR U2764 ( .A(n1803), .B(n1841), .Z(n1804) );
  AND U2765 ( .A(n1554), .B(n1031), .Z(n1841) );
  XNOR U2766 ( .A(n1845), .B(n1805), .Z(n1840) );
  NAND U2767 ( .A(n998), .B(n1593), .Z(n1805) );
  IV U2768 ( .A(n1807), .Z(n1845) );
  XOR U2769 ( .A(n1849), .B(n1850), .Z(n1810) );
  AND U2770 ( .A(n1851), .B(n1852), .Z(n1850) );
  XNOR U2771 ( .A(n1853), .B(n1854), .Z(n1852) );
  XOR U2772 ( .A(n1849), .B(n1855), .Z(n1854) );
  XOR U2773 ( .A(n1838), .B(n1856), .Z(n1851) );
  XNOR U2774 ( .A(n1849), .B(n1839), .Z(n1856) );
  XOR U2775 ( .A(n1820), .B(n1858), .Z(n1821) );
  AND U2776 ( .A(n1749), .B(n907), .Z(n1858) );
  XNOR U2777 ( .A(n1862), .B(n1822), .Z(n1857) );
  NAND U2778 ( .A(n880), .B(n1788), .Z(n1822) );
  IV U2779 ( .A(n1824), .Z(n1862) );
  XOR U2780 ( .A(n1863), .B(n1864), .Z(n1824) );
  AND U2781 ( .A(n1865), .B(n1866), .Z(n1864) );
  XNOR U2782 ( .A(n1863), .B(n1867), .Z(n1865) );
  XNOR U2783 ( .A(n1830), .B(n1831), .Z(n1826) );
  NAND U2784 ( .A(n846), .B(n1868), .Z(n1831) );
  XNOR U2785 ( .A(n1829), .B(n1869), .Z(n1830) );
  AND U2786 ( .A(n1827), .B(n864), .Z(n1869) );
  XOR U2787 ( .A(n1873), .B(n1848), .Z(n1838) );
  XNOR U2788 ( .A(n1835), .B(n1836), .Z(n1848) );
  NAND U2789 ( .A(n925), .B(n1710), .Z(n1836) );
  XNOR U2790 ( .A(n1834), .B(n1874), .Z(n1835) );
  AND U2791 ( .A(n1671), .B(n954), .Z(n1874) );
  XNOR U2792 ( .A(n1847), .B(n1837), .Z(n1873) );
  XOR U2793 ( .A(n1842), .B(n1882), .Z(n1843) );
  AND U2794 ( .A(n1593), .B(n1031), .Z(n1882) );
  XNOR U2795 ( .A(n1886), .B(n1844), .Z(n1881) );
  NAND U2796 ( .A(n998), .B(n1632), .Z(n1844) );
  IV U2797 ( .A(n1846), .Z(n1886) );
  XOR U2798 ( .A(n1890), .B(n1891), .Z(n1849) );
  AND U2799 ( .A(n1892), .B(n1893), .Z(n1891) );
  XNOR U2800 ( .A(n1894), .B(n1895), .Z(n1893) );
  XOR U2801 ( .A(n1890), .B(n1896), .Z(n1895) );
  XOR U2802 ( .A(n1879), .B(n1897), .Z(n1892) );
  XNOR U2803 ( .A(n1890), .B(n1880), .Z(n1897) );
  XOR U2804 ( .A(n1859), .B(n1899), .Z(n1860) );
  AND U2805 ( .A(n1788), .B(n907), .Z(n1899) );
  XNOR U2806 ( .A(n1903), .B(n1861), .Z(n1898) );
  NAND U2807 ( .A(n880), .B(n1827), .Z(n1861) );
  IV U2808 ( .A(n1863), .Z(n1903) );
  XNOR U2809 ( .A(n1871), .B(n1872), .Z(n1867) );
  NAND U2810 ( .A(n846), .B(n1907), .Z(n1872) );
  XNOR U2811 ( .A(n1870), .B(n1908), .Z(n1871) );
  AND U2812 ( .A(n1868), .B(n864), .Z(n1908) );
  XOR U2813 ( .A(n1912), .B(n1889), .Z(n1879) );
  XNOR U2814 ( .A(n1876), .B(n1877), .Z(n1889) );
  NAND U2815 ( .A(n925), .B(n1749), .Z(n1877) );
  XNOR U2816 ( .A(n1875), .B(n1913), .Z(n1876) );
  AND U2817 ( .A(n1710), .B(n954), .Z(n1913) );
  XNOR U2818 ( .A(n1888), .B(n1878), .Z(n1912) );
  XOR U2819 ( .A(n1883), .B(n1921), .Z(n1884) );
  AND U2820 ( .A(n1632), .B(n1031), .Z(n1921) );
  XNOR U2821 ( .A(n1925), .B(n1885), .Z(n1920) );
  NAND U2822 ( .A(n998), .B(n1671), .Z(n1885) );
  IV U2823 ( .A(n1887), .Z(n1925) );
  XOR U2824 ( .A(n1929), .B(n1930), .Z(n1890) );
  AND U2825 ( .A(n1931), .B(n1932), .Z(n1930) );
  XNOR U2826 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U2827 ( .A(n1929), .B(n1935), .Z(n1934) );
  XOR U2828 ( .A(n1918), .B(n1936), .Z(n1931) );
  XNOR U2829 ( .A(n1929), .B(n1919), .Z(n1936) );
  XOR U2830 ( .A(n1900), .B(n1938), .Z(n1901) );
  AND U2831 ( .A(n1827), .B(n907), .Z(n1938) );
  XNOR U2832 ( .A(n1942), .B(n1902), .Z(n1937) );
  NAND U2833 ( .A(n880), .B(n1868), .Z(n1902) );
  IV U2834 ( .A(n1904), .Z(n1942) );
  XNOR U2835 ( .A(n1910), .B(n1911), .Z(n1906) );
  NAND U2836 ( .A(n846), .B(n1946), .Z(n1911) );
  XNOR U2837 ( .A(n1909), .B(n1947), .Z(n1910) );
  AND U2838 ( .A(n1907), .B(n864), .Z(n1947) );
  XOR U2839 ( .A(n1951), .B(n1928), .Z(n1918) );
  XNOR U2840 ( .A(n1915), .B(n1916), .Z(n1928) );
  NAND U2841 ( .A(n925), .B(n1788), .Z(n1916) );
  XNOR U2842 ( .A(n1914), .B(n1952), .Z(n1915) );
  AND U2843 ( .A(n1749), .B(n954), .Z(n1952) );
  XNOR U2844 ( .A(n1927), .B(n1917), .Z(n1951) );
  XOR U2845 ( .A(n1922), .B(n1960), .Z(n1923) );
  AND U2846 ( .A(n1671), .B(n1031), .Z(n1960) );
  XNOR U2847 ( .A(n1964), .B(n1924), .Z(n1959) );
  NAND U2848 ( .A(n998), .B(n1710), .Z(n1924) );
  IV U2849 ( .A(n1926), .Z(n1964) );
  XOR U2850 ( .A(n1968), .B(n1969), .Z(n1929) );
  AND U2851 ( .A(n1970), .B(n1971), .Z(n1969) );
  XNOR U2852 ( .A(n1972), .B(n1973), .Z(n1971) );
  XOR U2853 ( .A(n1968), .B(n1974), .Z(n1973) );
  XOR U2854 ( .A(n1957), .B(n1975), .Z(n1970) );
  XNOR U2855 ( .A(n1968), .B(n1958), .Z(n1975) );
  XOR U2856 ( .A(n1939), .B(n1977), .Z(n1940) );
  AND U2857 ( .A(n1868), .B(n907), .Z(n1977) );
  XOR U2858 ( .A(n1978), .B(n1979), .Z(n1939) );
  AND U2859 ( .A(n1980), .B(n1981), .Z(n1979) );
  XNOR U2860 ( .A(n1982), .B(n1978), .Z(n1980) );
  XNOR U2861 ( .A(n1983), .B(n1941), .Z(n1976) );
  NAND U2862 ( .A(n880), .B(n1907), .Z(n1941) );
  IV U2863 ( .A(n1943), .Z(n1983) );
  XNOR U2864 ( .A(n1949), .B(n1950), .Z(n1945) );
  NAND U2865 ( .A(n846), .B(n1987), .Z(n1950) );
  XNOR U2866 ( .A(n1948), .B(n1988), .Z(n1949) );
  AND U2867 ( .A(n1946), .B(n864), .Z(n1988) );
  XOR U2868 ( .A(n1992), .B(n1967), .Z(n1957) );
  XNOR U2869 ( .A(n1954), .B(n1955), .Z(n1967) );
  NAND U2870 ( .A(n925), .B(n1827), .Z(n1955) );
  XNOR U2871 ( .A(n1953), .B(n1993), .Z(n1954) );
  AND U2872 ( .A(n1788), .B(n954), .Z(n1993) );
  XNOR U2873 ( .A(n1966), .B(n1956), .Z(n1992) );
  XOR U2874 ( .A(n1961), .B(n2001), .Z(n1962) );
  AND U2875 ( .A(n1710), .B(n1031), .Z(n2001) );
  XNOR U2876 ( .A(n2005), .B(n1963), .Z(n2000) );
  NAND U2877 ( .A(n998), .B(n1749), .Z(n1963) );
  IV U2878 ( .A(n1965), .Z(n2005) );
  XOR U2879 ( .A(n2009), .B(n2010), .Z(n1968) );
  AND U2880 ( .A(n2011), .B(n2012), .Z(n2010) );
  XNOR U2881 ( .A(n2013), .B(n2014), .Z(n2012) );
  XOR U2882 ( .A(n2009), .B(n2015), .Z(n2014) );
  XOR U2883 ( .A(n1998), .B(n2016), .Z(n2011) );
  XNOR U2884 ( .A(n2009), .B(n1999), .Z(n2016) );
  XOR U2885 ( .A(n1978), .B(n2018), .Z(n1981) );
  AND U2886 ( .A(n1907), .B(n907), .Z(n2018) );
  XNOR U2887 ( .A(n2022), .B(n1982), .Z(n2017) );
  NAND U2888 ( .A(n880), .B(n1946), .Z(n1982) );
  IV U2889 ( .A(n1984), .Z(n2022) );
  XOR U2890 ( .A(n2023), .B(n2024), .Z(n1984) );
  AND U2891 ( .A(n2025), .B(n2026), .Z(n2024) );
  XNOR U2892 ( .A(n2023), .B(n2027), .Z(n2025) );
  XNOR U2893 ( .A(n1990), .B(n1991), .Z(n1986) );
  NAND U2894 ( .A(n846), .B(n2028), .Z(n1991) );
  XNOR U2895 ( .A(n1989), .B(n2029), .Z(n1990) );
  AND U2896 ( .A(n1987), .B(n864), .Z(n2029) );
  XOR U2897 ( .A(n2030), .B(n2031), .Z(n1989) );
  ANDN U2898 ( .A(n2032), .B(n2033), .Z(n2031) );
  XNOR U2899 ( .A(n2034), .B(n2030), .Z(n2032) );
  XOR U2900 ( .A(n2035), .B(n2008), .Z(n1998) );
  XNOR U2901 ( .A(n1995), .B(n1996), .Z(n2008) );
  NAND U2902 ( .A(n925), .B(n1868), .Z(n1996) );
  XNOR U2903 ( .A(n1994), .B(n2036), .Z(n1995) );
  AND U2904 ( .A(n1827), .B(n954), .Z(n2036) );
  XNOR U2905 ( .A(n2007), .B(n1997), .Z(n2035) );
  XOR U2906 ( .A(n2002), .B(n2044), .Z(n2003) );
  AND U2907 ( .A(n1749), .B(n1031), .Z(n2044) );
  XNOR U2908 ( .A(n2048), .B(n2004), .Z(n2043) );
  NAND U2909 ( .A(n998), .B(n1788), .Z(n2004) );
  IV U2910 ( .A(n2006), .Z(n2048) );
  XOR U2911 ( .A(n2049), .B(n2050), .Z(n2006) );
  AND U2912 ( .A(n2051), .B(n2052), .Z(n2050) );
  XNOR U2913 ( .A(n2049), .B(n2053), .Z(n2052) );
  XOR U2914 ( .A(n2057), .B(n1411), .Z(n1404) );
  XNOR U2915 ( .A(n1401), .B(n1402), .Z(n1411) );
  NAND U2916 ( .A(n884), .B(n1334), .Z(n1402) );
  XNOR U2917 ( .A(n1400), .B(n2058), .Z(n1401) );
  AND U2918 ( .A(n1399), .B(n862), .Z(n2058) );
  XNOR U2919 ( .A(n1410), .B(n1403), .Z(n2057) );
  XOR U2920 ( .A(n1448), .B(n2064), .Z(n1449) );
  AND U2921 ( .A(n1256), .B(n945), .Z(n2064) );
  XNOR U2922 ( .A(n2068), .B(n1450), .Z(n2063) );
  NAND U2923 ( .A(n976), .B(n1206), .Z(n1450) );
  IV U2924 ( .A(n1452), .Z(n2068) );
  XNOR U2925 ( .A(n1457), .B(n1458), .Z(n1454) );
  NAND U2926 ( .A(n1048), .B(n1106), .Z(n1458) );
  XNOR U2927 ( .A(n1456), .B(n2072), .Z(n1457) );
  AND U2928 ( .A(n1158), .B(n1011), .Z(n2072) );
  XOR U2929 ( .A(n2076), .B(n2077), .Z(n1465) );
  XNOR U2930 ( .A(n2078), .B(n2062), .Z(n2076) );
  XOR U2931 ( .A(n2065), .B(n2081), .Z(n2066) );
  AND U2932 ( .A(n1256), .B(n976), .Z(n2081) );
  XNOR U2933 ( .A(n2085), .B(n2067), .Z(n2080) );
  NAND U2934 ( .A(n1011), .B(n1206), .Z(n2067) );
  IV U2935 ( .A(n2069), .Z(n2085) );
  XNOR U2936 ( .A(n2074), .B(n2075), .Z(n2071) );
  NAND U2937 ( .A(n1097), .B(n1106), .Z(n2075) );
  XNOR U2938 ( .A(n2073), .B(n2089), .Z(n2074) );
  AND U2939 ( .A(n1158), .B(n1048), .Z(n2089) );
  XOR U2940 ( .A(n2093), .B(n2094), .Z(n1504) );
  XNOR U2941 ( .A(n2095), .B(n2079), .Z(n2093) );
  XOR U2942 ( .A(n2082), .B(n2098), .Z(n2083) );
  AND U2943 ( .A(n1256), .B(n1011), .Z(n2098) );
  XNOR U2944 ( .A(n2102), .B(n2084), .Z(n2097) );
  NAND U2945 ( .A(n1048), .B(n1206), .Z(n2084) );
  IV U2946 ( .A(n2086), .Z(n2102) );
  XNOR U2947 ( .A(n2091), .B(n2092), .Z(n2088) );
  NAND U2948 ( .A(n1145), .B(n1106), .Z(n2092) );
  XNOR U2949 ( .A(n2090), .B(n2106), .Z(n2091) );
  AND U2950 ( .A(n1158), .B(n1097), .Z(n2106) );
  XOR U2951 ( .A(n2110), .B(n2111), .Z(n1543) );
  XNOR U2952 ( .A(n2112), .B(n2096), .Z(n2110) );
  XOR U2953 ( .A(n2099), .B(n2115), .Z(n2100) );
  AND U2954 ( .A(n1256), .B(n1048), .Z(n2115) );
  XNOR U2955 ( .A(n2119), .B(n2101), .Z(n2114) );
  NAND U2956 ( .A(n1097), .B(n1206), .Z(n2101) );
  IV U2957 ( .A(n2103), .Z(n2119) );
  XNOR U2958 ( .A(n2108), .B(n2109), .Z(n2105) );
  NAND U2959 ( .A(n1195), .B(n1106), .Z(n2109) );
  XNOR U2960 ( .A(n2107), .B(n2123), .Z(n2108) );
  AND U2961 ( .A(n1158), .B(n1145), .Z(n2123) );
  XOR U2962 ( .A(n2127), .B(n2128), .Z(n1582) );
  XNOR U2963 ( .A(n2129), .B(n2113), .Z(n2127) );
  XOR U2964 ( .A(n2116), .B(n2132), .Z(n2117) );
  AND U2965 ( .A(n1256), .B(n1097), .Z(n2132) );
  XNOR U2966 ( .A(n2136), .B(n2118), .Z(n2131) );
  NAND U2967 ( .A(n1145), .B(n1206), .Z(n2118) );
  IV U2968 ( .A(n2120), .Z(n2136) );
  XNOR U2969 ( .A(n2125), .B(n2126), .Z(n2122) );
  NAND U2970 ( .A(n1248), .B(n1106), .Z(n2126) );
  XNOR U2971 ( .A(n2124), .B(n2140), .Z(n2125) );
  AND U2972 ( .A(n1158), .B(n1195), .Z(n2140) );
  XOR U2973 ( .A(n2144), .B(n2145), .Z(n1621) );
  XNOR U2974 ( .A(n2146), .B(n2130), .Z(n2144) );
  XOR U2975 ( .A(n2133), .B(n2149), .Z(n2134) );
  AND U2976 ( .A(n1256), .B(n1145), .Z(n2149) );
  XNOR U2977 ( .A(n2153), .B(n2135), .Z(n2148) );
  NAND U2978 ( .A(n1195), .B(n1206), .Z(n2135) );
  IV U2979 ( .A(n2137), .Z(n2153) );
  XNOR U2980 ( .A(n2142), .B(n2143), .Z(n2139) );
  NAND U2981 ( .A(n1311), .B(n1106), .Z(n2143) );
  XNOR U2982 ( .A(n2141), .B(n2157), .Z(n2142) );
  AND U2983 ( .A(n1158), .B(n1248), .Z(n2157) );
  XOR U2984 ( .A(n2161), .B(n2162), .Z(n1660) );
  XNOR U2985 ( .A(n2163), .B(n2147), .Z(n2161) );
  XOR U2986 ( .A(n2150), .B(n2166), .Z(n2151) );
  AND U2987 ( .A(n1256), .B(n1195), .Z(n2166) );
  XNOR U2988 ( .A(n2170), .B(n2152), .Z(n2165) );
  NAND U2989 ( .A(n1248), .B(n1206), .Z(n2152) );
  IV U2990 ( .A(n2154), .Z(n2170) );
  XNOR U2991 ( .A(n2159), .B(n2160), .Z(n2156) );
  NAND U2992 ( .A(n1373), .B(n1106), .Z(n2160) );
  XNOR U2993 ( .A(n2158), .B(n2174), .Z(n2159) );
  AND U2994 ( .A(n1158), .B(n1311), .Z(n2174) );
  XOR U2995 ( .A(n2178), .B(n2179), .Z(n1699) );
  XNOR U2996 ( .A(n2180), .B(n2164), .Z(n2178) );
  XOR U2997 ( .A(n2167), .B(n2183), .Z(n2168) );
  AND U2998 ( .A(n1256), .B(n1248), .Z(n2183) );
  XNOR U2999 ( .A(n2187), .B(n2169), .Z(n2182) );
  NAND U3000 ( .A(n1311), .B(n1206), .Z(n2169) );
  IV U3001 ( .A(n2171), .Z(n2187) );
  XNOR U3002 ( .A(n2176), .B(n2177), .Z(n2173) );
  NAND U3003 ( .A(n1440), .B(n1106), .Z(n2177) );
  XNOR U3004 ( .A(n2175), .B(n2191), .Z(n2176) );
  AND U3005 ( .A(n1158), .B(n1373), .Z(n2191) );
  XOR U3006 ( .A(n2195), .B(n2196), .Z(n1738) );
  XNOR U3007 ( .A(n2197), .B(n2181), .Z(n2195) );
  XOR U3008 ( .A(n2184), .B(n2200), .Z(n2185) );
  AND U3009 ( .A(n1256), .B(n1311), .Z(n2200) );
  XNOR U3010 ( .A(n2204), .B(n2186), .Z(n2199) );
  NAND U3011 ( .A(n1373), .B(n1206), .Z(n2186) );
  IV U3012 ( .A(n2188), .Z(n2204) );
  XNOR U3013 ( .A(n2193), .B(n2194), .Z(n2190) );
  NAND U3014 ( .A(n1476), .B(n1106), .Z(n2194) );
  XNOR U3015 ( .A(n2192), .B(n2208), .Z(n2193) );
  AND U3016 ( .A(n1158), .B(n1440), .Z(n2208) );
  XOR U3017 ( .A(n2212), .B(n2213), .Z(n1777) );
  XNOR U3018 ( .A(n2214), .B(n2198), .Z(n2212) );
  XOR U3019 ( .A(n2201), .B(n2217), .Z(n2202) );
  AND U3020 ( .A(n1256), .B(n1373), .Z(n2217) );
  XNOR U3021 ( .A(n2221), .B(n2203), .Z(n2216) );
  NAND U3022 ( .A(n1440), .B(n1206), .Z(n2203) );
  IV U3023 ( .A(n2205), .Z(n2221) );
  XNOR U3024 ( .A(n2210), .B(n2211), .Z(n2207) );
  NAND U3025 ( .A(n1515), .B(n1106), .Z(n2211) );
  XNOR U3026 ( .A(n2209), .B(n2225), .Z(n2210) );
  AND U3027 ( .A(n1158), .B(n1476), .Z(n2225) );
  XOR U3028 ( .A(n2229), .B(n2230), .Z(n1816) );
  XNOR U3029 ( .A(n2231), .B(n2215), .Z(n2229) );
  XOR U3030 ( .A(n2218), .B(n2234), .Z(n2219) );
  AND U3031 ( .A(n1256), .B(n1440), .Z(n2234) );
  XNOR U3032 ( .A(n2238), .B(n2220), .Z(n2233) );
  NAND U3033 ( .A(n1476), .B(n1206), .Z(n2220) );
  IV U3034 ( .A(n2222), .Z(n2238) );
  XNOR U3035 ( .A(n2227), .B(n2228), .Z(n2224) );
  NAND U3036 ( .A(n1554), .B(n1106), .Z(n2228) );
  XNOR U3037 ( .A(n2226), .B(n2242), .Z(n2227) );
  AND U3038 ( .A(n1158), .B(n1515), .Z(n2242) );
  XOR U3039 ( .A(n2246), .B(n2247), .Z(n1855) );
  XNOR U3040 ( .A(n2248), .B(n2232), .Z(n2246) );
  XOR U3041 ( .A(n2235), .B(n2251), .Z(n2236) );
  AND U3042 ( .A(n1256), .B(n1476), .Z(n2251) );
  XNOR U3043 ( .A(n2255), .B(n2237), .Z(n2250) );
  NAND U3044 ( .A(n1515), .B(n1206), .Z(n2237) );
  IV U3045 ( .A(n2239), .Z(n2255) );
  XNOR U3046 ( .A(n2244), .B(n2245), .Z(n2241) );
  NAND U3047 ( .A(n1593), .B(n1106), .Z(n2245) );
  XNOR U3048 ( .A(n2243), .B(n2259), .Z(n2244) );
  AND U3049 ( .A(n1158), .B(n1554), .Z(n2259) );
  XOR U3050 ( .A(n2263), .B(n2264), .Z(n1896) );
  XNOR U3051 ( .A(n2265), .B(n2249), .Z(n2263) );
  XOR U3052 ( .A(n2252), .B(n2268), .Z(n2253) );
  AND U3053 ( .A(n1256), .B(n1515), .Z(n2268) );
  XNOR U3054 ( .A(n2272), .B(n2254), .Z(n2267) );
  NAND U3055 ( .A(n1554), .B(n1206), .Z(n2254) );
  IV U3056 ( .A(n2256), .Z(n2272) );
  XNOR U3057 ( .A(n2261), .B(n2262), .Z(n2258) );
  NAND U3058 ( .A(n1632), .B(n1106), .Z(n2262) );
  XNOR U3059 ( .A(n2260), .B(n2276), .Z(n2261) );
  AND U3060 ( .A(n1158), .B(n1593), .Z(n2276) );
  XOR U3061 ( .A(n2280), .B(n2281), .Z(n1935) );
  XNOR U3062 ( .A(n2282), .B(n2266), .Z(n2280) );
  XOR U3063 ( .A(n2269), .B(n2285), .Z(n2270) );
  AND U3064 ( .A(n1256), .B(n1554), .Z(n2285) );
  XNOR U3065 ( .A(n2289), .B(n2271), .Z(n2284) );
  NAND U3066 ( .A(n1593), .B(n1206), .Z(n2271) );
  IV U3067 ( .A(n2273), .Z(n2289) );
  XOR U3068 ( .A(n2290), .B(n2291), .Z(n2273) );
  AND U3069 ( .A(n2292), .B(n2293), .Z(n2291) );
  XNOR U3070 ( .A(n2290), .B(n2294), .Z(n2292) );
  XNOR U3071 ( .A(n2278), .B(n2279), .Z(n2275) );
  NAND U3072 ( .A(n1671), .B(n1106), .Z(n2279) );
  XNOR U3073 ( .A(n2277), .B(n2295), .Z(n2278) );
  AND U3074 ( .A(n1158), .B(n1632), .Z(n2295) );
  XOR U3075 ( .A(n2299), .B(n2300), .Z(n1974) );
  XNOR U3076 ( .A(n2301), .B(n2283), .Z(n2299) );
  XOR U3077 ( .A(n2286), .B(n2304), .Z(n2287) );
  AND U3078 ( .A(n1256), .B(n1593), .Z(n2304) );
  XNOR U3079 ( .A(n2308), .B(n2288), .Z(n2303) );
  NAND U3080 ( .A(n1632), .B(n1206), .Z(n2288) );
  IV U3081 ( .A(n2290), .Z(n2308) );
  XOR U3082 ( .A(n2309), .B(n2310), .Z(n2290) );
  AND U3083 ( .A(n2311), .B(n2312), .Z(n2310) );
  XNOR U3084 ( .A(n2309), .B(n2313), .Z(n2311) );
  XNOR U3085 ( .A(n2297), .B(n2298), .Z(n2294) );
  NAND U3086 ( .A(n1710), .B(n1106), .Z(n2298) );
  XNOR U3087 ( .A(n2296), .B(n2314), .Z(n2297) );
  AND U3088 ( .A(n1158), .B(n1671), .Z(n2314) );
  XOR U3089 ( .A(n2318), .B(n2319), .Z(n2015) );
  XNOR U3090 ( .A(n2320), .B(n2302), .Z(n2318) );
  XNOR U3091 ( .A(n2328), .B(n1408), .Z(n2324) );
  OR U3092 ( .A(n845), .B(n2329), .Z(n1408) );
  IV U3093 ( .A(n1409), .Z(n2328) );
  XNOR U3094 ( .A(n2060), .B(n2061), .Z(n2077) );
  NAND U3095 ( .A(n915), .B(n1334), .Z(n2061) );
  XNOR U3096 ( .A(n2059), .B(n2331), .Z(n2060) );
  AND U3097 ( .A(n1399), .B(n884), .Z(n2331) );
  XOR U3098 ( .A(n2325), .B(n2336), .Z(n2326) );
  NOR U3099 ( .A(n845), .B(n2337), .Z(n2336) );
  XNOR U3100 ( .A(n2341), .B(n2327), .Z(n2335) );
  NANDN U3101 ( .B(n2329), .A(n862), .Z(n2327) );
  IV U3102 ( .A(n2330), .Z(n2341) );
  XNOR U3103 ( .A(n2333), .B(n2334), .Z(n2094) );
  NAND U3104 ( .A(n945), .B(n1334), .Z(n2334) );
  XNOR U3105 ( .A(n2332), .B(n2343), .Z(n2333) );
  AND U3106 ( .A(n1399), .B(n915), .Z(n2343) );
  XOR U3107 ( .A(n2338), .B(n2348), .Z(n2339) );
  ANDN U3108 ( .A(n862), .B(n2337), .Z(n2348) );
  XNOR U3109 ( .A(n2352), .B(n2340), .Z(n2347) );
  NANDN U3110 ( .B(n2329), .A(n884), .Z(n2340) );
  IV U3111 ( .A(n2342), .Z(n2352) );
  XNOR U3112 ( .A(n2345), .B(n2346), .Z(n2111) );
  NAND U3113 ( .A(n976), .B(n1334), .Z(n2346) );
  XNOR U3114 ( .A(n2344), .B(n2354), .Z(n2345) );
  AND U3115 ( .A(n1399), .B(n945), .Z(n2354) );
  XOR U3116 ( .A(n2349), .B(n2359), .Z(n2350) );
  ANDN U3117 ( .A(n884), .B(n2337), .Z(n2359) );
  XNOR U3118 ( .A(n2363), .B(n2351), .Z(n2358) );
  NANDN U3119 ( .B(n2329), .A(n915), .Z(n2351) );
  IV U3120 ( .A(n2353), .Z(n2363) );
  XNOR U3121 ( .A(n2356), .B(n2357), .Z(n2128) );
  NAND U3122 ( .A(n1011), .B(n1334), .Z(n2357) );
  XNOR U3123 ( .A(n2355), .B(n2365), .Z(n2356) );
  AND U3124 ( .A(n1399), .B(n976), .Z(n2365) );
  XOR U3125 ( .A(n2360), .B(n2370), .Z(n2361) );
  ANDN U3126 ( .A(n915), .B(n2337), .Z(n2370) );
  XNOR U3127 ( .A(n2374), .B(n2362), .Z(n2369) );
  NANDN U3128 ( .B(n2329), .A(n945), .Z(n2362) );
  IV U3129 ( .A(n2364), .Z(n2374) );
  XNOR U3130 ( .A(n2367), .B(n2368), .Z(n2145) );
  NAND U3131 ( .A(n1048), .B(n1334), .Z(n2368) );
  XNOR U3132 ( .A(n2366), .B(n2376), .Z(n2367) );
  AND U3133 ( .A(n1399), .B(n1011), .Z(n2376) );
  XOR U3134 ( .A(n2371), .B(n2381), .Z(n2372) );
  ANDN U3135 ( .A(n945), .B(n2337), .Z(n2381) );
  XNOR U3136 ( .A(n2385), .B(n2373), .Z(n2380) );
  NANDN U3137 ( .B(n2329), .A(n976), .Z(n2373) );
  IV U3138 ( .A(n2375), .Z(n2385) );
  XNOR U3139 ( .A(n2378), .B(n2379), .Z(n2162) );
  NAND U3140 ( .A(n1097), .B(n1334), .Z(n2379) );
  XNOR U3141 ( .A(n2377), .B(n2387), .Z(n2378) );
  AND U3142 ( .A(n1399), .B(n1048), .Z(n2387) );
  XOR U3143 ( .A(n2382), .B(n2392), .Z(n2383) );
  ANDN U3144 ( .A(n976), .B(n2337), .Z(n2392) );
  XNOR U3145 ( .A(n2396), .B(n2384), .Z(n2391) );
  NANDN U3146 ( .B(n2329), .A(n1011), .Z(n2384) );
  IV U3147 ( .A(n2386), .Z(n2396) );
  XNOR U3148 ( .A(n2389), .B(n2390), .Z(n2179) );
  NAND U3149 ( .A(n1145), .B(n1334), .Z(n2390) );
  XNOR U3150 ( .A(n2388), .B(n2398), .Z(n2389) );
  AND U3151 ( .A(n1399), .B(n1097), .Z(n2398) );
  XOR U3152 ( .A(n2393), .B(n2403), .Z(n2394) );
  ANDN U3153 ( .A(n1011), .B(n2337), .Z(n2403) );
  XNOR U3154 ( .A(n2407), .B(n2395), .Z(n2402) );
  NANDN U3155 ( .B(n2329), .A(n1048), .Z(n2395) );
  IV U3156 ( .A(n2397), .Z(n2407) );
  XNOR U3157 ( .A(n2400), .B(n2401), .Z(n2196) );
  NAND U3158 ( .A(n1195), .B(n1334), .Z(n2401) );
  XNOR U3159 ( .A(n2399), .B(n2409), .Z(n2400) );
  AND U3160 ( .A(n1399), .B(n1145), .Z(n2409) );
  XOR U3161 ( .A(n2404), .B(n2414), .Z(n2405) );
  ANDN U3162 ( .A(n1048), .B(n2337), .Z(n2414) );
  XNOR U3163 ( .A(n2418), .B(n2406), .Z(n2413) );
  NANDN U3164 ( .B(n2329), .A(n1097), .Z(n2406) );
  IV U3165 ( .A(n2408), .Z(n2418) );
  XNOR U3166 ( .A(n2411), .B(n2412), .Z(n2213) );
  NAND U3167 ( .A(n1248), .B(n1334), .Z(n2412) );
  XNOR U3168 ( .A(n2410), .B(n2420), .Z(n2411) );
  AND U3169 ( .A(n1399), .B(n1195), .Z(n2420) );
  XOR U3170 ( .A(n2415), .B(n2425), .Z(n2416) );
  ANDN U3171 ( .A(n1097), .B(n2337), .Z(n2425) );
  XNOR U3172 ( .A(n2429), .B(n2417), .Z(n2424) );
  NANDN U3173 ( .B(n2329), .A(n1145), .Z(n2417) );
  IV U3174 ( .A(n2419), .Z(n2429) );
  XNOR U3175 ( .A(n2422), .B(n2423), .Z(n2230) );
  NAND U3176 ( .A(n1311), .B(n1334), .Z(n2423) );
  XNOR U3177 ( .A(n2421), .B(n2431), .Z(n2422) );
  AND U3178 ( .A(n1399), .B(n1248), .Z(n2431) );
  XOR U3179 ( .A(n2426), .B(n2436), .Z(n2427) );
  ANDN U3180 ( .A(n1145), .B(n2337), .Z(n2436) );
  XNOR U3181 ( .A(n2440), .B(n2428), .Z(n2435) );
  NANDN U3182 ( .B(n2329), .A(n1195), .Z(n2428) );
  IV U3183 ( .A(n2430), .Z(n2440) );
  XNOR U3184 ( .A(n2433), .B(n2434), .Z(n2247) );
  NAND U3185 ( .A(n1373), .B(n1334), .Z(n2434) );
  XNOR U3186 ( .A(n2432), .B(n2442), .Z(n2433) );
  AND U3187 ( .A(n1399), .B(n1311), .Z(n2442) );
  XOR U3188 ( .A(n2437), .B(n2447), .Z(n2438) );
  ANDN U3189 ( .A(n1195), .B(n2337), .Z(n2447) );
  XNOR U3190 ( .A(n2451), .B(n2439), .Z(n2446) );
  NANDN U3191 ( .B(n2329), .A(n1248), .Z(n2439) );
  IV U3192 ( .A(n2441), .Z(n2451) );
  XNOR U3193 ( .A(n2444), .B(n2445), .Z(n2264) );
  NAND U3194 ( .A(n1440), .B(n1334), .Z(n2445) );
  XNOR U3195 ( .A(n2443), .B(n2453), .Z(n2444) );
  AND U3196 ( .A(n1399), .B(n1373), .Z(n2453) );
  XOR U3197 ( .A(n2448), .B(n2458), .Z(n2449) );
  ANDN U3198 ( .A(n1248), .B(n2337), .Z(n2458) );
  XNOR U3199 ( .A(n2462), .B(n2450), .Z(n2457) );
  NANDN U3200 ( .B(n2329), .A(n1311), .Z(n2450) );
  IV U3201 ( .A(n2452), .Z(n2462) );
  XNOR U3202 ( .A(n2455), .B(n2456), .Z(n2281) );
  NAND U3203 ( .A(n1476), .B(n1334), .Z(n2456) );
  XNOR U3204 ( .A(n2454), .B(n2464), .Z(n2455) );
  AND U3205 ( .A(n1399), .B(n1440), .Z(n2464) );
  XOR U3206 ( .A(n2459), .B(n2469), .Z(n2460) );
  ANDN U3207 ( .A(n1311), .B(n2337), .Z(n2469) );
  XNOR U3208 ( .A(n2473), .B(n2461), .Z(n2468) );
  NANDN U3209 ( .B(n2329), .A(n1373), .Z(n2461) );
  IV U3210 ( .A(n2463), .Z(n2473) );
  XNOR U3211 ( .A(n2466), .B(n2467), .Z(n2300) );
  NAND U3212 ( .A(n1515), .B(n1334), .Z(n2467) );
  XNOR U3213 ( .A(n2465), .B(n2475), .Z(n2466) );
  AND U3214 ( .A(n1399), .B(n1476), .Z(n2475) );
  XOR U3215 ( .A(n2470), .B(n2480), .Z(n2471) );
  ANDN U3216 ( .A(n1373), .B(n2337), .Z(n2480) );
  XNOR U3217 ( .A(n2484), .B(n2472), .Z(n2479) );
  NANDN U3218 ( .B(n2329), .A(n1440), .Z(n2472) );
  IV U3219 ( .A(n2474), .Z(n2484) );
  XNOR U3220 ( .A(n2477), .B(n2478), .Z(n2319) );
  NAND U3221 ( .A(n1554), .B(n1334), .Z(n2478) );
  XNOR U3222 ( .A(n2476), .B(n2486), .Z(n2477) );
  AND U3223 ( .A(n1399), .B(n1515), .Z(n2486) );
  XOR U3224 ( .A(n2481), .B(n2491), .Z(n2482) );
  ANDN U3225 ( .A(n1440), .B(n2337), .Z(n2491) );
  XNOR U3226 ( .A(n2495), .B(n2483), .Z(n2490) );
  NANDN U3227 ( .B(n2329), .A(n1476), .Z(n2483) );
  IV U3228 ( .A(n2485), .Z(n2495) );
  XNOR U3229 ( .A(n2056), .B(n2055), .Z(n1412) );
  XOR U3230 ( .A(n2499), .B(n2323), .Z(n2055) );
  XOR U3231 ( .A(n2305), .B(n2501), .Z(n2306) );
  AND U3232 ( .A(n1256), .B(n1632), .Z(n2501) );
  XNOR U3233 ( .A(n2505), .B(n2307), .Z(n2500) );
  NAND U3234 ( .A(n1671), .B(n1206), .Z(n2307) );
  IV U3235 ( .A(n2309), .Z(n2505) );
  XNOR U3236 ( .A(n2316), .B(n2317), .Z(n2313) );
  NAND U3237 ( .A(n1749), .B(n1106), .Z(n2317) );
  XNOR U3238 ( .A(n2315), .B(n2509), .Z(n2316) );
  AND U3239 ( .A(n1158), .B(n1710), .Z(n2509) );
  XNOR U3240 ( .A(n2322), .B(n2054), .Z(n2499) );
  XOR U3241 ( .A(n2513), .B(n2514), .Z(n2054) );
  XOR U3242 ( .A(n2515), .B(n2498), .Z(n2322) );
  XNOR U3243 ( .A(n2488), .B(n2489), .Z(n2498) );
  NAND U3244 ( .A(n1593), .B(n1334), .Z(n2489) );
  XNOR U3245 ( .A(n2487), .B(n2516), .Z(n2488) );
  AND U3246 ( .A(n1399), .B(n1554), .Z(n2516) );
  XNOR U3247 ( .A(n2497), .B(n2321), .Z(n2515) );
  XOR U3248 ( .A(n2520), .B(n2521), .Z(n2321) );
  AND U3249 ( .A(n2522), .B(n2523), .Z(n2521) );
  XOR U3250 ( .A(n2524), .B(n2525), .Z(n2523) );
  XOR U3251 ( .A(n2520), .B(n2526), .Z(n2525) );
  XOR U3252 ( .A(n2507), .B(n2527), .Z(n2522) );
  XOR U3253 ( .A(n2520), .B(n2508), .Z(n2527) );
  NAND U3254 ( .A(n1106), .B(n1788), .Z(n2512) );
  XOR U3255 ( .A(n2510), .B(n2528), .Z(n2511) );
  AND U3256 ( .A(n1158), .B(n1749), .Z(n2528) );
  XOR U3257 ( .A(n2502), .B(n2533), .Z(n2503) );
  AND U3258 ( .A(n1256), .B(n1671), .Z(n2533) );
  XNOR U3259 ( .A(n2537), .B(n2504), .Z(n2532) );
  NAND U3260 ( .A(n1710), .B(n1206), .Z(n2504) );
  IV U3261 ( .A(n2506), .Z(n2537) );
  XOR U3262 ( .A(n2541), .B(n2542), .Z(n2520) );
  AND U3263 ( .A(n2543), .B(n2544), .Z(n2542) );
  XOR U3264 ( .A(n2545), .B(n2546), .Z(n2544) );
  XOR U3265 ( .A(n2541), .B(n2547), .Z(n2546) );
  XOR U3266 ( .A(n2539), .B(n2548), .Z(n2543) );
  XOR U3267 ( .A(n2541), .B(n2540), .Z(n2548) );
  NAND U3268 ( .A(n1106), .B(n1827), .Z(n2531) );
  XOR U3269 ( .A(n2529), .B(n2549), .Z(n2530) );
  AND U3270 ( .A(n1788), .B(n1158), .Z(n2549) );
  XOR U3271 ( .A(n2534), .B(n2554), .Z(n2535) );
  AND U3272 ( .A(n1256), .B(n1710), .Z(n2554) );
  XNOR U3273 ( .A(n2558), .B(n2536), .Z(n2553) );
  NAND U3274 ( .A(n1749), .B(n1206), .Z(n2536) );
  IV U3275 ( .A(n2538), .Z(n2558) );
  XOR U3276 ( .A(n2562), .B(n2563), .Z(n2541) );
  AND U3277 ( .A(n2564), .B(n2565), .Z(n2563) );
  XOR U3278 ( .A(n2566), .B(n2567), .Z(n2565) );
  XOR U3279 ( .A(n2562), .B(n2568), .Z(n2567) );
  XOR U3280 ( .A(n2560), .B(n2569), .Z(n2564) );
  XOR U3281 ( .A(n2562), .B(n2561), .Z(n2569) );
  NAND U3282 ( .A(n1106), .B(n1868), .Z(n2552) );
  XOR U3283 ( .A(n2550), .B(n2570), .Z(n2551) );
  AND U3284 ( .A(n1827), .B(n1158), .Z(n2570) );
  XOR U3285 ( .A(n2555), .B(n2575), .Z(n2556) );
  AND U3286 ( .A(n1256), .B(n1749), .Z(n2575) );
  XNOR U3287 ( .A(n2579), .B(n2557), .Z(n2574) );
  NAND U3288 ( .A(n1206), .B(n1788), .Z(n2557) );
  IV U3289 ( .A(n2559), .Z(n2579) );
  XOR U3290 ( .A(n2583), .B(n2584), .Z(n2562) );
  AND U3291 ( .A(n2585), .B(n2586), .Z(n2584) );
  XOR U3292 ( .A(n2587), .B(n2588), .Z(n2586) );
  XOR U3293 ( .A(n2583), .B(n2589), .Z(n2588) );
  XOR U3294 ( .A(n2581), .B(n2590), .Z(n2585) );
  XOR U3295 ( .A(n2583), .B(n2582), .Z(n2590) );
  NAND U3296 ( .A(n1106), .B(n1907), .Z(n2573) );
  XOR U3297 ( .A(n2571), .B(n2591), .Z(n2572) );
  AND U3298 ( .A(n1868), .B(n1158), .Z(n2591) );
  XOR U3299 ( .A(n2576), .B(n2596), .Z(n2577) );
  AND U3300 ( .A(n1788), .B(n1256), .Z(n2596) );
  XNOR U3301 ( .A(n2600), .B(n2578), .Z(n2595) );
  NAND U3302 ( .A(n1206), .B(n1827), .Z(n2578) );
  IV U3303 ( .A(n2580), .Z(n2600) );
  XOR U3304 ( .A(n2604), .B(n2605), .Z(n2583) );
  AND U3305 ( .A(n2606), .B(n2607), .Z(n2605) );
  XOR U3306 ( .A(n2608), .B(n2609), .Z(n2607) );
  XOR U3307 ( .A(n2604), .B(n2610), .Z(n2609) );
  XOR U3308 ( .A(n2602), .B(n2611), .Z(n2606) );
  XOR U3309 ( .A(n2604), .B(n2603), .Z(n2611) );
  NAND U3310 ( .A(n1106), .B(n1946), .Z(n2594) );
  XOR U3311 ( .A(n2592), .B(n2612), .Z(n2593) );
  AND U3312 ( .A(n1907), .B(n1158), .Z(n2612) );
  XOR U3313 ( .A(n2597), .B(n2617), .Z(n2598) );
  AND U3314 ( .A(n1827), .B(n1256), .Z(n2617) );
  XNOR U3315 ( .A(n2621), .B(n2599), .Z(n2616) );
  NAND U3316 ( .A(n1206), .B(n1868), .Z(n2599) );
  IV U3317 ( .A(n2601), .Z(n2621) );
  XOR U3318 ( .A(n2625), .B(n2626), .Z(n2604) );
  AND U3319 ( .A(n2627), .B(n2628), .Z(n2626) );
  XOR U3320 ( .A(n2629), .B(n2630), .Z(n2628) );
  XOR U3321 ( .A(n2625), .B(n2631), .Z(n2630) );
  XOR U3322 ( .A(n2623), .B(n2632), .Z(n2627) );
  XOR U3323 ( .A(n2625), .B(n2624), .Z(n2632) );
  NAND U3324 ( .A(n1106), .B(n1987), .Z(n2615) );
  XOR U3325 ( .A(n2613), .B(n2633), .Z(n2614) );
  AND U3326 ( .A(n1946), .B(n1158), .Z(n2633) );
  XOR U3327 ( .A(n2618), .B(n2638), .Z(n2619) );
  AND U3328 ( .A(n1868), .B(n1256), .Z(n2638) );
  XNOR U3329 ( .A(n2642), .B(n2620), .Z(n2637) );
  NAND U3330 ( .A(n1206), .B(n1907), .Z(n2620) );
  IV U3331 ( .A(n2622), .Z(n2642) );
  XOR U3332 ( .A(n2646), .B(n2647), .Z(n2625) );
  AND U3333 ( .A(n2648), .B(n2649), .Z(n2647) );
  XOR U3334 ( .A(n2650), .B(n2651), .Z(n2649) );
  XOR U3335 ( .A(n2646), .B(n2652), .Z(n2651) );
  XOR U3336 ( .A(n2644), .B(n2653), .Z(n2648) );
  XOR U3337 ( .A(n2646), .B(n2645), .Z(n2653) );
  NAND U3338 ( .A(n1106), .B(n2028), .Z(n2636) );
  XOR U3339 ( .A(n2634), .B(n2654), .Z(n2635) );
  AND U3340 ( .A(n1987), .B(n1158), .Z(n2654) );
  XOR U3341 ( .A(n2655), .B(n2656), .Z(n2634) );
  ANDN U3342 ( .A(n2657), .B(n2658), .Z(n2656) );
  XNOR U3343 ( .A(n2659), .B(n2655), .Z(n2657) );
  XOR U3344 ( .A(n2639), .B(n2661), .Z(n2640) );
  AND U3345 ( .A(n1907), .B(n1256), .Z(n2661) );
  XNOR U3346 ( .A(n2665), .B(n2641), .Z(n2660) );
  NAND U3347 ( .A(n1206), .B(n1946), .Z(n2641) );
  IV U3348 ( .A(n2643), .Z(n2665) );
  XNOR U3349 ( .A(n2670), .B(n2671), .Z(n2514) );
  XNOR U3350 ( .A(n2672), .B(n2669), .Z(n2670) );
  XOR U3351 ( .A(n2662), .B(n2674), .Z(n2663) );
  AND U3352 ( .A(n1946), .B(n1256), .Z(n2674) );
  XOR U3353 ( .A(n2677), .B(n2675), .Z(n2676) );
  AND U3354 ( .A(n1987), .B(n1256), .Z(n2677) );
  AND U3355 ( .A(n2028), .B(n1206), .Z(n2678) );
  XNOR U3356 ( .A(n2682), .B(n2664), .Z(n2673) );
  NAND U3357 ( .A(n1206), .B(n1987), .Z(n2664) );
  IV U3358 ( .A(n2666), .Z(n2682) );
  NAND U3359 ( .A(n1206), .B(n2683), .Z(n2681) );
  XOR U3360 ( .A(n2679), .B(n2684), .Z(n2680) );
  AND U3361 ( .A(n2028), .B(n1256), .Z(n2684) );
  ANDN U3362 ( .A(n2685), .B(n2686), .Z(n2679) );
  NANDN U3363 ( .B(n1206), .A(n2687), .Z(n2685) );
  NAND U3364 ( .A(n2683), .B(n1256), .Z(n2687) );
  XNOR U3365 ( .A(n2688), .B(e_input[4]), .Z(n1256) );
  NAND U3366 ( .A(e_input[31]), .B(n2689), .Z(n2688) );
  XOR U3367 ( .A(e_input[4]), .B(\_MAC/_MULT/X_[4] ), .Z(n2689) );
  XNOR U3368 ( .A(n2690), .B(e_input[5]), .Z(n1206) );
  NAND U3369 ( .A(e_input[31]), .B(n2691), .Z(n2690) );
  XOR U3370 ( .A(e_input[5]), .B(\_MAC/_MULT/X_[5] ), .Z(n2691) );
  XNOR U3371 ( .A(n2658), .B(n2659), .Z(n2668) );
  NAND U3372 ( .A(n1106), .B(n2683), .Z(n2659) );
  XNOR U3373 ( .A(n2655), .B(n2692), .Z(n2658) );
  AND U3374 ( .A(n2028), .B(n1158), .Z(n2692) );
  ANDN U3375 ( .A(n2693), .B(n2686), .Z(n2655) );
  NANDN U3376 ( .B(n1106), .A(n2694), .Z(n2693) );
  NAND U3377 ( .A(n2683), .B(n1158), .Z(n2694) );
  XNOR U3378 ( .A(n2695), .B(e_input[6]), .Z(n1158) );
  NAND U3379 ( .A(e_input[31]), .B(n2696), .Z(n2695) );
  XOR U3380 ( .A(e_input[6]), .B(\_MAC/_MULT/X_[6] ), .Z(n2696) );
  XNOR U3381 ( .A(n2697), .B(e_input[7]), .Z(n1106) );
  NAND U3382 ( .A(e_input[31]), .B(n2698), .Z(n2697) );
  XOR U3383 ( .A(e_input[7]), .B(\_MAC/_MULT/X_[7] ), .Z(n2698) );
  XOR U3384 ( .A(n2699), .B(n2700), .Z(n2669) );
  XOR U3385 ( .A(n2492), .B(n2702), .Z(n2493) );
  ANDN U3386 ( .A(n1476), .B(n2337), .Z(n2702) );
  XNOR U3387 ( .A(n2706), .B(n2494), .Z(n2701) );
  NANDN U3388 ( .B(n2329), .A(n1515), .Z(n2494) );
  IV U3389 ( .A(n2496), .Z(n2706) );
  NAND U3390 ( .A(n1632), .B(n1334), .Z(n2519) );
  XOR U3391 ( .A(n2517), .B(n2708), .Z(n2518) );
  AND U3392 ( .A(n1399), .B(n1593), .Z(n2708) );
  XOR U3393 ( .A(n2703), .B(n2713), .Z(n2704) );
  ANDN U3394 ( .A(n1515), .B(n2337), .Z(n2713) );
  XNOR U3395 ( .A(n2717), .B(n2705), .Z(n2712) );
  NANDN U3396 ( .B(n2329), .A(n1554), .Z(n2705) );
  IV U3397 ( .A(n2707), .Z(n2717) );
  NAND U3398 ( .A(n1671), .B(n1334), .Z(n2711) );
  XOR U3399 ( .A(n2709), .B(n2719), .Z(n2710) );
  AND U3400 ( .A(n1399), .B(n1632), .Z(n2719) );
  XOR U3401 ( .A(n2714), .B(n2724), .Z(n2715) );
  ANDN U3402 ( .A(n1554), .B(n2337), .Z(n2724) );
  XNOR U3403 ( .A(n2728), .B(n2716), .Z(n2723) );
  NANDN U3404 ( .B(n2329), .A(n1593), .Z(n2716) );
  IV U3405 ( .A(n2718), .Z(n2728) );
  NAND U3406 ( .A(n1710), .B(n1334), .Z(n2722) );
  XOR U3407 ( .A(n2720), .B(n2730), .Z(n2721) );
  AND U3408 ( .A(n1399), .B(n1671), .Z(n2730) );
  XOR U3409 ( .A(n2725), .B(n2735), .Z(n2726) );
  ANDN U3410 ( .A(n1593), .B(n2337), .Z(n2735) );
  XNOR U3411 ( .A(n2739), .B(n2727), .Z(n2734) );
  NANDN U3412 ( .B(n2329), .A(n1632), .Z(n2727) );
  IV U3413 ( .A(n2729), .Z(n2739) );
  NAND U3414 ( .A(n1749), .B(n1334), .Z(n2733) );
  XOR U3415 ( .A(n2731), .B(n2741), .Z(n2732) );
  AND U3416 ( .A(n1399), .B(n1710), .Z(n2741) );
  XOR U3417 ( .A(n2736), .B(n2746), .Z(n2737) );
  ANDN U3418 ( .A(n1632), .B(n2337), .Z(n2746) );
  XNOR U3419 ( .A(n2750), .B(n2738), .Z(n2745) );
  NANDN U3420 ( .B(n2329), .A(n1671), .Z(n2738) );
  IV U3421 ( .A(n2740), .Z(n2750) );
  NAND U3422 ( .A(n1788), .B(n1334), .Z(n2744) );
  XOR U3423 ( .A(n2742), .B(n2752), .Z(n2743) );
  AND U3424 ( .A(n1399), .B(n1749), .Z(n2752) );
  XOR U3425 ( .A(n2747), .B(n2757), .Z(n2748) );
  ANDN U3426 ( .A(n1671), .B(n2337), .Z(n2757) );
  XNOR U3427 ( .A(n2761), .B(n2749), .Z(n2756) );
  NANDN U3428 ( .B(n2329), .A(n1710), .Z(n2749) );
  IV U3429 ( .A(n2751), .Z(n2761) );
  NAND U3430 ( .A(n1827), .B(n1334), .Z(n2755) );
  XOR U3431 ( .A(n2753), .B(n2763), .Z(n2754) );
  AND U3432 ( .A(n1399), .B(n1788), .Z(n2763) );
  XOR U3433 ( .A(n2758), .B(n2768), .Z(n2759) );
  ANDN U3434 ( .A(n1710), .B(n2337), .Z(n2768) );
  XNOR U3435 ( .A(n2772), .B(n2760), .Z(n2767) );
  NANDN U3436 ( .B(n2329), .A(n1749), .Z(n2760) );
  IV U3437 ( .A(n2762), .Z(n2772) );
  NAND U3438 ( .A(n1868), .B(n1334), .Z(n2766) );
  XOR U3439 ( .A(n2764), .B(n2774), .Z(n2765) );
  AND U3440 ( .A(n1399), .B(n1827), .Z(n2774) );
  XOR U3441 ( .A(n2769), .B(n2779), .Z(n2770) );
  ANDN U3442 ( .A(n1749), .B(n2337), .Z(n2779) );
  XNOR U3443 ( .A(n2783), .B(n2771), .Z(n2778) );
  NANDN U3444 ( .B(n2329), .A(n1788), .Z(n2771) );
  IV U3445 ( .A(n2773), .Z(n2783) );
  XOR U3446 ( .A(n2784), .B(n2785), .Z(n2773) );
  AND U3447 ( .A(n2672), .B(n2786), .Z(n2785) );
  XNOR U3448 ( .A(n2784), .B(n2671), .Z(n2786) );
  XNOR U3449 ( .A(n2776), .B(n2777), .Z(n2671) );
  NAND U3450 ( .A(n1907), .B(n1334), .Z(n2777) );
  XNOR U3451 ( .A(n2775), .B(n2787), .Z(n2776) );
  AND U3452 ( .A(n1399), .B(n1868), .Z(n2787) );
  XNOR U3453 ( .A(n2791), .B(n2788), .Z(n2790) );
  XOR U3454 ( .A(n2780), .B(n2793), .Z(n2781) );
  ANDN U3455 ( .A(n1788), .B(n2337), .Z(n2793) );
  XNOR U3456 ( .A(n2797), .B(n2794), .Z(n2796) );
  XNOR U3457 ( .A(n2798), .B(n2782), .Z(n2792) );
  NANDN U3458 ( .B(n2329), .A(n1827), .Z(n2782) );
  IV U3459 ( .A(n2784), .Z(n2798) );
  XOR U3460 ( .A(n2799), .B(n2800), .Z(n2784) );
  AND U3461 ( .A(n2801), .B(n2802), .Z(n2800) );
  XOR U3462 ( .A(n2795), .B(n2803), .Z(n2802) );
  XNOR U3463 ( .A(n2797), .B(n2799), .Z(n2803) );
  NANDN U3464 ( .B(n2329), .A(n1868), .Z(n2797) );
  XOR U3465 ( .A(n2794), .B(n2804), .Z(n2795) );
  ANDN U3466 ( .A(n1827), .B(n2337), .Z(n2804) );
  XNOR U3467 ( .A(n2808), .B(n2805), .Z(n2807) );
  XOR U3468 ( .A(n2789), .B(n2809), .Z(n2801) );
  XNOR U3469 ( .A(n2791), .B(n2799), .Z(n2809) );
  NAND U3470 ( .A(n1334), .B(n1946), .Z(n2791) );
  XOR U3471 ( .A(n2788), .B(n2810), .Z(n2789) );
  AND U3472 ( .A(n1399), .B(n1907), .Z(n2810) );
  XNOR U3473 ( .A(n2814), .B(n2811), .Z(n2813) );
  XOR U3474 ( .A(n2815), .B(n2816), .Z(n2799) );
  AND U3475 ( .A(n2817), .B(n2818), .Z(n2816) );
  XOR U3476 ( .A(n2806), .B(n2819), .Z(n2818) );
  XNOR U3477 ( .A(n2808), .B(n2815), .Z(n2819) );
  NANDN U3478 ( .B(n2329), .A(n1907), .Z(n2808) );
  XOR U3479 ( .A(n2805), .B(n2820), .Z(n2806) );
  ANDN U3480 ( .A(n1868), .B(n2337), .Z(n2820) );
  XNOR U3481 ( .A(n2824), .B(n2821), .Z(n2823) );
  XOR U3482 ( .A(n2812), .B(n2825), .Z(n2817) );
  XNOR U3483 ( .A(n2814), .B(n2815), .Z(n2825) );
  NAND U3484 ( .A(n1334), .B(n1987), .Z(n2814) );
  XOR U3485 ( .A(n2811), .B(n2826), .Z(n2812) );
  AND U3486 ( .A(n1946), .B(n1399), .Z(n2826) );
  XNOR U3487 ( .A(n2830), .B(n2827), .Z(n2829) );
  XOR U3488 ( .A(n2831), .B(n2832), .Z(n2815) );
  AND U3489 ( .A(n2833), .B(n2834), .Z(n2832) );
  XOR U3490 ( .A(n2822), .B(n2835), .Z(n2834) );
  XNOR U3491 ( .A(n2824), .B(n2831), .Z(n2835) );
  NANDN U3492 ( .B(n2329), .A(n1946), .Z(n2824) );
  XOR U3493 ( .A(n2821), .B(n2836), .Z(n2822) );
  ANDN U3494 ( .A(n1907), .B(n2337), .Z(n2836) );
  XOR U3495 ( .A(n2828), .B(n2840), .Z(n2833) );
  XNOR U3496 ( .A(n2830), .B(n2831), .Z(n2840) );
  NAND U3497 ( .A(n1334), .B(n2028), .Z(n2830) );
  XOR U3498 ( .A(n2827), .B(n2841), .Z(n2828) );
  AND U3499 ( .A(n1987), .B(n1399), .Z(n2841) );
  XOR U3500 ( .A(n2842), .B(n2843), .Z(n2827) );
  AND U3501 ( .A(n2844), .B(n2845), .Z(n2843) );
  XNOR U3502 ( .A(n2846), .B(n2842), .Z(n2844) );
  NAND U3503 ( .A(n1334), .B(n2683), .Z(n2846) );
  XOR U3504 ( .A(n2842), .B(n2848), .Z(n2845) );
  AND U3505 ( .A(n2028), .B(n1399), .Z(n2848) );
  ANDN U3506 ( .A(n2849), .B(n2686), .Z(n2842) );
  NANDN U3507 ( .B(n1334), .A(n2850), .Z(n2849) );
  NAND U3508 ( .A(n2683), .B(n1399), .Z(n2850) );
  XNOR U3509 ( .A(n2851), .B(e_input[2]), .Z(n1399) );
  NAND U3510 ( .A(e_input[31]), .B(n2852), .Z(n2851) );
  XOR U3511 ( .A(e_input[2]), .B(\_MAC/_MULT/X_[2] ), .Z(n2852) );
  XNOR U3512 ( .A(n2853), .B(e_input[3]), .Z(n1334) );
  NAND U3513 ( .A(e_input[31]), .B(n2854), .Z(n2853) );
  XOR U3514 ( .A(e_input[3]), .B(\_MAC/_MULT/X_[3] ), .Z(n2854) );
  XOR U3515 ( .A(n2837), .B(n2856), .Z(n2838) );
  ANDN U3516 ( .A(n1946), .B(n2337), .Z(n2856) );
  XOR U3517 ( .A(n2859), .B(n2857), .Z(n2858) );
  ANDN U3518 ( .A(n1987), .B(n2337), .Z(n2859) );
  ANDN U3519 ( .A(n2028), .B(n2329), .Z(n2860) );
  XOR U3520 ( .A(n2861), .B(n2862), .Z(n2857) );
  AND U3521 ( .A(n2863), .B(n2864), .Z(n2862) );
  XNOR U3522 ( .A(n2865), .B(n2861), .Z(n2863) );
  XNOR U3523 ( .A(n2866), .B(n2839), .Z(n2855) );
  NANDN U3524 ( .B(n2329), .A(n1987), .Z(n2839) );
  IV U3525 ( .A(n2847), .Z(n2866) );
  NANDN U3526 ( .B(n2329), .A(n2683), .Z(n2865) );
  XOR U3527 ( .A(n2861), .B(n2867), .Z(n2864) );
  ANDN U3528 ( .A(n2028), .B(n2337), .Z(n2867) );
  ANDN U3529 ( .A(n2868), .B(n2686), .Z(n2861) );
  NAND U3530 ( .A(n2869), .B(n2329), .Z(n2868) );
  XOR U3531 ( .A(n2870), .B(e_input[1]), .Z(n2329) );
  NAND U3532 ( .A(e_input[31]), .B(n2871), .Z(n2870) );
  XOR U3533 ( .A(e_input[1]), .B(\_MAC/_MULT/X_[1] ), .Z(n2871) );
  NANDN U3534 ( .B(n2337), .A(n2683), .Z(n2869) );
  XOR U3535 ( .A(n2872), .B(e_input[0]), .Z(n2337) );
  NAND U3536 ( .A(e_input[31]), .B(n2873), .Z(n2872) );
  XOR U3537 ( .A(e_input[0]), .B(\_MAC/_MULT/X_[0] ), .Z(n2873) );
  XOR U3538 ( .A(n2874), .B(n2053), .Z(n2041) );
  XNOR U3539 ( .A(n2038), .B(n2039), .Z(n2053) );
  NAND U3540 ( .A(n925), .B(n1907), .Z(n2039) );
  XNOR U3541 ( .A(n2037), .B(n2875), .Z(n2038) );
  AND U3542 ( .A(n1868), .B(n954), .Z(n2875) );
  XNOR U3543 ( .A(n2879), .B(n2876), .Z(n2878) );
  XNOR U3544 ( .A(n2051), .B(n2040), .Z(n2874) );
  XOR U3545 ( .A(n2880), .B(n2881), .Z(n2040) );
  XOR U3546 ( .A(n2045), .B(n2883), .Z(n2046) );
  AND U3547 ( .A(n1788), .B(n1031), .Z(n2883) );
  XNOR U3548 ( .A(n2887), .B(n2884), .Z(n2886) );
  XNOR U3549 ( .A(n2888), .B(n2047), .Z(n2882) );
  NAND U3550 ( .A(n998), .B(n1827), .Z(n2047) );
  IV U3551 ( .A(n2049), .Z(n2888) );
  XOR U3552 ( .A(n2889), .B(n2890), .Z(n2049) );
  AND U3553 ( .A(n2891), .B(n2892), .Z(n2890) );
  XOR U3554 ( .A(n2885), .B(n2893), .Z(n2892) );
  XNOR U3555 ( .A(n2887), .B(n2889), .Z(n2893) );
  NAND U3556 ( .A(n998), .B(n1868), .Z(n2887) );
  XOR U3557 ( .A(n2884), .B(n2894), .Z(n2885) );
  AND U3558 ( .A(n1827), .B(n1031), .Z(n2894) );
  XNOR U3559 ( .A(n2898), .B(n2895), .Z(n2897) );
  XOR U3560 ( .A(n2877), .B(n2899), .Z(n2891) );
  XNOR U3561 ( .A(n2879), .B(n2889), .Z(n2899) );
  NAND U3562 ( .A(n925), .B(n1946), .Z(n2879) );
  XOR U3563 ( .A(n2876), .B(n2900), .Z(n2877) );
  AND U3564 ( .A(n1907), .B(n954), .Z(n2900) );
  XNOR U3565 ( .A(n2904), .B(n2901), .Z(n2903) );
  XOR U3566 ( .A(n2905), .B(n2906), .Z(n2889) );
  AND U3567 ( .A(n2907), .B(n2908), .Z(n2906) );
  XOR U3568 ( .A(n2896), .B(n2909), .Z(n2908) );
  XNOR U3569 ( .A(n2898), .B(n2905), .Z(n2909) );
  NAND U3570 ( .A(n998), .B(n1907), .Z(n2898) );
  XOR U3571 ( .A(n2895), .B(n2910), .Z(n2896) );
  AND U3572 ( .A(n1868), .B(n1031), .Z(n2910) );
  XNOR U3573 ( .A(n2914), .B(n2911), .Z(n2913) );
  XOR U3574 ( .A(n2902), .B(n2915), .Z(n2907) );
  XNOR U3575 ( .A(n2904), .B(n2905), .Z(n2915) );
  NAND U3576 ( .A(n925), .B(n1987), .Z(n2904) );
  XOR U3577 ( .A(n2901), .B(n2916), .Z(n2902) );
  AND U3578 ( .A(n1946), .B(n954), .Z(n2916) );
  XNOR U3579 ( .A(n2920), .B(n2917), .Z(n2919) );
  XOR U3580 ( .A(n2921), .B(n2922), .Z(n2905) );
  AND U3581 ( .A(n2923), .B(n2924), .Z(n2922) );
  XOR U3582 ( .A(n2912), .B(n2925), .Z(n2924) );
  XNOR U3583 ( .A(n2914), .B(n2921), .Z(n2925) );
  NAND U3584 ( .A(n998), .B(n1946), .Z(n2914) );
  XOR U3585 ( .A(n2911), .B(n2926), .Z(n2912) );
  AND U3586 ( .A(n1907), .B(n1031), .Z(n2926) );
  XOR U3587 ( .A(n2918), .B(n2930), .Z(n2923) );
  XNOR U3588 ( .A(n2920), .B(n2921), .Z(n2930) );
  NAND U3589 ( .A(n925), .B(n2028), .Z(n2920) );
  XOR U3590 ( .A(n2917), .B(n2931), .Z(n2918) );
  AND U3591 ( .A(n1987), .B(n954), .Z(n2931) );
  XOR U3592 ( .A(n2932), .B(n2933), .Z(n2917) );
  AND U3593 ( .A(n2934), .B(n2935), .Z(n2933) );
  XNOR U3594 ( .A(n2936), .B(n2932), .Z(n2934) );
  NAND U3595 ( .A(n925), .B(n2683), .Z(n2936) );
  XOR U3596 ( .A(n2932), .B(n2938), .Z(n2935) );
  AND U3597 ( .A(n2028), .B(n954), .Z(n2938) );
  ANDN U3598 ( .A(n2939), .B(n2686), .Z(n2932) );
  NANDN U3599 ( .B(n925), .A(n2940), .Z(n2939) );
  NAND U3600 ( .A(n2683), .B(n954), .Z(n2940) );
  XNOR U3601 ( .A(n2941), .B(e_input[10]), .Z(n954) );
  NAND U3602 ( .A(e_input[31]), .B(n2942), .Z(n2941) );
  XOR U3603 ( .A(e_input[10]), .B(\_MAC/_MULT/X_[10] ), .Z(n2942) );
  XNOR U3604 ( .A(n2943), .B(e_input[11]), .Z(n925) );
  NAND U3605 ( .A(e_input[31]), .B(n2944), .Z(n2943) );
  XOR U3606 ( .A(e_input[11]), .B(\_MAC/_MULT/X_[11] ), .Z(n2944) );
  XOR U3607 ( .A(n2927), .B(n2946), .Z(n2928) );
  AND U3608 ( .A(n1946), .B(n1031), .Z(n2946) );
  XOR U3609 ( .A(n2949), .B(n2947), .Z(n2948) );
  AND U3610 ( .A(n1987), .B(n1031), .Z(n2949) );
  AND U3611 ( .A(n2028), .B(n998), .Z(n2950) );
  XNOR U3612 ( .A(n2954), .B(n2929), .Z(n2945) );
  NAND U3613 ( .A(n998), .B(n1987), .Z(n2929) );
  IV U3614 ( .A(n2937), .Z(n2954) );
  NAND U3615 ( .A(n998), .B(n2683), .Z(n2953) );
  XOR U3616 ( .A(n2951), .B(n2955), .Z(n2952) );
  AND U3617 ( .A(n2028), .B(n1031), .Z(n2955) );
  ANDN U3618 ( .A(n2956), .B(n2686), .Z(n2951) );
  NANDN U3619 ( .B(n998), .A(n2957), .Z(n2956) );
  NAND U3620 ( .A(n2683), .B(n1031), .Z(n2957) );
  XNOR U3621 ( .A(n2958), .B(e_input[8]), .Z(n1031) );
  NAND U3622 ( .A(e_input[31]), .B(n2959), .Z(n2958) );
  XOR U3623 ( .A(e_input[8]), .B(\_MAC/_MULT/X_[8] ), .Z(n2959) );
  XNOR U3624 ( .A(n2960), .B(e_input[9]), .Z(n998) );
  NAND U3625 ( .A(e_input[31]), .B(n2961), .Z(n2960) );
  XOR U3626 ( .A(e_input[9]), .B(\_MAC/_MULT/X_[9] ), .Z(n2961) );
  XOR U3627 ( .A(n2019), .B(n2963), .Z(n2020) );
  AND U3628 ( .A(n1946), .B(n907), .Z(n2963) );
  XOR U3629 ( .A(n2966), .B(n2964), .Z(n2965) );
  AND U3630 ( .A(n1987), .B(n907), .Z(n2966) );
  AND U3631 ( .A(n2028), .B(n880), .Z(n2967) );
  XNOR U3632 ( .A(n2971), .B(n2021), .Z(n2962) );
  NAND U3633 ( .A(n880), .B(n1987), .Z(n2021) );
  IV U3634 ( .A(n2023), .Z(n2971) );
  NAND U3635 ( .A(n880), .B(n2683), .Z(n2970) );
  XOR U3636 ( .A(n2968), .B(n2972), .Z(n2969) );
  AND U3637 ( .A(n2028), .B(n907), .Z(n2972) );
  ANDN U3638 ( .A(n2973), .B(n2686), .Z(n2968) );
  NANDN U3639 ( .B(n880), .A(n2974), .Z(n2973) );
  NAND U3640 ( .A(n2683), .B(n907), .Z(n2974) );
  XNOR U3641 ( .A(n2975), .B(e_input[12]), .Z(n907) );
  NAND U3642 ( .A(e_input[31]), .B(n2976), .Z(n2975) );
  XOR U3643 ( .A(e_input[12]), .B(\_MAC/_MULT/X_[12] ), .Z(n2976) );
  XNOR U3644 ( .A(n2977), .B(e_input[13]), .Z(n880) );
  NAND U3645 ( .A(e_input[31]), .B(n2978), .Z(n2977) );
  XOR U3646 ( .A(e_input[13]), .B(\_MAC/_MULT/X_[13] ), .Z(n2978) );
  XNOR U3647 ( .A(n2033), .B(n2034), .Z(n2027) );
  NAND U3648 ( .A(n846), .B(n2683), .Z(n2034) );
  XNOR U3649 ( .A(n2030), .B(n2979), .Z(n2033) );
  AND U3650 ( .A(n2028), .B(n864), .Z(n2979) );
  ANDN U3651 ( .A(n2980), .B(n2686), .Z(n2030) );
  NANDN U3652 ( .B(n846), .A(n2981), .Z(n2980) );
  NAND U3653 ( .A(n2683), .B(n864), .Z(n2981) );
  XNOR U3654 ( .A(n2982), .B(e_input[14]), .Z(n864) );
  NAND U3655 ( .A(e_input[31]), .B(n2983), .Z(n2982) );
  XOR U3656 ( .A(e_input[14]), .B(\_MAC/_MULT/X_[14] ), .Z(n2983) );
  XNOR U3657 ( .A(n2984), .B(e_input[15]), .Z(n846) );
  NAND U3658 ( .A(e_input[31]), .B(n2985), .Z(n2984) );
  XOR U3659 ( .A(e_input[15]), .B(\_MAC/_MULT/X_[15] ), .Z(n2985) );
  XNOR U3660 ( .A(n2986), .B(n2987), .Z(\_MAC/_MULT/MULT/S[3][1][9] ) );
  XNOR U3661 ( .A(n2988), .B(n2989), .Z(\_MAC/_MULT/MULT/S[3][1][8] ) );
  XNOR U3662 ( .A(n2990), .B(n2991), .Z(\_MAC/_MULT/MULT/S[3][1][7] ) );
  XNOR U3663 ( .A(n2992), .B(n2993), .Z(\_MAC/_MULT/MULT/S[3][1][6] ) );
  XNOR U3664 ( .A(n2994), .B(n2995), .Z(\_MAC/_MULT/MULT/S[3][1][5] ) );
  XNOR U3665 ( .A(n2996), .B(n2997), .Z(\_MAC/_MULT/MULT/S[3][1][4] ) );
  XNOR U3666 ( .A(n2998), .B(n2999), .Z(\_MAC/_MULT/MULT/S[3][1][3] ) );
  XOR U3667 ( .A(n3000), .B(n3001), .Z(\_MAC/_MULT/MULT/S[3][1][31] ) );
  XOR U3668 ( .A(n3002), .B(n3003), .Z(n3001) );
  XNOR U3669 ( .A(n3004), .B(n3005), .Z(n3003) );
  AND U3670 ( .A(n3006), .B(n3007), .Z(n3005) );
  NAND U3671 ( .A(n3008), .B(n3009), .Z(n3007) );
  NANDN U3672 ( .B(n3010), .A(n3011), .Z(n3006) );
  XOR U3673 ( .A(n3012), .B(n3013), .Z(n3002) );
  AND U3674 ( .A(n3014), .B(\_MAC/_MULT/MULT/S[3][1][30] ), .Z(n3013) );
  ANDN U3675 ( .A(n3015), .B(n3004), .Z(n3012) );
  XOR U3676 ( .A(n3016), .B(n3009), .Z(n3000) );
  XOR U3677 ( .A(n3017), .B(n3014), .Z(n3016) );
  XOR U3678 ( .A(n3014), .B(n3018), .Z(\_MAC/_MULT/MULT/S[3][1][30] ) );
  OR U3679 ( .A(n3019), .B(n3020), .Z(n3004) );
  XOR U3680 ( .A(n3010), .B(n3017), .Z(n3015) );
  IV U3681 ( .A(n3011), .Z(n3017) );
  XNOR U3682 ( .A(n3009), .B(n3008), .Z(n3010) );
  NANDN U3683 ( .B(n845), .A(n3024), .Z(n3008) );
  XNOR U3684 ( .A(n3029), .B(n3030), .Z(\_MAC/_MULT/MULT/S[3][1][2] ) );
  XOR U3685 ( .A(n3028), .B(n3031), .Z(\_MAC/_MULT/MULT/S[3][1][29] ) );
  XOR U3686 ( .A(n3019), .B(n3020), .Z(n3031) );
  NANDN U3687 ( .B(n3032), .A(n3033), .Z(n3020) );
  XOR U3688 ( .A(n3021), .B(n3034), .Z(n3022) );
  ANDN U3689 ( .A(n3035), .B(n3036), .Z(n3034) );
  XNOR U3690 ( .A(n3026), .B(n3027), .Z(n3023) );
  NAND U3691 ( .A(n3024), .B(n862), .Z(n3027) );
  XNOR U3692 ( .A(n3025), .B(n3040), .Z(n3026) );
  ANDN U3693 ( .A(n3041), .B(n845), .Z(n3040) );
  XNOR U3694 ( .A(n3045), .B(n3046), .Z(\_MAC/_MULT/MULT/S[3][1][28] ) );
  XNOR U3695 ( .A(n3054), .B(n3036), .Z(n3050) );
  NANDN U3696 ( .B(n845), .A(n3055), .Z(n3036) );
  IV U3697 ( .A(n3037), .Z(n3054) );
  XNOR U3698 ( .A(n3043), .B(n3044), .Z(n3039) );
  NAND U3699 ( .A(n3024), .B(n884), .Z(n3044) );
  XNOR U3700 ( .A(n3042), .B(n3059), .Z(n3043) );
  AND U3701 ( .A(n862), .B(n3041), .Z(n3059) );
  XNOR U3702 ( .A(n3064), .B(n3063), .Z(\_MAC/_MULT/MULT/S[3][1][27] ) );
  OR U3703 ( .A(n3065), .B(n3066), .Z(n3063) );
  XNOR U3704 ( .A(n3049), .B(n3048), .Z(n3064) );
  XOR U3705 ( .A(n3067), .B(n3068), .Z(n3048) );
  XOR U3706 ( .A(n3069), .B(n3070), .Z(n3068) );
  AND U3707 ( .A(n3071), .B(n3072), .Z(n3069) );
  NAND U3708 ( .A(n3073), .B(n3074), .Z(n3072) );
  NANDN U3709 ( .B(n3075), .A(n3070), .Z(n3071) );
  XOR U3710 ( .A(n3051), .B(n3080), .Z(n3052) );
  ANDN U3711 ( .A(n3081), .B(n845), .Z(n3080) );
  XNOR U3712 ( .A(n3085), .B(n3053), .Z(n3079) );
  NAND U3713 ( .A(n3055), .B(n862), .Z(n3053) );
  IV U3714 ( .A(n3056), .Z(n3085) );
  XNOR U3715 ( .A(n3061), .B(n3062), .Z(n3058) );
  NAND U3716 ( .A(n3024), .B(n915), .Z(n3062) );
  XNOR U3717 ( .A(n3060), .B(n3089), .Z(n3061) );
  AND U3718 ( .A(n884), .B(n3041), .Z(n3089) );
  XOR U3719 ( .A(n3066), .B(n3065), .Z(\_MAC/_MULT/MULT/S[3][1][26] ) );
  OR U3720 ( .A(n3093), .B(n3094), .Z(n3065) );
  XNOR U3721 ( .A(n3095), .B(n3075), .Z(n3077) );
  XNOR U3722 ( .A(n3074), .B(n3073), .Z(n3075) );
  NANDN U3723 ( .B(n845), .A(n3096), .Z(n3073) );
  XNOR U3724 ( .A(n3070), .B(n3076), .Z(n3095) );
  XNOR U3725 ( .A(n3103), .B(n3106), .Z(n3105) );
  XOR U3726 ( .A(n3082), .B(n3108), .Z(n3083) );
  AND U3727 ( .A(n862), .B(n3081), .Z(n3108) );
  XNOR U3728 ( .A(n3112), .B(n3084), .Z(n3107) );
  NAND U3729 ( .A(n3055), .B(n884), .Z(n3084) );
  IV U3730 ( .A(n3086), .Z(n3112) );
  XOR U3731 ( .A(n3113), .B(n3114), .Z(n3086) );
  AND U3732 ( .A(n3115), .B(n3116), .Z(n3114) );
  XNOR U3733 ( .A(n3113), .B(n3117), .Z(n3115) );
  XNOR U3734 ( .A(n3091), .B(n3092), .Z(n3088) );
  NAND U3735 ( .A(n3024), .B(n945), .Z(n3092) );
  XNOR U3736 ( .A(n3090), .B(n3118), .Z(n3091) );
  AND U3737 ( .A(n915), .B(n3041), .Z(n3118) );
  XOR U3738 ( .A(n3093), .B(n3094), .Z(\_MAC/_MULT/MULT/S[3][1][25] ) );
  NANDN U3739 ( .B(n3122), .A(n3123), .Z(n3094) );
  XOR U3740 ( .A(n3124), .B(n3106), .Z(n3101) );
  XNOR U3741 ( .A(n3098), .B(n3099), .Z(n3106) );
  NAND U3742 ( .A(n3096), .B(n862), .Z(n3099) );
  XNOR U3743 ( .A(n3097), .B(n3125), .Z(n3098) );
  ANDN U3744 ( .A(n3126), .B(n845), .Z(n3125) );
  XNOR U3745 ( .A(n3104), .B(n3100), .Z(n3124) );
  XOR U3746 ( .A(n3103), .B(n3133), .Z(n3104) );
  ANDN U3747 ( .A(n3134), .B(n3135), .Z(n3133) );
  XOR U3748 ( .A(n3109), .B(n3140), .Z(n3110) );
  AND U3749 ( .A(n884), .B(n3081), .Z(n3140) );
  XNOR U3750 ( .A(n3144), .B(n3111), .Z(n3139) );
  NAND U3751 ( .A(n3055), .B(n915), .Z(n3111) );
  IV U3752 ( .A(n3113), .Z(n3144) );
  XNOR U3753 ( .A(n3120), .B(n3121), .Z(n3117) );
  NAND U3754 ( .A(n3024), .B(n976), .Z(n3121) );
  XNOR U3755 ( .A(n3119), .B(n3148), .Z(n3120) );
  AND U3756 ( .A(n945), .B(n3041), .Z(n3148) );
  XNOR U3757 ( .A(n3122), .B(n3123), .Z(\_MAC/_MULT/MULT/S[3][1][24] ) );
  XOR U3758 ( .A(n3155), .B(n3138), .Z(n3131) );
  XNOR U3759 ( .A(n3128), .B(n3129), .Z(n3138) );
  NAND U3760 ( .A(n3096), .B(n884), .Z(n3129) );
  XNOR U3761 ( .A(n3127), .B(n3156), .Z(n3128) );
  AND U3762 ( .A(n862), .B(n3126), .Z(n3156) );
  XNOR U3763 ( .A(n3137), .B(n3130), .Z(n3155) );
  XNOR U3764 ( .A(n3167), .B(n3135), .Z(n3163) );
  NANDN U3765 ( .B(n845), .A(n3168), .Z(n3135) );
  IV U3766 ( .A(n3136), .Z(n3167) );
  XOR U3767 ( .A(n3141), .B(n3173), .Z(n3142) );
  AND U3768 ( .A(n915), .B(n3081), .Z(n3173) );
  XNOR U3769 ( .A(n3177), .B(n3143), .Z(n3172) );
  NAND U3770 ( .A(n3055), .B(n945), .Z(n3143) );
  IV U3771 ( .A(n3145), .Z(n3177) );
  XNOR U3772 ( .A(n3150), .B(n3151), .Z(n3147) );
  NAND U3773 ( .A(n3024), .B(n1011), .Z(n3151) );
  XNOR U3774 ( .A(n3149), .B(n3181), .Z(n3150) );
  AND U3775 ( .A(n976), .B(n3041), .Z(n3181) );
  XNOR U3776 ( .A(n3154), .B(n3153), .Z(\_MAC/_MULT/MULT/S[3][1][23] ) );
  XOR U3777 ( .A(n3185), .B(n3186), .Z(n3153) );
  XOR U3778 ( .A(n3187), .B(n3188), .Z(n3186) );
  XOR U3779 ( .A(n3189), .B(n3190), .Z(n3188) );
  NOR U3780 ( .A(n3191), .B(n3192), .Z(n3190) );
  AND U3781 ( .A(n3193), .B(n3194), .Z(n3189) );
  NAND U3782 ( .A(n3195), .B(n3196), .Z(n3194) );
  NANDN U3783 ( .B(n3197), .A(n3187), .Z(n3193) );
  XOR U3784 ( .A(n3201), .B(n3171), .Z(n3161) );
  XNOR U3785 ( .A(n3158), .B(n3159), .Z(n3171) );
  NAND U3786 ( .A(n3096), .B(n915), .Z(n3159) );
  XNOR U3787 ( .A(n3157), .B(n3202), .Z(n3158) );
  AND U3788 ( .A(n884), .B(n3126), .Z(n3202) );
  XNOR U3789 ( .A(n3170), .B(n3160), .Z(n3201) );
  XOR U3790 ( .A(n3164), .B(n3210), .Z(n3165) );
  ANDN U3791 ( .A(n3211), .B(n845), .Z(n3210) );
  XNOR U3792 ( .A(n3215), .B(n3166), .Z(n3209) );
  NAND U3793 ( .A(n3168), .B(n862), .Z(n3166) );
  IV U3794 ( .A(n3169), .Z(n3215) );
  XOR U3795 ( .A(n3174), .B(n3220), .Z(n3175) );
  AND U3796 ( .A(n945), .B(n3081), .Z(n3220) );
  XNOR U3797 ( .A(n3224), .B(n3176), .Z(n3219) );
  NAND U3798 ( .A(n3055), .B(n976), .Z(n3176) );
  IV U3799 ( .A(n3178), .Z(n3224) );
  XNOR U3800 ( .A(n3183), .B(n3184), .Z(n3180) );
  NAND U3801 ( .A(n3024), .B(n1048), .Z(n3184) );
  XNOR U3802 ( .A(n3182), .B(n3228), .Z(n3183) );
  AND U3803 ( .A(n1011), .B(n3041), .Z(n3228) );
  XOR U3804 ( .A(n3200), .B(n3199), .Z(\_MAC/_MULT/MULT/S[3][1][22] ) );
  XNOR U3805 ( .A(n3232), .B(n3192), .Z(n3199) );
  XNOR U3806 ( .A(n3197), .B(n3187), .Z(n3192) );
  XNOR U3807 ( .A(n3196), .B(n3195), .Z(n3197) );
  NANDN U3808 ( .B(n845), .A(n3236), .Z(n3195) );
  OR U3809 ( .A(n3240), .B(n3241), .Z(n3191) );
  XOR U3810 ( .A(n3245), .B(n3218), .Z(n3207) );
  XNOR U3811 ( .A(n3204), .B(n3205), .Z(n3218) );
  NAND U3812 ( .A(n3096), .B(n945), .Z(n3205) );
  XNOR U3813 ( .A(n3203), .B(n3246), .Z(n3204) );
  AND U3814 ( .A(n915), .B(n3126), .Z(n3246) );
  XNOR U3815 ( .A(n3217), .B(n3206), .Z(n3245) );
  XOR U3816 ( .A(n3212), .B(n3254), .Z(n3213) );
  AND U3817 ( .A(n862), .B(n3211), .Z(n3254) );
  XNOR U3818 ( .A(n3258), .B(n3214), .Z(n3253) );
  NAND U3819 ( .A(n3168), .B(n884), .Z(n3214) );
  IV U3820 ( .A(n3216), .Z(n3258) );
  XOR U3821 ( .A(n3221), .B(n3263), .Z(n3222) );
  AND U3822 ( .A(n976), .B(n3081), .Z(n3263) );
  XNOR U3823 ( .A(n3267), .B(n3223), .Z(n3262) );
  NAND U3824 ( .A(n3055), .B(n1011), .Z(n3223) );
  IV U3825 ( .A(n3225), .Z(n3267) );
  XOR U3826 ( .A(n3268), .B(n3269), .Z(n3225) );
  AND U3827 ( .A(n3270), .B(n3271), .Z(n3269) );
  XNOR U3828 ( .A(n3268), .B(n3272), .Z(n3270) );
  XNOR U3829 ( .A(n3230), .B(n3231), .Z(n3227) );
  NAND U3830 ( .A(n3024), .B(n1097), .Z(n3231) );
  XNOR U3831 ( .A(n3229), .B(n3273), .Z(n3230) );
  AND U3832 ( .A(n1048), .B(n3041), .Z(n3273) );
  XNOR U3833 ( .A(n3244), .B(n3243), .Z(\_MAC/_MULT/MULT/S[3][1][21] ) );
  XOR U3834 ( .A(n3277), .B(n3241), .Z(n3243) );
  XOR U3835 ( .A(n3233), .B(n3278), .Z(n3234) );
  ANDN U3836 ( .A(n3279), .B(n3280), .Z(n3278) );
  XNOR U3837 ( .A(n3238), .B(n3239), .Z(n3235) );
  NAND U3838 ( .A(n3236), .B(n862), .Z(n3239) );
  XNOR U3839 ( .A(n3237), .B(n3284), .Z(n3238) );
  ANDN U3840 ( .A(n3285), .B(n845), .Z(n3284) );
  NANDN U3841 ( .B(n3289), .A(n3290), .Z(n3240) );
  XOR U3842 ( .A(n3294), .B(n3261), .Z(n3251) );
  XNOR U3843 ( .A(n3248), .B(n3249), .Z(n3261) );
  NAND U3844 ( .A(n3096), .B(n976), .Z(n3249) );
  XNOR U3845 ( .A(n3247), .B(n3295), .Z(n3248) );
  AND U3846 ( .A(n945), .B(n3126), .Z(n3295) );
  XNOR U3847 ( .A(n3260), .B(n3250), .Z(n3294) );
  XOR U3848 ( .A(n3255), .B(n3303), .Z(n3256) );
  AND U3849 ( .A(n884), .B(n3211), .Z(n3303) );
  XNOR U3850 ( .A(n3307), .B(n3257), .Z(n3302) );
  NAND U3851 ( .A(n3168), .B(n915), .Z(n3257) );
  IV U3852 ( .A(n3259), .Z(n3307) );
  XOR U3853 ( .A(n3264), .B(n3312), .Z(n3265) );
  AND U3854 ( .A(n1011), .B(n3081), .Z(n3312) );
  XNOR U3855 ( .A(n3316), .B(n3266), .Z(n3311) );
  NAND U3856 ( .A(n3055), .B(n1048), .Z(n3266) );
  IV U3857 ( .A(n3268), .Z(n3316) );
  XNOR U3858 ( .A(n3275), .B(n3276), .Z(n3272) );
  NAND U3859 ( .A(n3024), .B(n1145), .Z(n3276) );
  XNOR U3860 ( .A(n3274), .B(n3320), .Z(n3275) );
  AND U3861 ( .A(n1097), .B(n3041), .Z(n3320) );
  XNOR U3862 ( .A(n3293), .B(n3292), .Z(\_MAC/_MULT/MULT/S[3][1][20] ) );
  XOR U3863 ( .A(n3324), .B(n3289), .Z(n3292) );
  XNOR U3864 ( .A(n3329), .B(n3280), .Z(n3325) );
  NANDN U3865 ( .B(n845), .A(n3330), .Z(n3280) );
  IV U3866 ( .A(n3281), .Z(n3329) );
  XNOR U3867 ( .A(n3287), .B(n3288), .Z(n3283) );
  NAND U3868 ( .A(n3236), .B(n884), .Z(n3288) );
  XNOR U3869 ( .A(n3286), .B(n3334), .Z(n3287) );
  AND U3870 ( .A(n862), .B(n3285), .Z(n3334) );
  XNOR U3871 ( .A(n3290), .B(n3291), .Z(n3324) );
  XOR U3872 ( .A(n3344), .B(n3310), .Z(n3300) );
  XNOR U3873 ( .A(n3297), .B(n3298), .Z(n3310) );
  NAND U3874 ( .A(n3096), .B(n1011), .Z(n3298) );
  XNOR U3875 ( .A(n3296), .B(n3345), .Z(n3297) );
  AND U3876 ( .A(n976), .B(n3126), .Z(n3345) );
  XNOR U3877 ( .A(n3309), .B(n3299), .Z(n3344) );
  XOR U3878 ( .A(n3304), .B(n3353), .Z(n3305) );
  AND U3879 ( .A(n915), .B(n3211), .Z(n3353) );
  XNOR U3880 ( .A(n3357), .B(n3306), .Z(n3352) );
  NAND U3881 ( .A(n3168), .B(n945), .Z(n3306) );
  IV U3882 ( .A(n3308), .Z(n3357) );
  XOR U3883 ( .A(n3313), .B(n3362), .Z(n3314) );
  AND U3884 ( .A(n1048), .B(n3081), .Z(n3362) );
  XNOR U3885 ( .A(n3366), .B(n3315), .Z(n3361) );
  NAND U3886 ( .A(n3055), .B(n1097), .Z(n3315) );
  IV U3887 ( .A(n3317), .Z(n3366) );
  XNOR U3888 ( .A(n3322), .B(n3323), .Z(n3319) );
  NAND U3889 ( .A(n3024), .B(n1195), .Z(n3323) );
  XNOR U3890 ( .A(n3321), .B(n3370), .Z(n3322) );
  AND U3891 ( .A(n1145), .B(n3041), .Z(n3370) );
  XNOR U3892 ( .A(n3374), .B(n3375), .Z(\_MAC/_MULT/MULT/S[3][1][1] ) );
  XNOR U3893 ( .A(n3340), .B(n3339), .Z(\_MAC/_MULT/MULT/S[3][1][19] ) );
  XNOR U3894 ( .A(n3376), .B(n3343), .Z(n3339) );
  XOR U3895 ( .A(n3326), .B(n3378), .Z(n3327) );
  ANDN U3896 ( .A(n3379), .B(n845), .Z(n3378) );
  XNOR U3897 ( .A(n3383), .B(n3328), .Z(n3377) );
  NAND U3898 ( .A(n3330), .B(n862), .Z(n3328) );
  IV U3899 ( .A(n3331), .Z(n3383) );
  XNOR U3900 ( .A(n3336), .B(n3337), .Z(n3333) );
  NAND U3901 ( .A(n3236), .B(n915), .Z(n3337) );
  XNOR U3902 ( .A(n3335), .B(n3387), .Z(n3336) );
  AND U3903 ( .A(n884), .B(n3285), .Z(n3387) );
  XNOR U3904 ( .A(n3342), .B(n3338), .Z(n3376) );
  XNOR U3905 ( .A(n3394), .B(n3395), .Z(n3342) );
  XOR U3906 ( .A(n3396), .B(n3397), .Z(n3395) );
  AND U3907 ( .A(n3398), .B(n3399), .Z(n3396) );
  NAND U3908 ( .A(n3400), .B(n3401), .Z(n3399) );
  NANDN U3909 ( .B(n3402), .A(n3397), .Z(n3398) );
  XOR U3910 ( .A(n3406), .B(n3360), .Z(n3350) );
  XNOR U3911 ( .A(n3347), .B(n3348), .Z(n3360) );
  NAND U3912 ( .A(n3096), .B(n1048), .Z(n3348) );
  XNOR U3913 ( .A(n3346), .B(n3407), .Z(n3347) );
  AND U3914 ( .A(n1011), .B(n3126), .Z(n3407) );
  XNOR U3915 ( .A(n3359), .B(n3349), .Z(n3406) );
  XOR U3916 ( .A(n3354), .B(n3415), .Z(n3355) );
  AND U3917 ( .A(n945), .B(n3211), .Z(n3415) );
  XNOR U3918 ( .A(n3419), .B(n3356), .Z(n3414) );
  NAND U3919 ( .A(n3168), .B(n976), .Z(n3356) );
  IV U3920 ( .A(n3358), .Z(n3419) );
  XOR U3921 ( .A(n3363), .B(n3424), .Z(n3364) );
  AND U3922 ( .A(n1097), .B(n3081), .Z(n3424) );
  XNOR U3923 ( .A(n3428), .B(n3365), .Z(n3423) );
  NAND U3924 ( .A(n3055), .B(n1145), .Z(n3365) );
  IV U3925 ( .A(n3367), .Z(n3428) );
  XNOR U3926 ( .A(n3372), .B(n3373), .Z(n3369) );
  NAND U3927 ( .A(n3024), .B(n1248), .Z(n3373) );
  XNOR U3928 ( .A(n3371), .B(n3432), .Z(n3372) );
  AND U3929 ( .A(n1195), .B(n3041), .Z(n3432) );
  XNOR U3930 ( .A(n3393), .B(n3392), .Z(\_MAC/_MULT/MULT/S[3][1][18] ) );
  XOR U3931 ( .A(n3436), .B(n3405), .Z(n3392) );
  XOR U3932 ( .A(n3380), .B(n3438), .Z(n3381) );
  AND U3933 ( .A(n862), .B(n3379), .Z(n3438) );
  XNOR U3934 ( .A(n3442), .B(n3382), .Z(n3437) );
  NAND U3935 ( .A(n3330), .B(n884), .Z(n3382) );
  IV U3936 ( .A(n3384), .Z(n3442) );
  XNOR U3937 ( .A(n3389), .B(n3390), .Z(n3386) );
  NAND U3938 ( .A(n3236), .B(n945), .Z(n3390) );
  XNOR U3939 ( .A(n3388), .B(n3446), .Z(n3389) );
  AND U3940 ( .A(n915), .B(n3285), .Z(n3446) );
  XOR U3941 ( .A(n3404), .B(n3391), .Z(n3436) );
  XOR U3942 ( .A(n3453), .B(n3402), .Z(n3404) );
  XNOR U3943 ( .A(n3401), .B(n3400), .Z(n3402) );
  NANDN U3944 ( .B(n845), .A(n3454), .Z(n3400) );
  XNOR U3945 ( .A(n3397), .B(n3403), .Z(n3453) );
  XNOR U3946 ( .A(n3461), .B(n3464), .Z(n3463) );
  XOR U3947 ( .A(n3465), .B(n3422), .Z(n3412) );
  XNOR U3948 ( .A(n3409), .B(n3410), .Z(n3422) );
  NAND U3949 ( .A(n3096), .B(n1097), .Z(n3410) );
  XNOR U3950 ( .A(n3408), .B(n3466), .Z(n3409) );
  AND U3951 ( .A(n1048), .B(n3126), .Z(n3466) );
  XNOR U3952 ( .A(n3421), .B(n3411), .Z(n3465) );
  XOR U3953 ( .A(n3416), .B(n3474), .Z(n3417) );
  AND U3954 ( .A(n976), .B(n3211), .Z(n3474) );
  XNOR U3955 ( .A(n3478), .B(n3418), .Z(n3473) );
  NAND U3956 ( .A(n3168), .B(n1011), .Z(n3418) );
  IV U3957 ( .A(n3420), .Z(n3478) );
  XOR U3958 ( .A(n3425), .B(n3483), .Z(n3426) );
  AND U3959 ( .A(n1145), .B(n3081), .Z(n3483) );
  XNOR U3960 ( .A(n3487), .B(n3427), .Z(n3482) );
  NAND U3961 ( .A(n3055), .B(n1195), .Z(n3427) );
  IV U3962 ( .A(n3429), .Z(n3487) );
  XNOR U3963 ( .A(n3434), .B(n3435), .Z(n3431) );
  NAND U3964 ( .A(n3024), .B(n1311), .Z(n3435) );
  XNOR U3965 ( .A(n3433), .B(n3491), .Z(n3434) );
  AND U3966 ( .A(n1248), .B(n3041), .Z(n3491) );
  XNOR U3967 ( .A(n3452), .B(n3451), .Z(\_MAC/_MULT/MULT/S[3][1][17] ) );
  XOR U3968 ( .A(n3495), .B(n3460), .Z(n3451) );
  XOR U3969 ( .A(n3439), .B(n3497), .Z(n3440) );
  AND U3970 ( .A(n884), .B(n3379), .Z(n3497) );
  XNOR U3971 ( .A(n3501), .B(n3441), .Z(n3496) );
  NAND U3972 ( .A(n3330), .B(n915), .Z(n3441) );
  IV U3973 ( .A(n3443), .Z(n3501) );
  XOR U3974 ( .A(n3502), .B(n3503), .Z(n3443) );
  AND U3975 ( .A(n3504), .B(n3505), .Z(n3503) );
  XNOR U3976 ( .A(n3502), .B(n3506), .Z(n3504) );
  XNOR U3977 ( .A(n3448), .B(n3449), .Z(n3445) );
  NAND U3978 ( .A(n3236), .B(n976), .Z(n3449) );
  XNOR U3979 ( .A(n3447), .B(n3507), .Z(n3448) );
  AND U3980 ( .A(n945), .B(n3285), .Z(n3507) );
  XNOR U3981 ( .A(n3459), .B(n3450), .Z(n3495) );
  XOR U3982 ( .A(n3514), .B(n3464), .Z(n3459) );
  XNOR U3983 ( .A(n3456), .B(n3457), .Z(n3464) );
  NAND U3984 ( .A(n3454), .B(n862), .Z(n3457) );
  XNOR U3985 ( .A(n3455), .B(n3515), .Z(n3456) );
  ANDN U3986 ( .A(n3516), .B(n845), .Z(n3515) );
  XNOR U3987 ( .A(n3462), .B(n3458), .Z(n3514) );
  XOR U3988 ( .A(n3461), .B(n3523), .Z(n3462) );
  ANDN U3989 ( .A(n3524), .B(n3525), .Z(n3523) );
  XOR U3990 ( .A(n3529), .B(n3481), .Z(n3471) );
  XNOR U3991 ( .A(n3468), .B(n3469), .Z(n3481) );
  NAND U3992 ( .A(n3096), .B(n1145), .Z(n3469) );
  XNOR U3993 ( .A(n3467), .B(n3530), .Z(n3468) );
  AND U3994 ( .A(n1097), .B(n3126), .Z(n3530) );
  XNOR U3995 ( .A(n3480), .B(n3470), .Z(n3529) );
  XOR U3996 ( .A(n3475), .B(n3538), .Z(n3476) );
  AND U3997 ( .A(n1011), .B(n3211), .Z(n3538) );
  XNOR U3998 ( .A(n3542), .B(n3477), .Z(n3537) );
  NAND U3999 ( .A(n3168), .B(n1048), .Z(n3477) );
  IV U4000 ( .A(n3479), .Z(n3542) );
  XOR U4001 ( .A(n3484), .B(n3547), .Z(n3485) );
  AND U4002 ( .A(n1195), .B(n3081), .Z(n3547) );
  XNOR U4003 ( .A(n3551), .B(n3486), .Z(n3546) );
  NAND U4004 ( .A(n3055), .B(n1248), .Z(n3486) );
  IV U4005 ( .A(n3488), .Z(n3551) );
  XNOR U4006 ( .A(n3493), .B(n3494), .Z(n3490) );
  NAND U4007 ( .A(n3024), .B(n1373), .Z(n3494) );
  XNOR U4008 ( .A(n3492), .B(n3555), .Z(n3493) );
  AND U4009 ( .A(n1311), .B(n3041), .Z(n3555) );
  XNOR U4010 ( .A(n3513), .B(n3512), .Z(\_MAC/_MULT/MULT/S[3][1][16] ) );
  XOR U4011 ( .A(n3559), .B(n3522), .Z(n3512) );
  XOR U4012 ( .A(n3498), .B(n3561), .Z(n3499) );
  AND U4013 ( .A(n915), .B(n3379), .Z(n3561) );
  XNOR U4014 ( .A(n3565), .B(n3500), .Z(n3560) );
  NAND U4015 ( .A(n3330), .B(n945), .Z(n3500) );
  IV U4016 ( .A(n3502), .Z(n3565) );
  XNOR U4017 ( .A(n3509), .B(n3510), .Z(n3506) );
  NAND U4018 ( .A(n3236), .B(n1011), .Z(n3510) );
  XNOR U4019 ( .A(n3508), .B(n3569), .Z(n3509) );
  AND U4020 ( .A(n976), .B(n3285), .Z(n3569) );
  XNOR U4021 ( .A(n3521), .B(n3511), .Z(n3559) );
  XOR U4022 ( .A(n3576), .B(n3528), .Z(n3521) );
  XNOR U4023 ( .A(n3518), .B(n3519), .Z(n3528) );
  NAND U4024 ( .A(n3454), .B(n884), .Z(n3519) );
  XNOR U4025 ( .A(n3517), .B(n3577), .Z(n3518) );
  AND U4026 ( .A(n862), .B(n3516), .Z(n3577) );
  XNOR U4027 ( .A(n3527), .B(n3520), .Z(n3576) );
  XNOR U4028 ( .A(n3588), .B(n3525), .Z(n3584) );
  NANDN U4029 ( .B(n845), .A(n3589), .Z(n3525) );
  IV U4030 ( .A(n3526), .Z(n3588) );
  XOR U4031 ( .A(n3593), .B(n3545), .Z(n3535) );
  XNOR U4032 ( .A(n3532), .B(n3533), .Z(n3545) );
  NAND U4033 ( .A(n3096), .B(n1195), .Z(n3533) );
  XNOR U4034 ( .A(n3531), .B(n3594), .Z(n3532) );
  AND U4035 ( .A(n1145), .B(n3126), .Z(n3594) );
  XNOR U4036 ( .A(n3544), .B(n3534), .Z(n3593) );
  XOR U4037 ( .A(n3539), .B(n3602), .Z(n3540) );
  AND U4038 ( .A(n1048), .B(n3211), .Z(n3602) );
  XNOR U4039 ( .A(n3606), .B(n3541), .Z(n3601) );
  NAND U4040 ( .A(n3168), .B(n1097), .Z(n3541) );
  IV U4041 ( .A(n3543), .Z(n3606) );
  XOR U4042 ( .A(n3548), .B(n3611), .Z(n3549) );
  AND U4043 ( .A(n1248), .B(n3081), .Z(n3611) );
  XNOR U4044 ( .A(n3615), .B(n3550), .Z(n3610) );
  NAND U4045 ( .A(n3055), .B(n1311), .Z(n3550) );
  IV U4046 ( .A(n3552), .Z(n3615) );
  XNOR U4047 ( .A(n3557), .B(n3558), .Z(n3554) );
  NAND U4048 ( .A(n3024), .B(n1440), .Z(n3558) );
  XNOR U4049 ( .A(n3556), .B(n3619), .Z(n3557) );
  AND U4050 ( .A(n1373), .B(n3041), .Z(n3619) );
  XNOR U4051 ( .A(n3575), .B(n3574), .Z(\_MAC/_MULT/MULT/S[3][1][15] ) );
  XOR U4052 ( .A(n3623), .B(n3583), .Z(n3574) );
  XOR U4053 ( .A(n3562), .B(n3625), .Z(n3563) );
  AND U4054 ( .A(n945), .B(n3379), .Z(n3625) );
  XNOR U4055 ( .A(n3629), .B(n3564), .Z(n3624) );
  NAND U4056 ( .A(n3330), .B(n976), .Z(n3564) );
  IV U4057 ( .A(n3566), .Z(n3629) );
  XNOR U4058 ( .A(n3571), .B(n3572), .Z(n3568) );
  NAND U4059 ( .A(n3236), .B(n1048), .Z(n3572) );
  XNOR U4060 ( .A(n3570), .B(n3633), .Z(n3571) );
  AND U4061 ( .A(n1011), .B(n3285), .Z(n3633) );
  XNOR U4062 ( .A(n3582), .B(n3573), .Z(n3623) );
  XOR U4063 ( .A(n3640), .B(n3592), .Z(n3582) );
  XNOR U4064 ( .A(n3579), .B(n3580), .Z(n3592) );
  NAND U4065 ( .A(n3454), .B(n915), .Z(n3580) );
  XNOR U4066 ( .A(n3578), .B(n3641), .Z(n3579) );
  AND U4067 ( .A(n884), .B(n3516), .Z(n3641) );
  XNOR U4068 ( .A(n3591), .B(n3581), .Z(n3640) );
  XOR U4069 ( .A(n3585), .B(n3649), .Z(n3586) );
  ANDN U4070 ( .A(n3650), .B(n845), .Z(n3649) );
  NAND U4071 ( .A(\_MAC/_MULT/A_[31] ), .B(g_input[31]), .Z(n845) );
  XNOR U4072 ( .A(n3654), .B(n3587), .Z(n3648) );
  NAND U4073 ( .A(n3589), .B(n862), .Z(n3587) );
  IV U4074 ( .A(n3590), .Z(n3654) );
  XOR U4075 ( .A(n3658), .B(n3609), .Z(n3599) );
  XNOR U4076 ( .A(n3596), .B(n3597), .Z(n3609) );
  NAND U4077 ( .A(n3096), .B(n1248), .Z(n3597) );
  XNOR U4078 ( .A(n3595), .B(n3659), .Z(n3596) );
  AND U4079 ( .A(n1195), .B(n3126), .Z(n3659) );
  XNOR U4080 ( .A(n3608), .B(n3598), .Z(n3658) );
  XOR U4081 ( .A(n3603), .B(n3667), .Z(n3604) );
  AND U4082 ( .A(n1097), .B(n3211), .Z(n3667) );
  XNOR U4083 ( .A(n3671), .B(n3605), .Z(n3666) );
  NAND U4084 ( .A(n3168), .B(n1145), .Z(n3605) );
  IV U4085 ( .A(n3607), .Z(n3671) );
  XOR U4086 ( .A(n3612), .B(n3676), .Z(n3613) );
  AND U4087 ( .A(n1311), .B(n3081), .Z(n3676) );
  XNOR U4088 ( .A(n3680), .B(n3614), .Z(n3675) );
  NAND U4089 ( .A(n3055), .B(n1373), .Z(n3614) );
  IV U4090 ( .A(n3616), .Z(n3680) );
  XNOR U4091 ( .A(n3621), .B(n3622), .Z(n3618) );
  NAND U4092 ( .A(n3024), .B(n1476), .Z(n3622) );
  XNOR U4093 ( .A(n3620), .B(n3684), .Z(n3621) );
  AND U4094 ( .A(n1440), .B(n3041), .Z(n3684) );
  XNOR U4095 ( .A(n3639), .B(n3638), .Z(\_MAC/_MULT/MULT/S[3][1][14] ) );
  XOR U4096 ( .A(n3688), .B(n3647), .Z(n3638) );
  XOR U4097 ( .A(n3626), .B(n3690), .Z(n3627) );
  AND U4098 ( .A(n976), .B(n3379), .Z(n3690) );
  XNOR U4099 ( .A(n3694), .B(n3628), .Z(n3689) );
  NAND U4100 ( .A(n3330), .B(n1011), .Z(n3628) );
  IV U4101 ( .A(n3630), .Z(n3694) );
  XNOR U4102 ( .A(n3635), .B(n3636), .Z(n3632) );
  NAND U4103 ( .A(n3236), .B(n1097), .Z(n3636) );
  XNOR U4104 ( .A(n3634), .B(n3698), .Z(n3635) );
  AND U4105 ( .A(n1048), .B(n3285), .Z(n3698) );
  XNOR U4106 ( .A(n3646), .B(n3637), .Z(n3688) );
  XOR U4107 ( .A(n3705), .B(n3657), .Z(n3646) );
  XNOR U4108 ( .A(n3643), .B(n3644), .Z(n3657) );
  NAND U4109 ( .A(n3454), .B(n945), .Z(n3644) );
  XNOR U4110 ( .A(n3642), .B(n3706), .Z(n3643) );
  AND U4111 ( .A(n915), .B(n3516), .Z(n3706) );
  XNOR U4112 ( .A(n3656), .B(n3645), .Z(n3705) );
  XOR U4113 ( .A(n3651), .B(n3714), .Z(n3652) );
  AND U4114 ( .A(n862), .B(n3650), .Z(n3714) );
  XNOR U4115 ( .A(n3715), .B(g_input[30]), .Z(n862) );
  NAND U4116 ( .A(n3716), .B(g_input[31]), .Z(n3715) );
  XOR U4117 ( .A(g_input[30]), .B(\_MAC/_MULT/A_[30] ), .Z(n3716) );
  XNOR U4118 ( .A(n3720), .B(n3653), .Z(n3713) );
  NAND U4119 ( .A(n3589), .B(n884), .Z(n3653) );
  IV U4120 ( .A(n3655), .Z(n3720) );
  XOR U4121 ( .A(n3724), .B(n3674), .Z(n3664) );
  XNOR U4122 ( .A(n3661), .B(n3662), .Z(n3674) );
  NAND U4123 ( .A(n3096), .B(n1311), .Z(n3662) );
  XNOR U4124 ( .A(n3660), .B(n3725), .Z(n3661) );
  AND U4125 ( .A(n1248), .B(n3126), .Z(n3725) );
  XNOR U4126 ( .A(n3673), .B(n3663), .Z(n3724) );
  XOR U4127 ( .A(n3668), .B(n3733), .Z(n3669) );
  AND U4128 ( .A(n1145), .B(n3211), .Z(n3733) );
  XNOR U4129 ( .A(n3737), .B(n3670), .Z(n3732) );
  NAND U4130 ( .A(n3168), .B(n1195), .Z(n3670) );
  IV U4131 ( .A(n3672), .Z(n3737) );
  XOR U4132 ( .A(n3677), .B(n3742), .Z(n3678) );
  AND U4133 ( .A(n1373), .B(n3081), .Z(n3742) );
  XNOR U4134 ( .A(n3746), .B(n3679), .Z(n3741) );
  NAND U4135 ( .A(n3055), .B(n1440), .Z(n3679) );
  IV U4136 ( .A(n3681), .Z(n3746) );
  XNOR U4137 ( .A(n3686), .B(n3687), .Z(n3683) );
  NAND U4138 ( .A(n3024), .B(n1515), .Z(n3687) );
  XNOR U4139 ( .A(n3685), .B(n3750), .Z(n3686) );
  AND U4140 ( .A(n1476), .B(n3041), .Z(n3750) );
  XNOR U4141 ( .A(n3704), .B(n3703), .Z(\_MAC/_MULT/MULT/S[3][1][13] ) );
  XOR U4142 ( .A(n3754), .B(n3712), .Z(n3703) );
  XOR U4143 ( .A(n3691), .B(n3756), .Z(n3692) );
  AND U4144 ( .A(n1011), .B(n3379), .Z(n3756) );
  XNOR U4145 ( .A(n3760), .B(n3693), .Z(n3755) );
  NAND U4146 ( .A(n3330), .B(n1048), .Z(n3693) );
  IV U4147 ( .A(n3695), .Z(n3760) );
  XNOR U4148 ( .A(n3700), .B(n3701), .Z(n3697) );
  NAND U4149 ( .A(n3236), .B(n1145), .Z(n3701) );
  XNOR U4150 ( .A(n3699), .B(n3764), .Z(n3700) );
  AND U4151 ( .A(n1097), .B(n3285), .Z(n3764) );
  XNOR U4152 ( .A(n3711), .B(n3702), .Z(n3754) );
  XOR U4153 ( .A(n3771), .B(n3723), .Z(n3711) );
  XNOR U4154 ( .A(n3708), .B(n3709), .Z(n3723) );
  NAND U4155 ( .A(n3454), .B(n976), .Z(n3709) );
  XNOR U4156 ( .A(n3707), .B(n3772), .Z(n3708) );
  AND U4157 ( .A(n945), .B(n3516), .Z(n3772) );
  XNOR U4158 ( .A(n3722), .B(n3710), .Z(n3771) );
  XOR U4159 ( .A(n3717), .B(n3780), .Z(n3718) );
  AND U4160 ( .A(n884), .B(n3650), .Z(n3780) );
  XNOR U4161 ( .A(n3781), .B(g_input[29]), .Z(n884) );
  NAND U4162 ( .A(n3782), .B(g_input[31]), .Z(n3781) );
  XOR U4163 ( .A(g_input[29]), .B(\_MAC/_MULT/A_[29] ), .Z(n3782) );
  XNOR U4164 ( .A(n3786), .B(n3719), .Z(n3779) );
  NAND U4165 ( .A(n3589), .B(n915), .Z(n3719) );
  IV U4166 ( .A(n3721), .Z(n3786) );
  XOR U4167 ( .A(n3790), .B(n3740), .Z(n3730) );
  XNOR U4168 ( .A(n3727), .B(n3728), .Z(n3740) );
  NAND U4169 ( .A(n3096), .B(n1373), .Z(n3728) );
  XNOR U4170 ( .A(n3726), .B(n3791), .Z(n3727) );
  AND U4171 ( .A(n1311), .B(n3126), .Z(n3791) );
  XNOR U4172 ( .A(n3739), .B(n3729), .Z(n3790) );
  XOR U4173 ( .A(n3734), .B(n3799), .Z(n3735) );
  AND U4174 ( .A(n1195), .B(n3211), .Z(n3799) );
  XNOR U4175 ( .A(n3803), .B(n3736), .Z(n3798) );
  NAND U4176 ( .A(n3168), .B(n1248), .Z(n3736) );
  IV U4177 ( .A(n3738), .Z(n3803) );
  XOR U4178 ( .A(n3743), .B(n3808), .Z(n3744) );
  AND U4179 ( .A(n1440), .B(n3081), .Z(n3808) );
  XNOR U4180 ( .A(n3812), .B(n3745), .Z(n3807) );
  NAND U4181 ( .A(n3055), .B(n1476), .Z(n3745) );
  IV U4182 ( .A(n3747), .Z(n3812) );
  XNOR U4183 ( .A(n3752), .B(n3753), .Z(n3749) );
  NAND U4184 ( .A(n3024), .B(n1554), .Z(n3753) );
  XNOR U4185 ( .A(n3751), .B(n3816), .Z(n3752) );
  AND U4186 ( .A(n1515), .B(n3041), .Z(n3816) );
  XNOR U4187 ( .A(n3770), .B(n3769), .Z(\_MAC/_MULT/MULT/S[3][1][12] ) );
  XOR U4188 ( .A(n3820), .B(n3778), .Z(n3769) );
  XOR U4189 ( .A(n3757), .B(n3822), .Z(n3758) );
  AND U4190 ( .A(n1048), .B(n3379), .Z(n3822) );
  XNOR U4191 ( .A(n3826), .B(n3759), .Z(n3821) );
  NAND U4192 ( .A(n3330), .B(n1097), .Z(n3759) );
  IV U4193 ( .A(n3761), .Z(n3826) );
  XNOR U4194 ( .A(n3766), .B(n3767), .Z(n3763) );
  NAND U4195 ( .A(n3236), .B(n1195), .Z(n3767) );
  XNOR U4196 ( .A(n3765), .B(n3830), .Z(n3766) );
  AND U4197 ( .A(n1145), .B(n3285), .Z(n3830) );
  XNOR U4198 ( .A(n3777), .B(n3768), .Z(n3820) );
  XOR U4199 ( .A(n3837), .B(n3789), .Z(n3777) );
  XNOR U4200 ( .A(n3774), .B(n3775), .Z(n3789) );
  NAND U4201 ( .A(n3454), .B(n1011), .Z(n3775) );
  XNOR U4202 ( .A(n3773), .B(n3838), .Z(n3774) );
  AND U4203 ( .A(n976), .B(n3516), .Z(n3838) );
  XNOR U4204 ( .A(n3788), .B(n3776), .Z(n3837) );
  XOR U4205 ( .A(n3783), .B(n3846), .Z(n3784) );
  AND U4206 ( .A(n915), .B(n3650), .Z(n3846) );
  XNOR U4207 ( .A(n3847), .B(g_input[28]), .Z(n915) );
  NAND U4208 ( .A(n3848), .B(g_input[31]), .Z(n3847) );
  XOR U4209 ( .A(g_input[28]), .B(\_MAC/_MULT/A_[28] ), .Z(n3848) );
  XNOR U4210 ( .A(n3852), .B(n3785), .Z(n3845) );
  NAND U4211 ( .A(n3589), .B(n945), .Z(n3785) );
  IV U4212 ( .A(n3787), .Z(n3852) );
  XOR U4213 ( .A(n3856), .B(n3806), .Z(n3796) );
  XNOR U4214 ( .A(n3793), .B(n3794), .Z(n3806) );
  NAND U4215 ( .A(n3096), .B(n1440), .Z(n3794) );
  XNOR U4216 ( .A(n3792), .B(n3857), .Z(n3793) );
  AND U4217 ( .A(n1373), .B(n3126), .Z(n3857) );
  XNOR U4218 ( .A(n3805), .B(n3795), .Z(n3856) );
  XOR U4219 ( .A(n3800), .B(n3865), .Z(n3801) );
  AND U4220 ( .A(n1248), .B(n3211), .Z(n3865) );
  XNOR U4221 ( .A(n3869), .B(n3802), .Z(n3864) );
  NAND U4222 ( .A(n3168), .B(n1311), .Z(n3802) );
  IV U4223 ( .A(n3804), .Z(n3869) );
  XOR U4224 ( .A(n3809), .B(n3874), .Z(n3810) );
  AND U4225 ( .A(n1476), .B(n3081), .Z(n3874) );
  XNOR U4226 ( .A(n3878), .B(n3811), .Z(n3873) );
  NAND U4227 ( .A(n3055), .B(n1515), .Z(n3811) );
  IV U4228 ( .A(n3813), .Z(n3878) );
  XNOR U4229 ( .A(n3818), .B(n3819), .Z(n3815) );
  NAND U4230 ( .A(n3024), .B(n1593), .Z(n3819) );
  XNOR U4231 ( .A(n3817), .B(n3882), .Z(n3818) );
  AND U4232 ( .A(n1554), .B(n3041), .Z(n3882) );
  XNOR U4233 ( .A(n3836), .B(n3835), .Z(\_MAC/_MULT/MULT/S[3][1][11] ) );
  XOR U4234 ( .A(n3886), .B(n3844), .Z(n3835) );
  XOR U4235 ( .A(n3823), .B(n3888), .Z(n3824) );
  AND U4236 ( .A(n1097), .B(n3379), .Z(n3888) );
  XNOR U4237 ( .A(n3892), .B(n3825), .Z(n3887) );
  NAND U4238 ( .A(n3330), .B(n1145), .Z(n3825) );
  IV U4239 ( .A(n3827), .Z(n3892) );
  XNOR U4240 ( .A(n3832), .B(n3833), .Z(n3829) );
  NAND U4241 ( .A(n3236), .B(n1248), .Z(n3833) );
  XNOR U4242 ( .A(n3831), .B(n3896), .Z(n3832) );
  AND U4243 ( .A(n1195), .B(n3285), .Z(n3896) );
  XNOR U4244 ( .A(n3843), .B(n3834), .Z(n3886) );
  XOR U4245 ( .A(n3903), .B(n3855), .Z(n3843) );
  XNOR U4246 ( .A(n3840), .B(n3841), .Z(n3855) );
  NAND U4247 ( .A(n3454), .B(n1048), .Z(n3841) );
  XNOR U4248 ( .A(n3839), .B(n3904), .Z(n3840) );
  AND U4249 ( .A(n1011), .B(n3516), .Z(n3904) );
  XNOR U4250 ( .A(n3854), .B(n3842), .Z(n3903) );
  XOR U4251 ( .A(n3849), .B(n3912), .Z(n3850) );
  AND U4252 ( .A(n945), .B(n3650), .Z(n3912) );
  XNOR U4253 ( .A(n3913), .B(g_input[27]), .Z(n945) );
  NAND U4254 ( .A(n3914), .B(g_input[31]), .Z(n3913) );
  XOR U4255 ( .A(g_input[27]), .B(\_MAC/_MULT/A_[27] ), .Z(n3914) );
  XNOR U4256 ( .A(n3918), .B(n3851), .Z(n3911) );
  NAND U4257 ( .A(n3589), .B(n976), .Z(n3851) );
  IV U4258 ( .A(n3853), .Z(n3918) );
  XOR U4259 ( .A(n3922), .B(n3872), .Z(n3862) );
  XNOR U4260 ( .A(n3859), .B(n3860), .Z(n3872) );
  NAND U4261 ( .A(n3096), .B(n1476), .Z(n3860) );
  XNOR U4262 ( .A(n3858), .B(n3923), .Z(n3859) );
  AND U4263 ( .A(n1440), .B(n3126), .Z(n3923) );
  XNOR U4264 ( .A(n3871), .B(n3861), .Z(n3922) );
  XOR U4265 ( .A(n3866), .B(n3931), .Z(n3867) );
  AND U4266 ( .A(n1311), .B(n3211), .Z(n3931) );
  XNOR U4267 ( .A(n3935), .B(n3868), .Z(n3930) );
  NAND U4268 ( .A(n3168), .B(n1373), .Z(n3868) );
  IV U4269 ( .A(n3870), .Z(n3935) );
  XOR U4270 ( .A(n3875), .B(n3940), .Z(n3876) );
  AND U4271 ( .A(n1515), .B(n3081), .Z(n3940) );
  XNOR U4272 ( .A(n3944), .B(n3877), .Z(n3939) );
  NAND U4273 ( .A(n3055), .B(n1554), .Z(n3877) );
  IV U4274 ( .A(n3879), .Z(n3944) );
  XNOR U4275 ( .A(n3884), .B(n3885), .Z(n3881) );
  NAND U4276 ( .A(n3024), .B(n1632), .Z(n3885) );
  XNOR U4277 ( .A(n3883), .B(n3948), .Z(n3884) );
  AND U4278 ( .A(n1593), .B(n3041), .Z(n3948) );
  XNOR U4279 ( .A(n3902), .B(n3901), .Z(\_MAC/_MULT/MULT/S[3][1][10] ) );
  XOR U4280 ( .A(n3952), .B(n3910), .Z(n3901) );
  XOR U4281 ( .A(n3889), .B(n3954), .Z(n3890) );
  AND U4282 ( .A(n1145), .B(n3379), .Z(n3954) );
  XNOR U4283 ( .A(n3958), .B(n3891), .Z(n3953) );
  NAND U4284 ( .A(n3330), .B(n1195), .Z(n3891) );
  IV U4285 ( .A(n3893), .Z(n3958) );
  XNOR U4286 ( .A(n3898), .B(n3899), .Z(n3895) );
  NAND U4287 ( .A(n3236), .B(n1311), .Z(n3899) );
  XNOR U4288 ( .A(n3897), .B(n3962), .Z(n3898) );
  AND U4289 ( .A(n1248), .B(n3285), .Z(n3962) );
  XNOR U4290 ( .A(n3909), .B(n3900), .Z(n3952) );
  XOR U4291 ( .A(n3969), .B(n3970), .Z(n2987) );
  XNOR U4292 ( .A(n3971), .B(n3966), .Z(n3969) );
  XOR U4293 ( .A(n3975), .B(n3976), .Z(n2989) );
  XNOR U4294 ( .A(n3977), .B(n3972), .Z(n3975) );
  XOR U4295 ( .A(n3981), .B(n3982), .Z(n2991) );
  XNOR U4296 ( .A(n3983), .B(n3978), .Z(n3981) );
  XOR U4297 ( .A(n3987), .B(n3988), .Z(n2993) );
  XNOR U4298 ( .A(n3989), .B(n3984), .Z(n3987) );
  XOR U4299 ( .A(n3993), .B(n3994), .Z(n2995) );
  XNOR U4300 ( .A(n3995), .B(n3990), .Z(n3993) );
  XOR U4301 ( .A(n3999), .B(n4000), .Z(n2997) );
  XNOR U4302 ( .A(n4001), .B(n3996), .Z(n3999) );
  XOR U4303 ( .A(n4005), .B(n4006), .Z(n2999) );
  XNOR U4304 ( .A(n4007), .B(n4002), .Z(n4005) );
  XOR U4305 ( .A(n4011), .B(n4012), .Z(n3030) );
  XNOR U4306 ( .A(n4013), .B(n4008), .Z(n4011) );
  XOR U4307 ( .A(n4017), .B(n4018), .Z(n3375) );
  XNOR U4308 ( .A(n4019), .B(n4014), .Z(n4017) );
  XOR U4309 ( .A(n4023), .B(n3921), .Z(n3909) );
  XNOR U4310 ( .A(n3906), .B(n3907), .Z(n3921) );
  NAND U4311 ( .A(n3454), .B(n1097), .Z(n3907) );
  XNOR U4312 ( .A(n3905), .B(n4024), .Z(n3906) );
  AND U4313 ( .A(n1048), .B(n3516), .Z(n4024) );
  XNOR U4314 ( .A(n3920), .B(n3908), .Z(n4023) );
  XOR U4315 ( .A(n3955), .B(n4030), .Z(n3956) );
  AND U4316 ( .A(n1195), .B(n3379), .Z(n4030) );
  XNOR U4317 ( .A(n4034), .B(n3957), .Z(n4029) );
  NAND U4318 ( .A(n3330), .B(n1248), .Z(n3957) );
  IV U4319 ( .A(n3959), .Z(n4034) );
  XNOR U4320 ( .A(n3964), .B(n3965), .Z(n3961) );
  NAND U4321 ( .A(n3236), .B(n1373), .Z(n3965) );
  XNOR U4322 ( .A(n3963), .B(n4038), .Z(n3964) );
  AND U4323 ( .A(n1311), .B(n3285), .Z(n4038) );
  XOR U4324 ( .A(n4042), .B(n4043), .Z(n3971) );
  XNOR U4325 ( .A(n4044), .B(n4028), .Z(n4042) );
  XOR U4326 ( .A(n4031), .B(n4047), .Z(n4032) );
  AND U4327 ( .A(n1248), .B(n3379), .Z(n4047) );
  XNOR U4328 ( .A(n4051), .B(n4033), .Z(n4046) );
  NAND U4329 ( .A(n3330), .B(n1311), .Z(n4033) );
  IV U4330 ( .A(n4035), .Z(n4051) );
  XNOR U4331 ( .A(n4040), .B(n4041), .Z(n4037) );
  NAND U4332 ( .A(n3236), .B(n1440), .Z(n4041) );
  XNOR U4333 ( .A(n4039), .B(n4055), .Z(n4040) );
  AND U4334 ( .A(n1373), .B(n3285), .Z(n4055) );
  XOR U4335 ( .A(n4059), .B(n4060), .Z(n3977) );
  XNOR U4336 ( .A(n4061), .B(n4045), .Z(n4059) );
  XOR U4337 ( .A(n4048), .B(n4064), .Z(n4049) );
  AND U4338 ( .A(n1311), .B(n3379), .Z(n4064) );
  XNOR U4339 ( .A(n4068), .B(n4050), .Z(n4063) );
  NAND U4340 ( .A(n3330), .B(n1373), .Z(n4050) );
  IV U4341 ( .A(n4052), .Z(n4068) );
  XNOR U4342 ( .A(n4057), .B(n4058), .Z(n4054) );
  NAND U4343 ( .A(n3236), .B(n1476), .Z(n4058) );
  XNOR U4344 ( .A(n4056), .B(n4072), .Z(n4057) );
  AND U4345 ( .A(n1440), .B(n3285), .Z(n4072) );
  XOR U4346 ( .A(n4076), .B(n4077), .Z(n3983) );
  XNOR U4347 ( .A(n4078), .B(n4062), .Z(n4076) );
  XOR U4348 ( .A(n4065), .B(n4081), .Z(n4066) );
  AND U4349 ( .A(n1373), .B(n3379), .Z(n4081) );
  XNOR U4350 ( .A(n4085), .B(n4067), .Z(n4080) );
  NAND U4351 ( .A(n3330), .B(n1440), .Z(n4067) );
  IV U4352 ( .A(n4069), .Z(n4085) );
  XNOR U4353 ( .A(n4074), .B(n4075), .Z(n4071) );
  NAND U4354 ( .A(n3236), .B(n1515), .Z(n4075) );
  XNOR U4355 ( .A(n4073), .B(n4089), .Z(n4074) );
  AND U4356 ( .A(n1476), .B(n3285), .Z(n4089) );
  XOR U4357 ( .A(n4093), .B(n4094), .Z(n3989) );
  XNOR U4358 ( .A(n4095), .B(n4079), .Z(n4093) );
  XOR U4359 ( .A(n4082), .B(n4098), .Z(n4083) );
  AND U4360 ( .A(n1440), .B(n3379), .Z(n4098) );
  XNOR U4361 ( .A(n4102), .B(n4084), .Z(n4097) );
  NAND U4362 ( .A(n3330), .B(n1476), .Z(n4084) );
  IV U4363 ( .A(n4086), .Z(n4102) );
  XNOR U4364 ( .A(n4091), .B(n4092), .Z(n4088) );
  NAND U4365 ( .A(n3236), .B(n1554), .Z(n4092) );
  XNOR U4366 ( .A(n4090), .B(n4106), .Z(n4091) );
  AND U4367 ( .A(n1515), .B(n3285), .Z(n4106) );
  XOR U4368 ( .A(n4110), .B(n4111), .Z(n3995) );
  XNOR U4369 ( .A(n4112), .B(n4096), .Z(n4110) );
  XOR U4370 ( .A(n4099), .B(n4115), .Z(n4100) );
  AND U4371 ( .A(n1476), .B(n3379), .Z(n4115) );
  XNOR U4372 ( .A(n4119), .B(n4101), .Z(n4114) );
  NAND U4373 ( .A(n3330), .B(n1515), .Z(n4101) );
  IV U4374 ( .A(n4103), .Z(n4119) );
  XNOR U4375 ( .A(n4108), .B(n4109), .Z(n4105) );
  NAND U4376 ( .A(n3236), .B(n1593), .Z(n4109) );
  XNOR U4377 ( .A(n4107), .B(n4123), .Z(n4108) );
  AND U4378 ( .A(n1554), .B(n3285), .Z(n4123) );
  XOR U4379 ( .A(n4127), .B(n4128), .Z(n4001) );
  XNOR U4380 ( .A(n4129), .B(n4113), .Z(n4127) );
  XOR U4381 ( .A(n4116), .B(n4132), .Z(n4117) );
  AND U4382 ( .A(n1515), .B(n3379), .Z(n4132) );
  XNOR U4383 ( .A(n4136), .B(n4118), .Z(n4131) );
  NAND U4384 ( .A(n3330), .B(n1554), .Z(n4118) );
  IV U4385 ( .A(n4120), .Z(n4136) );
  XNOR U4386 ( .A(n4125), .B(n4126), .Z(n4122) );
  NAND U4387 ( .A(n3236), .B(n1632), .Z(n4126) );
  XNOR U4388 ( .A(n4124), .B(n4140), .Z(n4125) );
  AND U4389 ( .A(n1593), .B(n3285), .Z(n4140) );
  XOR U4390 ( .A(n4144), .B(n4145), .Z(n4007) );
  XNOR U4391 ( .A(n4146), .B(n4130), .Z(n4144) );
  XOR U4392 ( .A(n4133), .B(n4149), .Z(n4134) );
  AND U4393 ( .A(n1554), .B(n3379), .Z(n4149) );
  XNOR U4394 ( .A(n4153), .B(n4135), .Z(n4148) );
  NAND U4395 ( .A(n3330), .B(n1593), .Z(n4135) );
  IV U4396 ( .A(n4137), .Z(n4153) );
  XNOR U4397 ( .A(n4142), .B(n4143), .Z(n4139) );
  NAND U4398 ( .A(n3236), .B(n1671), .Z(n4143) );
  XNOR U4399 ( .A(n4141), .B(n4157), .Z(n4142) );
  AND U4400 ( .A(n1632), .B(n3285), .Z(n4157) );
  XOR U4401 ( .A(n4161), .B(n4162), .Z(n4013) );
  XNOR U4402 ( .A(n4163), .B(n4147), .Z(n4161) );
  XOR U4403 ( .A(n4150), .B(n4166), .Z(n4151) );
  AND U4404 ( .A(n1593), .B(n3379), .Z(n4166) );
  XNOR U4405 ( .A(n4170), .B(n4152), .Z(n4165) );
  NAND U4406 ( .A(n3330), .B(n1632), .Z(n4152) );
  IV U4407 ( .A(n4154), .Z(n4170) );
  XNOR U4408 ( .A(n4159), .B(n4160), .Z(n4156) );
  NAND U4409 ( .A(n3236), .B(n1710), .Z(n4160) );
  XNOR U4410 ( .A(n4158), .B(n4174), .Z(n4159) );
  AND U4411 ( .A(n1671), .B(n3285), .Z(n4174) );
  XOR U4412 ( .A(n4178), .B(n4179), .Z(n4019) );
  XNOR U4413 ( .A(n4180), .B(n4164), .Z(n4178) );
  XOR U4414 ( .A(n3915), .B(n4185), .Z(n3916) );
  AND U4415 ( .A(n976), .B(n3650), .Z(n4185) );
  XNOR U4416 ( .A(n4186), .B(g_input[26]), .Z(n976) );
  NAND U4417 ( .A(n4187), .B(g_input[31]), .Z(n4186) );
  XOR U4418 ( .A(g_input[26]), .B(\_MAC/_MULT/A_[26] ), .Z(n4187) );
  XNOR U4419 ( .A(n4191), .B(n3917), .Z(n4184) );
  NAND U4420 ( .A(n3589), .B(n1011), .Z(n3917) );
  IV U4421 ( .A(n3919), .Z(n4191) );
  XNOR U4422 ( .A(n4026), .B(n4027), .Z(n4043) );
  NAND U4423 ( .A(n3454), .B(n1145), .Z(n4027) );
  XNOR U4424 ( .A(n4025), .B(n4193), .Z(n4026) );
  AND U4425 ( .A(n1097), .B(n3516), .Z(n4193) );
  XOR U4426 ( .A(n4188), .B(n4198), .Z(n4189) );
  AND U4427 ( .A(n1011), .B(n3650), .Z(n4198) );
  XNOR U4428 ( .A(n4199), .B(g_input[25]), .Z(n1011) );
  NAND U4429 ( .A(n4200), .B(g_input[31]), .Z(n4199) );
  XOR U4430 ( .A(g_input[25]), .B(\_MAC/_MULT/A_[25] ), .Z(n4200) );
  XNOR U4431 ( .A(n4204), .B(n4190), .Z(n4197) );
  NAND U4432 ( .A(n3589), .B(n1048), .Z(n4190) );
  IV U4433 ( .A(n4192), .Z(n4204) );
  XNOR U4434 ( .A(n4195), .B(n4196), .Z(n4060) );
  NAND U4435 ( .A(n3454), .B(n1195), .Z(n4196) );
  XNOR U4436 ( .A(n4194), .B(n4206), .Z(n4195) );
  AND U4437 ( .A(n1145), .B(n3516), .Z(n4206) );
  XOR U4438 ( .A(n4201), .B(n4211), .Z(n4202) );
  AND U4439 ( .A(n1048), .B(n3650), .Z(n4211) );
  XNOR U4440 ( .A(n4212), .B(g_input[24]), .Z(n1048) );
  NAND U4441 ( .A(n4213), .B(g_input[31]), .Z(n4212) );
  XOR U4442 ( .A(g_input[24]), .B(\_MAC/_MULT/A_[24] ), .Z(n4213) );
  XNOR U4443 ( .A(n4217), .B(n4203), .Z(n4210) );
  NAND U4444 ( .A(n3589), .B(n1097), .Z(n4203) );
  IV U4445 ( .A(n4205), .Z(n4217) );
  XNOR U4446 ( .A(n4208), .B(n4209), .Z(n4077) );
  NAND U4447 ( .A(n3454), .B(n1248), .Z(n4209) );
  XNOR U4448 ( .A(n4207), .B(n4219), .Z(n4208) );
  AND U4449 ( .A(n1195), .B(n3516), .Z(n4219) );
  XOR U4450 ( .A(n4214), .B(n4224), .Z(n4215) );
  AND U4451 ( .A(n1097), .B(n3650), .Z(n4224) );
  XNOR U4452 ( .A(n4225), .B(g_input[23]), .Z(n1097) );
  NAND U4453 ( .A(n4226), .B(g_input[31]), .Z(n4225) );
  XOR U4454 ( .A(g_input[23]), .B(\_MAC/_MULT/A_[23] ), .Z(n4226) );
  XNOR U4455 ( .A(n4230), .B(n4216), .Z(n4223) );
  NAND U4456 ( .A(n3589), .B(n1145), .Z(n4216) );
  IV U4457 ( .A(n4218), .Z(n4230) );
  XNOR U4458 ( .A(n4221), .B(n4222), .Z(n4094) );
  NAND U4459 ( .A(n3454), .B(n1311), .Z(n4222) );
  XNOR U4460 ( .A(n4220), .B(n4232), .Z(n4221) );
  AND U4461 ( .A(n1248), .B(n3516), .Z(n4232) );
  XOR U4462 ( .A(n4227), .B(n4237), .Z(n4228) );
  AND U4463 ( .A(n1145), .B(n3650), .Z(n4237) );
  XNOR U4464 ( .A(n4238), .B(g_input[22]), .Z(n1145) );
  NAND U4465 ( .A(n4239), .B(g_input[31]), .Z(n4238) );
  XOR U4466 ( .A(g_input[22]), .B(\_MAC/_MULT/A_[22] ), .Z(n4239) );
  XNOR U4467 ( .A(n4243), .B(n4229), .Z(n4236) );
  NAND U4468 ( .A(n3589), .B(n1195), .Z(n4229) );
  IV U4469 ( .A(n4231), .Z(n4243) );
  XNOR U4470 ( .A(n4234), .B(n4235), .Z(n4111) );
  NAND U4471 ( .A(n3454), .B(n1373), .Z(n4235) );
  XNOR U4472 ( .A(n4233), .B(n4245), .Z(n4234) );
  AND U4473 ( .A(n1311), .B(n3516), .Z(n4245) );
  XOR U4474 ( .A(n4240), .B(n4250), .Z(n4241) );
  AND U4475 ( .A(n1195), .B(n3650), .Z(n4250) );
  XNOR U4476 ( .A(n4251), .B(g_input[21]), .Z(n1195) );
  NAND U4477 ( .A(n4252), .B(g_input[31]), .Z(n4251) );
  XOR U4478 ( .A(g_input[21]), .B(\_MAC/_MULT/A_[21] ), .Z(n4252) );
  XNOR U4479 ( .A(n4256), .B(n4242), .Z(n4249) );
  NAND U4480 ( .A(n3589), .B(n1248), .Z(n4242) );
  IV U4481 ( .A(n4244), .Z(n4256) );
  XNOR U4482 ( .A(n4247), .B(n4248), .Z(n4128) );
  NAND U4483 ( .A(n3454), .B(n1440), .Z(n4248) );
  XNOR U4484 ( .A(n4246), .B(n4258), .Z(n4247) );
  AND U4485 ( .A(n1373), .B(n3516), .Z(n4258) );
  XOR U4486 ( .A(n4253), .B(n4263), .Z(n4254) );
  AND U4487 ( .A(n1248), .B(n3650), .Z(n4263) );
  XNOR U4488 ( .A(n4264), .B(g_input[20]), .Z(n1248) );
  NAND U4489 ( .A(n4265), .B(g_input[31]), .Z(n4264) );
  XOR U4490 ( .A(g_input[20]), .B(\_MAC/_MULT/A_[20] ), .Z(n4265) );
  XNOR U4491 ( .A(n4269), .B(n4255), .Z(n4262) );
  NAND U4492 ( .A(n3589), .B(n1311), .Z(n4255) );
  IV U4493 ( .A(n4257), .Z(n4269) );
  XNOR U4494 ( .A(n4260), .B(n4261), .Z(n4145) );
  NAND U4495 ( .A(n3454), .B(n1476), .Z(n4261) );
  XNOR U4496 ( .A(n4259), .B(n4271), .Z(n4260) );
  AND U4497 ( .A(n1440), .B(n3516), .Z(n4271) );
  XOR U4498 ( .A(n4266), .B(n4276), .Z(n4267) );
  AND U4499 ( .A(n1311), .B(n3650), .Z(n4276) );
  XNOR U4500 ( .A(n4277), .B(g_input[19]), .Z(n1311) );
  NAND U4501 ( .A(n4278), .B(g_input[31]), .Z(n4277) );
  XOR U4502 ( .A(g_input[19]), .B(\_MAC/_MULT/A_[19] ), .Z(n4278) );
  XNOR U4503 ( .A(n4282), .B(n4268), .Z(n4275) );
  NAND U4504 ( .A(n3589), .B(n1373), .Z(n4268) );
  IV U4505 ( .A(n4270), .Z(n4282) );
  XNOR U4506 ( .A(n4273), .B(n4274), .Z(n4162) );
  NAND U4507 ( .A(n3454), .B(n1515), .Z(n4274) );
  XNOR U4508 ( .A(n4272), .B(n4284), .Z(n4273) );
  AND U4509 ( .A(n1476), .B(n3516), .Z(n4284) );
  XOR U4510 ( .A(n4279), .B(n4289), .Z(n4280) );
  AND U4511 ( .A(n1373), .B(n3650), .Z(n4289) );
  XNOR U4512 ( .A(n4293), .B(n4281), .Z(n4288) );
  NAND U4513 ( .A(n3589), .B(n1440), .Z(n4281) );
  IV U4514 ( .A(n4283), .Z(n4293) );
  XNOR U4515 ( .A(n4286), .B(n4287), .Z(n4179) );
  NAND U4516 ( .A(n3454), .B(n1554), .Z(n4287) );
  XNOR U4517 ( .A(n4285), .B(n4295), .Z(n4286) );
  AND U4518 ( .A(n1515), .B(n3516), .Z(n4295) );
  XOR U4519 ( .A(n4290), .B(n4300), .Z(n4291) );
  AND U4520 ( .A(n1440), .B(n3650), .Z(n4300) );
  XNOR U4521 ( .A(n4304), .B(n4292), .Z(n4299) );
  NAND U4522 ( .A(n3589), .B(n1476), .Z(n4292) );
  IV U4523 ( .A(n4294), .Z(n4304) );
  XOR U4524 ( .A(n4308), .B(n3938), .Z(n3928) );
  XNOR U4525 ( .A(n3925), .B(n3926), .Z(n3938) );
  NAND U4526 ( .A(n3096), .B(n1515), .Z(n3926) );
  XNOR U4527 ( .A(n3924), .B(n4309), .Z(n3925) );
  AND U4528 ( .A(n1476), .B(n3126), .Z(n4309) );
  XNOR U4529 ( .A(n3937), .B(n3927), .Z(n4308) );
  XOR U4530 ( .A(n4314), .B(n4315), .Z(n3968) );
  XNOR U4531 ( .A(n4316), .B(n4313), .Z(n4314) );
  XOR U4532 ( .A(n4320), .B(n4321), .Z(n3974) );
  XNOR U4533 ( .A(n4322), .B(n4319), .Z(n4320) );
  XOR U4534 ( .A(n4326), .B(n4327), .Z(n3980) );
  XNOR U4535 ( .A(n4328), .B(n4325), .Z(n4326) );
  XOR U4536 ( .A(n4332), .B(n4333), .Z(n3986) );
  XNOR U4537 ( .A(n4334), .B(n4331), .Z(n4332) );
  XOR U4538 ( .A(n4338), .B(n4339), .Z(n3992) );
  XNOR U4539 ( .A(n4340), .B(n4337), .Z(n4338) );
  XOR U4540 ( .A(n4344), .B(n4345), .Z(n3998) );
  XNOR U4541 ( .A(n4346), .B(n4343), .Z(n4344) );
  XOR U4542 ( .A(n4350), .B(n4351), .Z(n4004) );
  XNOR U4543 ( .A(n4352), .B(n4349), .Z(n4350) );
  XOR U4544 ( .A(n4356), .B(n4357), .Z(n4010) );
  XNOR U4545 ( .A(n4358), .B(n4355), .Z(n4356) );
  XOR U4546 ( .A(n4362), .B(n4363), .Z(n4016) );
  XNOR U4547 ( .A(n4364), .B(n4361), .Z(n4362) );
  XOR U4548 ( .A(n3932), .B(n4371), .Z(n3933) );
  AND U4549 ( .A(n1373), .B(n3211), .Z(n4371) );
  XNOR U4550 ( .A(n4372), .B(g_input[18]), .Z(n1373) );
  NAND U4551 ( .A(n4373), .B(g_input[31]), .Z(n4372) );
  XOR U4552 ( .A(g_input[18]), .B(\_MAC/_MULT/A_[18] ), .Z(n4373) );
  XNOR U4553 ( .A(n4377), .B(n3934), .Z(n4370) );
  NAND U4554 ( .A(n3168), .B(n1440), .Z(n3934) );
  IV U4555 ( .A(n3936), .Z(n4377) );
  XNOR U4556 ( .A(n4311), .B(n4312), .Z(n4315) );
  NAND U4557 ( .A(n3096), .B(n1554), .Z(n4312) );
  XNOR U4558 ( .A(n4310), .B(n4379), .Z(n4311) );
  AND U4559 ( .A(n1515), .B(n3126), .Z(n4379) );
  XOR U4560 ( .A(n4374), .B(n4384), .Z(n4375) );
  AND U4561 ( .A(n1440), .B(n3211), .Z(n4384) );
  XNOR U4562 ( .A(n4385), .B(g_input[17]), .Z(n1440) );
  NAND U4563 ( .A(n4386), .B(g_input[31]), .Z(n4385) );
  XOR U4564 ( .A(g_input[17]), .B(\_MAC/_MULT/A_[17] ), .Z(n4386) );
  XNOR U4565 ( .A(n4390), .B(n4376), .Z(n4383) );
  NAND U4566 ( .A(n3168), .B(n1476), .Z(n4376) );
  IV U4567 ( .A(n4378), .Z(n4390) );
  XNOR U4568 ( .A(n4381), .B(n4382), .Z(n4321) );
  NAND U4569 ( .A(n3096), .B(n1593), .Z(n4382) );
  XNOR U4570 ( .A(n4380), .B(n4392), .Z(n4381) );
  AND U4571 ( .A(n1554), .B(n3126), .Z(n4392) );
  XOR U4572 ( .A(n4387), .B(n4397), .Z(n4388) );
  AND U4573 ( .A(n1476), .B(n3211), .Z(n4397) );
  XNOR U4574 ( .A(n4401), .B(n4389), .Z(n4396) );
  NAND U4575 ( .A(n3168), .B(n1515), .Z(n4389) );
  IV U4576 ( .A(n4391), .Z(n4401) );
  XNOR U4577 ( .A(n4394), .B(n4395), .Z(n4327) );
  NAND U4578 ( .A(n3096), .B(n1632), .Z(n4395) );
  XNOR U4579 ( .A(n4393), .B(n4403), .Z(n4394) );
  AND U4580 ( .A(n1593), .B(n3126), .Z(n4403) );
  XOR U4581 ( .A(n4398), .B(n4408), .Z(n4399) );
  AND U4582 ( .A(n1515), .B(n3211), .Z(n4408) );
  XNOR U4583 ( .A(n4412), .B(n4400), .Z(n4407) );
  NAND U4584 ( .A(n3168), .B(n1554), .Z(n4400) );
  IV U4585 ( .A(n4402), .Z(n4412) );
  XNOR U4586 ( .A(n4405), .B(n4406), .Z(n4333) );
  NAND U4587 ( .A(n3096), .B(n1671), .Z(n4406) );
  XNOR U4588 ( .A(n4404), .B(n4414), .Z(n4405) );
  AND U4589 ( .A(n1632), .B(n3126), .Z(n4414) );
  XOR U4590 ( .A(n4409), .B(n4419), .Z(n4410) );
  AND U4591 ( .A(n1554), .B(n3211), .Z(n4419) );
  XNOR U4592 ( .A(n4423), .B(n4411), .Z(n4418) );
  NAND U4593 ( .A(n3168), .B(n1593), .Z(n4411) );
  IV U4594 ( .A(n4413), .Z(n4423) );
  XNOR U4595 ( .A(n4416), .B(n4417), .Z(n4339) );
  NAND U4596 ( .A(n3096), .B(n1710), .Z(n4417) );
  XNOR U4597 ( .A(n4415), .B(n4425), .Z(n4416) );
  AND U4598 ( .A(n1671), .B(n3126), .Z(n4425) );
  XOR U4599 ( .A(n4420), .B(n4430), .Z(n4421) );
  AND U4600 ( .A(n1593), .B(n3211), .Z(n4430) );
  XNOR U4601 ( .A(n4434), .B(n4422), .Z(n4429) );
  NAND U4602 ( .A(n3168), .B(n1632), .Z(n4422) );
  IV U4603 ( .A(n4424), .Z(n4434) );
  XNOR U4604 ( .A(n4427), .B(n4428), .Z(n4345) );
  NAND U4605 ( .A(n3096), .B(n1749), .Z(n4428) );
  XNOR U4606 ( .A(n4426), .B(n4436), .Z(n4427) );
  AND U4607 ( .A(n1710), .B(n3126), .Z(n4436) );
  XOR U4608 ( .A(n4431), .B(n4441), .Z(n4432) );
  AND U4609 ( .A(n1632), .B(n3211), .Z(n4441) );
  XNOR U4610 ( .A(n4445), .B(n4433), .Z(n4440) );
  NAND U4611 ( .A(n3168), .B(n1671), .Z(n4433) );
  IV U4612 ( .A(n4435), .Z(n4445) );
  XNOR U4613 ( .A(n4438), .B(n4439), .Z(n4351) );
  NAND U4614 ( .A(n3096), .B(n1788), .Z(n4439) );
  XNOR U4615 ( .A(n4437), .B(n4447), .Z(n4438) );
  AND U4616 ( .A(n1749), .B(n3126), .Z(n4447) );
  XOR U4617 ( .A(n4442), .B(n4452), .Z(n4443) );
  AND U4618 ( .A(n1671), .B(n3211), .Z(n4452) );
  XNOR U4619 ( .A(n4456), .B(n4444), .Z(n4451) );
  NAND U4620 ( .A(n3168), .B(n1710), .Z(n4444) );
  IV U4621 ( .A(n4446), .Z(n4456) );
  XNOR U4622 ( .A(n4449), .B(n4450), .Z(n4357) );
  NAND U4623 ( .A(n3096), .B(n1827), .Z(n4450) );
  XNOR U4624 ( .A(n4448), .B(n4458), .Z(n4449) );
  AND U4625 ( .A(n1788), .B(n3126), .Z(n4458) );
  XOR U4626 ( .A(n4453), .B(n4463), .Z(n4454) );
  AND U4627 ( .A(n1710), .B(n3211), .Z(n4463) );
  XOR U4628 ( .A(n4464), .B(n4465), .Z(n4453) );
  AND U4629 ( .A(n4466), .B(n4467), .Z(n4465) );
  XNOR U4630 ( .A(n4468), .B(n4464), .Z(n4466) );
  XNOR U4631 ( .A(n4469), .B(n4455), .Z(n4462) );
  NAND U4632 ( .A(n3168), .B(n1749), .Z(n4455) );
  IV U4633 ( .A(n4457), .Z(n4469) );
  XNOR U4634 ( .A(n4460), .B(n4461), .Z(n4363) );
  NAND U4635 ( .A(n3096), .B(n1868), .Z(n4461) );
  XNOR U4636 ( .A(n4459), .B(n4471), .Z(n4460) );
  AND U4637 ( .A(n1827), .B(n3126), .Z(n4471) );
  XOR U4638 ( .A(n4464), .B(n4476), .Z(n4467) );
  AND U4639 ( .A(n1749), .B(n3211), .Z(n4476) );
  XNOR U4640 ( .A(n4480), .B(n4468), .Z(n4475) );
  NAND U4641 ( .A(n3168), .B(n1788), .Z(n4468) );
  IV U4642 ( .A(n4470), .Z(n4480) );
  XOR U4643 ( .A(n3941), .B(n4485), .Z(n3942) );
  AND U4644 ( .A(n1554), .B(n3081), .Z(n4485) );
  XNOR U4645 ( .A(n4489), .B(n3943), .Z(n4484) );
  NAND U4646 ( .A(n3055), .B(n1593), .Z(n3943) );
  IV U4647 ( .A(n3945), .Z(n4489) );
  XOR U4648 ( .A(n4486), .B(n4492), .Z(n4487) );
  AND U4649 ( .A(n1593), .B(n3081), .Z(n4492) );
  XNOR U4650 ( .A(n4496), .B(n4488), .Z(n4491) );
  NAND U4651 ( .A(n3055), .B(n1632), .Z(n4488) );
  IV U4652 ( .A(n4490), .Z(n4496) );
  XNOR U4653 ( .A(n4497), .B(n4498), .Z(n4317) );
  XOR U4654 ( .A(n4499), .B(n4500), .Z(n4490) );
  AND U4655 ( .A(n4501), .B(n4324), .Z(n4500) );
  XOR U4656 ( .A(n4493), .B(n4503), .Z(n4494) );
  AND U4657 ( .A(n1632), .B(n3081), .Z(n4503) );
  XNOR U4658 ( .A(n4507), .B(n4495), .Z(n4502) );
  NAND U4659 ( .A(n3055), .B(n1671), .Z(n4495) );
  IV U4660 ( .A(n4499), .Z(n4507) );
  XNOR U4661 ( .A(n4499), .B(n4323), .Z(n4501) );
  XNOR U4662 ( .A(n4508), .B(n4509), .Z(n4323) );
  XOR U4663 ( .A(n4504), .B(n4512), .Z(n4505) );
  AND U4664 ( .A(n1671), .B(n3081), .Z(n4512) );
  XNOR U4665 ( .A(n4516), .B(n4506), .Z(n4511) );
  NAND U4666 ( .A(n3055), .B(n1710), .Z(n4506) );
  IV U4667 ( .A(n4510), .Z(n4516) );
  XNOR U4668 ( .A(n4517), .B(n4518), .Z(n4329) );
  XOR U4669 ( .A(n4513), .B(n4521), .Z(n4514) );
  AND U4670 ( .A(n1710), .B(n3081), .Z(n4521) );
  XNOR U4671 ( .A(n4525), .B(n4515), .Z(n4520) );
  NAND U4672 ( .A(n3055), .B(n1749), .Z(n4515) );
  IV U4673 ( .A(n4519), .Z(n4525) );
  XNOR U4674 ( .A(n4526), .B(n4527), .Z(n4335) );
  XOR U4675 ( .A(n4522), .B(n4530), .Z(n4523) );
  AND U4676 ( .A(n1749), .B(n3081), .Z(n4530) );
  XNOR U4677 ( .A(n4534), .B(n4524), .Z(n4529) );
  NAND U4678 ( .A(n3055), .B(n1788), .Z(n4524) );
  IV U4679 ( .A(n4528), .Z(n4534) );
  XNOR U4680 ( .A(n4535), .B(n4536), .Z(n4341) );
  XOR U4681 ( .A(n4531), .B(n4539), .Z(n4532) );
  AND U4682 ( .A(n1788), .B(n3081), .Z(n4539) );
  XNOR U4683 ( .A(n4543), .B(n4533), .Z(n4538) );
  NAND U4684 ( .A(n3055), .B(n1827), .Z(n4533) );
  IV U4685 ( .A(n4537), .Z(n4543) );
  XNOR U4686 ( .A(n4544), .B(n4545), .Z(n4347) );
  XOR U4687 ( .A(n4546), .B(n4547), .Z(n4537) );
  AND U4688 ( .A(n4548), .B(n4354), .Z(n4547) );
  XOR U4689 ( .A(n4540), .B(n4550), .Z(n4541) );
  AND U4690 ( .A(n1827), .B(n3081), .Z(n4550) );
  XNOR U4691 ( .A(n4554), .B(n4542), .Z(n4549) );
  NAND U4692 ( .A(n3055), .B(n1868), .Z(n4542) );
  IV U4693 ( .A(n4546), .Z(n4554) );
  XNOR U4694 ( .A(n4546), .B(n4353), .Z(n4548) );
  XNOR U4695 ( .A(n4555), .B(n4556), .Z(n4353) );
  XOR U4696 ( .A(n4551), .B(n4559), .Z(n4552) );
  AND U4697 ( .A(n1868), .B(n3081), .Z(n4559) );
  XNOR U4698 ( .A(n4563), .B(n4553), .Z(n4558) );
  NAND U4699 ( .A(n3055), .B(n1907), .Z(n4553) );
  IV U4700 ( .A(n4557), .Z(n4563) );
  XNOR U4701 ( .A(n4564), .B(n4565), .Z(n4359) );
  XOR U4702 ( .A(n4560), .B(n4568), .Z(n4561) );
  AND U4703 ( .A(n1907), .B(n3081), .Z(n4568) );
  XNOR U4704 ( .A(n4572), .B(n4562), .Z(n4567) );
  NAND U4705 ( .A(n3055), .B(n1946), .Z(n4562) );
  IV U4706 ( .A(n4566), .Z(n4572) );
  XNOR U4707 ( .A(n4573), .B(n4574), .Z(n4365) );
  XNOR U4708 ( .A(n3950), .B(n3951), .Z(n3947) );
  NAND U4709 ( .A(n3024), .B(n1671), .Z(n3951) );
  XNOR U4710 ( .A(n3949), .B(n4578), .Z(n3950) );
  AND U4711 ( .A(n1632), .B(n3041), .Z(n4578) );
  XNOR U4712 ( .A(n4579), .B(n4580), .Z(n4497) );
  AND U4713 ( .A(n1671), .B(n3041), .Z(n4580) );
  NAND U4714 ( .A(n3024), .B(n1710), .Z(n4498) );
  XNOR U4715 ( .A(n4581), .B(n4582), .Z(n4508) );
  AND U4716 ( .A(n1710), .B(n3041), .Z(n4582) );
  NAND U4717 ( .A(n3024), .B(n1749), .Z(n4509) );
  XNOR U4718 ( .A(n4583), .B(n4584), .Z(n4517) );
  AND U4719 ( .A(n1749), .B(n3041), .Z(n4584) );
  NAND U4720 ( .A(n3024), .B(n1788), .Z(n4518) );
  XNOR U4721 ( .A(n4585), .B(n4586), .Z(n4526) );
  AND U4722 ( .A(n1788), .B(n3041), .Z(n4586) );
  NAND U4723 ( .A(n3024), .B(n1827), .Z(n4527) );
  XNOR U4724 ( .A(n4587), .B(n4588), .Z(n4535) );
  AND U4725 ( .A(n1827), .B(n3041), .Z(n4588) );
  NAND U4726 ( .A(n3024), .B(n1868), .Z(n4536) );
  XNOR U4727 ( .A(n4589), .B(n4590), .Z(n4544) );
  AND U4728 ( .A(n1868), .B(n3041), .Z(n4590) );
  NAND U4729 ( .A(n3024), .B(n1907), .Z(n4545) );
  XNOR U4730 ( .A(n4591), .B(n4592), .Z(n4555) );
  AND U4731 ( .A(n1907), .B(n3041), .Z(n4592) );
  NAND U4732 ( .A(n3024), .B(n1946), .Z(n4556) );
  XNOR U4733 ( .A(n4593), .B(n4594), .Z(n4564) );
  AND U4734 ( .A(n1946), .B(n3041), .Z(n4594) );
  NAND U4735 ( .A(n3024), .B(n1987), .Z(n4565) );
  XNOR U4736 ( .A(n4595), .B(n4596), .Z(n4573) );
  AND U4737 ( .A(n1987), .B(n3041), .Z(n4596) );
  NAND U4738 ( .A(n3024), .B(n2028), .Z(n4574) );
  XNOR U4739 ( .A(n4022), .B(n4021), .Z(\_MAC/_MULT/MULT/S[3][1][0] ) );
  XOR U4740 ( .A(n4600), .B(n4183), .Z(n4021) );
  XOR U4741 ( .A(n4167), .B(n4602), .Z(n4168) );
  AND U4742 ( .A(n1632), .B(n3379), .Z(n4602) );
  XNOR U4743 ( .A(n4606), .B(n4169), .Z(n4601) );
  NAND U4744 ( .A(n3330), .B(n1671), .Z(n4169) );
  IV U4745 ( .A(n4171), .Z(n4606) );
  XNOR U4746 ( .A(n4176), .B(n4177), .Z(n4173) );
  NAND U4747 ( .A(n3236), .B(n1749), .Z(n4177) );
  XNOR U4748 ( .A(n4175), .B(n4610), .Z(n4176) );
  AND U4749 ( .A(n1710), .B(n3285), .Z(n4610) );
  XNOR U4750 ( .A(n4182), .B(n4020), .Z(n4600) );
  XOR U4751 ( .A(n4614), .B(n4615), .Z(n4020) );
  XOR U4752 ( .A(n4616), .B(n4307), .Z(n4182) );
  XNOR U4753 ( .A(n4297), .B(n4298), .Z(n4307) );
  NAND U4754 ( .A(n3454), .B(n1593), .Z(n4298) );
  XNOR U4755 ( .A(n4296), .B(n4617), .Z(n4297) );
  AND U4756 ( .A(n1554), .B(n3516), .Z(n4617) );
  XNOR U4757 ( .A(n4306), .B(n4181), .Z(n4616) );
  XOR U4758 ( .A(n4621), .B(n4622), .Z(n4181) );
  AND U4759 ( .A(n4623), .B(n4624), .Z(n4622) );
  XOR U4760 ( .A(n4625), .B(n4626), .Z(n4624) );
  XOR U4761 ( .A(n4621), .B(n4627), .Z(n4626) );
  XOR U4762 ( .A(n4608), .B(n4628), .Z(n4623) );
  XOR U4763 ( .A(n4621), .B(n4609), .Z(n4628) );
  NAND U4764 ( .A(n3236), .B(n1788), .Z(n4613) );
  XOR U4765 ( .A(n4611), .B(n4629), .Z(n4612) );
  AND U4766 ( .A(n1749), .B(n3285), .Z(n4629) );
  XOR U4767 ( .A(n4603), .B(n4634), .Z(n4604) );
  AND U4768 ( .A(n1671), .B(n3379), .Z(n4634) );
  XNOR U4769 ( .A(n4638), .B(n4605), .Z(n4633) );
  NAND U4770 ( .A(n3330), .B(n1710), .Z(n4605) );
  IV U4771 ( .A(n4607), .Z(n4638) );
  XOR U4772 ( .A(n4642), .B(n4643), .Z(n4621) );
  AND U4773 ( .A(n4644), .B(n4645), .Z(n4643) );
  XOR U4774 ( .A(n4646), .B(n4647), .Z(n4645) );
  XOR U4775 ( .A(n4642), .B(n4648), .Z(n4647) );
  XOR U4776 ( .A(n4640), .B(n4649), .Z(n4644) );
  XOR U4777 ( .A(n4642), .B(n4641), .Z(n4649) );
  NAND U4778 ( .A(n3236), .B(n1827), .Z(n4632) );
  XOR U4779 ( .A(n4630), .B(n4650), .Z(n4631) );
  AND U4780 ( .A(n1788), .B(n3285), .Z(n4650) );
  XOR U4781 ( .A(n4635), .B(n4655), .Z(n4636) );
  AND U4782 ( .A(n1710), .B(n3379), .Z(n4655) );
  XNOR U4783 ( .A(n4659), .B(n4637), .Z(n4654) );
  NAND U4784 ( .A(n3330), .B(n1749), .Z(n4637) );
  IV U4785 ( .A(n4639), .Z(n4659) );
  XOR U4786 ( .A(n4663), .B(n4664), .Z(n4642) );
  AND U4787 ( .A(n4665), .B(n4666), .Z(n4664) );
  XOR U4788 ( .A(n4667), .B(n4668), .Z(n4666) );
  XOR U4789 ( .A(n4663), .B(n4669), .Z(n4668) );
  XOR U4790 ( .A(n4661), .B(n4670), .Z(n4665) );
  XOR U4791 ( .A(n4663), .B(n4662), .Z(n4670) );
  NAND U4792 ( .A(n3236), .B(n1868), .Z(n4653) );
  XOR U4793 ( .A(n4651), .B(n4671), .Z(n4652) );
  AND U4794 ( .A(n1827), .B(n3285), .Z(n4671) );
  XOR U4795 ( .A(n4656), .B(n4676), .Z(n4657) );
  AND U4796 ( .A(n1749), .B(n3379), .Z(n4676) );
  XNOR U4797 ( .A(n4680), .B(n4658), .Z(n4675) );
  NAND U4798 ( .A(n3330), .B(n1788), .Z(n4658) );
  IV U4799 ( .A(n4660), .Z(n4680) );
  XOR U4800 ( .A(n4684), .B(n4685), .Z(n4663) );
  AND U4801 ( .A(n4686), .B(n4687), .Z(n4685) );
  XOR U4802 ( .A(n4688), .B(n4689), .Z(n4687) );
  XOR U4803 ( .A(n4684), .B(n4690), .Z(n4689) );
  XOR U4804 ( .A(n4682), .B(n4691), .Z(n4686) );
  XOR U4805 ( .A(n4684), .B(n4683), .Z(n4691) );
  NAND U4806 ( .A(n3236), .B(n1907), .Z(n4674) );
  XOR U4807 ( .A(n4672), .B(n4692), .Z(n4673) );
  AND U4808 ( .A(n1868), .B(n3285), .Z(n4692) );
  XOR U4809 ( .A(n4677), .B(n4697), .Z(n4678) );
  AND U4810 ( .A(n1788), .B(n3379), .Z(n4697) );
  XNOR U4811 ( .A(n4701), .B(n4679), .Z(n4696) );
  NAND U4812 ( .A(n3330), .B(n1827), .Z(n4679) );
  IV U4813 ( .A(n4681), .Z(n4701) );
  XOR U4814 ( .A(n4705), .B(n4706), .Z(n4684) );
  AND U4815 ( .A(n4707), .B(n4708), .Z(n4706) );
  XOR U4816 ( .A(n4709), .B(n4710), .Z(n4708) );
  XOR U4817 ( .A(n4705), .B(n4711), .Z(n4710) );
  XOR U4818 ( .A(n4703), .B(n4712), .Z(n4707) );
  XOR U4819 ( .A(n4705), .B(n4704), .Z(n4712) );
  NAND U4820 ( .A(n3236), .B(n1946), .Z(n4695) );
  XOR U4821 ( .A(n4693), .B(n4713), .Z(n4694) );
  AND U4822 ( .A(n1907), .B(n3285), .Z(n4713) );
  XOR U4823 ( .A(n4698), .B(n4718), .Z(n4699) );
  AND U4824 ( .A(n1827), .B(n3379), .Z(n4718) );
  XNOR U4825 ( .A(n4722), .B(n4700), .Z(n4717) );
  NAND U4826 ( .A(n3330), .B(n1868), .Z(n4700) );
  IV U4827 ( .A(n4702), .Z(n4722) );
  XOR U4828 ( .A(n4726), .B(n4727), .Z(n4705) );
  AND U4829 ( .A(n4728), .B(n4729), .Z(n4727) );
  XOR U4830 ( .A(n4730), .B(n4731), .Z(n4729) );
  XOR U4831 ( .A(n4726), .B(n4732), .Z(n4731) );
  XOR U4832 ( .A(n4724), .B(n4733), .Z(n4728) );
  XOR U4833 ( .A(n4726), .B(n4725), .Z(n4733) );
  NAND U4834 ( .A(n3236), .B(n1987), .Z(n4716) );
  XOR U4835 ( .A(n4714), .B(n4734), .Z(n4715) );
  AND U4836 ( .A(n1946), .B(n3285), .Z(n4734) );
  XOR U4837 ( .A(n4719), .B(n4739), .Z(n4720) );
  AND U4838 ( .A(n1868), .B(n3379), .Z(n4739) );
  XNOR U4839 ( .A(n4743), .B(n4721), .Z(n4738) );
  NAND U4840 ( .A(n3330), .B(n1907), .Z(n4721) );
  IV U4841 ( .A(n4723), .Z(n4743) );
  XOR U4842 ( .A(n4747), .B(n4748), .Z(n4726) );
  AND U4843 ( .A(n4749), .B(n4750), .Z(n4748) );
  XOR U4844 ( .A(n4751), .B(n4752), .Z(n4750) );
  XOR U4845 ( .A(n4747), .B(n4753), .Z(n4752) );
  XOR U4846 ( .A(n4745), .B(n4754), .Z(n4749) );
  XOR U4847 ( .A(n4747), .B(n4746), .Z(n4754) );
  NAND U4848 ( .A(n3236), .B(n2028), .Z(n4737) );
  XOR U4849 ( .A(n4735), .B(n4755), .Z(n4736) );
  AND U4850 ( .A(n1987), .B(n3285), .Z(n4755) );
  XOR U4851 ( .A(n4756), .B(n4757), .Z(n4735) );
  ANDN U4852 ( .A(n4758), .B(n4759), .Z(n4757) );
  XNOR U4853 ( .A(n4760), .B(n4756), .Z(n4758) );
  XOR U4854 ( .A(n4740), .B(n4762), .Z(n4741) );
  AND U4855 ( .A(n1907), .B(n3379), .Z(n4762) );
  XNOR U4856 ( .A(n4766), .B(n4742), .Z(n4761) );
  NAND U4857 ( .A(n3330), .B(n1946), .Z(n4742) );
  IV U4858 ( .A(n4744), .Z(n4766) );
  XOR U4859 ( .A(n4771), .B(n4772), .Z(n4615) );
  XNOR U4860 ( .A(n4773), .B(n4770), .Z(n4771) );
  XOR U4861 ( .A(n4763), .B(n4775), .Z(n4764) );
  AND U4862 ( .A(n1946), .B(n3379), .Z(n4775) );
  XOR U4863 ( .A(n4778), .B(n4776), .Z(n4777) );
  AND U4864 ( .A(n1987), .B(n3379), .Z(n4778) );
  AND U4865 ( .A(n2028), .B(n3330), .Z(n4779) );
  XNOR U4866 ( .A(n4783), .B(n4765), .Z(n4774) );
  NAND U4867 ( .A(n3330), .B(n1987), .Z(n4765) );
  IV U4868 ( .A(n4767), .Z(n4783) );
  NAND U4869 ( .A(n3330), .B(n2683), .Z(n4782) );
  XOR U4870 ( .A(n4780), .B(n4784), .Z(n4781) );
  AND U4871 ( .A(n2028), .B(n3379), .Z(n4784) );
  ANDN U4872 ( .A(n4785), .B(n2686), .Z(n4780) );
  NANDN U4873 ( .B(n3330), .A(n4786), .Z(n4785) );
  NAND U4874 ( .A(n2683), .B(n3379), .Z(n4786) );
  XNOR U4875 ( .A(n4787), .B(e_input[20]), .Z(n3379) );
  NAND U4876 ( .A(e_input[31]), .B(n4788), .Z(n4787) );
  XOR U4877 ( .A(e_input[20]), .B(\_MAC/_MULT/X_[20] ), .Z(n4788) );
  XNOR U4878 ( .A(n4789), .B(e_input[21]), .Z(n3330) );
  NAND U4879 ( .A(e_input[31]), .B(n4790), .Z(n4789) );
  XOR U4880 ( .A(e_input[21]), .B(\_MAC/_MULT/X_[21] ), .Z(n4790) );
  XNOR U4881 ( .A(n4759), .B(n4760), .Z(n4769) );
  NAND U4882 ( .A(n3236), .B(n2683), .Z(n4760) );
  XNOR U4883 ( .A(n4756), .B(n4791), .Z(n4759) );
  AND U4884 ( .A(n2028), .B(n3285), .Z(n4791) );
  ANDN U4885 ( .A(n4792), .B(n2686), .Z(n4756) );
  NANDN U4886 ( .B(n3236), .A(n4793), .Z(n4792) );
  NAND U4887 ( .A(n2683), .B(n3285), .Z(n4793) );
  XNOR U4888 ( .A(n4794), .B(e_input[22]), .Z(n3285) );
  NAND U4889 ( .A(e_input[31]), .B(n4795), .Z(n4794) );
  XOR U4890 ( .A(e_input[22]), .B(\_MAC/_MULT/X_[22] ), .Z(n4795) );
  XNOR U4891 ( .A(n4796), .B(e_input[23]), .Z(n3236) );
  NAND U4892 ( .A(e_input[31]), .B(n4797), .Z(n4796) );
  XOR U4893 ( .A(e_input[23]), .B(\_MAC/_MULT/X_[23] ), .Z(n4797) );
  XOR U4894 ( .A(n4798), .B(n4799), .Z(n4770) );
  XOR U4895 ( .A(n4301), .B(n4801), .Z(n4302) );
  AND U4896 ( .A(n1476), .B(n3650), .Z(n4801) );
  XNOR U4897 ( .A(n4802), .B(g_input[16]), .Z(n1476) );
  NAND U4898 ( .A(n4803), .B(g_input[31]), .Z(n4802) );
  XOR U4899 ( .A(g_input[16]), .B(\_MAC/_MULT/A_[16] ), .Z(n4803) );
  XNOR U4900 ( .A(n4807), .B(n4303), .Z(n4800) );
  NAND U4901 ( .A(n3589), .B(n1515), .Z(n4303) );
  IV U4902 ( .A(n4305), .Z(n4807) );
  NAND U4903 ( .A(n3454), .B(n1632), .Z(n4620) );
  XOR U4904 ( .A(n4618), .B(n4809), .Z(n4619) );
  AND U4905 ( .A(n1593), .B(n3516), .Z(n4809) );
  XOR U4906 ( .A(n4804), .B(n4814), .Z(n4805) );
  AND U4907 ( .A(n1515), .B(n3650), .Z(n4814) );
  XNOR U4908 ( .A(n4815), .B(g_input[15]), .Z(n1515) );
  NAND U4909 ( .A(n4816), .B(g_input[31]), .Z(n4815) );
  XOR U4910 ( .A(g_input[15]), .B(\_MAC/_MULT/A_[15] ), .Z(n4816) );
  XNOR U4911 ( .A(n4820), .B(n4806), .Z(n4813) );
  NAND U4912 ( .A(n3589), .B(n1554), .Z(n4806) );
  IV U4913 ( .A(n4808), .Z(n4820) );
  NAND U4914 ( .A(n3454), .B(n1671), .Z(n4812) );
  XOR U4915 ( .A(n4810), .B(n4822), .Z(n4811) );
  AND U4916 ( .A(n1632), .B(n3516), .Z(n4822) );
  XOR U4917 ( .A(n4817), .B(n4827), .Z(n4818) );
  AND U4918 ( .A(n1554), .B(n3650), .Z(n4827) );
  XNOR U4919 ( .A(n4828), .B(g_input[14]), .Z(n1554) );
  NAND U4920 ( .A(n4829), .B(g_input[31]), .Z(n4828) );
  XOR U4921 ( .A(g_input[14]), .B(\_MAC/_MULT/A_[14] ), .Z(n4829) );
  XNOR U4922 ( .A(n4833), .B(n4819), .Z(n4826) );
  NAND U4923 ( .A(n3589), .B(n1593), .Z(n4819) );
  IV U4924 ( .A(n4821), .Z(n4833) );
  NAND U4925 ( .A(n3454), .B(n1710), .Z(n4825) );
  XOR U4926 ( .A(n4823), .B(n4835), .Z(n4824) );
  AND U4927 ( .A(n1671), .B(n3516), .Z(n4835) );
  XOR U4928 ( .A(n4830), .B(n4840), .Z(n4831) );
  AND U4929 ( .A(n1593), .B(n3650), .Z(n4840) );
  XNOR U4930 ( .A(n4841), .B(g_input[13]), .Z(n1593) );
  NAND U4931 ( .A(n4842), .B(g_input[31]), .Z(n4841) );
  XOR U4932 ( .A(g_input[13]), .B(\_MAC/_MULT/A_[13] ), .Z(n4842) );
  XNOR U4933 ( .A(n4846), .B(n4832), .Z(n4839) );
  NAND U4934 ( .A(n3589), .B(n1632), .Z(n4832) );
  IV U4935 ( .A(n4834), .Z(n4846) );
  NAND U4936 ( .A(n3454), .B(n1749), .Z(n4838) );
  XOR U4937 ( .A(n4836), .B(n4848), .Z(n4837) );
  AND U4938 ( .A(n1710), .B(n3516), .Z(n4848) );
  XOR U4939 ( .A(n4843), .B(n4853), .Z(n4844) );
  AND U4940 ( .A(n1632), .B(n3650), .Z(n4853) );
  XNOR U4941 ( .A(n4854), .B(g_input[12]), .Z(n1632) );
  NAND U4942 ( .A(n4855), .B(g_input[31]), .Z(n4854) );
  XOR U4943 ( .A(g_input[12]), .B(\_MAC/_MULT/A_[12] ), .Z(n4855) );
  XNOR U4944 ( .A(n4859), .B(n4845), .Z(n4852) );
  NAND U4945 ( .A(n3589), .B(n1671), .Z(n4845) );
  IV U4946 ( .A(n4847), .Z(n4859) );
  NAND U4947 ( .A(n3454), .B(n1788), .Z(n4851) );
  XOR U4948 ( .A(n4849), .B(n4861), .Z(n4850) );
  AND U4949 ( .A(n1749), .B(n3516), .Z(n4861) );
  XOR U4950 ( .A(n4856), .B(n4866), .Z(n4857) );
  AND U4951 ( .A(n1671), .B(n3650), .Z(n4866) );
  XNOR U4952 ( .A(n4867), .B(g_input[11]), .Z(n1671) );
  NAND U4953 ( .A(n4868), .B(g_input[31]), .Z(n4867) );
  XOR U4954 ( .A(g_input[11]), .B(\_MAC/_MULT/A_[11] ), .Z(n4868) );
  XNOR U4955 ( .A(n4872), .B(n4858), .Z(n4865) );
  NAND U4956 ( .A(n3589), .B(n1710), .Z(n4858) );
  IV U4957 ( .A(n4860), .Z(n4872) );
  NAND U4958 ( .A(n3454), .B(n1827), .Z(n4864) );
  XOR U4959 ( .A(n4862), .B(n4874), .Z(n4863) );
  AND U4960 ( .A(n1788), .B(n3516), .Z(n4874) );
  XOR U4961 ( .A(n4869), .B(n4879), .Z(n4870) );
  AND U4962 ( .A(n1710), .B(n3650), .Z(n4879) );
  XNOR U4963 ( .A(n4880), .B(g_input[10]), .Z(n1710) );
  NAND U4964 ( .A(n4881), .B(g_input[31]), .Z(n4880) );
  XOR U4965 ( .A(g_input[10]), .B(\_MAC/_MULT/A_[10] ), .Z(n4881) );
  XNOR U4966 ( .A(n4885), .B(n4871), .Z(n4878) );
  NAND U4967 ( .A(n3589), .B(n1749), .Z(n4871) );
  IV U4968 ( .A(n4873), .Z(n4885) );
  NAND U4969 ( .A(n3454), .B(n1868), .Z(n4877) );
  XOR U4970 ( .A(n4875), .B(n4887), .Z(n4876) );
  AND U4971 ( .A(n1827), .B(n3516), .Z(n4887) );
  XOR U4972 ( .A(n4882), .B(n4892), .Z(n4883) );
  AND U4973 ( .A(n1749), .B(n3650), .Z(n4892) );
  XNOR U4974 ( .A(n4893), .B(g_input[9]), .Z(n1749) );
  NAND U4975 ( .A(n4894), .B(g_input[31]), .Z(n4893) );
  XOR U4976 ( .A(g_input[9]), .B(\_MAC/_MULT/A_[9] ), .Z(n4894) );
  XNOR U4977 ( .A(n4898), .B(n4884), .Z(n4891) );
  NAND U4978 ( .A(n3589), .B(n1788), .Z(n4884) );
  IV U4979 ( .A(n4886), .Z(n4898) );
  NAND U4980 ( .A(n3454), .B(n1907), .Z(n4890) );
  XOR U4981 ( .A(n4888), .B(n4900), .Z(n4889) );
  AND U4982 ( .A(n1868), .B(n3516), .Z(n4900) );
  XNOR U4983 ( .A(n4904), .B(n4901), .Z(n4903) );
  XOR U4984 ( .A(n4895), .B(n4906), .Z(n4896) );
  AND U4985 ( .A(n1788), .B(n3650), .Z(n4906) );
  XNOR U4986 ( .A(n4910), .B(n4907), .Z(n4909) );
  XNOR U4987 ( .A(n4911), .B(n4897), .Z(n4905) );
  NAND U4988 ( .A(n3589), .B(n1827), .Z(n4897) );
  IV U4989 ( .A(n4899), .Z(n4911) );
  XOR U4990 ( .A(n4912), .B(n4913), .Z(n4899) );
  AND U4991 ( .A(n4914), .B(n4915), .Z(n4913) );
  XOR U4992 ( .A(n4908), .B(n4916), .Z(n4915) );
  XNOR U4993 ( .A(n4910), .B(n4912), .Z(n4916) );
  NAND U4994 ( .A(n3589), .B(n1868), .Z(n4910) );
  XOR U4995 ( .A(n4907), .B(n4917), .Z(n4908) );
  AND U4996 ( .A(n1827), .B(n3650), .Z(n4917) );
  XNOR U4997 ( .A(n4921), .B(n4918), .Z(n4920) );
  XOR U4998 ( .A(n4902), .B(n4922), .Z(n4914) );
  XNOR U4999 ( .A(n4904), .B(n4912), .Z(n4922) );
  NAND U5000 ( .A(n3454), .B(n1946), .Z(n4904) );
  XOR U5001 ( .A(n4901), .B(n4923), .Z(n4902) );
  AND U5002 ( .A(n1907), .B(n3516), .Z(n4923) );
  XNOR U5003 ( .A(n4927), .B(n4924), .Z(n4926) );
  XOR U5004 ( .A(n4928), .B(n4929), .Z(n4912) );
  AND U5005 ( .A(n4930), .B(n4931), .Z(n4929) );
  XOR U5006 ( .A(n4919), .B(n4932), .Z(n4931) );
  XNOR U5007 ( .A(n4921), .B(n4928), .Z(n4932) );
  NAND U5008 ( .A(n3589), .B(n1907), .Z(n4921) );
  XOR U5009 ( .A(n4918), .B(n4933), .Z(n4919) );
  AND U5010 ( .A(n1868), .B(n3650), .Z(n4933) );
  XNOR U5011 ( .A(n4937), .B(n4934), .Z(n4936) );
  XOR U5012 ( .A(n4925), .B(n4938), .Z(n4930) );
  XNOR U5013 ( .A(n4927), .B(n4928), .Z(n4938) );
  NAND U5014 ( .A(n3454), .B(n1987), .Z(n4927) );
  XOR U5015 ( .A(n4924), .B(n4939), .Z(n4925) );
  AND U5016 ( .A(n1946), .B(n3516), .Z(n4939) );
  XNOR U5017 ( .A(n4943), .B(n4940), .Z(n4942) );
  XOR U5018 ( .A(n4944), .B(n4945), .Z(n4928) );
  AND U5019 ( .A(n4946), .B(n4947), .Z(n4945) );
  XOR U5020 ( .A(n4935), .B(n4948), .Z(n4947) );
  XNOR U5021 ( .A(n4937), .B(n4944), .Z(n4948) );
  NAND U5022 ( .A(n3589), .B(n1946), .Z(n4937) );
  XOR U5023 ( .A(n4934), .B(n4949), .Z(n4935) );
  AND U5024 ( .A(n1907), .B(n3650), .Z(n4949) );
  XOR U5025 ( .A(n4941), .B(n4953), .Z(n4946) );
  XNOR U5026 ( .A(n4943), .B(n4944), .Z(n4953) );
  NAND U5027 ( .A(n3454), .B(n2028), .Z(n4943) );
  XOR U5028 ( .A(n4940), .B(n4954), .Z(n4941) );
  AND U5029 ( .A(n1987), .B(n3516), .Z(n4954) );
  XOR U5030 ( .A(n4955), .B(n4956), .Z(n4940) );
  AND U5031 ( .A(n4957), .B(n4958), .Z(n4956) );
  XNOR U5032 ( .A(n4959), .B(n4955), .Z(n4957) );
  NAND U5033 ( .A(n3454), .B(n2683), .Z(n4959) );
  XOR U5034 ( .A(n4955), .B(n4961), .Z(n4958) );
  AND U5035 ( .A(n2028), .B(n3516), .Z(n4961) );
  ANDN U5036 ( .A(n4962), .B(n2686), .Z(n4955) );
  NANDN U5037 ( .B(n3454), .A(n4963), .Z(n4962) );
  NAND U5038 ( .A(n2683), .B(n3516), .Z(n4963) );
  XNOR U5039 ( .A(n4964), .B(e_input[18]), .Z(n3516) );
  NAND U5040 ( .A(e_input[31]), .B(n4965), .Z(n4964) );
  XOR U5041 ( .A(e_input[18]), .B(\_MAC/_MULT/X_[18] ), .Z(n4965) );
  XNOR U5042 ( .A(n4966), .B(e_input[19]), .Z(n3454) );
  NAND U5043 ( .A(e_input[31]), .B(n4967), .Z(n4966) );
  XOR U5044 ( .A(e_input[19]), .B(\_MAC/_MULT/X_[19] ), .Z(n4967) );
  XOR U5045 ( .A(n4950), .B(n4969), .Z(n4951) );
  AND U5046 ( .A(n1946), .B(n3650), .Z(n4969) );
  XOR U5047 ( .A(n4972), .B(n4970), .Z(n4971) );
  AND U5048 ( .A(n1987), .B(n3650), .Z(n4972) );
  AND U5049 ( .A(n2028), .B(n3589), .Z(n4973) );
  XNOR U5050 ( .A(n4977), .B(n4952), .Z(n4968) );
  NAND U5051 ( .A(n3589), .B(n1987), .Z(n4952) );
  IV U5052 ( .A(n4960), .Z(n4977) );
  NAND U5053 ( .A(n3589), .B(n2683), .Z(n4976) );
  XOR U5054 ( .A(n4974), .B(n4978), .Z(n4975) );
  AND U5055 ( .A(n2028), .B(n3650), .Z(n4978) );
  ANDN U5056 ( .A(n4979), .B(n2686), .Z(n4974) );
  NANDN U5057 ( .B(n3589), .A(n4980), .Z(n4979) );
  NAND U5058 ( .A(n2683), .B(n3650), .Z(n4980) );
  XNOR U5059 ( .A(n4981), .B(e_input[16]), .Z(n3650) );
  NAND U5060 ( .A(e_input[31]), .B(n4982), .Z(n4981) );
  XOR U5061 ( .A(e_input[16]), .B(\_MAC/_MULT/X_[16] ), .Z(n4982) );
  XNOR U5062 ( .A(n4983), .B(e_input[17]), .Z(n3589) );
  NAND U5063 ( .A(e_input[31]), .B(n4984), .Z(n4983) );
  XOR U5064 ( .A(e_input[17]), .B(\_MAC/_MULT/X_[17] ), .Z(n4984) );
  XOR U5065 ( .A(n4985), .B(n4483), .Z(n4368) );
  XNOR U5066 ( .A(n4473), .B(n4474), .Z(n4483) );
  NAND U5067 ( .A(n3096), .B(n1907), .Z(n4474) );
  XNOR U5068 ( .A(n4472), .B(n4986), .Z(n4473) );
  AND U5069 ( .A(n1868), .B(n3126), .Z(n4986) );
  XNOR U5070 ( .A(n4990), .B(n4987), .Z(n4989) );
  XNOR U5071 ( .A(n4482), .B(n4367), .Z(n4985) );
  XOR U5072 ( .A(n4991), .B(n4992), .Z(n4367) );
  XOR U5073 ( .A(n4477), .B(n4994), .Z(n4478) );
  AND U5074 ( .A(n1788), .B(n3211), .Z(n4994) );
  XNOR U5075 ( .A(n4995), .B(g_input[8]), .Z(n1788) );
  NAND U5076 ( .A(n4996), .B(g_input[31]), .Z(n4995) );
  XOR U5077 ( .A(g_input[8]), .B(\_MAC/_MULT/A_[8] ), .Z(n4996) );
  XNOR U5078 ( .A(n5000), .B(n4997), .Z(n4999) );
  XNOR U5079 ( .A(n5001), .B(n4479), .Z(n4993) );
  NAND U5080 ( .A(n3168), .B(n1827), .Z(n4479) );
  IV U5081 ( .A(n4481), .Z(n5001) );
  XOR U5082 ( .A(n5002), .B(n5003), .Z(n4481) );
  AND U5083 ( .A(n5004), .B(n5005), .Z(n5003) );
  XOR U5084 ( .A(n4998), .B(n5006), .Z(n5005) );
  XNOR U5085 ( .A(n5000), .B(n5002), .Z(n5006) );
  NAND U5086 ( .A(n3168), .B(n1868), .Z(n5000) );
  XOR U5087 ( .A(n4997), .B(n5007), .Z(n4998) );
  AND U5088 ( .A(n1827), .B(n3211), .Z(n5007) );
  XNOR U5089 ( .A(n5008), .B(g_input[7]), .Z(n1827) );
  NAND U5090 ( .A(n5009), .B(g_input[31]), .Z(n5008) );
  XOR U5091 ( .A(g_input[7]), .B(\_MAC/_MULT/A_[7] ), .Z(n5009) );
  XNOR U5092 ( .A(n5013), .B(n5010), .Z(n5012) );
  XOR U5093 ( .A(n4988), .B(n5014), .Z(n5004) );
  XNOR U5094 ( .A(n4990), .B(n5002), .Z(n5014) );
  NAND U5095 ( .A(n3096), .B(n1946), .Z(n4990) );
  XOR U5096 ( .A(n4987), .B(n5015), .Z(n4988) );
  AND U5097 ( .A(n1907), .B(n3126), .Z(n5015) );
  XNOR U5098 ( .A(n5019), .B(n5016), .Z(n5018) );
  XOR U5099 ( .A(n5020), .B(n5021), .Z(n5002) );
  AND U5100 ( .A(n5022), .B(n5023), .Z(n5021) );
  XOR U5101 ( .A(n5011), .B(n5024), .Z(n5023) );
  XNOR U5102 ( .A(n5013), .B(n5020), .Z(n5024) );
  NAND U5103 ( .A(n3168), .B(n1907), .Z(n5013) );
  XOR U5104 ( .A(n5010), .B(n5025), .Z(n5011) );
  AND U5105 ( .A(n1868), .B(n3211), .Z(n5025) );
  XNOR U5106 ( .A(n5026), .B(g_input[6]), .Z(n1868) );
  NAND U5107 ( .A(n5027), .B(g_input[31]), .Z(n5026) );
  XOR U5108 ( .A(g_input[6]), .B(\_MAC/_MULT/A_[6] ), .Z(n5027) );
  XNOR U5109 ( .A(n5031), .B(n5028), .Z(n5030) );
  XOR U5110 ( .A(n5017), .B(n5032), .Z(n5022) );
  XNOR U5111 ( .A(n5019), .B(n5020), .Z(n5032) );
  NAND U5112 ( .A(n3096), .B(n1987), .Z(n5019) );
  XOR U5113 ( .A(n5016), .B(n5033), .Z(n5017) );
  AND U5114 ( .A(n1946), .B(n3126), .Z(n5033) );
  XNOR U5115 ( .A(n5037), .B(n5034), .Z(n5036) );
  XOR U5116 ( .A(n5038), .B(n5039), .Z(n5020) );
  AND U5117 ( .A(n5040), .B(n5041), .Z(n5039) );
  XOR U5118 ( .A(n5029), .B(n5042), .Z(n5041) );
  XNOR U5119 ( .A(n5031), .B(n5038), .Z(n5042) );
  NAND U5120 ( .A(n3168), .B(n1946), .Z(n5031) );
  XOR U5121 ( .A(n5028), .B(n5043), .Z(n5029) );
  AND U5122 ( .A(n1907), .B(n3211), .Z(n5043) );
  XNOR U5123 ( .A(n5044), .B(g_input[5]), .Z(n1907) );
  NAND U5124 ( .A(n5045), .B(g_input[31]), .Z(n5044) );
  XOR U5125 ( .A(g_input[5]), .B(\_MAC/_MULT/A_[5] ), .Z(n5045) );
  XOR U5126 ( .A(n5035), .B(n5049), .Z(n5040) );
  XNOR U5127 ( .A(n5037), .B(n5038), .Z(n5049) );
  NAND U5128 ( .A(n3096), .B(n2028), .Z(n5037) );
  XOR U5129 ( .A(n5034), .B(n5050), .Z(n5035) );
  AND U5130 ( .A(n1987), .B(n3126), .Z(n5050) );
  NAND U5131 ( .A(n3096), .B(n2683), .Z(n5053) );
  XOR U5132 ( .A(n5051), .B(n5055), .Z(n5052) );
  AND U5133 ( .A(n2028), .B(n3126), .Z(n5055) );
  ANDN U5134 ( .A(n5056), .B(n2686), .Z(n5051) );
  NANDN U5135 ( .B(n3096), .A(n5057), .Z(n5056) );
  NAND U5136 ( .A(n2683), .B(n3126), .Z(n5057) );
  XNOR U5137 ( .A(n5058), .B(e_input[26]), .Z(n3126) );
  NAND U5138 ( .A(e_input[31]), .B(n5059), .Z(n5058) );
  XOR U5139 ( .A(e_input[26]), .B(\_MAC/_MULT/X_[26] ), .Z(n5059) );
  XNOR U5140 ( .A(n5060), .B(e_input[27]), .Z(n3096) );
  NAND U5141 ( .A(e_input[31]), .B(n5061), .Z(n5060) );
  XOR U5142 ( .A(e_input[27]), .B(\_MAC/_MULT/X_[27] ), .Z(n5061) );
  XOR U5143 ( .A(n5046), .B(n5063), .Z(n5047) );
  AND U5144 ( .A(n1946), .B(n3211), .Z(n5063) );
  XOR U5145 ( .A(n5066), .B(n5064), .Z(n5065) );
  AND U5146 ( .A(n1987), .B(n3211), .Z(n5066) );
  AND U5147 ( .A(n2028), .B(n3168), .Z(n5067) );
  XNOR U5148 ( .A(n5071), .B(n5048), .Z(n5062) );
  NAND U5149 ( .A(n3168), .B(n1987), .Z(n5048) );
  IV U5150 ( .A(n5054), .Z(n5071) );
  NAND U5151 ( .A(n3168), .B(n2683), .Z(n5070) );
  XOR U5152 ( .A(n5068), .B(n5072), .Z(n5069) );
  AND U5153 ( .A(n2028), .B(n3211), .Z(n5072) );
  ANDN U5154 ( .A(n5073), .B(n2686), .Z(n5068) );
  NANDN U5155 ( .B(n3168), .A(n5074), .Z(n5073) );
  NAND U5156 ( .A(n2683), .B(n3211), .Z(n5074) );
  XNOR U5157 ( .A(n5075), .B(e_input[24]), .Z(n3211) );
  NAND U5158 ( .A(e_input[31]), .B(n5076), .Z(n5075) );
  XOR U5159 ( .A(e_input[24]), .B(\_MAC/_MULT/X_[24] ), .Z(n5076) );
  XNOR U5160 ( .A(n5077), .B(e_input[25]), .Z(n3168) );
  NAND U5161 ( .A(e_input[31]), .B(n5078), .Z(n5077) );
  XOR U5162 ( .A(e_input[25]), .B(\_MAC/_MULT/X_[25] ), .Z(n5078) );
  XOR U5163 ( .A(n4569), .B(n5080), .Z(n4570) );
  AND U5164 ( .A(n1946), .B(n3081), .Z(n5080) );
  XNOR U5165 ( .A(n5081), .B(g_input[4]), .Z(n1946) );
  NAND U5166 ( .A(n5082), .B(g_input[31]), .Z(n5081) );
  XOR U5167 ( .A(g_input[4]), .B(\_MAC/_MULT/A_[4] ), .Z(n5082) );
  XOR U5168 ( .A(n5085), .B(n5083), .Z(n5084) );
  AND U5169 ( .A(n1987), .B(n3081), .Z(n5085) );
  AND U5170 ( .A(n2028), .B(n3055), .Z(n5086) );
  XNOR U5171 ( .A(n5090), .B(n4571), .Z(n5079) );
  NAND U5172 ( .A(n3055), .B(n1987), .Z(n4571) );
  XNOR U5173 ( .A(n5091), .B(g_input[3]), .Z(n1987) );
  NAND U5174 ( .A(n5092), .B(g_input[31]), .Z(n5091) );
  XOR U5175 ( .A(g_input[3]), .B(\_MAC/_MULT/A_[3] ), .Z(n5092) );
  IV U5176 ( .A(n4575), .Z(n5090) );
  NAND U5177 ( .A(n3055), .B(n2683), .Z(n5089) );
  XOR U5178 ( .A(n5087), .B(n5093), .Z(n5088) );
  AND U5179 ( .A(n2028), .B(n3081), .Z(n5093) );
  ANDN U5180 ( .A(n5094), .B(n2686), .Z(n5087) );
  NANDN U5181 ( .B(n3055), .A(n5095), .Z(n5094) );
  NAND U5182 ( .A(n2683), .B(n3081), .Z(n5095) );
  XNOR U5183 ( .A(n5096), .B(e_input[28]), .Z(n3081) );
  NAND U5184 ( .A(e_input[31]), .B(n5097), .Z(n5096) );
  XOR U5185 ( .A(e_input[28]), .B(\_MAC/_MULT/X_[28] ), .Z(n5097) );
  XNOR U5186 ( .A(n5098), .B(e_input[29]), .Z(n3055) );
  NAND U5187 ( .A(e_input[31]), .B(n5099), .Z(n5098) );
  XOR U5188 ( .A(e_input[29]), .B(\_MAC/_MULT/X_[29] ), .Z(n5099) );
  XNOR U5189 ( .A(n4598), .B(n4599), .Z(n4577) );
  NAND U5190 ( .A(n3024), .B(n2683), .Z(n4599) );
  XNOR U5191 ( .A(n4597), .B(n5100), .Z(n4598) );
  AND U5192 ( .A(n2028), .B(n3041), .Z(n5100) );
  XNOR U5193 ( .A(n5101), .B(g_input[2]), .Z(n2028) );
  NAND U5194 ( .A(n5102), .B(g_input[31]), .Z(n5101) );
  XOR U5195 ( .A(g_input[2]), .B(\_MAC/_MULT/A_[2] ), .Z(n5102) );
  ANDN U5196 ( .A(n5103), .B(n2686), .Z(n4597) );
  XOR U5197 ( .A(n5104), .B(g_input[0]), .Z(n2686) );
  NAND U5198 ( .A(n5105), .B(g_input[31]), .Z(n5104) );
  XOR U5199 ( .A(g_input[0]), .B(\_MAC/_MULT/A_[0] ), .Z(n5105) );
  NANDN U5200 ( .B(n3024), .A(n5106), .Z(n5103) );
  NAND U5201 ( .A(n2683), .B(n3041), .Z(n5106) );
  XNOR U5202 ( .A(n5107), .B(e_input[30]), .Z(n3041) );
  NAND U5203 ( .A(e_input[31]), .B(n5108), .Z(n5107) );
  XOR U5204 ( .A(e_input[30]), .B(\_MAC/_MULT/X_[30] ), .Z(n5108) );
  XNOR U5205 ( .A(n5109), .B(g_input[1]), .Z(n2683) );
  NAND U5206 ( .A(n5110), .B(g_input[31]), .Z(n5109) );
  XOR U5207 ( .A(g_input[1]), .B(\_MAC/_MULT/A_[1] ), .Z(n5110) );
  ANDN U5208 ( .A(\_MAC/_MULT/X_[31] ), .B(n5111), .Z(n3024) );
  IV U5209 ( .A(e_input[31]), .Z(n5111) );
endmodule

