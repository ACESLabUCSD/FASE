
module MAC_TG_N16 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MAC/AX[15] , \_MAC/AX[14] , \_MAC/AX[13] , \_MAC/AX[12] ,
         \_MAC/AX[11] , \_MAC/AX[10] , \_MAC/AX[9] , \_MAC/AX[8] ,
         \_MAC/AX[7] , \_MAC/AX[6] , \_MAC/AX[5] , \_MAC/AX[4] , \_MAC/AX[3] ,
         \_MAC/AX[2] , \_MAC/AX[1] , \_MAC/AX[0] , \_MAC/_MULT/AX__[15] ,
         \_MAC/_MULT/AX__[14] , \_MAC/_MULT/AX__[13] , \_MAC/_MULT/AX__[12] ,
         \_MAC/_MULT/AX__[11] , \_MAC/_MULT/AX__[10] , \_MAC/_MULT/AX__[9] ,
         \_MAC/_MULT/AX__[8] , \_MAC/_MULT/AX__[7] , \_MAC/_MULT/AX__[6] ,
         \_MAC/_MULT/AX__[5] , \_MAC/_MULT/AX__[4] , \_MAC/_MULT/AX__[3] ,
         \_MAC/_MULT/AX__[2] , \_MAC/_MULT/AX__[1] , \_MAC/_MULT/AX__[0] ,
         \_MAC/_MULT/AX_[0] , \_MAC/_MULT/AX_[1] , \_MAC/_MULT/AX_[2] ,
         \_MAC/_MULT/AX_[3] , \_MAC/_MULT/AX_[4] , \_MAC/_MULT/AX_[5] ,
         \_MAC/_MULT/AX_[6] , \_MAC/_MULT/AX_[7] , \_MAC/_MULT/AX_[8] ,
         \_MAC/_MULT/AX_[9] , \_MAC/_MULT/AX_[10] , \_MAC/_MULT/AX_[11] ,
         \_MAC/_MULT/AX_[12] , \_MAC/_MULT/AX_[13] , \_MAC/_MULT/AX_[14] ,
         \_MAC/_MULT/AX_[15] , \_MAC/_MULT/X_[15] , \_MAC/_MULT/X_[14] ,
         \_MAC/_MULT/X_[13] , \_MAC/_MULT/X_[12] , \_MAC/_MULT/X_[11] ,
         \_MAC/_MULT/X_[10] , \_MAC/_MULT/X_[9] , \_MAC/_MULT/X_[8] ,
         \_MAC/_MULT/X_[7] , \_MAC/_MULT/X_[6] , \_MAC/_MULT/X_[5] ,
         \_MAC/_MULT/X_[4] , \_MAC/_MULT/X_[3] , \_MAC/_MULT/X_[2] ,
         \_MAC/_MULT/X_[1] , \_MAC/_MULT/X_[0] , \_MAC/_MULT/A_[15] ,
         \_MAC/_MULT/A_[14] , \_MAC/_MULT/A_[13] , \_MAC/_MULT/A_[12] ,
         \_MAC/_MULT/A_[11] , \_MAC/_MULT/A_[10] , \_MAC/_MULT/A_[9] ,
         \_MAC/_MULT/A_[8] , \_MAC/_MULT/A_[7] , \_MAC/_MULT/A_[6] ,
         \_MAC/_MULT/A_[5] , \_MAC/_MULT/A_[4] , \_MAC/_MULT/A_[3] ,
         \_MAC/_MULT/A_[2] , \_MAC/_MULT/A_[1] , \_MAC/_MULT/A_[0] ,
         \_MAC/_MULT/MULT/S[2][1][0] , \_MAC/_MULT/MULT/S[2][1][1] ,
         \_MAC/_MULT/MULT/S[2][1][2] , \_MAC/_MULT/MULT/S[2][1][3] ,
         \_MAC/_MULT/MULT/S[2][1][4] , \_MAC/_MULT/MULT/S[2][1][5] ,
         \_MAC/_MULT/MULT/S[2][1][6] , \_MAC/_MULT/MULT/S[2][1][7] ,
         \_MAC/_MULT/MULT/S[2][1][8] , \_MAC/_MULT/MULT/S[2][1][9] ,
         \_MAC/_MULT/MULT/S[2][1][10] , \_MAC/_MULT/MULT/S[2][1][11] ,
         \_MAC/_MULT/MULT/S[2][1][12] , \_MAC/_MULT/MULT/S[2][1][13] ,
         \_MAC/_MULT/MULT/S[2][1][14] , \_MAC/_MULT/MULT/S[2][1][15] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[15] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[14] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[13] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[12] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[11] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[10] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[9] ,
         \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[8] , n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266;
  wire   [15:0] o_reg;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFF \o_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[0])
         );
  DFF \o_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[1])
         );
  DFF \o_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[2])
         );
  DFF \o_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[3])
         );
  DFF \o_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[4])
         );
  DFF \o_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[5])
         );
  DFF \o_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[6])
         );
  DFF \o_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[7])
         );
  DFF \o_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[8])
         );
  DFF \o_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[9])
         );
  DFF \o_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[10]) );
  DFF \o_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[11]) );
  DFF \o_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[12]) );
  DFF \o_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[13]) );
  DFF \o_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[14]) );
  DFF \o_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[15]) );
  ADD_ \_MAC/_ADD  ( .A({\_MAC/AX[15] , \_MAC/AX[14] , \_MAC/AX[13] , 
        \_MAC/AX[12] , \_MAC/AX[11] , \_MAC/AX[10] , \_MAC/AX[9] , 
        \_MAC/AX[8] , \_MAC/AX[7] , \_MAC/AX[6] , \_MAC/AX[5] , \_MAC/AX[4] , 
        \_MAC/AX[3] , \_MAC/AX[2] , \_MAC/AX[1] , \_MAC/AX[0] }), .B(o_reg), 
        .O({o, SYNOPSYS_UNCONNECTED__0}) );
  TwosComplement \_MAC/_MULT/TwosComplement_O  ( .A({\_MAC/_MULT/AX_[15] , 
        \_MAC/_MULT/AX_[14] , \_MAC/_MULT/AX_[13] , \_MAC/_MULT/AX_[12] , 
        \_MAC/_MULT/AX_[11] , \_MAC/_MULT/AX_[10] , \_MAC/_MULT/AX_[9] , 
        \_MAC/_MULT/AX_[8] , \_MAC/_MULT/AX_[7] , \_MAC/_MULT/AX_[6] , 
        \_MAC/_MULT/AX_[5] , \_MAC/_MULT/AX_[4] , \_MAC/_MULT/AX_[3] , 
        \_MAC/_MULT/AX_[2] , \_MAC/_MULT/AX_[1] , \_MAC/_MULT/AX_[0] }), .O({
        \_MAC/_MULT/AX__[15] , \_MAC/_MULT/AX__[14] , \_MAC/_MULT/AX__[13] , 
        \_MAC/_MULT/AX__[12] , \_MAC/_MULT/AX__[11] , \_MAC/_MULT/AX__[10] , 
        \_MAC/_MULT/AX__[9] , \_MAC/_MULT/AX__[8] , \_MAC/_MULT/AX__[7] , 
        \_MAC/_MULT/AX__[6] , \_MAC/_MULT/AX__[5] , \_MAC/_MULT/AX__[4] , 
        \_MAC/_MULT/AX__[3] , \_MAC/_MULT/AX__[2] , \_MAC/_MULT/AX__[1] , 
        \_MAC/_MULT/AX__[0] }) );
  TwosComplement \_MAC/_MULT/TwosComplement_B  ( .A(e_input), .O({
        \_MAC/_MULT/X_[15] , \_MAC/_MULT/X_[14] , \_MAC/_MULT/X_[13] , 
        \_MAC/_MULT/X_[12] , \_MAC/_MULT/X_[11] , \_MAC/_MULT/X_[10] , 
        \_MAC/_MULT/X_[9] , \_MAC/_MULT/X_[8] , \_MAC/_MULT/X_[7] , 
        \_MAC/_MULT/X_[6] , \_MAC/_MULT/X_[5] , \_MAC/_MULT/X_[4] , 
        \_MAC/_MULT/X_[3] , \_MAC/_MULT/X_[2] , \_MAC/_MULT/X_[1] , 
        \_MAC/_MULT/X_[0] }) );
  TwosComplement \_MAC/_MULT/TwosComplement_A  ( .A(g_input), .O({
        \_MAC/_MULT/A_[15] , \_MAC/_MULT/A_[14] , \_MAC/_MULT/A_[13] , 
        \_MAC/_MULT/A_[12] , \_MAC/_MULT/A_[11] , \_MAC/_MULT/A_[10] , 
        \_MAC/_MULT/A_[9] , \_MAC/_MULT/A_[8] , \_MAC/_MULT/A_[7] , 
        \_MAC/_MULT/A_[6] , \_MAC/_MULT/A_[5] , \_MAC/_MULT/A_[4] , 
        \_MAC/_MULT/A_[3] , \_MAC/_MULT/A_[2] , \_MAC/_MULT/A_[1] , 
        \_MAC/_MULT/A_[0] }) );
  XOR \_MAC/_MULT/MUX_O/U46  ( .A(\_MAC/_MULT/AX_[0] ), .B(n1266), .Z(
        \_MAC/AX[0] ) );
  XOR \_MAC/_MULT/MUX_O/U43  ( .A(\_MAC/_MULT/AX_[10] ), .B(n1265), .Z(
        \_MAC/AX[10] ) );
  XOR \_MAC/_MULT/MUX_O/U40  ( .A(\_MAC/_MULT/AX_[11] ), .B(n1264), .Z(
        \_MAC/AX[11] ) );
  XOR \_MAC/_MULT/MUX_O/U37  ( .A(\_MAC/_MULT/AX_[12] ), .B(n1263), .Z(
        \_MAC/AX[12] ) );
  XOR \_MAC/_MULT/MUX_O/U34  ( .A(\_MAC/_MULT/AX_[13] ), .B(n1262), .Z(
        \_MAC/AX[13] ) );
  XOR \_MAC/_MULT/MUX_O/U31  ( .A(\_MAC/_MULT/AX_[14] ), .B(n1261), .Z(
        \_MAC/AX[14] ) );
  XOR \_MAC/_MULT/MUX_O/U28  ( .A(\_MAC/_MULT/AX_[15] ), .B(n1260), .Z(
        \_MAC/AX[15] ) );
  XOR \_MAC/_MULT/MUX_O/U25  ( .A(\_MAC/_MULT/AX_[1] ), .B(n1259), .Z(
        \_MAC/AX[1] ) );
  XOR \_MAC/_MULT/MUX_O/U22  ( .A(\_MAC/_MULT/AX_[2] ), .B(n1258), .Z(
        \_MAC/AX[2] ) );
  XOR \_MAC/_MULT/MUX_O/U19  ( .A(\_MAC/_MULT/AX_[3] ), .B(n1257), .Z(
        \_MAC/AX[3] ) );
  XOR \_MAC/_MULT/MUX_O/U16  ( .A(\_MAC/_MULT/AX_[4] ), .B(n1256), .Z(
        \_MAC/AX[4] ) );
  XOR \_MAC/_MULT/MUX_O/U13  ( .A(\_MAC/_MULT/AX_[5] ), .B(n1255), .Z(
        \_MAC/AX[5] ) );
  XOR \_MAC/_MULT/MUX_O/U10  ( .A(\_MAC/_MULT/AX_[6] ), .B(n1254), .Z(
        \_MAC/AX[6] ) );
  XOR \_MAC/_MULT/MUX_O/U7  ( .A(\_MAC/_MULT/AX_[7] ), .B(n1253), .Z(
        \_MAC/AX[7] ) );
  XOR \_MAC/_MULT/MUX_O/U4  ( .A(\_MAC/_MULT/AX_[8] ), .B(n1252), .Z(
        \_MAC/AX[8] ) );
  XOR \_MAC/_MULT/MUX_O/U1  ( .A(\_MAC/_MULT/AX_[9] ), .B(n1251), .Z(
        \_MAC/AX[9] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[15].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][15] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[15] ), .Z(
        \_MAC/_MULT/AX_[15] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[14].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][14] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[14] ), .Z(
        \_MAC/_MULT/AX_[14] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[13].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][13] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[13] ), .Z(
        \_MAC/_MULT/AX_[13] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[12].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][12] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[12] ), .Z(
        \_MAC/_MULT/AX_[12] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[11].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][11] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[11] ), .Z(
        \_MAC/_MULT/AX_[11] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[10].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][10] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[10] ), .Z(
        \_MAC/_MULT/AX_[10] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[9].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][9] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[9] ), .Z(
        \_MAC/_MULT/AX_[9] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[8].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][8] ), .B(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[8] ), .Z(
        \_MAC/_MULT/AX_[8] ) );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[7].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][7] ), .B(n1250), .Z(\_MAC/_MULT/AX_[7] )
         );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[6].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][6] ), .B(n1249), .Z(\_MAC/_MULT/AX_[6] )
         );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[5].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][5] ), .B(n1248), .Z(\_MAC/_MULT/AX_[5] )
         );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[4].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][4] ), .B(n1247), .Z(\_MAC/_MULT/AX_[4] )
         );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[3].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][3] ), .B(n1246), .Z(\_MAC/_MULT/AX_[3] )
         );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[2].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][2] ), .B(n1245), .Z(\_MAC/_MULT/AX_[2] )
         );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[1].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][1] ), .B(n1244), .Z(\_MAC/_MULT/AX_[1] )
         );
  XOR \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/FA_IF2.FAINST[0].FA_/U2  ( 
        .A(\_MAC/_MULT/MULT/S[2][1][0] ), .B(n1243), .Z(\_MAC/_MULT/AX_[0] )
         );
  MUX U19 ( .IN0(n569), .IN1(n572), .SEL(n570), .F(n564) );
  MUX U20 ( .IN0(n17), .IN1(n395), .SEL(n396), .F(n380) );
  IV U21 ( .A(n397), .Z(n17) );
  XOR U22 ( .A(n390), .B(n391), .Z(n319) );
  MUX U23 ( .IN0(n18), .IN1(n674), .SEL(n675), .F(n670) );
  IV U24 ( .A(n676), .Z(n18) );
  MUX U25 ( .IN0(n1134), .IN1(n1152), .SEL(n1136), .F(n1103) );
  MUX U26 ( .IN0(n19), .IN1(n923), .SEL(n924), .F(n912) );
  IV U27 ( .A(n925), .Z(n19) );
  MUX U28 ( .IN0(n20), .IN1(n777), .SEL(n778), .F(n750) );
  IV U29 ( .A(n779), .Z(n20) );
  MUX U30 ( .IN0(n613), .IN1(n628), .SEL(n615), .F(n597) );
  XOR U31 ( .A(n376), .B(n377), .Z(n311) );
  MUX U32 ( .IN0(n670), .IN1(n673), .SEL(n671), .F(n538) );
  MUX U33 ( .IN0(n21), .IN1(n912), .SEL(n913), .F(n901) );
  IV U34 ( .A(n914), .Z(n21) );
  XNOR U35 ( .A(n1220), .B(n1221), .Z(n1067) );
  MUX U36 ( .IN0(n1153), .IN1(n1171), .SEL(n1155), .F(n1134) );
  XOR U37 ( .A(n378), .B(n370), .Z(n305) );
  MUX U38 ( .IN0(n22), .IN1(n364), .SEL(n365), .F(n352) );
  IV U39 ( .A(n366), .Z(n22) );
  XOR U40 ( .A(n475), .B(n469), .Z(n299) );
  MUX U41 ( .IN0(n23), .IN1(n1094), .SEL(n1054), .F(n1092) );
  IV U42 ( .A(n1055), .Z(n23) );
  MUX U43 ( .IN0(n24), .IN1(n901), .SEL(n902), .F(n890) );
  IV U44 ( .A(n903), .Z(n24) );
  MUX U45 ( .IN0(n752), .IN1(n25), .SEL(n751), .F(n736) );
  IV U46 ( .A(n750), .Z(n25) );
  MUX U47 ( .IN0(n619), .IN1(n635), .SEL(n621), .F(n603) );
  XOR U48 ( .A(n367), .B(n359), .Z(n297) );
  MUX U49 ( .IN0(n1103), .IN1(n1133), .SEL(n1105), .F(n942) );
  MUX U50 ( .IN0(n26), .IN1(n457), .SEL(n458), .F(n266) );
  IV U51 ( .A(n459), .Z(n26) );
  MUX U52 ( .IN0(n27), .IN1(n1098), .SEL(n1099), .F(n1096) );
  IV U53 ( .A(n1100), .Z(n27) );
  MUX U54 ( .IN0(n28), .IN1(n890), .SEL(n891), .F(n879) );
  IV U55 ( .A(n892), .Z(n28) );
  XNOR U56 ( .A(n1207), .B(n1062), .Z(n1068) );
  MUX U57 ( .IN0(n29), .IN1(n573), .SEL(n574), .F(n569) );
  IV U58 ( .A(n575), .Z(n29) );
  MUX U59 ( .IN0(n30), .IN1(n380), .SEL(n381), .F(n369) );
  IV U60 ( .A(n382), .Z(n30) );
  XOR U61 ( .A(n365), .B(n366), .Z(n303) );
  MUX U62 ( .IN0(n31), .IN1(n942), .SEL(n943), .F(n929) );
  IV U63 ( .A(n944), .Z(n31) );
  MUX U64 ( .IN0(n32), .IN1(n1096), .SEL(n1065), .F(n1094) );
  IV U65 ( .A(n1066), .Z(n32) );
  MUX U66 ( .IN0(n33), .IN1(n235), .SEL(n236), .F(n207) );
  IV U67 ( .A(n237), .Z(n33) );
  XOR U68 ( .A(n1185), .B(n1168), .Z(n1108) );
  XNOR U69 ( .A(n1057), .B(n1051), .Z(n843) );
  MUX U70 ( .IN0(n561), .IN1(n563), .SEL(n562), .F(n558) );
  MUX U71 ( .IN0(n34), .IN1(n358), .SEL(n359), .F(n345) );
  IV U72 ( .A(n360), .Z(n34) );
  XOR U73 ( .A(n464), .B(n458), .Z(n291) );
  MUX U74 ( .IN0(n35), .IN1(n282), .SEL(n283), .F(n252) );
  IV U75 ( .A(n284), .Z(n35) );
  MUX U76 ( .IN0(n36), .IN1(n873), .SEL(n874), .F(n862) );
  IV U77 ( .A(n875), .Z(n36) );
  MUX U78 ( .IN0(n37), .IN1(n1077), .SEL(n988), .F(n1073) );
  IV U79 ( .A(n989), .Z(n37) );
  MUX U80 ( .IN0(n812), .IN1(n1001), .SEL(n813), .F(n990) );
  MUX U81 ( .IN0(n868), .IN1(n38), .SEL(n867), .F(n858) );
  IV U82 ( .A(n866), .Z(n38) );
  XNOR U83 ( .A(n1046), .B(n1040), .Z(n837) );
  MUX U84 ( .IN0(n39), .IN1(n352), .SEL(n353), .F(n282) );
  IV U85 ( .A(n354), .Z(n39) );
  MUX U86 ( .IN0(n549), .IN1(n551), .SEL(n550), .F(n275) );
  XOR U87 ( .A(n355), .B(n346), .Z(n289) );
  MUX U88 ( .IN0(n40), .IN1(n1092), .SEL(n1043), .F(n1090) );
  IV U89 ( .A(n1044), .Z(n40) );
  MUX U90 ( .IN0(n41), .IN1(n207), .SEL(n208), .F(n177) );
  IV U91 ( .A(n209), .Z(n41) );
  MUX U92 ( .IN0(n42), .IN1(n862), .SEL(n863), .F(n854) );
  IV U93 ( .A(n864), .Z(n42) );
  MUX U94 ( .IN0(n894), .IN1(n821), .SEL(n822), .F(n883) );
  MUX U95 ( .IN0(n803), .IN1(n979), .SEL(n804), .F(n966) );
  XOR U96 ( .A(n1109), .B(n950), .Z(n954) );
  XNOR U97 ( .A(n1035), .B(n1029), .Z(n831) );
  MUX U98 ( .IN0(n43), .IN1(n275), .SEL(n276), .F(n244) );
  IV U99 ( .A(n277), .Z(n43) );
  MUX U100 ( .IN0(n44), .IN1(n266), .SEL(n267), .F(n235) );
  IV U101 ( .A(n268), .Z(n44) );
  MUX U102 ( .IN0(n45), .IN1(n929), .SEL(n930), .F(n918) );
  IV U103 ( .A(n931), .Z(n45) );
  MUX U104 ( .IN0(n46), .IN1(n1090), .SEL(n1032), .F(n1088) );
  IV U105 ( .A(n1033), .Z(n46) );
  MUX U106 ( .IN0(n461), .IN1(n292), .SEL(n291), .F(n270) );
  MUX U107 ( .IN0(n347), .IN1(n47), .SEL(n346), .F(n259) );
  IV U108 ( .A(n345), .Z(n47) );
  XOR U109 ( .A(n283), .B(n284), .Z(n287) );
  MUX U110 ( .IN0(n883), .IN1(n815), .SEL(n816), .F(n871) );
  MUX U111 ( .IN0(n184), .IN1(n182), .SEL(n183), .F(n162) );
  MUX U112 ( .IN0(n797), .IN1(n966), .SEL(n798), .F(n781) );
  XOR U113 ( .A(n945), .B(n937), .Z(n846) );
  XNOR U114 ( .A(n1024), .B(n1018), .Z(n825) );
  MUX U115 ( .IN0(n48), .IN1(n341), .SEL(n342), .F(n333) );
  IV U116 ( .A(n343), .Z(n48) );
  MUX U117 ( .IN0(n558), .IN1(n560), .SEL(n559), .F(n555) );
  MUX U118 ( .IN0(n49), .IN1(n369), .SEL(n370), .F(n358) );
  IV U119 ( .A(n371), .Z(n49) );
  MUX U120 ( .IN0(n50), .IN1(n918), .SEL(n919), .F(n907) );
  IV U121 ( .A(n920), .Z(n50) );
  MUX U122 ( .IN0(n51), .IN1(n1088), .SEL(n1021), .F(n1086) );
  IV U123 ( .A(n1022), .Z(n51) );
  MUX U124 ( .IN0(n52), .IN1(n252), .SEL(n253), .F(n223) );
  IV U125 ( .A(n254), .Z(n52) );
  MUX U126 ( .IN0(n213), .IN1(n211), .SEL(n212), .F(n182) );
  MUX U127 ( .IN0(n179), .IN1(n53), .SEL(n178), .F(n160) );
  IV U128 ( .A(n177), .Z(n53) );
  MUX U129 ( .IN0(n871), .IN1(n54), .SEL(n808), .F(n860) );
  IV U130 ( .A(n807), .Z(n54) );
  MUX U131 ( .IN0(n783), .IN1(n781), .SEL(n782), .F(n755) );
  XOR U132 ( .A(n932), .B(n924), .Z(n840) );
  XNOR U133 ( .A(n1013), .B(n1007), .Z(n819) );
  XNOR U134 ( .A(n675), .B(n676), .Z(n545) );
  MUX U135 ( .IN0(n55), .IN1(n1086), .SEL(n1010), .F(n1081) );
  IV U136 ( .A(n1011), .Z(n55) );
  MUX U137 ( .IN0(n241), .IN1(n239), .SEL(n240), .F(n211) );
  MUX U138 ( .IN0(n56), .IN1(n187), .SEL(n188), .F(n168) );
  IV U139 ( .A(n189), .Z(n56) );
  MUX U140 ( .IN0(n57), .IN1(n854), .SEL(n855), .F(n790) );
  IV U141 ( .A(n856), .Z(n57) );
  MUX U142 ( .IN0(n757), .IN1(n755), .SEL(n756), .F(n738) );
  XOR U143 ( .A(n344), .B(n259), .Z(n262) );
  MUX U144 ( .IN0(n58), .IN1(n223), .SEL(n224), .F(n199) );
  IV U145 ( .A(n225), .Z(n58) );
  XOR U146 ( .A(n910), .B(n902), .Z(n828) );
  XNOR U147 ( .A(n1002), .B(n998), .Z(n813) );
  MUX U148 ( .IN0(n59), .IN1(n805), .SEL(n697), .F(n799) );
  IV U149 ( .A(n696), .Z(n59) );
  MUX U150 ( .IN0(n333), .IN1(n338), .SEL(n334), .F(n325) );
  MUX U151 ( .IN0(n597), .IN1(n612), .SEL(n599), .F(n586) );
  MUX U152 ( .IN0(n552), .IN1(n554), .SEL(n553), .F(n549) );
  XOR U153 ( .A(n353), .B(n354), .Z(n295) );
  MUX U154 ( .IN0(n60), .IN1(n879), .SEL(n880), .F(n866) );
  IV U155 ( .A(n881), .Z(n60) );
  MUX U156 ( .IN0(n61), .IN1(n1073), .SEL(n977), .F(n785) );
  IV U157 ( .A(n978), .Z(n61) );
  XNOR U158 ( .A(n668), .B(n541), .Z(n546) );
  MUX U159 ( .IN0(n272), .IN1(n270), .SEL(n271), .F(n239) );
  MUX U160 ( .IN0(n830), .IN1(n1034), .SEL(n831), .F(n1023) );
  MUX U161 ( .IN0(n916), .IN1(n833), .SEL(n834), .F(n905) );
  MUX U162 ( .IN0(n990), .IN1(n809), .SEL(n810), .F(n979) );
  MUX U163 ( .IN0(n841), .IN1(n62), .SEL(n709), .F(n835) );
  IV U164 ( .A(n708), .Z(n62) );
  MUX U165 ( .IN0(n817), .IN1(n63), .SEL(n701), .F(n811) );
  IV U166 ( .A(n700), .Z(n63) );
  XOR U167 ( .A(n863), .B(n864), .Z(n807) );
  MUX U168 ( .IN0(n164), .IN1(n162), .SEL(n163), .F(n64) );
  IV U169 ( .A(n64), .Z(n147) );
  MUX U170 ( .IN0(n793), .IN1(n65), .SEL(n693), .F(n771) );
  IV U171 ( .A(n692), .Z(n65) );
  XNOR U172 ( .A(n774), .B(n751), .Z(n756) );
  XOR U173 ( .A(n173), .B(n199), .Z(n192) );
  MUX U174 ( .IN0(n547), .IN1(n545), .SEL(n546), .F(n532) );
  MUX U175 ( .IN0(n452), .IN1(n454), .SEL(n453), .F(n434) );
  MUX U176 ( .IN0(n66), .IN1(n636), .SEL(n637), .F(n619) );
  IV U177 ( .A(n638), .Z(n66) );
  MUX U178 ( .IN0(n325), .IN1(n330), .SEL(n326), .F(n317) );
  MUX U179 ( .IN0(n651), .IN1(n654), .SEL(n652), .F(n629) );
  MUX U180 ( .IN0(n483), .IN1(n308), .SEL(n307), .F(n472) );
  MUX U181 ( .IN0(n373), .IN1(n67), .SEL(n305), .F(n362) );
  IV U182 ( .A(n303), .Z(n67) );
  MUX U183 ( .IN0(n68), .IN1(n244), .SEL(n245), .F(n216) );
  IV U184 ( .A(n246), .Z(n68) );
  MUX U185 ( .IN0(n69), .IN1(n907), .SEL(n908), .F(n896) );
  IV U186 ( .A(n909), .Z(n69) );
  MUX U187 ( .IN0(n1069), .IN1(n1067), .SEL(n1068), .F(n1056) );
  MUX U188 ( .IN0(n953), .IN1(n955), .SEL(n954), .F(n940) );
  MUX U189 ( .IN0(n818), .IN1(n1012), .SEL(n819), .F(n1001) );
  MUX U190 ( .IN0(n70), .IN1(n785), .SEL(n786), .F(n759) );
  IV U191 ( .A(n787), .Z(n70) );
  MUX U192 ( .IN0(n285), .IN1(n290), .SEL(n286), .F(n255) );
  XNOR U193 ( .A(n233), .B(n208), .Z(n212) );
  MUX U194 ( .IN0(n835), .IN1(n71), .SEL(n707), .F(n829) );
  IV U195 ( .A(n706), .Z(n71) );
  XOR U196 ( .A(n876), .B(n867), .Z(n808) );
  XNOR U197 ( .A(n967), .B(n963), .Z(n798) );
  MUX U198 ( .IN0(n799), .IN1(n72), .SEL(n695), .F(n793) );
  IV U199 ( .A(n694), .Z(n72) );
  MUX U200 ( .IN0(n850), .IN1(n857), .SEL(n851), .F(n765) );
  MUX U201 ( .IN0(n740), .IN1(n738), .SEL(n739), .F(n73) );
  IV U202 ( .A(n73), .Z(n726) );
  MUX U203 ( .IN0(n171), .IN1(\_MAC/_MULT/MULT/S[2][1][4] ), .SEL(n1247), .F(
        n155) );
  MUX U204 ( .IN0(n149), .IN1(n74), .SEL(n148), .F(n141) );
  IV U205 ( .A(n147), .Z(n74) );
  MUX U206 ( .IN0(n532), .IN1(n340), .SEL(n339), .F(n519) );
  MUX U207 ( .IN0(n434), .IN1(n75), .SEL(n337), .F(n416) );
  IV U208 ( .A(n335), .Z(n75) );
  MUX U209 ( .IN0(n317), .IN1(n322), .SEL(n318), .F(n309) );
  MUX U210 ( .IN0(n603), .IN1(n618), .SEL(n605), .F(n578) );
  XNOR U211 ( .A(n658), .B(n659), .Z(n639) );
  MUX U212 ( .IN0(n362), .IN1(n76), .SEL(n297), .F(n350) );
  IV U213 ( .A(n295), .Z(n76) );
  MUX U214 ( .IN0(n77), .IN1(n896), .SEL(n897), .F(n885) );
  IV U215 ( .A(n898), .Z(n77) );
  MUX U216 ( .IN0(n842), .IN1(n1056), .SEL(n843), .F(n1045) );
  MUX U217 ( .IN0(n927), .IN1(n839), .SEL(n840), .F(n916) );
  XNOR U218 ( .A(n455), .B(n267), .Z(n271) );
  MUX U219 ( .IN0(n226), .IN1(n78), .SEL(n227), .F(n201) );
  IV U220 ( .A(n228), .Z(n78) );
  MUX U221 ( .IN0(n829), .IN1(n79), .SEL(n705), .F(n823) );
  IV U222 ( .A(n704), .Z(n79) );
  XOR U223 ( .A(n888), .B(n880), .Z(n816) );
  XOR U224 ( .A(n993), .B(n985), .Z(n810) );
  MUX U225 ( .IN0(n80), .IN1(n773), .SEL(n772), .F(n746) );
  IV U226 ( .A(n771), .Z(n80) );
  MUX U227 ( .IN0(n81), .IN1(n759), .SEL(n760), .F(n743) );
  IV U228 ( .A(n761), .Z(n81) );
  MUX U229 ( .IN0(n278), .IN1(\_MAC/_MULT/MULT/S[2][1][0] ), .SEL(n1243), .F(
        n247) );
  XNOR U230 ( .A(n184), .B(n183), .Z(n175) );
  MUX U231 ( .IN0(n155), .IN1(\_MAC/_MULT/MULT/S[2][1][5] ), .SEL(n1248), .F(
        n143) );
  MUX U232 ( .IN0(n82), .IN1(n152), .SEL(n153), .F(n132) );
  IV U233 ( .A(n154), .Z(n82) );
  XNOR U234 ( .A(n728), .B(n727), .Z(n725) );
  MUX U235 ( .IN0(n519), .IN1(n332), .SEL(n331), .F(n507) );
  MUX U236 ( .IN0(n416), .IN1(n83), .SEL(n329), .F(n399) );
  IV U237 ( .A(n327), .Z(n83) );
  MUX U238 ( .IN0(n84), .IN1(n1107), .SEL(n1108), .F(n1157) );
  IV U239 ( .A(n1177), .Z(n84) );
  MUX U240 ( .IN0(n309), .IN1(n314), .SEL(n310), .F(n301) );
  MUX U241 ( .IN0(n586), .IN1(n596), .SEL(n588), .F(n446) );
  MUX U242 ( .IN0(n472), .IN1(n300), .SEL(n299), .F(n461) );
  XOR U243 ( .A(n637), .B(n638), .Z(n582) );
  MUX U244 ( .IN0(n1081), .IN1(n1083), .SEL(n1082), .F(n1077) );
  MUX U245 ( .IN0(n350), .IN1(n85), .SEL(n289), .F(n261) );
  IV U246 ( .A(n287), .Z(n85) );
  MUX U247 ( .IN0(n836), .IN1(n1045), .SEL(n837), .F(n1034) );
  MUX U248 ( .IN0(n860), .IN1(n801), .SEL(n802), .F(n86) );
  IV U249 ( .A(n86), .Z(n850) );
  MUX U250 ( .IN0(n255), .IN1(n87), .SEL(n256), .F(n226) );
  IV U251 ( .A(n257), .Z(n87) );
  XOR U252 ( .A(n921), .B(n913), .Z(n834) );
  XNOR U253 ( .A(n176), .B(n160), .Z(n163) );
  MUX U254 ( .IN0(n823), .IN1(n88), .SEL(n703), .F(n817) );
  IV U255 ( .A(n702), .Z(n88) );
  MUX U256 ( .IN0(n89), .IN1(n168), .SEL(n169), .F(n152) );
  IV U257 ( .A(n170), .Z(n89) );
  XNOR U258 ( .A(n980), .B(n974), .Z(n804) );
  MUX U259 ( .IN0(n90), .IN1(n790), .SEL(n791), .F(n769) );
  IV U260 ( .A(n792), .Z(n90) );
  MUX U261 ( .IN0(n247), .IN1(\_MAC/_MULT/MULT/S[2][1][1] ), .SEL(n1244), .F(
        n219) );
  MUX U262 ( .IN0(n175), .IN1(n173), .SEL(n174), .F(n91) );
  IV U263 ( .A(n91), .Z(n158) );
  MUX U264 ( .IN0(n143), .IN1(\_MAC/_MULT/MULT/S[2][1][6] ), .SEL(n1249), .F(
        n92) );
  IV U265 ( .A(n92), .Z(n128) );
  XNOR U266 ( .A(n797), .B(n798), .Z(n692) );
  XNOR U267 ( .A(n783), .B(n782), .Z(n773) );
  XNOR U268 ( .A(n757), .B(n756), .Z(n748) );
  XNOR U269 ( .A(n740), .B(n739), .Z(n733) );
  MUX U270 ( .IN0(n728), .IN1(n93), .SEL(n727), .F(n723) );
  IV U271 ( .A(n726), .Z(n93) );
  MUX U272 ( .IN0(n507), .IN1(n324), .SEL(n323), .F(n495) );
  MUX U273 ( .IN0(n399), .IN1(n94), .SEL(n321), .F(n384) );
  IV U274 ( .A(n319), .Z(n94) );
  MUX U275 ( .IN0(n95), .IN1(n375), .SEL(n376), .F(n364) );
  IV U276 ( .A(n377), .Z(n95) );
  MUX U277 ( .IN0(n301), .IN1(n306), .SEL(n302), .F(n293) );
  XOR U278 ( .A(n649), .B(n632), .Z(n583) );
  MUX U279 ( .IN0(n96), .IN1(n885), .SEL(n886), .F(n873) );
  IV U280 ( .A(n887), .Z(n96) );
  MUX U281 ( .IN0(n97), .IN1(n216), .SEL(n217), .F(n187) );
  IV U282 ( .A(n218), .Z(n97) );
  MUX U283 ( .IN0(n261), .IN1(n263), .SEL(n262), .F(n98) );
  IV U284 ( .A(n98), .Z(n229) );
  MUX U285 ( .IN0(n824), .IN1(n1023), .SEL(n825), .F(n1012) );
  MUX U286 ( .IN0(n905), .IN1(n827), .SEL(n828), .F(n894) );
  MUX U287 ( .IN0(n847), .IN1(n99), .SEL(n848), .F(n841) );
  IV U288 ( .A(n849), .Z(n99) );
  XNOR U289 ( .A(n264), .B(n236), .Z(n240) );
  MUX U290 ( .IN0(n100), .IN1(n203), .SEL(n202), .F(n173) );
  IV U291 ( .A(n201), .Z(n100) );
  MUX U292 ( .IN0(n811), .IN1(n101), .SEL(n699), .F(n805) );
  IV U293 ( .A(n698), .Z(n101) );
  XOR U294 ( .A(n865), .B(n858), .Z(n802) );
  XNOR U295 ( .A(n956), .B(n778), .Z(n782) );
  XNOR U296 ( .A(n830), .B(n831), .Z(n704) );
  MUX U297 ( .IN0(n219), .IN1(\_MAC/_MULT/MULT/S[2][1][2] ), .SEL(n1245), .F(
        n102) );
  IV U298 ( .A(n102), .Z(n190) );
  XNOR U299 ( .A(n164), .B(n163), .Z(n157) );
  MUX U300 ( .IN0(n746), .IN1(n748), .SEL(n747), .F(n103) );
  IV U301 ( .A(n103), .Z(n734) );
  XNOR U302 ( .A(n128), .B(n141), .Z(n129) );
  MUX U303 ( .IN0(n104), .IN1(n730), .SEL(n731), .F(n710) );
  IV U304 ( .A(n732), .Z(n104) );
  MUX U305 ( .IN0(n105), .IN1(n582), .SEL(n583), .F(n623) );
  IV U306 ( .A(n639), .Z(n105) );
  MUX U307 ( .IN0(n555), .IN1(n557), .SEL(n556), .F(n552) );
  MUX U308 ( .IN0(n495), .IN1(n316), .SEL(n315), .F(n483) );
  MUX U309 ( .IN0(n384), .IN1(n106), .SEL(n313), .F(n373) );
  IV U310 ( .A(n311), .Z(n106) );
  MUX U311 ( .IN0(n578), .IN1(n602), .SEL(n580), .F(n438) );
  XOR U312 ( .A(n1175), .B(n1176), .Z(n1107) );
  MUX U313 ( .IN0(n293), .IN1(n298), .SEL(n294), .F(n285) );
  XOR U314 ( .A(n584), .B(n449), .Z(n453) );
  MUX U315 ( .IN0(n940), .IN1(n845), .SEL(n846), .F(n927) );
  XNOR U316 ( .A(n547), .B(n546), .Z(n343) );
  MUX U317 ( .IN0(n229), .IN1(n258), .SEL(n231), .F(n195) );
  XNOR U318 ( .A(n204), .B(n178), .Z(n183) );
  XOR U319 ( .A(n899), .B(n891), .Z(n822) );
  XNOR U320 ( .A(n749), .B(n736), .Z(n739) );
  XNOR U321 ( .A(n1069), .B(n1068), .Z(n849) );
  XNOR U322 ( .A(n272), .B(n271), .Z(n257) );
  XNOR U323 ( .A(n842), .B(n843), .Z(n708) );
  XNOR U324 ( .A(n241), .B(n240), .Z(n228) );
  XNOR U325 ( .A(n836), .B(n837), .Z(n706) );
  XNOR U326 ( .A(n213), .B(n212), .Z(n203) );
  XNOR U327 ( .A(n824), .B(n825), .Z(n702) );
  MUX U328 ( .IN0(n107), .IN1(\_MAC/_MULT/MULT/S[2][1][3] ), .SEL(n1246), .F(
        n171) );
  IV U329 ( .A(n190), .Z(n107) );
  XNOR U330 ( .A(n818), .B(n819), .Z(n700) );
  XNOR U331 ( .A(n149), .B(n148), .Z(n145) );
  XNOR U332 ( .A(n812), .B(n813), .Z(n698) );
  XNOR U333 ( .A(n803), .B(n804), .Z(n694) );
  XOR U334 ( .A(n746), .B(n769), .Z(n762) );
  MUX U335 ( .IN0(n108), .IN1(n743), .SEL(n744), .F(n730) );
  IV U336 ( .A(n745), .Z(n108) );
  MUX U337 ( .IN0(n109), .IN1(\_MAC/_MULT/MULT/S[2][1][7] ), .SEL(n1250), .F(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[8] ) );
  IV U338 ( .A(n128), .Z(n109) );
  XNOR U339 ( .A(n718), .B(n714), .Z(\_MAC/_MULT/MULT/S[2][1][14] ) );
  AND U340 ( .A(n110), .B(n111), .Z(n1255) );
  XOR U341 ( .A(\_MAC/_MULT/AX__[5] ), .B(\_MAC/_MULT/AX_[5] ), .Z(n111) );
  AND U342 ( .A(n110), .B(n112), .Z(n1254) );
  XOR U343 ( .A(\_MAC/_MULT/AX__[6] ), .B(\_MAC/_MULT/AX_[6] ), .Z(n112) );
  AND U344 ( .A(n110), .B(n113), .Z(n1253) );
  XOR U345 ( .A(\_MAC/_MULT/AX__[7] ), .B(\_MAC/_MULT/AX_[7] ), .Z(n113) );
  AND U346 ( .A(n110), .B(n114), .Z(n1266) );
  XOR U347 ( .A(\_MAC/_MULT/AX__[0] ), .B(\_MAC/_MULT/AX_[0] ), .Z(n114) );
  AND U348 ( .A(n110), .B(n115), .Z(n1252) );
  XOR U349 ( .A(\_MAC/_MULT/AX__[8] ), .B(\_MAC/_MULT/AX_[8] ), .Z(n115) );
  AND U350 ( .A(n110), .B(n116), .Z(n1265) );
  XOR U351 ( .A(\_MAC/_MULT/AX__[10] ), .B(\_MAC/_MULT/AX_[10] ), .Z(n116) );
  AND U352 ( .A(n110), .B(n117), .Z(n1264) );
  XOR U353 ( .A(\_MAC/_MULT/AX__[11] ), .B(\_MAC/_MULT/AX_[11] ), .Z(n117) );
  AND U354 ( .A(n110), .B(n118), .Z(n1263) );
  XOR U355 ( .A(\_MAC/_MULT/AX__[12] ), .B(\_MAC/_MULT/AX_[12] ), .Z(n118) );
  AND U356 ( .A(n110), .B(n119), .Z(n1262) );
  XOR U357 ( .A(\_MAC/_MULT/AX__[13] ), .B(\_MAC/_MULT/AX_[13] ), .Z(n119) );
  AND U358 ( .A(n110), .B(n120), .Z(n1261) );
  XOR U359 ( .A(\_MAC/_MULT/AX__[14] ), .B(\_MAC/_MULT/AX_[14] ), .Z(n120) );
  AND U360 ( .A(n110), .B(n121), .Z(n1260) );
  XOR U361 ( .A(\_MAC/_MULT/AX__[15] ), .B(\_MAC/_MULT/AX_[15] ), .Z(n121) );
  AND U362 ( .A(n110), .B(n122), .Z(n1259) );
  XOR U363 ( .A(\_MAC/_MULT/AX__[1] ), .B(\_MAC/_MULT/AX_[1] ), .Z(n122) );
  AND U364 ( .A(n110), .B(n123), .Z(n1258) );
  XOR U365 ( .A(\_MAC/_MULT/AX__[2] ), .B(\_MAC/_MULT/AX_[2] ), .Z(n123) );
  AND U366 ( .A(n110), .B(n124), .Z(n1257) );
  XOR U367 ( .A(\_MAC/_MULT/AX__[3] ), .B(\_MAC/_MULT/AX_[3] ), .Z(n124) );
  AND U368 ( .A(n110), .B(n125), .Z(n1256) );
  XOR U369 ( .A(\_MAC/_MULT/AX__[4] ), .B(\_MAC/_MULT/AX_[4] ), .Z(n125) );
  AND U370 ( .A(n110), .B(n126), .Z(n1251) );
  XOR U371 ( .A(\_MAC/_MULT/AX__[9] ), .B(\_MAC/_MULT/AX_[9] ), .Z(n126) );
  XNOR U372 ( .A(n127), .B(g_input[15]), .Z(n110) );
  AND U373 ( .A(\_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[14] ), .B(
        \_MAC/_MULT/MULT/S[2][1][14] ), .Z(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[15] ) );
  AND U374 ( .A(\_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[13] ), .B(
        \_MAC/_MULT/MULT/S[2][1][13] ), .Z(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[14] ) );
  AND U375 ( .A(\_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[12] ), .B(
        \_MAC/_MULT/MULT/S[2][1][12] ), .Z(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[13] ) );
  AND U376 ( .A(\_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[11] ), .B(
        \_MAC/_MULT/MULT/S[2][1][11] ), .Z(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[12] ) );
  AND U377 ( .A(\_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[10] ), .B(
        \_MAC/_MULT/MULT/S[2][1][10] ), .Z(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[11] ) );
  AND U378 ( .A(\_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[9] ), .B(
        \_MAC/_MULT/MULT/S[2][1][9] ), .Z(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[10] ) );
  AND U379 ( .A(\_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[8] ), .B(
        \_MAC/_MULT/MULT/S[2][1][8] ), .Z(
        \_MAC/_MULT/MULT/col[2].row[0]._SHIFT_ADD/_ADD/C[9] ) );
  XOR U380 ( .A(n129), .B(n130), .Z(n1250) );
  XOR U381 ( .A(n131), .B(n132), .Z(n130) );
  AND U382 ( .A(n133), .B(n134), .Z(n131) );
  OR U383 ( .A(n135), .B(n136), .Z(n134) );
  AND U384 ( .A(n137), .B(n138), .Z(n133) );
  NAND U385 ( .A(n139), .B(n132), .Z(n138) );
  OR U386 ( .A(n140), .B(n141), .Z(n137) );
  XNOR U387 ( .A(n144), .B(n143), .Z(n1249) );
  XNOR U388 ( .A(n136), .B(n135), .Z(n144) );
  OR U389 ( .A(n145), .B(n146), .Z(n135) );
  XNOR U390 ( .A(n140), .B(n142), .Z(n136) );
  IV U391 ( .A(n141), .Z(n142) );
  XNOR U392 ( .A(n132), .B(n139), .Z(n140) );
  NANDN U393 ( .B(n150), .A(n151), .Z(n139) );
  XNOR U394 ( .A(n156), .B(n155), .Z(n1248) );
  XNOR U395 ( .A(n145), .B(n146), .Z(n156) );
  NANDN U396 ( .B(n157), .A(n158), .Z(n146) );
  XNOR U397 ( .A(n147), .B(n159), .Z(n148) );
  NOR U398 ( .A(n160), .B(n161), .Z(n159) );
  XNOR U399 ( .A(n153), .B(n154), .Z(n149) );
  NAND U400 ( .A(n151), .B(n165), .Z(n154) );
  XNOR U401 ( .A(n152), .B(n166), .Z(n153) );
  NOR U402 ( .A(n150), .B(n167), .Z(n166) );
  XNOR U403 ( .A(n172), .B(n171), .Z(n1247) );
  XOR U404 ( .A(n157), .B(n158), .Z(n172) );
  XOR U405 ( .A(n180), .B(n161), .Z(n176) );
  NANDN U406 ( .B(n150), .A(n181), .Z(n161) );
  IV U407 ( .A(n162), .Z(n180) );
  XNOR U408 ( .A(n169), .B(n170), .Z(n164) );
  NAND U409 ( .A(n151), .B(n185), .Z(n170) );
  XNOR U410 ( .A(n168), .B(n186), .Z(n169) );
  ANDN U411 ( .A(n165), .B(n167), .Z(n186) );
  XNOR U412 ( .A(n191), .B(n190), .Z(n1246) );
  XOR U413 ( .A(n175), .B(n174), .Z(n191) );
  XNOR U414 ( .A(n192), .B(n193), .Z(n174) );
  XOR U415 ( .A(n194), .B(n195), .Z(n193) );
  AND U416 ( .A(n196), .B(n197), .Z(n194) );
  NAND U417 ( .A(n198), .B(n199), .Z(n197) );
  NANDN U418 ( .B(n200), .A(n195), .Z(n196) );
  XNOR U419 ( .A(n177), .B(n205), .Z(n178) );
  ANDN U420 ( .A(n206), .B(n150), .Z(n205) );
  XOR U421 ( .A(n210), .B(n179), .Z(n204) );
  NAND U422 ( .A(n181), .B(n165), .Z(n179) );
  IV U423 ( .A(n182), .Z(n210) );
  XNOR U424 ( .A(n188), .B(n189), .Z(n184) );
  NAND U425 ( .A(n151), .B(n214), .Z(n189) );
  XNOR U426 ( .A(n187), .B(n215), .Z(n188) );
  ANDN U427 ( .A(n185), .B(n167), .Z(n215) );
  XNOR U428 ( .A(n220), .B(n219), .Z(n1245) );
  XOR U429 ( .A(n203), .B(n202), .Z(n220) );
  XNOR U430 ( .A(n221), .B(n200), .Z(n202) );
  XNOR U431 ( .A(n199), .B(n198), .Z(n200) );
  NANDN U432 ( .B(n150), .A(n222), .Z(n198) );
  XNOR U433 ( .A(n195), .B(n201), .Z(n221) );
  XNOR U434 ( .A(n229), .B(n232), .Z(n231) );
  XNOR U435 ( .A(n207), .B(n234), .Z(n208) );
  AND U436 ( .A(n165), .B(n206), .Z(n234) );
  XOR U437 ( .A(n238), .B(n209), .Z(n233) );
  NAND U438 ( .A(n181), .B(n185), .Z(n209) );
  IV U439 ( .A(n211), .Z(n238) );
  XNOR U440 ( .A(n217), .B(n218), .Z(n213) );
  NAND U441 ( .A(n151), .B(n242), .Z(n218) );
  XNOR U442 ( .A(n216), .B(n243), .Z(n217) );
  ANDN U443 ( .A(n214), .B(n167), .Z(n243) );
  XNOR U444 ( .A(n248), .B(n247), .Z(n1244) );
  XOR U445 ( .A(n228), .B(n227), .Z(n248) );
  XOR U446 ( .A(n249), .B(n232), .Z(n227) );
  XNOR U447 ( .A(n224), .B(n225), .Z(n232) );
  NAND U448 ( .A(n222), .B(n165), .Z(n225) );
  XNOR U449 ( .A(n223), .B(n250), .Z(n224) );
  ANDN U450 ( .A(n251), .B(n150), .Z(n250) );
  XNOR U451 ( .A(n230), .B(n226), .Z(n249) );
  XOR U452 ( .A(n229), .B(n258), .Z(n230) );
  NOR U453 ( .A(n259), .B(n260), .Z(n258) );
  XNOR U454 ( .A(n235), .B(n265), .Z(n236) );
  AND U455 ( .A(n185), .B(n206), .Z(n265) );
  XOR U456 ( .A(n269), .B(n237), .Z(n264) );
  NAND U457 ( .A(n181), .B(n214), .Z(n237) );
  IV U458 ( .A(n239), .Z(n269) );
  XNOR U459 ( .A(n245), .B(n246), .Z(n241) );
  NANDN U460 ( .B(n273), .A(n151), .Z(n246) );
  XNOR U461 ( .A(n244), .B(n274), .Z(n245) );
  ANDN U462 ( .A(n242), .B(n167), .Z(n274) );
  XNOR U463 ( .A(n279), .B(n278), .Z(n1243) );
  XOR U464 ( .A(n257), .B(n256), .Z(n279) );
  XOR U465 ( .A(n280), .B(n263), .Z(n256) );
  XNOR U466 ( .A(n253), .B(n254), .Z(n263) );
  NAND U467 ( .A(n222), .B(n185), .Z(n254) );
  XNOR U468 ( .A(n252), .B(n281), .Z(n253) );
  AND U469 ( .A(n165), .B(n251), .Z(n281) );
  XNOR U470 ( .A(n262), .B(n255), .Z(n280) );
  XOR U471 ( .A(n287), .B(n288), .Z(n286) );
  XOR U472 ( .A(n285), .B(n289), .Z(n288) );
  XNOR U473 ( .A(n291), .B(n292), .Z(n290) );
  XOR U474 ( .A(n295), .B(n296), .Z(n294) );
  XOR U475 ( .A(n293), .B(n297), .Z(n296) );
  XNOR U476 ( .A(n299), .B(n300), .Z(n298) );
  XOR U477 ( .A(n303), .B(n304), .Z(n302) );
  XOR U478 ( .A(n301), .B(n305), .Z(n304) );
  XNOR U479 ( .A(n307), .B(n308), .Z(n306) );
  XOR U480 ( .A(n311), .B(n312), .Z(n310) );
  XOR U481 ( .A(n309), .B(n313), .Z(n312) );
  XNOR U482 ( .A(n315), .B(n316), .Z(n314) );
  XOR U483 ( .A(n319), .B(n320), .Z(n318) );
  XOR U484 ( .A(n317), .B(n321), .Z(n320) );
  XNOR U485 ( .A(n323), .B(n324), .Z(n322) );
  XOR U486 ( .A(n327), .B(n328), .Z(n326) );
  XOR U487 ( .A(n325), .B(n329), .Z(n328) );
  XNOR U488 ( .A(n331), .B(n332), .Z(n330) );
  XOR U489 ( .A(n335), .B(n336), .Z(n334) );
  XOR U490 ( .A(n333), .B(n337), .Z(n336) );
  XNOR U491 ( .A(n339), .B(n340), .Z(n338) );
  XOR U492 ( .A(n348), .B(n260), .Z(n344) );
  NANDN U493 ( .B(n150), .A(n349), .Z(n260) );
  IV U494 ( .A(n261), .Z(n348) );
  NAND U495 ( .A(n222), .B(n214), .Z(n284) );
  XNOR U496 ( .A(n282), .B(n351), .Z(n283) );
  AND U497 ( .A(n185), .B(n251), .Z(n351) );
  XNOR U498 ( .A(n345), .B(n356), .Z(n346) );
  ANDN U499 ( .A(n357), .B(n150), .Z(n356) );
  XOR U500 ( .A(n361), .B(n347), .Z(n355) );
  NAND U501 ( .A(n349), .B(n165), .Z(n347) );
  IV U502 ( .A(n350), .Z(n361) );
  NAND U503 ( .A(n222), .B(n242), .Z(n354) );
  XNOR U504 ( .A(n352), .B(n363), .Z(n353) );
  AND U505 ( .A(n214), .B(n251), .Z(n363) );
  XNOR U506 ( .A(n358), .B(n368), .Z(n359) );
  AND U507 ( .A(n165), .B(n357), .Z(n368) );
  XOR U508 ( .A(n372), .B(n360), .Z(n367) );
  NAND U509 ( .A(n349), .B(n185), .Z(n360) );
  IV U510 ( .A(n362), .Z(n372) );
  NANDN U511 ( .B(n273), .A(n222), .Z(n366) );
  XNOR U512 ( .A(n364), .B(n374), .Z(n365) );
  AND U513 ( .A(n242), .B(n251), .Z(n374) );
  XNOR U514 ( .A(n369), .B(n379), .Z(n370) );
  AND U515 ( .A(n185), .B(n357), .Z(n379) );
  XOR U516 ( .A(n383), .B(n371), .Z(n378) );
  NAND U517 ( .A(n349), .B(n214), .Z(n371) );
  IV U518 ( .A(n373), .Z(n383) );
  NANDN U519 ( .B(n385), .A(n222), .Z(n377) );
  XNOR U520 ( .A(n375), .B(n386), .Z(n376) );
  ANDN U521 ( .A(n251), .B(n273), .Z(n386) );
  XOR U522 ( .A(n387), .B(n388), .Z(n375) );
  ANDN U523 ( .A(n389), .B(n390), .Z(n388) );
  XNOR U524 ( .A(n391), .B(n387), .Z(n389) );
  XNOR U525 ( .A(n392), .B(n393), .Z(n313) );
  IV U526 ( .A(n381), .Z(n393) );
  XNOR U527 ( .A(n380), .B(n394), .Z(n381) );
  AND U528 ( .A(n214), .B(n357), .Z(n394) );
  XOR U529 ( .A(n398), .B(n382), .Z(n392) );
  NAND U530 ( .A(n349), .B(n242), .Z(n382) );
  IV U531 ( .A(n384), .Z(n398) );
  NAND U532 ( .A(n222), .B(n400), .Z(n391) );
  XNOR U533 ( .A(n387), .B(n401), .Z(n390) );
  ANDN U534 ( .A(n251), .B(n385), .Z(n401) );
  XOR U535 ( .A(n402), .B(n403), .Z(n387) );
  ANDN U536 ( .A(n404), .B(n405), .Z(n403) );
  XNOR U537 ( .A(n406), .B(n402), .Z(n404) );
  XNOR U538 ( .A(n407), .B(n408), .Z(n321) );
  IV U539 ( .A(n396), .Z(n408) );
  XNOR U540 ( .A(n395), .B(n409), .Z(n396) );
  AND U541 ( .A(n242), .B(n357), .Z(n409) );
  XOR U542 ( .A(n410), .B(n411), .Z(n395) );
  ANDN U543 ( .A(n412), .B(n413), .Z(n411) );
  XNOR U544 ( .A(n414), .B(n410), .Z(n412) );
  XOR U545 ( .A(n415), .B(n397), .Z(n407) );
  NANDN U546 ( .B(n273), .A(n349), .Z(n397) );
  IV U547 ( .A(n399), .Z(n415) );
  XNOR U548 ( .A(n417), .B(n406), .Z(n327) );
  NAND U549 ( .A(n222), .B(n418), .Z(n406) );
  IV U550 ( .A(n405), .Z(n417) );
  XNOR U551 ( .A(n402), .B(n419), .Z(n405) );
  AND U552 ( .A(n400), .B(n251), .Z(n419) );
  XOR U553 ( .A(n420), .B(n421), .Z(n402) );
  ANDN U554 ( .A(n422), .B(n423), .Z(n421) );
  XNOR U555 ( .A(n424), .B(n420), .Z(n422) );
  XNOR U556 ( .A(n425), .B(n426), .Z(n329) );
  IV U557 ( .A(n413), .Z(n426) );
  XNOR U558 ( .A(n410), .B(n427), .Z(n413) );
  ANDN U559 ( .A(n357), .B(n273), .Z(n427) );
  XOR U560 ( .A(n428), .B(n429), .Z(n410) );
  ANDN U561 ( .A(n430), .B(n431), .Z(n429) );
  XNOR U562 ( .A(n432), .B(n428), .Z(n430) );
  XOR U563 ( .A(n433), .B(n414), .Z(n425) );
  NANDN U564 ( .B(n385), .A(n349), .Z(n414) );
  IV U565 ( .A(n416), .Z(n433) );
  XNOR U566 ( .A(n435), .B(n424), .Z(n335) );
  NAND U567 ( .A(n222), .B(n436), .Z(n424) );
  IV U568 ( .A(n423), .Z(n435) );
  XNOR U569 ( .A(n420), .B(n437), .Z(n423) );
  AND U570 ( .A(n418), .B(n251), .Z(n437) );
  XOR U571 ( .A(n438), .B(n439), .Z(n420) );
  ANDN U572 ( .A(n440), .B(n441), .Z(n439) );
  XNOR U573 ( .A(n442), .B(n438), .Z(n440) );
  XNOR U574 ( .A(n443), .B(n444), .Z(n337) );
  IV U575 ( .A(n431), .Z(n444) );
  XNOR U576 ( .A(n428), .B(n445), .Z(n431) );
  ANDN U577 ( .A(n357), .B(n385), .Z(n445) );
  XOR U578 ( .A(n446), .B(n447), .Z(n428) );
  ANDN U579 ( .A(n448), .B(n449), .Z(n447) );
  XNOR U580 ( .A(n450), .B(n446), .Z(n448) );
  XOR U581 ( .A(n451), .B(n432), .Z(n443) );
  NAND U582 ( .A(n349), .B(n400), .Z(n432) );
  IV U583 ( .A(n434), .Z(n451) );
  XNOR U584 ( .A(n266), .B(n456), .Z(n267) );
  AND U585 ( .A(n214), .B(n206), .Z(n456) );
  XOR U586 ( .A(n460), .B(n268), .Z(n455) );
  NAND U587 ( .A(n181), .B(n242), .Z(n268) );
  IV U588 ( .A(n270), .Z(n460) );
  XOR U589 ( .A(n462), .B(n463), .Z(n292) );
  XNOR U590 ( .A(n457), .B(n465), .Z(n458) );
  AND U591 ( .A(n242), .B(n206), .Z(n465) );
  XOR U592 ( .A(n466), .B(n467), .Z(n457) );
  ANDN U593 ( .A(n468), .B(n469), .Z(n467) );
  XNOR U594 ( .A(n470), .B(n466), .Z(n468) );
  XOR U595 ( .A(n471), .B(n459), .Z(n464) );
  NANDN U596 ( .B(n273), .A(n181), .Z(n459) );
  IV U597 ( .A(n461), .Z(n471) );
  XOR U598 ( .A(n473), .B(n474), .Z(n300) );
  XNOR U599 ( .A(n466), .B(n476), .Z(n469) );
  ANDN U600 ( .A(n206), .B(n273), .Z(n476) );
  XOR U601 ( .A(n477), .B(n478), .Z(n466) );
  ANDN U602 ( .A(n479), .B(n480), .Z(n478) );
  XNOR U603 ( .A(n481), .B(n477), .Z(n479) );
  XOR U604 ( .A(n482), .B(n470), .Z(n475) );
  NANDN U605 ( .B(n385), .A(n181), .Z(n470) );
  IV U606 ( .A(n472), .Z(n482) );
  XOR U607 ( .A(n484), .B(n485), .Z(n308) );
  XNOR U608 ( .A(n486), .B(n487), .Z(n307) );
  IV U609 ( .A(n480), .Z(n487) );
  XNOR U610 ( .A(n477), .B(n488), .Z(n480) );
  ANDN U611 ( .A(n206), .B(n385), .Z(n488) );
  XOR U612 ( .A(n489), .B(n490), .Z(n477) );
  ANDN U613 ( .A(n491), .B(n492), .Z(n490) );
  XNOR U614 ( .A(n493), .B(n489), .Z(n491) );
  XOR U615 ( .A(n494), .B(n481), .Z(n486) );
  NAND U616 ( .A(n181), .B(n400), .Z(n481) );
  IV U617 ( .A(n483), .Z(n494) );
  XOR U618 ( .A(n496), .B(n497), .Z(n316) );
  XNOR U619 ( .A(n498), .B(n499), .Z(n315) );
  IV U620 ( .A(n492), .Z(n499) );
  XNOR U621 ( .A(n489), .B(n500), .Z(n492) );
  AND U622 ( .A(n400), .B(n206), .Z(n500) );
  XOR U623 ( .A(n501), .B(n502), .Z(n489) );
  ANDN U624 ( .A(n503), .B(n504), .Z(n502) );
  XNOR U625 ( .A(n505), .B(n501), .Z(n503) );
  XOR U626 ( .A(n506), .B(n493), .Z(n498) );
  NAND U627 ( .A(n181), .B(n418), .Z(n493) );
  IV U628 ( .A(n495), .Z(n506) );
  XOR U629 ( .A(n508), .B(n509), .Z(n324) );
  XNOR U630 ( .A(n510), .B(n511), .Z(n323) );
  IV U631 ( .A(n504), .Z(n511) );
  XNOR U632 ( .A(n501), .B(n512), .Z(n504) );
  AND U633 ( .A(n418), .B(n206), .Z(n512) );
  XOR U634 ( .A(n513), .B(n514), .Z(n501) );
  ANDN U635 ( .A(n515), .B(n516), .Z(n514) );
  XNOR U636 ( .A(n517), .B(n513), .Z(n515) );
  XOR U637 ( .A(n518), .B(n505), .Z(n510) );
  NAND U638 ( .A(n181), .B(n436), .Z(n505) );
  IV U639 ( .A(n507), .Z(n518) );
  XOR U640 ( .A(n520), .B(n521), .Z(n332) );
  XNOR U641 ( .A(n522), .B(n523), .Z(n331) );
  IV U642 ( .A(n516), .Z(n523) );
  XNOR U643 ( .A(n513), .B(n524), .Z(n516) );
  AND U644 ( .A(n436), .B(n206), .Z(n524) );
  XOR U645 ( .A(n525), .B(n526), .Z(n513) );
  ANDN U646 ( .A(n527), .B(n528), .Z(n526) );
  XNOR U647 ( .A(n529), .B(n525), .Z(n527) );
  XOR U648 ( .A(n530), .B(n517), .Z(n522) );
  NAND U649 ( .A(n181), .B(n531), .Z(n517) );
  IV U650 ( .A(n519), .Z(n530) );
  XOR U651 ( .A(n533), .B(n534), .Z(n340) );
  XNOR U652 ( .A(n535), .B(n536), .Z(n339) );
  IV U653 ( .A(n528), .Z(n536) );
  XNOR U654 ( .A(n525), .B(n537), .Z(n528) );
  AND U655 ( .A(n531), .B(n206), .Z(n537) );
  XOR U656 ( .A(n538), .B(n539), .Z(n525) );
  ANDN U657 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U658 ( .A(n542), .B(n538), .Z(n540) );
  XOR U659 ( .A(n543), .B(n529), .Z(n535) );
  NAND U660 ( .A(n181), .B(n544), .Z(n529) );
  IV U661 ( .A(n532), .Z(n543) );
  XNOR U662 ( .A(n276), .B(n277), .Z(n272) );
  NANDN U663 ( .B(n385), .A(n151), .Z(n277) );
  XNOR U664 ( .A(n275), .B(n548), .Z(n276) );
  NOR U665 ( .A(n167), .B(n273), .Z(n548) );
  XNOR U666 ( .A(n463), .B(n549), .Z(n550) );
  NAND U667 ( .A(n151), .B(n400), .Z(n463) );
  XOR U668 ( .A(n549), .B(n551), .Z(n462) );
  NOR U669 ( .A(n167), .B(n385), .Z(n551) );
  XNOR U670 ( .A(n474), .B(n552), .Z(n553) );
  NAND U671 ( .A(n151), .B(n418), .Z(n474) );
  XOR U672 ( .A(n552), .B(n554), .Z(n473) );
  ANDN U673 ( .A(n400), .B(n167), .Z(n554) );
  XNOR U674 ( .A(n485), .B(n555), .Z(n556) );
  NAND U675 ( .A(n151), .B(n436), .Z(n485) );
  XOR U676 ( .A(n555), .B(n557), .Z(n484) );
  ANDN U677 ( .A(n418), .B(n167), .Z(n557) );
  XNOR U678 ( .A(n497), .B(n558), .Z(n559) );
  NAND U679 ( .A(n151), .B(n531), .Z(n497) );
  XOR U680 ( .A(n558), .B(n560), .Z(n496) );
  ANDN U681 ( .A(n436), .B(n167), .Z(n560) );
  XNOR U682 ( .A(n509), .B(n561), .Z(n562) );
  NAND U683 ( .A(n151), .B(n544), .Z(n509) );
  XOR U684 ( .A(n561), .B(n563), .Z(n508) );
  ANDN U685 ( .A(n531), .B(n167), .Z(n563) );
  XOR U686 ( .A(n564), .B(n565), .Z(n561) );
  AND U687 ( .A(n520), .B(n566), .Z(n565) );
  XNOR U688 ( .A(n521), .B(n564), .Z(n566) );
  NAND U689 ( .A(n151), .B(n567), .Z(n521) );
  XOR U690 ( .A(n564), .B(n568), .Z(n520) );
  ANDN U691 ( .A(n544), .B(n167), .Z(n568) );
  XNOR U692 ( .A(n534), .B(n569), .Z(n570) );
  NANDN U693 ( .B(n571), .A(n151), .Z(n534) );
  XOR U694 ( .A(n569), .B(n572), .Z(n533) );
  ANDN U695 ( .A(n567), .B(n167), .Z(n572) );
  XOR U696 ( .A(n343), .B(n342), .Z(n278) );
  XNOR U697 ( .A(n576), .B(n454), .Z(n342) );
  XNOR U698 ( .A(n441), .B(n442), .Z(n454) );
  NAND U699 ( .A(n222), .B(n531), .Z(n442) );
  XNOR U700 ( .A(n438), .B(n577), .Z(n441) );
  AND U701 ( .A(n436), .B(n251), .Z(n577) );
  XNOR U702 ( .A(n581), .B(n578), .Z(n580) );
  XNOR U703 ( .A(n453), .B(n341), .Z(n576) );
  XOR U704 ( .A(n582), .B(n583), .Z(n341) );
  XNOR U705 ( .A(n446), .B(n585), .Z(n449) );
  AND U706 ( .A(n400), .B(n357), .Z(n585) );
  XNOR U707 ( .A(n589), .B(n586), .Z(n588) );
  XOR U708 ( .A(n590), .B(n450), .Z(n584) );
  NAND U709 ( .A(n349), .B(n418), .Z(n450) );
  IV U710 ( .A(n452), .Z(n590) );
  XNOR U711 ( .A(n591), .B(n592), .Z(n452) );
  AND U712 ( .A(n593), .B(n594), .Z(n592) );
  XOR U713 ( .A(n587), .B(n595), .Z(n594) );
  XNOR U714 ( .A(n589), .B(n591), .Z(n595) );
  NAND U715 ( .A(n349), .B(n436), .Z(n589) );
  XOR U716 ( .A(n586), .B(n596), .Z(n587) );
  AND U717 ( .A(n418), .B(n357), .Z(n596) );
  XNOR U718 ( .A(n600), .B(n597), .Z(n599) );
  XOR U719 ( .A(n579), .B(n601), .Z(n593) );
  XNOR U720 ( .A(n581), .B(n591), .Z(n601) );
  NAND U721 ( .A(n222), .B(n544), .Z(n581) );
  XOR U722 ( .A(n578), .B(n602), .Z(n579) );
  AND U723 ( .A(n531), .B(n251), .Z(n602) );
  XNOR U724 ( .A(n606), .B(n603), .Z(n605) );
  XOR U725 ( .A(n607), .B(n608), .Z(n591) );
  AND U726 ( .A(n609), .B(n610), .Z(n608) );
  XOR U727 ( .A(n598), .B(n611), .Z(n610) );
  XNOR U728 ( .A(n600), .B(n607), .Z(n611) );
  NAND U729 ( .A(n349), .B(n531), .Z(n600) );
  XOR U730 ( .A(n597), .B(n612), .Z(n598) );
  AND U731 ( .A(n436), .B(n357), .Z(n612) );
  XNOR U732 ( .A(n616), .B(n613), .Z(n615) );
  XOR U733 ( .A(n604), .B(n617), .Z(n609) );
  XNOR U734 ( .A(n606), .B(n607), .Z(n617) );
  NAND U735 ( .A(n222), .B(n567), .Z(n606) );
  XOR U736 ( .A(n603), .B(n618), .Z(n604) );
  AND U737 ( .A(n544), .B(n251), .Z(n618) );
  XNOR U738 ( .A(n622), .B(n619), .Z(n621) );
  XOR U739 ( .A(n623), .B(n624), .Z(n607) );
  AND U740 ( .A(n625), .B(n626), .Z(n624) );
  XOR U741 ( .A(n614), .B(n627), .Z(n626) );
  XNOR U742 ( .A(n616), .B(n623), .Z(n627) );
  NAND U743 ( .A(n349), .B(n544), .Z(n616) );
  XOR U744 ( .A(n613), .B(n628), .Z(n614) );
  AND U745 ( .A(n531), .B(n357), .Z(n628) );
  XOR U746 ( .A(n629), .B(n630), .Z(n613) );
  ANDN U747 ( .A(n631), .B(n632), .Z(n630) );
  XNOR U748 ( .A(n633), .B(n629), .Z(n631) );
  XOR U749 ( .A(n620), .B(n634), .Z(n625) );
  XNOR U750 ( .A(n622), .B(n623), .Z(n634) );
  NANDN U751 ( .B(n571), .A(n222), .Z(n622) );
  XOR U752 ( .A(n619), .B(n635), .Z(n620) );
  AND U753 ( .A(n567), .B(n251), .Z(n635) );
  NAND U754 ( .A(n222), .B(n640), .Z(n638) );
  XNOR U755 ( .A(n636), .B(n641), .Z(n637) );
  ANDN U756 ( .A(n251), .B(n571), .Z(n641) );
  ANDN U757 ( .A(n642), .B(n643), .Z(n636) );
  NANDN U758 ( .B(n222), .A(n644), .Z(n642) );
  NAND U759 ( .A(n640), .B(n251), .Z(n644) );
  XNOR U760 ( .A(n645), .B(e_input[2]), .Z(n251) );
  NANDN U761 ( .B(n127), .A(n646), .Z(n645) );
  XOR U762 ( .A(e_input[2]), .B(\_MAC/_MULT/X_[2] ), .Z(n646) );
  XNOR U763 ( .A(n647), .B(e_input[3]), .Z(n222) );
  NANDN U764 ( .B(n127), .A(n648), .Z(n647) );
  XOR U765 ( .A(e_input[3]), .B(\_MAC/_MULT/X_[3] ), .Z(n648) );
  XNOR U766 ( .A(n629), .B(n650), .Z(n632) );
  AND U767 ( .A(n544), .B(n357), .Z(n650) );
  XOR U768 ( .A(n653), .B(n651), .Z(n652) );
  AND U769 ( .A(n567), .B(n357), .Z(n653) );
  ANDN U770 ( .A(n349), .B(n571), .Z(n654) );
  XOR U771 ( .A(n655), .B(n656), .Z(n651) );
  ANDN U772 ( .A(n657), .B(n658), .Z(n656) );
  XNOR U773 ( .A(n659), .B(n655), .Z(n657) );
  XOR U774 ( .A(n660), .B(n633), .Z(n649) );
  NAND U775 ( .A(n349), .B(n567), .Z(n633) );
  IV U776 ( .A(n639), .Z(n660) );
  NAND U777 ( .A(n349), .B(n640), .Z(n659) );
  XNOR U778 ( .A(n655), .B(n661), .Z(n658) );
  ANDN U779 ( .A(n357), .B(n571), .Z(n661) );
  ANDN U780 ( .A(n662), .B(n643), .Z(n655) );
  NANDN U781 ( .B(n349), .A(n663), .Z(n662) );
  NAND U782 ( .A(n640), .B(n357), .Z(n663) );
  XNOR U783 ( .A(n664), .B(e_input[0]), .Z(n357) );
  NANDN U784 ( .B(n127), .A(n665), .Z(n664) );
  XOR U785 ( .A(e_input[0]), .B(\_MAC/_MULT/X_[0] ), .Z(n665) );
  XNOR U786 ( .A(n666), .B(e_input[1]), .Z(n349) );
  NANDN U787 ( .B(n127), .A(n667), .Z(n666) );
  XOR U788 ( .A(e_input[1]), .B(\_MAC/_MULT/X_[1] ), .Z(n667) );
  XNOR U789 ( .A(n538), .B(n669), .Z(n541) );
  AND U790 ( .A(n544), .B(n206), .Z(n669) );
  XOR U791 ( .A(n672), .B(n670), .Z(n671) );
  AND U792 ( .A(n567), .B(n206), .Z(n672) );
  ANDN U793 ( .A(n181), .B(n571), .Z(n673) );
  XOR U794 ( .A(n677), .B(n542), .Z(n668) );
  NAND U795 ( .A(n181), .B(n567), .Z(n542) );
  IV U796 ( .A(n545), .Z(n677) );
  NAND U797 ( .A(n181), .B(n640), .Z(n676) );
  XNOR U798 ( .A(n674), .B(n678), .Z(n675) );
  ANDN U799 ( .A(n206), .B(n571), .Z(n678) );
  ANDN U800 ( .A(n679), .B(n643), .Z(n674) );
  NANDN U801 ( .B(n181), .A(n680), .Z(n679) );
  NAND U802 ( .A(n640), .B(n206), .Z(n680) );
  XNOR U803 ( .A(n681), .B(e_input[4]), .Z(n206) );
  NANDN U804 ( .B(n127), .A(n682), .Z(n681) );
  XOR U805 ( .A(e_input[4]), .B(\_MAC/_MULT/X_[4] ), .Z(n682) );
  XNOR U806 ( .A(n683), .B(e_input[5]), .Z(n181) );
  NANDN U807 ( .B(n127), .A(n684), .Z(n683) );
  XOR U808 ( .A(e_input[5]), .B(\_MAC/_MULT/X_[5] ), .Z(n684) );
  XNOR U809 ( .A(n574), .B(n575), .Z(n547) );
  NAND U810 ( .A(n151), .B(n640), .Z(n575) );
  XNOR U811 ( .A(n573), .B(n685), .Z(n574) );
  NOR U812 ( .A(n167), .B(n571), .Z(n685) );
  ANDN U813 ( .A(n686), .B(n643), .Z(n573) );
  NANDN U814 ( .B(n151), .A(n687), .Z(n686) );
  NANDN U815 ( .B(n167), .A(n640), .Z(n687) );
  XOR U816 ( .A(n688), .B(e_input[6]), .Z(n167) );
  NANDN U817 ( .B(n127), .A(n689), .Z(n688) );
  XOR U818 ( .A(e_input[6]), .B(\_MAC/_MULT/X_[6] ), .Z(n689) );
  XNOR U819 ( .A(n690), .B(e_input[7]), .Z(n151) );
  NANDN U820 ( .B(n127), .A(n691), .Z(n690) );
  XOR U821 ( .A(e_input[7]), .B(\_MAC/_MULT/X_[7] ), .Z(n691) );
  XNOR U822 ( .A(n692), .B(n693), .Z(\_MAC/_MULT/MULT/S[2][1][9] ) );
  XNOR U823 ( .A(n694), .B(n695), .Z(\_MAC/_MULT/MULT/S[2][1][8] ) );
  XOR U824 ( .A(n696), .B(n697), .Z(\_MAC/_MULT/MULT/S[2][1][7] ) );
  XNOR U825 ( .A(n698), .B(n699), .Z(\_MAC/_MULT/MULT/S[2][1][6] ) );
  XNOR U826 ( .A(n700), .B(n701), .Z(\_MAC/_MULT/MULT/S[2][1][5] ) );
  XNOR U827 ( .A(n702), .B(n703), .Z(\_MAC/_MULT/MULT/S[2][1][4] ) );
  XNOR U828 ( .A(n704), .B(n705), .Z(\_MAC/_MULT/MULT/S[2][1][3] ) );
  XNOR U829 ( .A(n706), .B(n707), .Z(\_MAC/_MULT/MULT/S[2][1][2] ) );
  XNOR U830 ( .A(n708), .B(n709), .Z(\_MAC/_MULT/MULT/S[2][1][1] ) );
  XOR U831 ( .A(n710), .B(n711), .Z(\_MAC/_MULT/MULT/S[2][1][15] ) );
  XOR U832 ( .A(n712), .B(n713), .Z(n711) );
  ANDN U833 ( .A(n714), .B(n715), .Z(n713) );
  AND U834 ( .A(n716), .B(n717), .Z(n712) );
  OR U835 ( .A(n714), .B(n718), .Z(n717) );
  AND U836 ( .A(n719), .B(n720), .Z(n716) );
  NAND U837 ( .A(n721), .B(n710), .Z(n720) );
  OR U838 ( .A(n722), .B(n723), .Z(n719) );
  OR U839 ( .A(n724), .B(n725), .Z(n714) );
  XOR U840 ( .A(n722), .B(n715), .Z(n718) );
  IV U841 ( .A(n723), .Z(n715) );
  XNOR U842 ( .A(n710), .B(n721), .Z(n722) );
  NANDN U843 ( .B(n150), .A(n729), .Z(n721) );
  XOR U844 ( .A(n725), .B(n724), .Z(\_MAC/_MULT/MULT/S[2][1][13] ) );
  NANDN U845 ( .B(n733), .A(n734), .Z(n724) );
  XNOR U846 ( .A(n726), .B(n735), .Z(n727) );
  NOR U847 ( .A(n736), .B(n737), .Z(n735) );
  XNOR U848 ( .A(n731), .B(n732), .Z(n728) );
  NAND U849 ( .A(n729), .B(n165), .Z(n732) );
  XNOR U850 ( .A(n730), .B(n741), .Z(n731) );
  ANDN U851 ( .A(n742), .B(n150), .Z(n741) );
  XNOR U852 ( .A(n733), .B(n734), .Z(\_MAC/_MULT/MULT/S[2][1][12] ) );
  XOR U853 ( .A(n753), .B(n737), .Z(n749) );
  NANDN U854 ( .B(n150), .A(n754), .Z(n737) );
  IV U855 ( .A(n738), .Z(n753) );
  XNOR U856 ( .A(n744), .B(n745), .Z(n740) );
  NAND U857 ( .A(n729), .B(n185), .Z(n745) );
  XNOR U858 ( .A(n743), .B(n758), .Z(n744) );
  AND U859 ( .A(n165), .B(n742), .Z(n758) );
  XNOR U860 ( .A(n748), .B(n747), .Z(\_MAC/_MULT/MULT/S[2][1][11] ) );
  XOR U861 ( .A(n762), .B(n763), .Z(n747) );
  XOR U862 ( .A(n764), .B(n765), .Z(n763) );
  AND U863 ( .A(n766), .B(n767), .Z(n764) );
  NAND U864 ( .A(n768), .B(n769), .Z(n767) );
  NANDN U865 ( .B(n770), .A(n765), .Z(n766) );
  XNOR U866 ( .A(n750), .B(n775), .Z(n751) );
  ANDN U867 ( .A(n776), .B(n150), .Z(n775) );
  XOR U868 ( .A(n780), .B(n752), .Z(n774) );
  NAND U869 ( .A(n754), .B(n165), .Z(n752) );
  IV U870 ( .A(n755), .Z(n780) );
  XNOR U871 ( .A(n760), .B(n761), .Z(n757) );
  NAND U872 ( .A(n729), .B(n214), .Z(n761) );
  XNOR U873 ( .A(n759), .B(n784), .Z(n760) );
  AND U874 ( .A(n185), .B(n742), .Z(n784) );
  XNOR U875 ( .A(n773), .B(n772), .Z(\_MAC/_MULT/MULT/S[2][1][10] ) );
  XNOR U876 ( .A(n788), .B(n770), .Z(n772) );
  XNOR U877 ( .A(n769), .B(n768), .Z(n770) );
  NANDN U878 ( .B(n150), .A(n789), .Z(n768) );
  XNOR U879 ( .A(n765), .B(n771), .Z(n788) );
  XOR U880 ( .A(n794), .B(n795), .Z(n693) );
  XNOR U881 ( .A(n796), .B(n793), .Z(n794) );
  XOR U882 ( .A(n800), .B(n801), .Z(n695) );
  XNOR U883 ( .A(n802), .B(n799), .Z(n800) );
  XOR U884 ( .A(n806), .B(n807), .Z(n697) );
  XNOR U885 ( .A(n808), .B(n805), .Z(n806) );
  XOR U886 ( .A(n809), .B(n810), .Z(n696) );
  XOR U887 ( .A(n814), .B(n815), .Z(n699) );
  XNOR U888 ( .A(n816), .B(n811), .Z(n814) );
  XOR U889 ( .A(n820), .B(n821), .Z(n701) );
  XNOR U890 ( .A(n822), .B(n817), .Z(n820) );
  XOR U891 ( .A(n826), .B(n827), .Z(n703) );
  XNOR U892 ( .A(n828), .B(n823), .Z(n826) );
  XOR U893 ( .A(n832), .B(n833), .Z(n705) );
  XNOR U894 ( .A(n834), .B(n829), .Z(n832) );
  XOR U895 ( .A(n838), .B(n839), .Z(n707) );
  XNOR U896 ( .A(n840), .B(n835), .Z(n838) );
  XOR U897 ( .A(n844), .B(n845), .Z(n709) );
  XNOR U898 ( .A(n846), .B(n841), .Z(n844) );
  XNOR U899 ( .A(n850), .B(n795), .Z(n851) );
  XNOR U900 ( .A(n791), .B(n792), .Z(n795) );
  NAND U901 ( .A(n789), .B(n165), .Z(n792) );
  XNOR U902 ( .A(n790), .B(n852), .Z(n791) );
  ANDN U903 ( .A(n853), .B(n150), .Z(n852) );
  XOR U904 ( .A(n850), .B(n857), .Z(n796) );
  NOR U905 ( .A(n858), .B(n859), .Z(n857) );
  XNOR U906 ( .A(n855), .B(n856), .Z(n801) );
  NAND U907 ( .A(n789), .B(n185), .Z(n856) );
  XNOR U908 ( .A(n854), .B(n861), .Z(n855) );
  AND U909 ( .A(n165), .B(n853), .Z(n861) );
  XOR U910 ( .A(n869), .B(n859), .Z(n865) );
  NANDN U911 ( .B(n150), .A(n870), .Z(n859) );
  IV U912 ( .A(n860), .Z(n869) );
  NAND U913 ( .A(n789), .B(n214), .Z(n864) );
  XNOR U914 ( .A(n862), .B(n872), .Z(n863) );
  AND U915 ( .A(n185), .B(n853), .Z(n872) );
  XNOR U916 ( .A(n866), .B(n877), .Z(n867) );
  ANDN U917 ( .A(n878), .B(n150), .Z(n877) );
  NAND U918 ( .A(\_MAC/_MULT/A_[15] ), .B(g_input[15]), .Z(n150) );
  XOR U919 ( .A(n882), .B(n868), .Z(n876) );
  NAND U920 ( .A(n870), .B(n165), .Z(n868) );
  IV U921 ( .A(n871), .Z(n882) );
  XNOR U922 ( .A(n874), .B(n875), .Z(n815) );
  NAND U923 ( .A(n789), .B(n242), .Z(n875) );
  XNOR U924 ( .A(n873), .B(n884), .Z(n874) );
  AND U925 ( .A(n214), .B(n853), .Z(n884) );
  XNOR U926 ( .A(n879), .B(n889), .Z(n880) );
  AND U927 ( .A(n165), .B(n878), .Z(n889) );
  XOR U928 ( .A(n893), .B(n881), .Z(n888) );
  NAND U929 ( .A(n870), .B(n185), .Z(n881) );
  IV U930 ( .A(n883), .Z(n893) );
  XNOR U931 ( .A(n886), .B(n887), .Z(n821) );
  NANDN U932 ( .B(n273), .A(n789), .Z(n887) );
  XNOR U933 ( .A(n885), .B(n895), .Z(n886) );
  AND U934 ( .A(n242), .B(n853), .Z(n895) );
  XNOR U935 ( .A(n890), .B(n900), .Z(n891) );
  AND U936 ( .A(n185), .B(n878), .Z(n900) );
  XOR U937 ( .A(n904), .B(n892), .Z(n899) );
  NAND U938 ( .A(n870), .B(n214), .Z(n892) );
  IV U939 ( .A(n894), .Z(n904) );
  XNOR U940 ( .A(n897), .B(n898), .Z(n827) );
  NANDN U941 ( .B(n385), .A(n789), .Z(n898) );
  XNOR U942 ( .A(n896), .B(n906), .Z(n897) );
  ANDN U943 ( .A(n853), .B(n273), .Z(n906) );
  XNOR U944 ( .A(n901), .B(n911), .Z(n902) );
  AND U945 ( .A(n214), .B(n878), .Z(n911) );
  XOR U946 ( .A(n915), .B(n903), .Z(n910) );
  NAND U947 ( .A(n870), .B(n242), .Z(n903) );
  IV U948 ( .A(n905), .Z(n915) );
  XNOR U949 ( .A(n908), .B(n909), .Z(n833) );
  NAND U950 ( .A(n789), .B(n400), .Z(n909) );
  XNOR U951 ( .A(n907), .B(n917), .Z(n908) );
  ANDN U952 ( .A(n853), .B(n385), .Z(n917) );
  XNOR U953 ( .A(n912), .B(n922), .Z(n913) );
  AND U954 ( .A(n242), .B(n878), .Z(n922) );
  XOR U955 ( .A(n926), .B(n914), .Z(n921) );
  NANDN U956 ( .B(n273), .A(n870), .Z(n914) );
  IV U957 ( .A(n916), .Z(n926) );
  XNOR U958 ( .A(n919), .B(n920), .Z(n839) );
  NAND U959 ( .A(n789), .B(n418), .Z(n920) );
  XNOR U960 ( .A(n918), .B(n928), .Z(n919) );
  AND U961 ( .A(n400), .B(n853), .Z(n928) );
  XNOR U962 ( .A(n923), .B(n933), .Z(n924) );
  ANDN U963 ( .A(n878), .B(n273), .Z(n933) );
  XOR U964 ( .A(n934), .B(n935), .Z(n923) );
  ANDN U965 ( .A(n936), .B(n937), .Z(n935) );
  XNOR U966 ( .A(n938), .B(n934), .Z(n936) );
  XOR U967 ( .A(n939), .B(n925), .Z(n932) );
  NANDN U968 ( .B(n385), .A(n870), .Z(n925) );
  IV U969 ( .A(n927), .Z(n939) );
  XNOR U970 ( .A(n930), .B(n931), .Z(n845) );
  NAND U971 ( .A(n789), .B(n436), .Z(n931) );
  XNOR U972 ( .A(n929), .B(n941), .Z(n930) );
  AND U973 ( .A(n418), .B(n853), .Z(n941) );
  XNOR U974 ( .A(n934), .B(n946), .Z(n937) );
  ANDN U975 ( .A(n878), .B(n385), .Z(n946) );
  XOR U976 ( .A(n947), .B(n948), .Z(n934) );
  ANDN U977 ( .A(n949), .B(n950), .Z(n948) );
  XNOR U978 ( .A(n951), .B(n947), .Z(n949) );
  XOR U979 ( .A(n952), .B(n938), .Z(n945) );
  NAND U980 ( .A(n870), .B(n400), .Z(n938) );
  IV U981 ( .A(n940), .Z(n952) );
  XNOR U982 ( .A(n777), .B(n957), .Z(n778) );
  AND U983 ( .A(n165), .B(n776), .Z(n957) );
  XNOR U984 ( .A(n958), .B(g_input[14]), .Z(n165) );
  NAND U985 ( .A(n959), .B(g_input[15]), .Z(n958) );
  XOR U986 ( .A(g_input[14]), .B(\_MAC/_MULT/A_[14] ), .Z(n959) );
  XOR U987 ( .A(n960), .B(n961), .Z(n777) );
  ANDN U988 ( .A(n962), .B(n963), .Z(n961) );
  XNOR U989 ( .A(n964), .B(n960), .Z(n962) );
  XOR U990 ( .A(n965), .B(n779), .Z(n956) );
  NAND U991 ( .A(n754), .B(n185), .Z(n779) );
  IV U992 ( .A(n781), .Z(n965) );
  XNOR U993 ( .A(n960), .B(n968), .Z(n963) );
  AND U994 ( .A(n185), .B(n776), .Z(n968) );
  XNOR U995 ( .A(n969), .B(g_input[13]), .Z(n185) );
  NAND U996 ( .A(n970), .B(g_input[15]), .Z(n969) );
  XOR U997 ( .A(g_input[13]), .B(\_MAC/_MULT/A_[13] ), .Z(n970) );
  XOR U998 ( .A(n971), .B(n972), .Z(n960) );
  ANDN U999 ( .A(n973), .B(n974), .Z(n972) );
  XNOR U1000 ( .A(n975), .B(n971), .Z(n973) );
  XOR U1001 ( .A(n976), .B(n964), .Z(n967) );
  NAND U1002 ( .A(n754), .B(n214), .Z(n964) );
  IV U1003 ( .A(n966), .Z(n976) );
  XNOR U1004 ( .A(n977), .B(n978), .Z(n797) );
  XNOR U1005 ( .A(n971), .B(n981), .Z(n974) );
  AND U1006 ( .A(n214), .B(n776), .Z(n981) );
  XOR U1007 ( .A(n982), .B(n983), .Z(n971) );
  ANDN U1008 ( .A(n984), .B(n985), .Z(n983) );
  XNOR U1009 ( .A(n986), .B(n982), .Z(n984) );
  XOR U1010 ( .A(n987), .B(n975), .Z(n980) );
  NAND U1011 ( .A(n754), .B(n242), .Z(n975) );
  IV U1012 ( .A(n979), .Z(n987) );
  XNOR U1013 ( .A(n988), .B(n989), .Z(n803) );
  XOR U1014 ( .A(n991), .B(n992), .Z(n809) );
  XNOR U1015 ( .A(n982), .B(n994), .Z(n985) );
  AND U1016 ( .A(n242), .B(n776), .Z(n994) );
  XOR U1017 ( .A(n995), .B(n996), .Z(n982) );
  ANDN U1018 ( .A(n997), .B(n998), .Z(n996) );
  XNOR U1019 ( .A(n999), .B(n995), .Z(n997) );
  XOR U1020 ( .A(n1000), .B(n986), .Z(n993) );
  NANDN U1021 ( .B(n273), .A(n754), .Z(n986) );
  IV U1022 ( .A(n990), .Z(n1000) );
  XNOR U1023 ( .A(n995), .B(n1003), .Z(n998) );
  ANDN U1024 ( .A(n776), .B(n273), .Z(n1003) );
  XOR U1025 ( .A(n1004), .B(n1005), .Z(n995) );
  ANDN U1026 ( .A(n1006), .B(n1007), .Z(n1005) );
  XNOR U1027 ( .A(n1008), .B(n1004), .Z(n1006) );
  XOR U1028 ( .A(n1009), .B(n999), .Z(n1002) );
  NANDN U1029 ( .B(n385), .A(n754), .Z(n999) );
  IV U1030 ( .A(n1001), .Z(n1009) );
  XNOR U1031 ( .A(n1010), .B(n1011), .Z(n812) );
  XNOR U1032 ( .A(n1004), .B(n1014), .Z(n1007) );
  ANDN U1033 ( .A(n776), .B(n385), .Z(n1014) );
  XOR U1034 ( .A(n1015), .B(n1016), .Z(n1004) );
  ANDN U1035 ( .A(n1017), .B(n1018), .Z(n1016) );
  XNOR U1036 ( .A(n1019), .B(n1015), .Z(n1017) );
  XOR U1037 ( .A(n1020), .B(n1008), .Z(n1013) );
  NAND U1038 ( .A(n754), .B(n400), .Z(n1008) );
  IV U1039 ( .A(n1012), .Z(n1020) );
  XNOR U1040 ( .A(n1021), .B(n1022), .Z(n818) );
  XNOR U1041 ( .A(n1015), .B(n1025), .Z(n1018) );
  AND U1042 ( .A(n400), .B(n776), .Z(n1025) );
  XOR U1043 ( .A(n1026), .B(n1027), .Z(n1015) );
  ANDN U1044 ( .A(n1028), .B(n1029), .Z(n1027) );
  XNOR U1045 ( .A(n1030), .B(n1026), .Z(n1028) );
  XOR U1046 ( .A(n1031), .B(n1019), .Z(n1024) );
  NAND U1047 ( .A(n754), .B(n418), .Z(n1019) );
  IV U1048 ( .A(n1023), .Z(n1031) );
  XNOR U1049 ( .A(n1032), .B(n1033), .Z(n824) );
  XNOR U1050 ( .A(n1026), .B(n1036), .Z(n1029) );
  AND U1051 ( .A(n418), .B(n776), .Z(n1036) );
  XOR U1052 ( .A(n1037), .B(n1038), .Z(n1026) );
  ANDN U1053 ( .A(n1039), .B(n1040), .Z(n1038) );
  XNOR U1054 ( .A(n1041), .B(n1037), .Z(n1039) );
  XOR U1055 ( .A(n1042), .B(n1030), .Z(n1035) );
  NAND U1056 ( .A(n754), .B(n436), .Z(n1030) );
  IV U1057 ( .A(n1034), .Z(n1042) );
  XNOR U1058 ( .A(n1043), .B(n1044), .Z(n830) );
  XNOR U1059 ( .A(n1037), .B(n1047), .Z(n1040) );
  AND U1060 ( .A(n436), .B(n776), .Z(n1047) );
  XOR U1061 ( .A(n1048), .B(n1049), .Z(n1037) );
  ANDN U1062 ( .A(n1050), .B(n1051), .Z(n1049) );
  XNOR U1063 ( .A(n1052), .B(n1048), .Z(n1050) );
  XOR U1064 ( .A(n1053), .B(n1041), .Z(n1046) );
  NAND U1065 ( .A(n754), .B(n531), .Z(n1041) );
  IV U1066 ( .A(n1045), .Z(n1053) );
  XNOR U1067 ( .A(n1054), .B(n1055), .Z(n836) );
  XNOR U1068 ( .A(n1048), .B(n1058), .Z(n1051) );
  AND U1069 ( .A(n531), .B(n776), .Z(n1058) );
  XOR U1070 ( .A(n1059), .B(n1060), .Z(n1048) );
  ANDN U1071 ( .A(n1061), .B(n1062), .Z(n1060) );
  XNOR U1072 ( .A(n1063), .B(n1059), .Z(n1061) );
  XOR U1073 ( .A(n1064), .B(n1052), .Z(n1057) );
  NAND U1074 ( .A(n754), .B(n544), .Z(n1052) );
  IV U1075 ( .A(n1056), .Z(n1064) );
  XNOR U1076 ( .A(n1065), .B(n1066), .Z(n842) );
  XNOR U1077 ( .A(n786), .B(n787), .Z(n783) );
  NAND U1078 ( .A(n729), .B(n242), .Z(n787) );
  XNOR U1079 ( .A(n785), .B(n1070), .Z(n786) );
  AND U1080 ( .A(n214), .B(n742), .Z(n1070) );
  XNOR U1081 ( .A(n1071), .B(g_input[12]), .Z(n214) );
  NAND U1082 ( .A(n1072), .B(g_input[15]), .Z(n1071) );
  XOR U1083 ( .A(g_input[12]), .B(\_MAC/_MULT/A_[12] ), .Z(n1072) );
  XNOR U1084 ( .A(n1073), .B(n1074), .Z(n977) );
  AND U1085 ( .A(n242), .B(n742), .Z(n1074) );
  XNOR U1086 ( .A(n1075), .B(g_input[11]), .Z(n242) );
  NAND U1087 ( .A(n1076), .B(g_input[15]), .Z(n1075) );
  XOR U1088 ( .A(g_input[11]), .B(\_MAC/_MULT/A_[11] ), .Z(n1076) );
  NANDN U1089 ( .B(n273), .A(n729), .Z(n978) );
  XNOR U1090 ( .A(n1077), .B(n1078), .Z(n988) );
  ANDN U1091 ( .A(n742), .B(n273), .Z(n1078) );
  XOR U1092 ( .A(n1079), .B(g_input[10]), .Z(n273) );
  NAND U1093 ( .A(n1080), .B(g_input[15]), .Z(n1079) );
  XOR U1094 ( .A(g_input[10]), .B(\_MAC/_MULT/A_[10] ), .Z(n1080) );
  NANDN U1095 ( .B(n385), .A(n729), .Z(n989) );
  XNOR U1096 ( .A(n992), .B(n1081), .Z(n1082) );
  NAND U1097 ( .A(n729), .B(n400), .Z(n992) );
  XOR U1098 ( .A(n1081), .B(n1083), .Z(n991) );
  ANDN U1099 ( .A(n742), .B(n385), .Z(n1083) );
  XOR U1100 ( .A(n1084), .B(g_input[9]), .Z(n385) );
  NAND U1101 ( .A(n1085), .B(g_input[15]), .Z(n1084) );
  XOR U1102 ( .A(g_input[9]), .B(\_MAC/_MULT/A_[9] ), .Z(n1085) );
  XNOR U1103 ( .A(n1086), .B(n1087), .Z(n1010) );
  AND U1104 ( .A(n400), .B(n742), .Z(n1087) );
  NAND U1105 ( .A(n729), .B(n418), .Z(n1011) );
  XNOR U1106 ( .A(n1088), .B(n1089), .Z(n1021) );
  AND U1107 ( .A(n418), .B(n742), .Z(n1089) );
  NAND U1108 ( .A(n729), .B(n436), .Z(n1022) );
  XNOR U1109 ( .A(n1090), .B(n1091), .Z(n1032) );
  AND U1110 ( .A(n436), .B(n742), .Z(n1091) );
  NAND U1111 ( .A(n729), .B(n531), .Z(n1033) );
  XNOR U1112 ( .A(n1092), .B(n1093), .Z(n1043) );
  AND U1113 ( .A(n531), .B(n742), .Z(n1093) );
  NAND U1114 ( .A(n729), .B(n544), .Z(n1044) );
  XNOR U1115 ( .A(n1094), .B(n1095), .Z(n1054) );
  AND U1116 ( .A(n544), .B(n742), .Z(n1095) );
  NAND U1117 ( .A(n729), .B(n567), .Z(n1055) );
  XNOR U1118 ( .A(n1096), .B(n1097), .Z(n1065) );
  AND U1119 ( .A(n567), .B(n742), .Z(n1097) );
  NANDN U1120 ( .B(n571), .A(n729), .Z(n1066) );
  XNOR U1121 ( .A(n849), .B(n848), .Z(\_MAC/_MULT/MULT/S[2][1][0] ) );
  XOR U1122 ( .A(n1101), .B(n955), .Z(n848) );
  XNOR U1123 ( .A(n943), .B(n944), .Z(n955) );
  NAND U1124 ( .A(n789), .B(n531), .Z(n944) );
  XNOR U1125 ( .A(n942), .B(n1102), .Z(n943) );
  AND U1126 ( .A(n436), .B(n853), .Z(n1102) );
  XNOR U1127 ( .A(n1106), .B(n1103), .Z(n1105) );
  XNOR U1128 ( .A(n954), .B(n847), .Z(n1101) );
  XOR U1129 ( .A(n1107), .B(n1108), .Z(n847) );
  XNOR U1130 ( .A(n947), .B(n1110), .Z(n950) );
  AND U1131 ( .A(n400), .B(n878), .Z(n1110) );
  XNOR U1132 ( .A(n1111), .B(g_input[8]), .Z(n400) );
  NAND U1133 ( .A(n1112), .B(g_input[15]), .Z(n1111) );
  XOR U1134 ( .A(g_input[8]), .B(\_MAC/_MULT/A_[8] ), .Z(n1112) );
  XOR U1135 ( .A(n1113), .B(n1114), .Z(n947) );
  AND U1136 ( .A(n1115), .B(n1116), .Z(n1114) );
  XNOR U1137 ( .A(n1117), .B(n1113), .Z(n1116) );
  XOR U1138 ( .A(n1118), .B(n951), .Z(n1109) );
  NAND U1139 ( .A(n870), .B(n418), .Z(n951) );
  IV U1140 ( .A(n953), .Z(n1118) );
  XNOR U1141 ( .A(n1119), .B(n1120), .Z(n953) );
  AND U1142 ( .A(n1121), .B(n1122), .Z(n1120) );
  XOR U1143 ( .A(n1115), .B(n1123), .Z(n1122) );
  XNOR U1144 ( .A(n1117), .B(n1119), .Z(n1123) );
  NAND U1145 ( .A(n870), .B(n436), .Z(n1117) );
  XOR U1146 ( .A(n1113), .B(n1124), .Z(n1115) );
  AND U1147 ( .A(n418), .B(n878), .Z(n1124) );
  XNOR U1148 ( .A(n1125), .B(g_input[7]), .Z(n418) );
  NAND U1149 ( .A(n1126), .B(g_input[15]), .Z(n1125) );
  XOR U1150 ( .A(g_input[7]), .B(\_MAC/_MULT/A_[7] ), .Z(n1126) );
  XOR U1151 ( .A(n1127), .B(n1128), .Z(n1113) );
  AND U1152 ( .A(n1129), .B(n1130), .Z(n1128) );
  XNOR U1153 ( .A(n1131), .B(n1127), .Z(n1130) );
  XOR U1154 ( .A(n1104), .B(n1132), .Z(n1121) );
  XNOR U1155 ( .A(n1106), .B(n1119), .Z(n1132) );
  NAND U1156 ( .A(n789), .B(n544), .Z(n1106) );
  XOR U1157 ( .A(n1103), .B(n1133), .Z(n1104) );
  AND U1158 ( .A(n531), .B(n853), .Z(n1133) );
  XNOR U1159 ( .A(n1137), .B(n1134), .Z(n1136) );
  XOR U1160 ( .A(n1138), .B(n1139), .Z(n1119) );
  AND U1161 ( .A(n1140), .B(n1141), .Z(n1139) );
  XOR U1162 ( .A(n1129), .B(n1142), .Z(n1141) );
  XNOR U1163 ( .A(n1131), .B(n1138), .Z(n1142) );
  NAND U1164 ( .A(n870), .B(n531), .Z(n1131) );
  XOR U1165 ( .A(n1127), .B(n1143), .Z(n1129) );
  AND U1166 ( .A(n436), .B(n878), .Z(n1143) );
  XNOR U1167 ( .A(n1144), .B(g_input[6]), .Z(n436) );
  NAND U1168 ( .A(n1145), .B(g_input[15]), .Z(n1144) );
  XOR U1169 ( .A(g_input[6]), .B(\_MAC/_MULT/A_[6] ), .Z(n1145) );
  XOR U1170 ( .A(n1146), .B(n1147), .Z(n1127) );
  AND U1171 ( .A(n1148), .B(n1149), .Z(n1147) );
  XNOR U1172 ( .A(n1150), .B(n1146), .Z(n1149) );
  XOR U1173 ( .A(n1135), .B(n1151), .Z(n1140) );
  XNOR U1174 ( .A(n1137), .B(n1138), .Z(n1151) );
  NAND U1175 ( .A(n789), .B(n567), .Z(n1137) );
  XOR U1176 ( .A(n1134), .B(n1152), .Z(n1135) );
  AND U1177 ( .A(n544), .B(n853), .Z(n1152) );
  XNOR U1178 ( .A(n1156), .B(n1153), .Z(n1155) );
  XOR U1179 ( .A(n1157), .B(n1158), .Z(n1138) );
  AND U1180 ( .A(n1159), .B(n1160), .Z(n1158) );
  XOR U1181 ( .A(n1148), .B(n1161), .Z(n1160) );
  XNOR U1182 ( .A(n1150), .B(n1157), .Z(n1161) );
  NAND U1183 ( .A(n870), .B(n544), .Z(n1150) );
  XOR U1184 ( .A(n1146), .B(n1162), .Z(n1148) );
  AND U1185 ( .A(n531), .B(n878), .Z(n1162) );
  XNOR U1186 ( .A(n1163), .B(g_input[5]), .Z(n531) );
  NAND U1187 ( .A(n1164), .B(g_input[15]), .Z(n1163) );
  XOR U1188 ( .A(g_input[5]), .B(\_MAC/_MULT/A_[5] ), .Z(n1164) );
  XOR U1189 ( .A(n1165), .B(n1166), .Z(n1146) );
  ANDN U1190 ( .A(n1167), .B(n1168), .Z(n1166) );
  XNOR U1191 ( .A(n1169), .B(n1165), .Z(n1167) );
  XOR U1192 ( .A(n1154), .B(n1170), .Z(n1159) );
  XNOR U1193 ( .A(n1156), .B(n1157), .Z(n1170) );
  NANDN U1194 ( .B(n571), .A(n789), .Z(n1156) );
  XOR U1195 ( .A(n1153), .B(n1171), .Z(n1154) );
  AND U1196 ( .A(n567), .B(n853), .Z(n1171) );
  XOR U1197 ( .A(n1172), .B(n1173), .Z(n1153) );
  ANDN U1198 ( .A(n1174), .B(n1175), .Z(n1173) );
  XNOR U1199 ( .A(n1176), .B(n1172), .Z(n1174) );
  NAND U1200 ( .A(n789), .B(n640), .Z(n1176) );
  XNOR U1201 ( .A(n1172), .B(n1178), .Z(n1175) );
  ANDN U1202 ( .A(n853), .B(n571), .Z(n1178) );
  ANDN U1203 ( .A(n1179), .B(n643), .Z(n1172) );
  NANDN U1204 ( .B(n789), .A(n1180), .Z(n1179) );
  NAND U1205 ( .A(n640), .B(n853), .Z(n1180) );
  XNOR U1206 ( .A(n1181), .B(e_input[10]), .Z(n853) );
  NANDN U1207 ( .B(n127), .A(n1182), .Z(n1181) );
  XOR U1208 ( .A(e_input[10]), .B(\_MAC/_MULT/X_[10] ), .Z(n1182) );
  XNOR U1209 ( .A(n1183), .B(e_input[11]), .Z(n789) );
  NANDN U1210 ( .B(n127), .A(n1184), .Z(n1183) );
  XOR U1211 ( .A(e_input[11]), .B(\_MAC/_MULT/X_[11] ), .Z(n1184) );
  XNOR U1212 ( .A(n1165), .B(n1186), .Z(n1168) );
  AND U1213 ( .A(n544), .B(n878), .Z(n1186) );
  XOR U1214 ( .A(n1187), .B(n1188), .Z(n1165) );
  AND U1215 ( .A(n1189), .B(n1190), .Z(n1188) );
  XOR U1216 ( .A(n1191), .B(n1187), .Z(n1190) );
  AND U1217 ( .A(n567), .B(n878), .Z(n1191) );
  XOR U1218 ( .A(n1192), .B(n1187), .Z(n1189) );
  ANDN U1219 ( .A(n870), .B(n571), .Z(n1192) );
  XOR U1220 ( .A(n1193), .B(n1194), .Z(n1187) );
  ANDN U1221 ( .A(n1195), .B(n1196), .Z(n1194) );
  XNOR U1222 ( .A(n1197), .B(n1193), .Z(n1195) );
  XOR U1223 ( .A(n1198), .B(n1169), .Z(n1185) );
  NAND U1224 ( .A(n870), .B(n567), .Z(n1169) );
  IV U1225 ( .A(n1177), .Z(n1198) );
  XOR U1226 ( .A(n1199), .B(n1197), .Z(n1177) );
  NAND U1227 ( .A(n870), .B(n640), .Z(n1197) );
  IV U1228 ( .A(n1196), .Z(n1199) );
  XNOR U1229 ( .A(n1193), .B(n1200), .Z(n1196) );
  ANDN U1230 ( .A(n878), .B(n571), .Z(n1200) );
  ANDN U1231 ( .A(n1201), .B(n643), .Z(n1193) );
  NANDN U1232 ( .B(n870), .A(n1202), .Z(n1201) );
  NAND U1233 ( .A(n640), .B(n878), .Z(n1202) );
  XNOR U1234 ( .A(n1203), .B(e_input[8]), .Z(n878) );
  NANDN U1235 ( .B(n127), .A(n1204), .Z(n1203) );
  XOR U1236 ( .A(e_input[8]), .B(\_MAC/_MULT/X_[8] ), .Z(n1204) );
  XNOR U1237 ( .A(n1205), .B(e_input[9]), .Z(n870) );
  NANDN U1238 ( .B(n127), .A(n1206), .Z(n1205) );
  XOR U1239 ( .A(e_input[9]), .B(\_MAC/_MULT/X_[9] ), .Z(n1206) );
  XNOR U1240 ( .A(n1059), .B(n1208), .Z(n1062) );
  AND U1241 ( .A(n544), .B(n776), .Z(n1208) );
  XNOR U1242 ( .A(n1209), .B(g_input[4]), .Z(n544) );
  NAND U1243 ( .A(n1210), .B(g_input[15]), .Z(n1209) );
  XOR U1244 ( .A(g_input[4]), .B(\_MAC/_MULT/A_[4] ), .Z(n1210) );
  XOR U1245 ( .A(n1211), .B(n1212), .Z(n1059) );
  AND U1246 ( .A(n1213), .B(n1214), .Z(n1212) );
  XOR U1247 ( .A(n1215), .B(n1211), .Z(n1214) );
  AND U1248 ( .A(n567), .B(n776), .Z(n1215) );
  XOR U1249 ( .A(n1216), .B(n1211), .Z(n1213) );
  ANDN U1250 ( .A(n754), .B(n571), .Z(n1216) );
  XOR U1251 ( .A(n1217), .B(n1218), .Z(n1211) );
  ANDN U1252 ( .A(n1219), .B(n1220), .Z(n1218) );
  XNOR U1253 ( .A(n1221), .B(n1217), .Z(n1219) );
  XOR U1254 ( .A(n1222), .B(n1063), .Z(n1207) );
  NAND U1255 ( .A(n754), .B(n567), .Z(n1063) );
  XNOR U1256 ( .A(n1223), .B(g_input[3]), .Z(n567) );
  NAND U1257 ( .A(n1224), .B(g_input[15]), .Z(n1223) );
  XOR U1258 ( .A(g_input[3]), .B(\_MAC/_MULT/A_[3] ), .Z(n1224) );
  IV U1259 ( .A(n1067), .Z(n1222) );
  NAND U1260 ( .A(n754), .B(n640), .Z(n1221) );
  XNOR U1261 ( .A(n1217), .B(n1225), .Z(n1220) );
  ANDN U1262 ( .A(n776), .B(n571), .Z(n1225) );
  ANDN U1263 ( .A(n1226), .B(n643), .Z(n1217) );
  NANDN U1264 ( .B(n754), .A(n1227), .Z(n1226) );
  NAND U1265 ( .A(n640), .B(n776), .Z(n1227) );
  XNOR U1266 ( .A(n1228), .B(e_input[12]), .Z(n776) );
  NANDN U1267 ( .B(n127), .A(n1229), .Z(n1228) );
  XOR U1268 ( .A(e_input[12]), .B(\_MAC/_MULT/X_[12] ), .Z(n1229) );
  XNOR U1269 ( .A(n1230), .B(e_input[13]), .Z(n754) );
  NANDN U1270 ( .B(n127), .A(n1231), .Z(n1230) );
  XOR U1271 ( .A(e_input[13]), .B(\_MAC/_MULT/X_[13] ), .Z(n1231) );
  XNOR U1272 ( .A(n1099), .B(n1100), .Z(n1069) );
  NAND U1273 ( .A(n729), .B(n640), .Z(n1100) );
  XNOR U1274 ( .A(n1098), .B(n1232), .Z(n1099) );
  ANDN U1275 ( .A(n742), .B(n571), .Z(n1232) );
  XOR U1276 ( .A(n1233), .B(g_input[2]), .Z(n571) );
  NAND U1277 ( .A(n1234), .B(g_input[15]), .Z(n1233) );
  XOR U1278 ( .A(g_input[2]), .B(\_MAC/_MULT/A_[2] ), .Z(n1234) );
  ANDN U1279 ( .A(n1235), .B(n643), .Z(n1098) );
  XOR U1280 ( .A(n1236), .B(g_input[0]), .Z(n643) );
  NAND U1281 ( .A(n1237), .B(g_input[15]), .Z(n1236) );
  XOR U1282 ( .A(g_input[0]), .B(\_MAC/_MULT/A_[0] ), .Z(n1237) );
  NANDN U1283 ( .B(n729), .A(n1238), .Z(n1235) );
  NAND U1284 ( .A(n640), .B(n742), .Z(n1238) );
  XNOR U1285 ( .A(n1239), .B(e_input[14]), .Z(n742) );
  NANDN U1286 ( .B(n127), .A(n1240), .Z(n1239) );
  XOR U1287 ( .A(e_input[14]), .B(\_MAC/_MULT/X_[14] ), .Z(n1240) );
  IV U1288 ( .A(e_input[15]), .Z(n127) );
  XNOR U1289 ( .A(n1241), .B(g_input[1]), .Z(n640) );
  NAND U1290 ( .A(n1242), .B(g_input[15]), .Z(n1241) );
  XOR U1291 ( .A(g_input[1]), .B(\_MAC/_MULT/A_[1] ), .Z(n1242) );
  AND U1292 ( .A(\_MAC/_MULT/X_[15] ), .B(e_input[15]), .Z(n729) );
endmodule

