
module MxM_TG_W16_N10000 ( clk, rst, g_input, e_input, o );
  input [15:0] g_input;
  input [15:0] e_input;
  output [15:0] o;
  input clk, rst;
  wire   \_MxM/n262 , \_MxM/n261 , \_MxM/n260 , \_MxM/n259 , \_MxM/n258 ,
         \_MxM/n257 , \_MxM/n256 , \_MxM/n255 , \_MxM/n254 , \_MxM/n253 ,
         \_MxM/n252 , \_MxM/n251 , \_MxM/n250 , \_MxM/n249 , \_MxM/n248 ,
         \_MxM/n247 , \_MxM/n246 , \_MxM/n245 , \_MxM/n244 , \_MxM/n243 ,
         \_MxM/n242 , \_MxM/n241 , \_MxM/n240 , \_MxM/n239 , \_MxM/n238 ,
         \_MxM/n237 , \_MxM/n236 , \_MxM/n235 , \_MxM/n234 , \_MxM/n233 ,
         \_MxM/n232 , \_MxM/n231 , \_MxM/n230 , \_MxM/n229 , \_MxM/n228 ,
         \_MxM/n227 , \_MxM/n226 , \_MxM/n225 , \_MxM/n224 , \_MxM/n223 ,
         \_MxM/n222 , \_MxM/n221 , \_MxM/n220 , \_MxM/n219 , \_MxM/n218 ,
         \_MxM/n217 , \_MxM/N19 , \_MxM/N18 , \_MxM/N17 , \_MxM/N16 ,
         \_MxM/N15 , \_MxM/N14 , \_MxM/N13 , \_MxM/N12 , \_MxM/N11 ,
         \_MxM/N10 , \_MxM/N9 , \_MxM/N8 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/n[7] , \_MxM/n[8] , \_MxM/n[9] , \_MxM/n[10] , \_MxM/n[11] ,
         \_MxM/n[12] , \_MxM/n[13] , \_MxM/Y0[0] , \_MxM/Y0[1] , \_MxM/Y0[2] ,
         \_MxM/Y0[3] , \_MxM/Y0[4] , \_MxM/Y0[5] , \_MxM/Y0[6] , \_MxM/Y0[7] ,
         \_MxM/Y0[8] , \_MxM/Y0[9] , \_MxM/Y0[10] , \_MxM/Y0[11] ,
         \_MxM/Y0[12] , \_MxM/Y0[13] , \_MxM/Y0[14] , \_MxM/Y0[15] ,
         \_MxM/add_39/carry[13] , \_MxM/add_39/carry[12] ,
         \_MxM/add_39/carry[11] , \_MxM/add_39/carry[10] ,
         \_MxM/add_39/carry[9] , \_MxM/add_39/carry[8] ,
         \_MxM/add_39/carry[7] , \_MxM/add_39/carry[6] ,
         \_MxM/add_39/carry[5] , \_MxM/add_39/carry[4] ,
         \_MxM/add_39/carry[3] , \_MxM/add_39/carry[2] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498;

  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n217 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n218 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n219 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n220 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n221 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n222 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n223 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n224 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n225 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n226 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n227 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n228 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n229 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n230 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n231 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n232 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/n233 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/n234 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/n235 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/n236 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/n237 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/n238 ), .CLK(clk), .RST(1'b0), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/n239 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/n240 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/n241 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/n242 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/n243 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/n244 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/n245 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/n246 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/n247 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/n248 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[13]  ( .D(\_MxM/n249 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[13] ) );
  DFF \_MxM/n_reg[12]  ( .D(\_MxM/n250 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[12] ) );
  DFF \_MxM/n_reg[11]  ( .D(\_MxM/n251 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[11] ) );
  DFF \_MxM/n_reg[10]  ( .D(\_MxM/n252 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[10] ) );
  DFF \_MxM/n_reg[9]  ( .D(\_MxM/n253 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[9] ) );
  DFF \_MxM/n_reg[8]  ( .D(\_MxM/n254 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[8] ) );
  DFF \_MxM/n_reg[7]  ( .D(\_MxM/n255 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[7] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/n256 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/n257 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/n258 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/n259 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/n260 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/n261 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/n262 ), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_39/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_39/carry[2] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_39/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_39/carry[2] ), .COUT(\_MxM/add_39/carry[3] ), .SUM(\_MxM/N9 ) );
  HADDER \_MxM/add_39/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_39/carry[3] ), .COUT(\_MxM/add_39/carry[4] ), .SUM(\_MxM/N10 ) );
  HADDER \_MxM/add_39/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_39/carry[4] ), .COUT(\_MxM/add_39/carry[5] ), .SUM(\_MxM/N11 ) );
  HADDER \_MxM/add_39/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_39/carry[5] ), .COUT(\_MxM/add_39/carry[6] ), .SUM(\_MxM/N12 ) );
  HADDER \_MxM/add_39/U1_1_6  ( .IN0(\_MxM/n[6] ), .IN1(\_MxM/add_39/carry[6] ), .COUT(\_MxM/add_39/carry[7] ), .SUM(\_MxM/N13 ) );
  HADDER \_MxM/add_39/U1_1_7  ( .IN0(\_MxM/n[7] ), .IN1(\_MxM/add_39/carry[7] ), .COUT(\_MxM/add_39/carry[8] ), .SUM(\_MxM/N14 ) );
  HADDER \_MxM/add_39/U1_1_8  ( .IN0(\_MxM/n[8] ), .IN1(\_MxM/add_39/carry[8] ), .COUT(\_MxM/add_39/carry[9] ), .SUM(\_MxM/N15 ) );
  HADDER \_MxM/add_39/U1_1_9  ( .IN0(\_MxM/n[9] ), .IN1(\_MxM/add_39/carry[9] ), .COUT(\_MxM/add_39/carry[10] ), .SUM(\_MxM/N16 ) );
  HADDER \_MxM/add_39/U1_1_10  ( .IN0(\_MxM/n[10] ), .IN1(
        \_MxM/add_39/carry[10] ), .COUT(\_MxM/add_39/carry[11] ), .SUM(
        \_MxM/N17 ) );
  HADDER \_MxM/add_39/U1_1_11  ( .IN0(\_MxM/n[11] ), .IN1(
        \_MxM/add_39/carry[11] ), .COUT(\_MxM/add_39/carry[12] ), .SUM(
        \_MxM/N18 ) );
  HADDER \_MxM/add_39/U1_1_12  ( .IN0(\_MxM/n[12] ), .IN1(
        \_MxM/add_39/carry[12] ), .COUT(\_MxM/add_39/carry[13] ), .SUM(
        \_MxM/N19 ) );
  MUX U1 ( .IN0(n1), .IN1(n1321), .SEL(n1322), .F(n1305) );
  IV U2 ( .A(n1323), .Z(n1) );
  MUX U3 ( .IN0(n2), .IN1(n988), .SEL(n989), .F(n965) );
  IV U4 ( .A(n990), .Z(n2) );
  MUX U5 ( .IN0(n1396), .IN1(n1414), .SEL(n1398), .F(n1377) );
  XOR U6 ( .A(n1179), .B(n1169), .Z(n985) );
  XOR U7 ( .A(n991), .B(n973), .Z(n977) );
  MUX U8 ( .IN0(n3), .IN1(n738), .SEL(n739), .F(n668) );
  IV U9 ( .A(n740), .Z(n3) );
  MUX U10 ( .IN0(n4), .IN1(n899), .SEL(n900), .F(n824) );
  IV U11 ( .A(n901), .Z(n4) );
  MUX U12 ( .IN0(n5), .IN1(n965), .SEL(n966), .F(n942) );
  IV U13 ( .A(n967), .Z(n5) );
  MUX U14 ( .IN0(n6), .IN1(n1161), .SEL(n1162), .F(n1151) );
  IV U15 ( .A(n1163), .Z(n6) );
  XOR U16 ( .A(n1164), .B(n1156), .Z(n962) );
  MUX U17 ( .IN0(n1116), .IN1(n1119), .SEL(n1117), .F(n1101) );
  MUX U18 ( .IN0(n7), .IN1(n463), .SEL(n464), .F(n412) );
  IV U19 ( .A(n465), .Z(n7) );
  MUX U20 ( .IN0(n8), .IN1(n815), .SEL(n816), .F(n738) );
  IV U21 ( .A(n817), .Z(n8) );
  XNOR U22 ( .A(n1459), .B(n1460), .Z(n903) );
  XOR U23 ( .A(n966), .B(n967), .Z(n978) );
  MUX U24 ( .IN0(n9), .IN1(n915), .SEL(n916), .F(n853) );
  IV U25 ( .A(n917), .Z(n9) );
  XOR U26 ( .A(n1152), .B(n1153), .Z(n960) );
  MUX U27 ( .IN0(n10), .IN1(n592), .SEL(n593), .F(n527) );
  IV U28 ( .A(n594), .Z(n10) );
  MUX U29 ( .IN0(e_input[8]), .IN1(n1444), .SEL(e_input[15]), .F(n475) );
  MUX U30 ( .IN0(n1157), .IN1(n11), .SEL(n1156), .F(n1148) );
  IV U31 ( .A(n1155), .Z(n11) );
  MUX U32 ( .IN0(e_input[13]), .IN1(n1470), .SEL(e_input[15]), .F(n257) );
  MUX U33 ( .IN0(n1332), .IN1(n1335), .SEL(n1333), .F(n1316) );
  MUX U34 ( .IN0(n12), .IN1(n942), .SEL(n943), .F(n923) );
  IV U35 ( .A(n944), .Z(n12) );
  MUX U36 ( .IN0(n13), .IN1(n1151), .SEL(n1152), .F(n930) );
  IV U37 ( .A(n1153), .Z(n13) );
  XOR U38 ( .A(n968), .B(n950), .Z(n954) );
  MUX U39 ( .IN0(e_input[9]), .IN1(n1445), .SEL(e_input[15]), .F(n421) );
  MUX U40 ( .IN0(n298), .IN1(n14), .SEL(n297), .F(n259) );
  IV U41 ( .A(n296), .Z(n14) );
  MUX U42 ( .IN0(e_input[11]), .IN1(n1425), .SEL(e_input[15]), .F(n327) );
  MUX U43 ( .IN0(n388), .IN1(n386), .SEL(n387), .F(n341) );
  MUX U44 ( .IN0(n15), .IN1(n181), .SEL(n180), .F(n189) );
  IV U45 ( .A(n192), .Z(n15) );
  MUX U46 ( .IN0(n16), .IN1(n1336), .SEL(n1337), .F(n1332) );
  IV U47 ( .A(n1338), .Z(n16) );
  XOR U48 ( .A(n1162), .B(n1163), .Z(n983) );
  MUX U49 ( .IN0(n17), .IN1(n719), .SEL(n720), .F(n650) );
  IV U50 ( .A(n721), .Z(n17) );
  MUX U51 ( .IN0(n18), .IN1(n778), .SEL(n779), .F(n715) );
  IV U52 ( .A(n780), .Z(n18) );
  MUX U53 ( .IN0(e_input[10]), .IN1(n1424), .SEL(e_input[15]), .F(n368) );
  MUX U54 ( .IN0(n478), .IN1(n19), .SEL(n477), .F(n423) );
  IV U55 ( .A(n476), .Z(n19) );
  MUX U56 ( .IN0(n554), .IN1(n552), .SEL(n553), .F(n487) );
  XNOR U57 ( .A(n1446), .B(n900), .Z(n904) );
  XOR U58 ( .A(n190), .B(n211), .Z(n209) );
  MUX U59 ( .IN0(n1377), .IN1(n1395), .SEL(n1379), .F(n1346) );
  MUX U60 ( .IN0(n1265), .IN1(n1287), .SEL(n1267), .F(n1247) );
  MUX U61 ( .IN0(n20), .IN1(n923), .SEL(n924), .F(n861) );
  IV U62 ( .A(n925), .Z(n20) );
  MUX U63 ( .IN0(n21), .IN1(n1168), .SEL(n1169), .F(n1155) );
  IV U64 ( .A(n1170), .Z(n21) );
  MUX U65 ( .IN0(n22), .IN1(n890), .SEL(n891), .F(n815) );
  IV U66 ( .A(n892), .Z(n22) );
  MUX U67 ( .IN0(g_input[11]), .IN1(n1199), .SEL(g_input[15]), .F(n344) );
  MUX U68 ( .IN0(n426), .IN1(n27), .SEL(n425), .F(n375) );
  MUX U69 ( .IN0(n687), .IN1(n685), .SEL(n686), .F(n617) );
  MUX U70 ( .IN0(n717), .IN1(n23), .SEL(n716), .F(n645) );
  IV U71 ( .A(n715), .Z(n23) );
  NAND U72 ( .A(n259), .B(n294), .Z(n293) );
  XOR U73 ( .A(n237), .B(n245), .Z(n243) );
  MUX U74 ( .IN0(n24), .IN1(n1183), .SEL(n1184), .F(n1168) );
  IV U75 ( .A(n1185), .Z(n24) );
  MUX U76 ( .IN0(n25), .IN1(n730), .SEL(n731), .F(n660) );
  IV U77 ( .A(n732), .Z(n25) );
  MUX U78 ( .IN0(n26), .IN1(n786), .SEL(n787), .F(n719) );
  IV U79 ( .A(n788), .Z(n26) );
  MUX U80 ( .IN0(e_input[4]), .IN1(n1130), .SEL(e_input[15]), .F(n714) );
  XOR U81 ( .A(n1426), .B(n1411), .Z(n1351) );
  MUX U82 ( .IN0(n470), .IN1(n472), .SEL(n471), .F(n27) );
  IV U83 ( .A(n27), .Z(n424) );
  MUX U84 ( .IN0(n648), .IN1(n28), .SEL(n647), .F(n575) );
  IV U85 ( .A(n646), .Z(n28) );
  MUX U86 ( .IN0(n755), .IN1(n753), .SEL(n754), .F(n685) );
  MUX U87 ( .IN0(n873), .IN1(n29), .SEL(n872), .F(n796) );
  IV U88 ( .A(n871), .Z(n29) );
  XNOR U89 ( .A(n378), .B(n338), .Z(n342) );
  XOR U90 ( .A(n268), .B(n276), .Z(n274) );
  XOR U91 ( .A(n943), .B(n944), .Z(n955) );
  MUX U92 ( .IN0(n1271), .IN1(n1281), .SEL(n1273), .F(n1257) );
  MUX U93 ( .IN0(n1346), .IN1(n1376), .SEL(n1348), .F(n882) );
  XNOR U94 ( .A(n1123), .B(n1124), .Z(n1107) );
  MUX U95 ( .IN0(g_input[9]), .IN1(n1237), .SEL(g_input[15]), .F(n438) );
  MUX U96 ( .IN0(g_input[12]), .IN1(n1181), .SEL(g_input[15]), .F(n299) );
  XOR U97 ( .A(n347), .B(n390), .Z(n348) );
  MUX U98 ( .IN0(n742), .IN1(n744), .SEL(n743), .F(n674) );
  MUX U99 ( .IN0(n784), .IN1(n782), .SEL(n783), .F(n709) );
  XOR U100 ( .A(n872), .B(n873), .Z(n879) );
  XNOR U101 ( .A(n375), .B(n418), .Z(n376) );
  XNOR U102 ( .A(n479), .B(n432), .Z(n436) );
  MUX U103 ( .IN0(n30), .IN1(n663), .SEL(n664), .F(n595) );
  IV U104 ( .A(n665), .Z(n30) );
  MUX U105 ( .IN0(n522), .IN1(n524), .SEL(n523), .F(n31) );
  IV U106 ( .A(n31), .Z(n458) );
  XOR U107 ( .A(n305), .B(n313), .Z(n311) );
  MUX U108 ( .IN0(n1263), .IN1(n32), .SEL(n1113), .F(n1244) );
  IV U109 ( .A(n1112), .Z(n32) );
  MUX U110 ( .IN0(n1109), .IN1(n1107), .SEL(n1108), .F(n1080) );
  XOR U111 ( .A(n1154), .B(n1148), .Z(n939) );
  MUX U112 ( .IN0(n33), .IN1(n882), .SEL(n883), .F(n807) );
  IV U113 ( .A(n884), .Z(n33) );
  MUX U114 ( .IN0(n34), .IN1(n930), .SEL(n931), .F(n871) );
  IV U115 ( .A(n932), .Z(n34) );
  XOR U116 ( .A(n945), .B(n916), .Z(n920) );
  MUX U117 ( .IN0(n606), .IN1(n608), .SEL(n607), .F(n541) );
  MUX U118 ( .IN0(n832), .IN1(n830), .SEL(n831), .F(n753) );
  XOR U119 ( .A(n1352), .B(n891), .Z(n895) );
  XNOR U120 ( .A(n427), .B(n383), .Z(n387) );
  MUX U121 ( .IN0(n35), .IN1(n466), .SEL(n467), .F(n415) );
  IV U122 ( .A(n468), .Z(n35) );
  MUX U123 ( .IN0(n36), .IN1(n581), .SEL(n582), .F(n521) );
  IV U124 ( .A(n583), .Z(n36) );
  NAND U125 ( .A(n645), .B(n713), .Z(n712) );
  MUX U126 ( .IN0(n587), .IN1(n589), .SEL(n588), .F(n522) );
  MUX U127 ( .IN0(n37), .IN1(n561), .SEL(n562), .F(n496) );
  IV U128 ( .A(\_MxM/Y0[5] ), .Z(n37) );
  XOR U129 ( .A(n350), .B(n358), .Z(n356) );
  MUX U130 ( .IN0(n38), .IN1(n1316), .SEL(n1317), .F(n1299) );
  IV U131 ( .A(n1318), .Z(n38) );
  MUX U132 ( .IN0(g_input[1]), .IN1(n1472), .SEL(g_input[15]), .F(n1126) );
  MUX U133 ( .IN0(n39), .IN1(n527), .SEL(n528), .F(n463) );
  IV U134 ( .A(n529), .Z(n39) );
  MUX U135 ( .IN0(g_input[6]), .IN1(n1368), .SEL(g_input[15]), .F(n620) );
  MUX U136 ( .IN0(g_input[7]), .IN1(n1355), .SEL(g_input[15]), .F(n555) );
  MUX U137 ( .IN0(g_input[5]), .IN1(n1388), .SEL(g_input[15]), .F(n688) );
  MUX U138 ( .IN0(n40), .IN1(n861), .SEL(n862), .F(n786) );
  IV U139 ( .A(n863), .Z(n40) );
  XOR U140 ( .A(n931), .B(n932), .Z(n937) );
  MUX U141 ( .IN0(n674), .IN1(n676), .SEL(n675), .F(n606) );
  XNOR U142 ( .A(n913), .B(n854), .Z(n858) );
  XOR U143 ( .A(n265), .B(n300), .Z(n266) );
  MUX U144 ( .IN0(n41), .IN1(n330), .SEL(n331), .F(n283) );
  IV U145 ( .A(n332), .Z(n41) );
  NAND U146 ( .A(n423), .B(n474), .Z(n473) );
  MUX U147 ( .IN0(n577), .IN1(n575), .SEL(n576), .F(n519) );
  XNOR U148 ( .A(n609), .B(n549), .Z(n553) );
  MUX U149 ( .IN0(n42), .IN1(n810), .SEL(n811), .F(n733) );
  IV U150 ( .A(n812), .Z(n42) );
  MUX U151 ( .IN0(n43), .IN1(n657), .SEL(n656), .F(n587) );
  IV U152 ( .A(n655), .Z(n43) );
  MUX U153 ( .IN0(n44), .IN1(n626), .SEL(n627), .F(n561) );
  IV U154 ( .A(\_MxM/Y0[4] ), .Z(n44) );
  XOR U155 ( .A(n395), .B(n403), .Z(n401) );
  MUX U156 ( .IN0(n1080), .IN1(n45), .SEL(n1081), .F(n1053) );
  IV U157 ( .A(n1082), .Z(n45) );
  MUX U158 ( .IN0(n1172), .IN1(n46), .SEL(n985), .F(n1159) );
  IV U159 ( .A(n983), .Z(n46) );
  XNOR U160 ( .A(n1337), .B(n1338), .Z(n1324) );
  MUX U161 ( .IN0(n47), .IN1(n660), .SEL(n661), .F(n592) );
  IV U162 ( .A(n662), .Z(n47) );
  MUX U163 ( .IN0(g_input[3]), .IN1(n1449), .SEL(g_input[15]), .F(n48) );
  IV U164 ( .A(n48), .Z(n833) );
  MUX U165 ( .IN0(g_input[4]), .IN1(n1406), .SEL(g_input[15]), .F(n49) );
  IV U166 ( .A(n49), .Z(n756) );
  MUX U167 ( .IN0(n919), .IN1(n50), .SEL(n920), .F(n857) );
  IV U168 ( .A(n921), .Z(n50) );
  XOR U169 ( .A(n1250), .B(n1251), .Z(n1112) );
  MUX U170 ( .IN0(n343), .IN1(n341), .SEL(n342), .F(n288) );
  MUX U171 ( .IN0(n51), .IN1(n650), .SEL(n651), .F(n581) );
  IV U172 ( .A(n652), .Z(n51) );
  XOR U173 ( .A(n558), .B(n621), .Z(n559) );
  MUX U174 ( .IN0(n819), .IN1(n821), .SEL(n820), .F(n742) );
  MUX U175 ( .IN0(n905), .IN1(n903), .SEL(n904), .F(n830) );
  MUX U176 ( .IN0(n52), .IN1(n372), .SEL(n373), .F(n330) );
  IV U177 ( .A(n374), .Z(n52) );
  XOR U178 ( .A(n533), .B(n477), .Z(n471) );
  XNOR U179 ( .A(n544), .B(n484), .Z(n488) );
  MUX U180 ( .IN0(n53), .IN1(n595), .SEL(n596), .F(n530) );
  IV U181 ( .A(n597), .Z(n53) );
  XOR U182 ( .A(n708), .B(n646), .Z(n647) );
  MUX U183 ( .IN0(n804), .IN1(n54), .SEL(n803), .F(n725) );
  IV U184 ( .A(n802), .Z(n54) );
  MUX U185 ( .IN0(n722), .IN1(n55), .SEL(n723), .F(n655) );
  IV U186 ( .A(n724), .Z(n55) );
  MUX U187 ( .IN0(n56), .IN1(n694), .SEL(n695), .F(n626) );
  IV U188 ( .A(\_MxM/Y0[3] ), .Z(n56) );
  XOR U189 ( .A(n450), .B(n456), .Z(n445) );
  MUX U190 ( .IN0(n57), .IN1(n1110), .SEL(n927), .F(n1083) );
  IV U191 ( .A(n926), .Z(n57) );
  MUX U192 ( .IN0(n1026), .IN1(n58), .SEL(n1027), .F(n999) );
  IV U193 ( .A(n1028), .Z(n58) );
  MUX U194 ( .IN0(e_input[1]), .IN1(n59), .SEL(e_input[15]), .F(n1143) );
  IV U195 ( .A(n1343), .Z(n59) );
  MUX U196 ( .IN0(e_input[6]), .IN1(n1135), .SEL(e_input[15]), .F(n580) );
  MUX U197 ( .IN0(e_input[3]), .IN1(n1329), .SEL(e_input[15]), .F(n799) );
  MUX U198 ( .IN0(n894), .IN1(n896), .SEL(n895), .F(n819) );
  MUX U199 ( .IN0(e_input[14]), .IN1(n1475), .SEL(e_input[15]), .F(n226) );
  NAND U200 ( .A(n324), .B(n367), .Z(n366) );
  XOR U201 ( .A(n598), .B(n538), .Z(n542) );
  XNOR U202 ( .A(n677), .B(n614), .Z(n618) );
  MUX U203 ( .IN0(n60), .IN1(n733), .SEL(n734), .F(n663) );
  IV U204 ( .A(n735), .Z(n60) );
  XNOR U205 ( .A(n776), .B(n716), .Z(n710) );
  MUX U206 ( .IN0(n789), .IN1(n61), .SEL(n790), .F(n722) );
  IV U207 ( .A(n791), .Z(n61) );
  MUX U208 ( .IN0(n62), .IN1(n268), .SEL(n269), .F(n237) );
  IV U209 ( .A(\_MxM/Y0[11] ), .Z(n62) );
  XOR U210 ( .A(n496), .B(n504), .Z(n502) );
  MUX U211 ( .IN0(n1244), .IN1(n63), .SEL(n1089), .F(n1225) );
  IV U212 ( .A(n1087), .Z(n63) );
  MUX U213 ( .IN0(n1299), .IN1(n1315), .SEL(n1301), .F(n1282) );
  MUX U214 ( .IN0(n976), .IN1(n64), .SEL(n977), .F(n953) );
  IV U215 ( .A(n978), .Z(n64) );
  XOR U216 ( .A(n924), .B(n925), .Z(n921) );
  XOR U217 ( .A(n1322), .B(n1323), .Z(n1137) );
  MUX U218 ( .IN0(n65), .IN1(n807), .SEL(n808), .F(n730) );
  IV U219 ( .A(n809), .Z(n65) );
  MUX U220 ( .IN0(g_input[10]), .IN1(n1217), .SEL(g_input[15]), .F(n389) );
  XNOR U221 ( .A(n1114), .B(n1104), .Z(n1108) );
  XOR U222 ( .A(n441), .B(n491), .Z(n442) );
  MUX U223 ( .IN0(n489), .IN1(n487), .SEL(n488), .F(n435) );
  MUX U224 ( .IN0(n711), .IN1(n709), .SEL(n710), .F(n646) );
  MUX U225 ( .IN0(g_input[13]), .IN1(n1167), .SEL(g_input[15]), .F(n262) );
  MUX U226 ( .IN0(n66), .IN1(n530), .SEL(n531), .F(n466) );
  IV U227 ( .A(n532), .Z(n66) );
  XOR U228 ( .A(n666), .B(n603), .Z(n607) );
  XNOR U229 ( .A(n822), .B(n750), .Z(n754) );
  MUX U230 ( .IN0(n67), .IN1(n885), .SEL(n886), .F(n810) );
  IV U231 ( .A(n887), .Z(n67) );
  MUX U232 ( .IN0(n68), .IN1(n874), .SEL(n875), .F(n802) );
  IV U233 ( .A(n876), .Z(n68) );
  MUX U234 ( .IN0(g_input[14]), .IN1(n1144), .SEL(g_input[15]), .F(n227) );
  MUX U235 ( .IN0(n285), .IN1(n69), .SEL(n284), .F(n253) );
  IV U236 ( .A(n283), .Z(n69) );
  XNOR U237 ( .A(n587), .B(n586), .Z(n639) );
  MUX U238 ( .IN0(\_MxM/Y0[13] ), .IN1(n70), .SEL(n191), .F(n183) );
  IV U239 ( .A(n190), .Z(n70) );
  MUX U240 ( .IN0(n71), .IN1(n350), .SEL(n351), .F(n305) );
  IV U241 ( .A(\_MxM/Y0[9] ), .Z(n71) );
  MUX U242 ( .IN0(n72), .IN1(n839), .SEL(n840), .F(n762) );
  IV U243 ( .A(\_MxM/Y0[1] ), .Z(n72) );
  XOR U244 ( .A(n561), .B(n569), .Z(n567) );
  MUX U245 ( .IN0(n1225), .IN1(n73), .SEL(n1062), .F(n1206) );
  IV U246 ( .A(n1060), .Z(n73) );
  MUX U247 ( .IN0(n999), .IN1(n74), .SEL(n1000), .F(n976) );
  IV U248 ( .A(n1001), .Z(n74) );
  MUX U249 ( .IN0(n1282), .IN1(n1298), .SEL(n1284), .F(n1271) );
  MUX U250 ( .IN0(n1159), .IN1(n75), .SEL(n962), .F(n1149) );
  IV U251 ( .A(n960), .Z(n75) );
  MUX U252 ( .IN0(g_input[8]), .IN1(n1255), .SEL(g_input[15]), .F(n490) );
  MUX U253 ( .IN0(g_input[2]), .IN1(n1462), .SEL(g_input[15]), .F(n906) );
  MUX U254 ( .IN0(n76), .IN1(n853), .SEL(n854), .F(n778) );
  IV U255 ( .A(n855), .Z(n76) );
  MUX U256 ( .IN0(n77), .IN1(n412), .SEL(n413), .F(n369) );
  IV U257 ( .A(n414), .Z(n77) );
  MUX U258 ( .IN0(n541), .IN1(n543), .SEL(n542), .F(n470) );
  MUX U259 ( .IN0(n619), .IN1(n617), .SEL(n618), .F(n552) );
  XOR U260 ( .A(n836), .B(n907), .Z(n837) );
  MUX U261 ( .IN0(n859), .IN1(n857), .SEL(n858), .F(n782) );
  XNOR U262 ( .A(n288), .B(n289), .Z(n287) );
  MUX U263 ( .IN0(n78), .IN1(n415), .SEL(n416), .F(n372) );
  IV U264 ( .A(n417), .Z(n78) );
  XOR U265 ( .A(n582), .B(n583), .Z(n577) );
  XOR U266 ( .A(n813), .B(n739), .Z(n743) );
  XNOR U267 ( .A(n897), .B(n827), .Z(n831) );
  NAND U268 ( .A(n796), .B(n869), .Z(n868) );
  XNOR U269 ( .A(n292), .B(n291), .Z(n285) );
  XNOR U270 ( .A(n687), .B(n686), .Z(n665) );
  MUX U271 ( .IN0(n727), .IN1(n725), .SEL(n726), .F(n79) );
  IV U272 ( .A(n79), .Z(n654) );
  MUX U273 ( .IN0(n864), .IN1(n80), .SEL(n865), .F(n789) );
  IV U274 ( .A(n866), .Z(n80) );
  MUX U275 ( .IN0(n458), .IN1(n81), .SEL(n459), .F(n409) );
  IV U276 ( .A(n460), .Z(n81) );
  MUX U277 ( .IN0(n82), .IN1(n237), .SEL(n238), .F(n190) );
  IV U278 ( .A(\_MxM/Y0[12] ), .Z(n82) );
  MUX U279 ( .IN0(n83), .IN1(n395), .SEL(n396), .F(n350) );
  IV U280 ( .A(\_MxM/Y0[8] ), .Z(n83) );
  XOR U281 ( .A(n626), .B(n634), .Z(n632) );
  MUX U282 ( .IN0(n1206), .IN1(n84), .SEL(n1035), .F(n1187) );
  IV U283 ( .A(n1033), .Z(n84) );
  MUX U284 ( .IN0(n85), .IN1(n1350), .SEL(n1351), .F(n1400) );
  IV U285 ( .A(n1420), .Z(n85) );
  NOR U286 ( .A(g_input[0]), .B(n1472), .Z(n1463) );
  XOR U287 ( .A(n1330), .B(n1317), .Z(n1138) );
  MUX U288 ( .IN0(n1149), .IN1(n86), .SEL(n939), .F(n877) );
  IV U289 ( .A(n937), .Z(n86) );
  MUX U290 ( .IN0(n437), .IN1(n435), .SEL(n436), .F(n386) );
  XOR U291 ( .A(n691), .B(n757), .Z(n692) );
  MUX U292 ( .IN0(n371), .IN1(n87), .SEL(n370), .F(n324) );
  IV U293 ( .A(n369), .Z(n87) );
  MUX U294 ( .IN0(e_input[7]), .IN1(n1136), .SEL(e_input[15]), .F(n513) );
  XNOR U295 ( .A(n745), .B(n682), .Z(n686) );
  XOR U296 ( .A(n736), .B(n671), .Z(n675) );
  XNOR U297 ( .A(n851), .B(n779), .Z(n783) );
  XNOR U298 ( .A(n905), .B(n904), .Z(n887) );
  MUX U299 ( .IN0(n261), .IN1(n287), .SEL(n260), .F(n232) );
  XNOR U300 ( .A(n343), .B(n342), .Z(n332) );
  XNOR U301 ( .A(n554), .B(n553), .Z(n532) );
  XNOR U302 ( .A(n619), .B(n618), .Z(n597) );
  XNOR U303 ( .A(n725), .B(n792), .Z(n726) );
  XNOR U304 ( .A(n468), .B(n467), .Z(n460) );
  XOR U305 ( .A(n574), .B(n515), .Z(n523) );
  XNOR U306 ( .A(n735), .B(n734), .Z(n724) );
  XNOR U307 ( .A(n812), .B(n811), .Z(n791) );
  XNOR U308 ( .A(n251), .B(n250), .Z(n275) );
  MUX U309 ( .IN0(n88), .IN1(n444), .SEL(n445), .F(n395) );
  IV U310 ( .A(\_MxM/Y0[7] ), .Z(n88) );
  MUX U311 ( .IN0(\_MxM/Y0[14] ), .IN1(n183), .SEL(n184), .F(n173) );
  XOR U312 ( .A(n694), .B(n702), .Z(n700) );
  MUX U313 ( .IN0(n1053), .IN1(n89), .SEL(n1054), .F(n1026) );
  IV U314 ( .A(n1055), .Z(n89) );
  MUX U315 ( .IN0(n90), .IN1(n1137), .SEL(n1138), .F(n1310) );
  IV U316 ( .A(n1324), .Z(n90) );
  MUX U317 ( .IN0(n1187), .IN1(n91), .SEL(n1008), .F(n1172) );
  IV U318 ( .A(n1006), .Z(n91) );
  XOR U319 ( .A(n1448), .B(g_input[3]), .Z(n1449) );
  MUX U320 ( .IN0(n953), .IN1(n92), .SEL(n954), .F(n919) );
  IV U321 ( .A(n955), .Z(n92) );
  XOR U322 ( .A(n1418), .B(n1419), .Z(n1350) );
  XOR U323 ( .A(n1269), .B(n1260), .Z(n1113) );
  MUX U324 ( .IN0(e_input[5]), .IN1(n1131), .SEL(e_input[15]), .F(n643) );
  MUX U325 ( .IN0(e_input[2]), .IN1(n1328), .SEL(e_input[15]), .F(n870) );
  XNOR U326 ( .A(n1109), .B(n1108), .Z(n926) );
  XNOR U327 ( .A(n333), .B(n297), .Z(n291) );
  MUX U328 ( .IN0(n377), .IN1(n375), .SEL(n376), .F(n93) );
  IV U329 ( .A(n93), .Z(n329) );
  XOR U330 ( .A(n651), .B(n652), .Z(n648) );
  XOR U331 ( .A(n888), .B(n816), .Z(n820) );
  MUX U332 ( .IN0(n879), .IN1(n1139), .SEL(n878), .F(n801) );
  XNOR U333 ( .A(n859), .B(n858), .Z(n876) );
  AND U334 ( .A(n221), .B(n198), .Z(n220) );
  XNOR U335 ( .A(n388), .B(n387), .Z(n374) );
  XNOR U336 ( .A(n437), .B(n436), .Z(n417) );
  XNOR U337 ( .A(n489), .B(n488), .Z(n468) );
  XNOR U338 ( .A(n711), .B(n710), .Z(n727) );
  XNOR U339 ( .A(n755), .B(n754), .Z(n735) );
  XNOR U340 ( .A(n832), .B(n831), .Z(n812) );
  XNOR U341 ( .A(n784), .B(n783), .Z(n804) );
  XNOR U342 ( .A(n887), .B(n886), .Z(n866) );
  XNOR U343 ( .A(n252), .B(n253), .Z(n251) );
  XNOR U344 ( .A(n532), .B(n531), .Z(n524) );
  XNOR U345 ( .A(n597), .B(n596), .Z(n589) );
  XNOR U346 ( .A(n665), .B(n664), .Z(n657) );
  MUX U347 ( .IN0(n94), .IN1(n305), .SEL(n306), .F(n268) );
  IV U348 ( .A(\_MxM/Y0[10] ), .Z(n94) );
  MUX U349 ( .IN0(n95), .IN1(n496), .SEL(n497), .F(n444) );
  IV U350 ( .A(\_MxM/Y0[6] ), .Z(n95) );
  MUX U351 ( .IN0(n96), .IN1(n762), .SEL(n763), .F(n694) );
  IV U352 ( .A(\_MxM/Y0[2] ), .Z(n96) );
  MUX U353 ( .IN0(\_MxM/Y0[15] ), .IN1(n173), .SEL(n174), .F(n97) );
  IV U354 ( .A(n97), .Z(n170) );
  XOR U355 ( .A(n840), .B(\_MxM/Y0[1] ), .Z(n115) );
  ANDN U356 ( .A(n98), .B(\_MxM/n[0] ), .Z(\_MxM/n262 ) );
  AND U357 ( .A(\_MxM/N8 ), .B(n98), .Z(\_MxM/n261 ) );
  AND U358 ( .A(\_MxM/N9 ), .B(n98), .Z(\_MxM/n260 ) );
  AND U359 ( .A(\_MxM/N10 ), .B(n98), .Z(\_MxM/n259 ) );
  AND U360 ( .A(\_MxM/N11 ), .B(n98), .Z(\_MxM/n258 ) );
  AND U361 ( .A(\_MxM/N12 ), .B(n98), .Z(\_MxM/n257 ) );
  AND U362 ( .A(\_MxM/N13 ), .B(n98), .Z(\_MxM/n256 ) );
  AND U363 ( .A(\_MxM/N14 ), .B(n98), .Z(\_MxM/n255 ) );
  AND U364 ( .A(\_MxM/N15 ), .B(n98), .Z(\_MxM/n254 ) );
  AND U365 ( .A(\_MxM/N16 ), .B(n98), .Z(\_MxM/n253 ) );
  AND U366 ( .A(\_MxM/N17 ), .B(n98), .Z(\_MxM/n252 ) );
  AND U367 ( .A(\_MxM/N18 ), .B(n98), .Z(\_MxM/n251 ) );
  AND U368 ( .A(\_MxM/N19 ), .B(n98), .Z(\_MxM/n250 ) );
  AND U369 ( .A(n98), .B(n99), .Z(\_MxM/n249 ) );
  XOR U370 ( .A(\_MxM/n[13] ), .B(\_MxM/add_39/carry[13] ), .Z(n99) );
  ANDN U371 ( .A(n100), .B(rst), .Z(n98) );
  NAND U372 ( .A(n101), .B(n102), .Z(n100) );
  AND U373 ( .A(n103), .B(n104), .Z(n102) );
  ANDN U374 ( .A(n105), .B(n106), .Z(n104) );
  NOR U375 ( .A(n107), .B(n108), .Z(n105) );
  AND U376 ( .A(n109), .B(\_MxM/n[13] ), .Z(n103) );
  AND U377 ( .A(\_MxM/n[10] ), .B(\_MxM/n[0] ), .Z(n109) );
  AND U378 ( .A(n110), .B(n111), .Z(n101) );
  AND U379 ( .A(\_MxM/n[3] ), .B(n112), .Z(n111) );
  AND U380 ( .A(\_MxM/n[2] ), .B(\_MxM/n[1] ), .Z(n112) );
  AND U381 ( .A(\_MxM/n[9] ), .B(\_MxM/n[8] ), .Z(n110) );
  NAND U382 ( .A(n113), .B(n114), .Z(\_MxM/n248 ) );
  OR U383 ( .A(n115), .B(n116), .Z(n114) );
  NANDN U384 ( .B(n117), .A(\_MxM/Y0[0] ), .Z(n113) );
  NAND U385 ( .A(n118), .B(n119), .Z(\_MxM/n247 ) );
  NANDN U386 ( .B(n116), .A(n120), .Z(n119) );
  NANDN U387 ( .B(n121), .A(rst), .Z(n118) );
  NAND U388 ( .A(n122), .B(n123), .Z(\_MxM/n246 ) );
  NANDN U389 ( .B(n116), .A(n124), .Z(n123) );
  NANDN U390 ( .B(n117), .A(\_MxM/Y0[2] ), .Z(n122) );
  NAND U391 ( .A(n125), .B(n126), .Z(\_MxM/n245 ) );
  NANDN U392 ( .B(n116), .A(n127), .Z(n126) );
  NANDN U393 ( .B(n117), .A(\_MxM/Y0[3] ), .Z(n125) );
  NAND U394 ( .A(n128), .B(n129), .Z(\_MxM/n244 ) );
  NANDN U395 ( .B(n116), .A(n130), .Z(n129) );
  NANDN U396 ( .B(n117), .A(\_MxM/Y0[4] ), .Z(n128) );
  NAND U397 ( .A(n131), .B(n132), .Z(\_MxM/n243 ) );
  NANDN U398 ( .B(n116), .A(n133), .Z(n132) );
  NANDN U399 ( .B(n117), .A(\_MxM/Y0[5] ), .Z(n131) );
  NAND U400 ( .A(n134), .B(n135), .Z(\_MxM/n242 ) );
  NANDN U401 ( .B(n116), .A(n136), .Z(n135) );
  NANDN U402 ( .B(n117), .A(\_MxM/Y0[6] ), .Z(n134) );
  NAND U403 ( .A(n137), .B(n138), .Z(\_MxM/n241 ) );
  NANDN U404 ( .B(n116), .A(n139), .Z(n138) );
  NANDN U405 ( .B(n117), .A(\_MxM/Y0[7] ), .Z(n137) );
  NAND U406 ( .A(n140), .B(n141), .Z(\_MxM/n240 ) );
  NANDN U407 ( .B(n116), .A(n142), .Z(n141) );
  NANDN U408 ( .B(n117), .A(\_MxM/Y0[8] ), .Z(n140) );
  NAND U409 ( .A(n143), .B(n144), .Z(\_MxM/n239 ) );
  NANDN U410 ( .B(n116), .A(n145), .Z(n144) );
  NANDN U411 ( .B(n117), .A(\_MxM/Y0[9] ), .Z(n143) );
  NAND U412 ( .A(n146), .B(n147), .Z(\_MxM/n238 ) );
  NANDN U413 ( .B(n116), .A(n148), .Z(n147) );
  NANDN U414 ( .B(n117), .A(\_MxM/Y0[10] ), .Z(n146) );
  NAND U415 ( .A(n149), .B(n150), .Z(\_MxM/n237 ) );
  NANDN U416 ( .B(n116), .A(n151), .Z(n150) );
  NANDN U417 ( .B(n117), .A(\_MxM/Y0[11] ), .Z(n149) );
  NAND U418 ( .A(n152), .B(n153), .Z(\_MxM/n236 ) );
  NANDN U419 ( .B(n116), .A(n154), .Z(n153) );
  NANDN U420 ( .B(n117), .A(\_MxM/Y0[12] ), .Z(n152) );
  NAND U421 ( .A(n155), .B(n156), .Z(\_MxM/n235 ) );
  NANDN U422 ( .B(n116), .A(n157), .Z(n156) );
  NANDN U423 ( .B(n117), .A(\_MxM/Y0[13] ), .Z(n155) );
  NAND U424 ( .A(n158), .B(n159), .Z(\_MxM/n234 ) );
  OR U425 ( .A(n160), .B(n116), .Z(n159) );
  NANDN U426 ( .B(n117), .A(\_MxM/Y0[14] ), .Z(n158) );
  NAND U427 ( .A(n161), .B(n162), .Z(\_MxM/n233 ) );
  OR U428 ( .A(n116), .B(n163), .Z(n162) );
  NANDN U429 ( .B(n164), .A(n117), .Z(n116) );
  NANDN U430 ( .B(n117), .A(\_MxM/Y0[15] ), .Z(n161) );
  NAND U431 ( .A(n165), .B(n166), .Z(\_MxM/n232 ) );
  NANDN U432 ( .B(n117), .A(o[15]), .Z(n166) );
  AND U433 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U434 ( .B(n164), .A(o[15]), .Z(n168) );
  OR U435 ( .A(n163), .B(n169), .Z(n167) );
  XOR U436 ( .A(n170), .B(n171), .Z(n163) );
  XNOR U437 ( .A(\_MxM/Y0[15] ), .B(n172), .Z(n171) );
  NAND U438 ( .A(n175), .B(n176), .Z(\_MxM/n231 ) );
  NANDN U439 ( .B(n117), .A(o[14]), .Z(n176) );
  AND U440 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U441 ( .B(n164), .A(o[14]), .Z(n178) );
  OR U442 ( .A(n160), .B(n169), .Z(n177) );
  XOR U443 ( .A(n174), .B(\_MxM/Y0[15] ), .Z(n160) );
  XOR U444 ( .A(n173), .B(n172), .Z(n174) );
  NAND U445 ( .A(n179), .B(n180), .Z(n172) );
  OR U446 ( .A(n181), .B(n182), .Z(n179) );
  NAND U447 ( .A(n185), .B(n186), .Z(\_MxM/n230 ) );
  NANDN U448 ( .B(n117), .A(o[13]), .Z(n186) );
  AND U449 ( .A(n187), .B(n188), .Z(n185) );
  NANDN U450 ( .B(n164), .A(o[13]), .Z(n188) );
  NANDN U451 ( .B(n169), .A(n157), .Z(n187) );
  XNOR U452 ( .A(n184), .B(\_MxM/Y0[14] ), .Z(n157) );
  XNOR U453 ( .A(n189), .B(n183), .Z(n184) );
  XNOR U454 ( .A(n182), .B(n192), .Z(n181) );
  OR U455 ( .A(n193), .B(n194), .Z(n182) );
  AND U456 ( .A(n195), .B(n196), .Z(n192) );
  OR U457 ( .A(n197), .B(n198), .Z(n196) );
  AND U458 ( .A(n199), .B(n200), .Z(n195) );
  OR U459 ( .A(n201), .B(n202), .Z(n200) );
  OR U460 ( .A(n203), .B(n204), .Z(n199) );
  NAND U461 ( .A(n205), .B(n206), .Z(\_MxM/n229 ) );
  NANDN U462 ( .B(n117), .A(o[12]), .Z(n206) );
  AND U463 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U464 ( .B(n164), .A(o[12]), .Z(n208) );
  NANDN U465 ( .B(n169), .A(n154), .Z(n207) );
  XNOR U466 ( .A(n191), .B(\_MxM/Y0[13] ), .Z(n154) );
  XNOR U467 ( .A(n209), .B(n210), .Z(n191) );
  AND U468 ( .A(n180), .B(n212), .Z(n211) );
  XOR U469 ( .A(n193), .B(n213), .Z(n212) );
  XOR U470 ( .A(n213), .B(n194), .Z(n193) );
  OR U471 ( .A(n214), .B(n215), .Z(n194) );
  IV U472 ( .A(n210), .Z(n213) );
  XNOR U473 ( .A(n204), .B(n203), .Z(n210) );
  OR U474 ( .A(n216), .B(n217), .Z(n203) );
  AND U475 ( .A(n218), .B(n219), .Z(n204) );
  XNOR U476 ( .A(n197), .B(n220), .Z(n219) );
  NAND U477 ( .A(n222), .B(n223), .Z(n198) );
  NANDN U478 ( .B(n224), .A(n225), .Z(n222) );
  NANDN U479 ( .B(n201), .A(n226), .Z(n221) );
  NANDN U480 ( .B(n202), .A(n227), .Z(n197) );
  AND U481 ( .A(n228), .B(n229), .Z(n218) );
  OR U482 ( .A(n230), .B(n231), .Z(n229) );
  XNOR U483 ( .A(n232), .B(n233), .Z(n228) );
  ANDN U484 ( .A(n234), .B(n235), .Z(n233) );
  XOR U485 ( .A(n232), .B(n236), .Z(n234) );
  NAND U486 ( .A(n239), .B(n240), .Z(\_MxM/n228 ) );
  NANDN U487 ( .B(n117), .A(o[11]), .Z(n240) );
  AND U488 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U489 ( .B(n164), .A(o[11]), .Z(n242) );
  NANDN U490 ( .B(n169), .A(n151), .Z(n241) );
  XNOR U491 ( .A(n238), .B(\_MxM/Y0[12] ), .Z(n151) );
  XNOR U492 ( .A(n243), .B(n244), .Z(n238) );
  AND U493 ( .A(n180), .B(n246), .Z(n245) );
  XOR U494 ( .A(n214), .B(n247), .Z(n246) );
  XOR U495 ( .A(n247), .B(n215), .Z(n214) );
  OR U496 ( .A(n248), .B(n249), .Z(n215) );
  IV U497 ( .A(n244), .Z(n247) );
  XNOR U498 ( .A(n217), .B(n216), .Z(n244) );
  OR U499 ( .A(n250), .B(n251), .Z(n216) );
  XNOR U500 ( .A(n231), .B(n230), .Z(n217) );
  OR U501 ( .A(n252), .B(n253), .Z(n230) );
  XOR U502 ( .A(n236), .B(n235), .Z(n231) );
  XOR U503 ( .A(n232), .B(n254), .Z(n235) );
  AND U504 ( .A(n255), .B(n256), .Z(n254) );
  NANDN U505 ( .B(n201), .A(n257), .Z(n256) );
  OR U506 ( .A(n258), .B(n259), .Z(n255) );
  XOR U507 ( .A(n224), .B(n225), .Z(n236) );
  NANDN U508 ( .B(n202), .A(n262), .Z(n225) );
  XNOR U509 ( .A(n223), .B(n263), .Z(n224) );
  AND U510 ( .A(n227), .B(n226), .Z(n263) );
  ANDN U511 ( .A(n264), .B(n265), .Z(n223) );
  NANDN U512 ( .B(n266), .A(n267), .Z(n264) );
  NAND U513 ( .A(n270), .B(n271), .Z(\_MxM/n227 ) );
  NANDN U514 ( .B(n117), .A(o[10]), .Z(n271) );
  AND U515 ( .A(n272), .B(n273), .Z(n270) );
  NANDN U516 ( .B(n164), .A(o[10]), .Z(n273) );
  NANDN U517 ( .B(n169), .A(n148), .Z(n272) );
  XNOR U518 ( .A(n269), .B(\_MxM/Y0[11] ), .Z(n148) );
  XNOR U519 ( .A(n274), .B(n275), .Z(n269) );
  AND U520 ( .A(n180), .B(n277), .Z(n276) );
  XOR U521 ( .A(n248), .B(n278), .Z(n277) );
  XOR U522 ( .A(n278), .B(n249), .Z(n248) );
  OR U523 ( .A(n279), .B(n280), .Z(n249) );
  IV U524 ( .A(n275), .Z(n278) );
  OR U525 ( .A(n281), .B(n282), .Z(n250) );
  XOR U526 ( .A(n261), .B(n260), .Z(n252) );
  XNOR U527 ( .A(n286), .B(n287), .Z(n260) );
  ANDN U528 ( .A(n290), .B(n291), .Z(n289) );
  XOR U529 ( .A(n288), .B(n292), .Z(n290) );
  XNOR U530 ( .A(n293), .B(n258), .Z(n286) );
  NAND U531 ( .A(n257), .B(n227), .Z(n258) );
  NANDN U532 ( .B(n201), .A(n295), .Z(n294) );
  XOR U533 ( .A(n266), .B(n267), .Z(n261) );
  NANDN U534 ( .B(n202), .A(n299), .Z(n267) );
  AND U535 ( .A(n262), .B(n226), .Z(n300) );
  NAND U536 ( .A(n301), .B(n302), .Z(n265) );
  NANDN U537 ( .B(n303), .A(n304), .Z(n301) );
  NAND U538 ( .A(n307), .B(n308), .Z(\_MxM/n226 ) );
  NANDN U539 ( .B(n117), .A(o[9]), .Z(n308) );
  AND U540 ( .A(n309), .B(n310), .Z(n307) );
  NANDN U541 ( .B(n164), .A(o[9]), .Z(n310) );
  NANDN U542 ( .B(n169), .A(n145), .Z(n309) );
  XNOR U543 ( .A(n306), .B(\_MxM/Y0[10] ), .Z(n145) );
  XNOR U544 ( .A(n311), .B(n312), .Z(n306) );
  AND U545 ( .A(n180), .B(n314), .Z(n313) );
  XOR U546 ( .A(n279), .B(n315), .Z(n314) );
  XOR U547 ( .A(n315), .B(n280), .Z(n279) );
  OR U548 ( .A(n316), .B(n317), .Z(n280) );
  IV U549 ( .A(n312), .Z(n315) );
  XNOR U550 ( .A(n282), .B(n281), .Z(n312) );
  OR U551 ( .A(n318), .B(n319), .Z(n281) );
  XNOR U552 ( .A(n285), .B(n284), .Z(n282) );
  XOR U553 ( .A(n283), .B(n320), .Z(n284) );
  AND U554 ( .A(n321), .B(n322), .Z(n320) );
  OR U555 ( .A(n323), .B(n324), .Z(n322) );
  AND U556 ( .A(n325), .B(n326), .Z(n321) );
  NANDN U557 ( .B(n201), .A(n327), .Z(n326) );
  NAND U558 ( .A(n328), .B(n329), .Z(n325) );
  XNOR U559 ( .A(n296), .B(n334), .Z(n297) );
  AND U560 ( .A(n227), .B(n295), .Z(n334) );
  XOR U561 ( .A(n335), .B(n336), .Z(n296) );
  ANDN U562 ( .A(n337), .B(n338), .Z(n336) );
  XNOR U563 ( .A(n339), .B(n335), .Z(n337) );
  XOR U564 ( .A(n340), .B(n298), .Z(n333) );
  NAND U565 ( .A(n257), .B(n262), .Z(n298) );
  IV U566 ( .A(n288), .Z(n340) );
  XNOR U567 ( .A(n303), .B(n304), .Z(n292) );
  NANDN U568 ( .B(n202), .A(n344), .Z(n304) );
  XNOR U569 ( .A(n302), .B(n345), .Z(n303) );
  AND U570 ( .A(n299), .B(n226), .Z(n345) );
  ANDN U571 ( .A(n346), .B(n347), .Z(n302) );
  NANDN U572 ( .B(n348), .A(n349), .Z(n346) );
  NAND U573 ( .A(n352), .B(n353), .Z(\_MxM/n225 ) );
  NANDN U574 ( .B(n117), .A(o[8]), .Z(n353) );
  AND U575 ( .A(n354), .B(n355), .Z(n352) );
  NANDN U576 ( .B(n164), .A(o[8]), .Z(n355) );
  NANDN U577 ( .B(n169), .A(n142), .Z(n354) );
  XNOR U578 ( .A(n351), .B(\_MxM/Y0[9] ), .Z(n142) );
  XNOR U579 ( .A(n356), .B(n357), .Z(n351) );
  AND U580 ( .A(n180), .B(n359), .Z(n358) );
  XOR U581 ( .A(n316), .B(n360), .Z(n359) );
  XOR U582 ( .A(n360), .B(n317), .Z(n316) );
  OR U583 ( .A(n361), .B(n362), .Z(n317) );
  IV U584 ( .A(n357), .Z(n360) );
  XNOR U585 ( .A(n319), .B(n318), .Z(n357) );
  OR U586 ( .A(n363), .B(n364), .Z(n318) );
  XNOR U587 ( .A(n332), .B(n331), .Z(n319) );
  XOR U588 ( .A(n365), .B(n328), .Z(n331) );
  XNOR U589 ( .A(n366), .B(n323), .Z(n328) );
  NAND U590 ( .A(n327), .B(n227), .Z(n323) );
  NANDN U591 ( .B(n201), .A(n368), .Z(n367) );
  XNOR U592 ( .A(n329), .B(n330), .Z(n365) );
  XNOR U593 ( .A(n335), .B(n379), .Z(n338) );
  AND U594 ( .A(n262), .B(n295), .Z(n379) );
  XOR U595 ( .A(n380), .B(n381), .Z(n335) );
  ANDN U596 ( .A(n382), .B(n383), .Z(n381) );
  XNOR U597 ( .A(n384), .B(n380), .Z(n382) );
  XOR U598 ( .A(n385), .B(n339), .Z(n378) );
  NAND U599 ( .A(n257), .B(n299), .Z(n339) );
  IV U600 ( .A(n341), .Z(n385) );
  XNOR U601 ( .A(n348), .B(n349), .Z(n343) );
  NANDN U602 ( .B(n202), .A(n389), .Z(n349) );
  AND U603 ( .A(n344), .B(n226), .Z(n390) );
  NAND U604 ( .A(n391), .B(n392), .Z(n347) );
  NANDN U605 ( .B(n393), .A(n394), .Z(n391) );
  NAND U606 ( .A(n397), .B(n398), .Z(\_MxM/n224 ) );
  NANDN U607 ( .B(n117), .A(o[7]), .Z(n398) );
  AND U608 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U609 ( .B(n164), .A(o[7]), .Z(n400) );
  NANDN U610 ( .B(n169), .A(n139), .Z(n399) );
  XNOR U611 ( .A(n396), .B(\_MxM/Y0[8] ), .Z(n139) );
  XNOR U612 ( .A(n401), .B(n402), .Z(n396) );
  AND U613 ( .A(n180), .B(n404), .Z(n403) );
  XOR U614 ( .A(n361), .B(n405), .Z(n404) );
  XOR U615 ( .A(n405), .B(n362), .Z(n361) );
  OR U616 ( .A(n406), .B(n407), .Z(n362) );
  IV U617 ( .A(n402), .Z(n405) );
  XNOR U618 ( .A(n364), .B(n363), .Z(n402) );
  NANDN U619 ( .B(n408), .A(n409), .Z(n363) );
  XNOR U620 ( .A(n374), .B(n373), .Z(n364) );
  XOR U621 ( .A(n410), .B(n377), .Z(n373) );
  XNOR U622 ( .A(n370), .B(n371), .Z(n377) );
  NAND U623 ( .A(n327), .B(n262), .Z(n371) );
  XNOR U624 ( .A(n369), .B(n411), .Z(n370) );
  AND U625 ( .A(n227), .B(n368), .Z(n411) );
  XNOR U626 ( .A(n376), .B(n372), .Z(n410) );
  AND U627 ( .A(n419), .B(n420), .Z(n418) );
  NANDN U628 ( .B(n201), .A(n421), .Z(n420) );
  OR U629 ( .A(n422), .B(n423), .Z(n419) );
  XNOR U630 ( .A(n380), .B(n428), .Z(n383) );
  AND U631 ( .A(n299), .B(n295), .Z(n428) );
  XOR U632 ( .A(n429), .B(n430), .Z(n380) );
  ANDN U633 ( .A(n431), .B(n432), .Z(n430) );
  XNOR U634 ( .A(n433), .B(n429), .Z(n431) );
  XOR U635 ( .A(n434), .B(n384), .Z(n427) );
  NAND U636 ( .A(n257), .B(n344), .Z(n384) );
  IV U637 ( .A(n386), .Z(n434) );
  XNOR U638 ( .A(n393), .B(n394), .Z(n388) );
  NANDN U639 ( .B(n202), .A(n438), .Z(n394) );
  XNOR U640 ( .A(n392), .B(n439), .Z(n393) );
  AND U641 ( .A(n389), .B(n226), .Z(n439) );
  ANDN U642 ( .A(n440), .B(n441), .Z(n392) );
  NANDN U643 ( .B(n442), .A(n443), .Z(n440) );
  NAND U644 ( .A(n446), .B(n447), .Z(\_MxM/n223 ) );
  NANDN U645 ( .B(n117), .A(o[6]), .Z(n447) );
  AND U646 ( .A(n448), .B(n449), .Z(n446) );
  NANDN U647 ( .B(n164), .A(o[6]), .Z(n449) );
  NANDN U648 ( .B(n169), .A(n136), .Z(n448) );
  XNOR U649 ( .A(n445), .B(\_MxM/Y0[7] ), .Z(n136) );
  XNOR U650 ( .A(n451), .B(n452), .Z(n450) );
  AND U651 ( .A(n180), .B(n453), .Z(n452) );
  XOR U652 ( .A(n406), .B(n456), .Z(n453) );
  XOR U653 ( .A(n456), .B(n407), .Z(n406) );
  OR U654 ( .A(n454), .B(n455), .Z(n407) );
  XNOR U655 ( .A(n408), .B(n409), .Z(n456) );
  XNOR U656 ( .A(n417), .B(n416), .Z(n408) );
  XOR U657 ( .A(n461), .B(n426), .Z(n416) );
  XNOR U658 ( .A(n413), .B(n414), .Z(n426) );
  NAND U659 ( .A(n327), .B(n299), .Z(n414) );
  XNOR U660 ( .A(n412), .B(n462), .Z(n413) );
  AND U661 ( .A(n262), .B(n368), .Z(n462) );
  XNOR U662 ( .A(n425), .B(n415), .Z(n461) );
  XNOR U663 ( .A(n469), .B(n424), .Z(n425) );
  XNOR U664 ( .A(n473), .B(n422), .Z(n469) );
  NAND U665 ( .A(n421), .B(n227), .Z(n422) );
  NANDN U666 ( .B(n201), .A(n475), .Z(n474) );
  XNOR U667 ( .A(n429), .B(n480), .Z(n432) );
  AND U668 ( .A(n344), .B(n295), .Z(n480) );
  XOR U669 ( .A(n481), .B(n482), .Z(n429) );
  ANDN U670 ( .A(n483), .B(n484), .Z(n482) );
  XNOR U671 ( .A(n485), .B(n481), .Z(n483) );
  XOR U672 ( .A(n486), .B(n433), .Z(n479) );
  NAND U673 ( .A(n257), .B(n389), .Z(n433) );
  IV U674 ( .A(n435), .Z(n486) );
  XNOR U675 ( .A(n442), .B(n443), .Z(n437) );
  NANDN U676 ( .B(n202), .A(n490), .Z(n443) );
  AND U677 ( .A(n438), .B(n226), .Z(n491) );
  NAND U678 ( .A(n492), .B(n493), .Z(n441) );
  NANDN U679 ( .B(n494), .A(n495), .Z(n492) );
  IV U680 ( .A(n444), .Z(n451) );
  NAND U681 ( .A(n498), .B(n499), .Z(\_MxM/n222 ) );
  NANDN U682 ( .B(n117), .A(o[5]), .Z(n499) );
  AND U683 ( .A(n500), .B(n501), .Z(n498) );
  NANDN U684 ( .B(n164), .A(o[5]), .Z(n501) );
  NANDN U685 ( .B(n169), .A(n133), .Z(n500) );
  XNOR U686 ( .A(n497), .B(\_MxM/Y0[6] ), .Z(n133) );
  XNOR U687 ( .A(n502), .B(n503), .Z(n497) );
  AND U688 ( .A(n180), .B(n505), .Z(n504) );
  XOR U689 ( .A(n454), .B(n506), .Z(n505) );
  XOR U690 ( .A(n506), .B(n455), .Z(n454) );
  OR U691 ( .A(n507), .B(n508), .Z(n455) );
  IV U692 ( .A(n503), .Z(n506) );
  XOR U693 ( .A(n460), .B(n459), .Z(n503) );
  XNOR U694 ( .A(n458), .B(n509), .Z(n459) );
  AND U695 ( .A(n457), .B(n510), .Z(n509) );
  AND U696 ( .A(n511), .B(n512), .Z(n510) );
  NANDN U697 ( .B(n201), .A(n513), .Z(n512) );
  OR U698 ( .A(n514), .B(n515), .Z(n511) );
  AND U699 ( .A(n516), .B(n517), .Z(n457) );
  NANDN U700 ( .B(n518), .A(n519), .Z(n517) );
  NANDN U701 ( .B(n520), .A(n521), .Z(n516) );
  XNOR U702 ( .A(n525), .B(n472), .Z(n467) );
  XNOR U703 ( .A(n464), .B(n465), .Z(n472) );
  NAND U704 ( .A(n327), .B(n344), .Z(n465) );
  XNOR U705 ( .A(n463), .B(n526), .Z(n464) );
  AND U706 ( .A(n299), .B(n368), .Z(n526) );
  XNOR U707 ( .A(n471), .B(n466), .Z(n525) );
  XNOR U708 ( .A(n476), .B(n534), .Z(n477) );
  AND U709 ( .A(n227), .B(n475), .Z(n534) );
  XOR U710 ( .A(n535), .B(n536), .Z(n476) );
  ANDN U711 ( .A(n537), .B(n538), .Z(n536) );
  XNOR U712 ( .A(n539), .B(n535), .Z(n537) );
  XOR U713 ( .A(n540), .B(n478), .Z(n533) );
  NAND U714 ( .A(n421), .B(n262), .Z(n478) );
  IV U715 ( .A(n470), .Z(n540) );
  XNOR U716 ( .A(n481), .B(n545), .Z(n484) );
  AND U717 ( .A(n389), .B(n295), .Z(n545) );
  XOR U718 ( .A(n546), .B(n547), .Z(n481) );
  ANDN U719 ( .A(n548), .B(n549), .Z(n547) );
  XNOR U720 ( .A(n550), .B(n546), .Z(n548) );
  XOR U721 ( .A(n551), .B(n485), .Z(n544) );
  NAND U722 ( .A(n257), .B(n438), .Z(n485) );
  IV U723 ( .A(n487), .Z(n551) );
  XNOR U724 ( .A(n494), .B(n495), .Z(n489) );
  NANDN U725 ( .B(n202), .A(n555), .Z(n495) );
  XNOR U726 ( .A(n493), .B(n556), .Z(n494) );
  AND U727 ( .A(n490), .B(n226), .Z(n556) );
  ANDN U728 ( .A(n557), .B(n558), .Z(n493) );
  NANDN U729 ( .B(n559), .A(n560), .Z(n557) );
  NAND U730 ( .A(n563), .B(n564), .Z(\_MxM/n221 ) );
  NANDN U731 ( .B(n117), .A(o[4]), .Z(n564) );
  AND U732 ( .A(n565), .B(n566), .Z(n563) );
  NANDN U733 ( .B(n164), .A(o[4]), .Z(n566) );
  NANDN U734 ( .B(n169), .A(n130), .Z(n565) );
  XNOR U735 ( .A(n562), .B(\_MxM/Y0[5] ), .Z(n130) );
  XNOR U736 ( .A(n567), .B(n568), .Z(n562) );
  AND U737 ( .A(n180), .B(n570), .Z(n569) );
  XOR U738 ( .A(n507), .B(n571), .Z(n570) );
  XOR U739 ( .A(n571), .B(n508), .Z(n507) );
  OR U740 ( .A(n572), .B(n573), .Z(n508) );
  IV U741 ( .A(n568), .Z(n571) );
  XOR U742 ( .A(n524), .B(n523), .Z(n568) );
  XOR U743 ( .A(n518), .B(n519), .Z(n515) );
  XOR U744 ( .A(n578), .B(n520), .Z(n518) );
  NAND U745 ( .A(n227), .B(n513), .Z(n520) );
  NANDN U746 ( .B(n521), .A(n579), .Z(n578) );
  NANDN U747 ( .B(n201), .A(n580), .Z(n579) );
  XOR U748 ( .A(n584), .B(n514), .Z(n574) );
  OR U749 ( .A(n585), .B(n586), .Z(n514) );
  IV U750 ( .A(n522), .Z(n584) );
  XNOR U751 ( .A(n590), .B(n543), .Z(n531) );
  XNOR U752 ( .A(n528), .B(n529), .Z(n543) );
  NAND U753 ( .A(n327), .B(n389), .Z(n529) );
  XNOR U754 ( .A(n527), .B(n591), .Z(n528) );
  AND U755 ( .A(n344), .B(n368), .Z(n591) );
  XNOR U756 ( .A(n542), .B(n530), .Z(n590) );
  XNOR U757 ( .A(n535), .B(n599), .Z(n538) );
  AND U758 ( .A(n262), .B(n475), .Z(n599) );
  XOR U759 ( .A(n600), .B(n601), .Z(n535) );
  ANDN U760 ( .A(n602), .B(n603), .Z(n601) );
  XNOR U761 ( .A(n604), .B(n600), .Z(n602) );
  XOR U762 ( .A(n605), .B(n539), .Z(n598) );
  NAND U763 ( .A(n421), .B(n299), .Z(n539) );
  IV U764 ( .A(n541), .Z(n605) );
  XNOR U765 ( .A(n546), .B(n610), .Z(n549) );
  AND U766 ( .A(n438), .B(n295), .Z(n610) );
  XOR U767 ( .A(n611), .B(n612), .Z(n546) );
  ANDN U768 ( .A(n613), .B(n614), .Z(n612) );
  XNOR U769 ( .A(n615), .B(n611), .Z(n613) );
  XOR U770 ( .A(n616), .B(n550), .Z(n609) );
  NAND U771 ( .A(n257), .B(n490), .Z(n550) );
  IV U772 ( .A(n552), .Z(n616) );
  XNOR U773 ( .A(n559), .B(n560), .Z(n554) );
  NANDN U774 ( .B(n202), .A(n620), .Z(n560) );
  AND U775 ( .A(n555), .B(n226), .Z(n621) );
  NAND U776 ( .A(n622), .B(n623), .Z(n558) );
  NANDN U777 ( .B(n624), .A(n625), .Z(n622) );
  NAND U778 ( .A(n628), .B(n629), .Z(\_MxM/n220 ) );
  NANDN U779 ( .B(n117), .A(o[3]), .Z(n629) );
  AND U780 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U781 ( .B(n164), .A(o[3]), .Z(n631) );
  NANDN U782 ( .B(n169), .A(n127), .Z(n630) );
  XNOR U783 ( .A(n627), .B(\_MxM/Y0[4] ), .Z(n127) );
  XNOR U784 ( .A(n632), .B(n633), .Z(n627) );
  AND U785 ( .A(n180), .B(n635), .Z(n634) );
  XOR U786 ( .A(n572), .B(n636), .Z(n635) );
  XOR U787 ( .A(n636), .B(n573), .Z(n572) );
  OR U788 ( .A(n637), .B(n638), .Z(n573) );
  IV U789 ( .A(n633), .Z(n636) );
  XOR U790 ( .A(n589), .B(n588), .Z(n633) );
  XOR U791 ( .A(n639), .B(n585), .Z(n588) );
  XOR U792 ( .A(n577), .B(n576), .Z(n585) );
  XOR U793 ( .A(n575), .B(n640), .Z(n576) );
  AND U794 ( .A(n641), .B(n642), .Z(n640) );
  NANDN U795 ( .B(n201), .A(n643), .Z(n642) );
  OR U796 ( .A(n644), .B(n645), .Z(n641) );
  NAND U797 ( .A(n262), .B(n513), .Z(n583) );
  XNOR U798 ( .A(n581), .B(n649), .Z(n582) );
  AND U799 ( .A(n580), .B(n227), .Z(n649) );
  NANDN U800 ( .B(n653), .A(n654), .Z(n586) );
  XNOR U801 ( .A(n658), .B(n608), .Z(n596) );
  XNOR U802 ( .A(n593), .B(n594), .Z(n608) );
  NAND U803 ( .A(n327), .B(n438), .Z(n594) );
  XNOR U804 ( .A(n592), .B(n659), .Z(n593) );
  AND U805 ( .A(n389), .B(n368), .Z(n659) );
  XNOR U806 ( .A(n607), .B(n595), .Z(n658) );
  XNOR U807 ( .A(n600), .B(n667), .Z(n603) );
  AND U808 ( .A(n299), .B(n475), .Z(n667) );
  XOR U809 ( .A(n668), .B(n669), .Z(n600) );
  ANDN U810 ( .A(n670), .B(n671), .Z(n669) );
  XNOR U811 ( .A(n672), .B(n668), .Z(n670) );
  XOR U812 ( .A(n673), .B(n604), .Z(n666) );
  NAND U813 ( .A(n421), .B(n344), .Z(n604) );
  IV U814 ( .A(n606), .Z(n673) );
  XNOR U815 ( .A(n611), .B(n678), .Z(n614) );
  AND U816 ( .A(n490), .B(n295), .Z(n678) );
  XOR U817 ( .A(n679), .B(n680), .Z(n611) );
  ANDN U818 ( .A(n681), .B(n682), .Z(n680) );
  XNOR U819 ( .A(n683), .B(n679), .Z(n681) );
  XOR U820 ( .A(n684), .B(n615), .Z(n677) );
  NAND U821 ( .A(n257), .B(n555), .Z(n615) );
  IV U822 ( .A(n617), .Z(n684) );
  XNOR U823 ( .A(n624), .B(n625), .Z(n619) );
  NANDN U824 ( .B(n202), .A(n688), .Z(n625) );
  XNOR U825 ( .A(n623), .B(n689), .Z(n624) );
  AND U826 ( .A(n620), .B(n226), .Z(n689) );
  ANDN U827 ( .A(n690), .B(n691), .Z(n623) );
  NANDN U828 ( .B(n692), .A(n693), .Z(n690) );
  NAND U829 ( .A(n696), .B(n697), .Z(\_MxM/n219 ) );
  NANDN U830 ( .B(n117), .A(o[2]), .Z(n697) );
  AND U831 ( .A(n698), .B(n699), .Z(n696) );
  NANDN U832 ( .B(n164), .A(o[2]), .Z(n699) );
  NANDN U833 ( .B(n169), .A(n124), .Z(n698) );
  XNOR U834 ( .A(n695), .B(\_MxM/Y0[3] ), .Z(n124) );
  XNOR U835 ( .A(n700), .B(n701), .Z(n695) );
  AND U836 ( .A(n180), .B(n703), .Z(n702) );
  XOR U837 ( .A(n637), .B(n704), .Z(n703) );
  XOR U838 ( .A(n704), .B(n638), .Z(n637) );
  OR U839 ( .A(n705), .B(n706), .Z(n638) );
  IV U840 ( .A(n701), .Z(n704) );
  XOR U841 ( .A(n657), .B(n656), .Z(n701) );
  XOR U842 ( .A(n707), .B(n653), .Z(n656) );
  XOR U843 ( .A(n648), .B(n647), .Z(n653) );
  XNOR U844 ( .A(n712), .B(n644), .Z(n708) );
  NAND U845 ( .A(n227), .B(n643), .Z(n644) );
  NANDN U846 ( .B(n201), .A(n714), .Z(n713) );
  NAND U847 ( .A(n299), .B(n513), .Z(n652) );
  XNOR U848 ( .A(n650), .B(n718), .Z(n651) );
  AND U849 ( .A(n580), .B(n262), .Z(n718) );
  XNOR U850 ( .A(n654), .B(n655), .Z(n707) );
  XNOR U851 ( .A(n728), .B(n676), .Z(n664) );
  XNOR U852 ( .A(n661), .B(n662), .Z(n676) );
  NAND U853 ( .A(n327), .B(n490), .Z(n662) );
  XNOR U854 ( .A(n660), .B(n729), .Z(n661) );
  AND U855 ( .A(n438), .B(n368), .Z(n729) );
  XNOR U856 ( .A(n675), .B(n663), .Z(n728) );
  XNOR U857 ( .A(n668), .B(n737), .Z(n671) );
  AND U858 ( .A(n344), .B(n475), .Z(n737) );
  XOR U859 ( .A(n741), .B(n672), .Z(n736) );
  NAND U860 ( .A(n421), .B(n389), .Z(n672) );
  IV U861 ( .A(n674), .Z(n741) );
  XNOR U862 ( .A(n679), .B(n746), .Z(n682) );
  AND U863 ( .A(n555), .B(n295), .Z(n746) );
  XOR U864 ( .A(n747), .B(n748), .Z(n679) );
  ANDN U865 ( .A(n749), .B(n750), .Z(n748) );
  XNOR U866 ( .A(n751), .B(n747), .Z(n749) );
  XOR U867 ( .A(n752), .B(n683), .Z(n745) );
  NAND U868 ( .A(n257), .B(n620), .Z(n683) );
  IV U869 ( .A(n685), .Z(n752) );
  XNOR U870 ( .A(n692), .B(n693), .Z(n687) );
  OR U871 ( .A(n756), .B(n202), .Z(n693) );
  AND U872 ( .A(n688), .B(n226), .Z(n757) );
  NAND U873 ( .A(n758), .B(n759), .Z(n691) );
  NANDN U874 ( .B(n760), .A(n761), .Z(n758) );
  NAND U875 ( .A(n764), .B(n765), .Z(\_MxM/n218 ) );
  NANDN U876 ( .B(n117), .A(o[1]), .Z(n765) );
  AND U877 ( .A(n766), .B(n767), .Z(n764) );
  NANDN U878 ( .B(n164), .A(o[1]), .Z(n767) );
  NANDN U879 ( .B(n169), .A(n120), .Z(n766) );
  XNOR U880 ( .A(n763), .B(\_MxM/Y0[2] ), .Z(n120) );
  XNOR U881 ( .A(n768), .B(n769), .Z(n763) );
  XOR U882 ( .A(n762), .B(n770), .Z(n768) );
  AND U883 ( .A(n180), .B(n771), .Z(n770) );
  XOR U884 ( .A(n705), .B(n772), .Z(n771) );
  XOR U885 ( .A(n772), .B(n706), .Z(n705) );
  NANDN U886 ( .B(n773), .A(n774), .Z(n706) );
  IV U887 ( .A(n769), .Z(n772) );
  XOR U888 ( .A(n724), .B(n723), .Z(n769) );
  XNOR U889 ( .A(n775), .B(n727), .Z(n723) );
  XNOR U890 ( .A(n715), .B(n777), .Z(n716) );
  AND U891 ( .A(n714), .B(n227), .Z(n777) );
  XOR U892 ( .A(n781), .B(n717), .Z(n776) );
  NAND U893 ( .A(n262), .B(n643), .Z(n717) );
  IV U894 ( .A(n709), .Z(n781) );
  XNOR U895 ( .A(n720), .B(n721), .Z(n711) );
  NAND U896 ( .A(n344), .B(n513), .Z(n721) );
  XNOR U897 ( .A(n719), .B(n785), .Z(n720) );
  AND U898 ( .A(n580), .B(n299), .Z(n785) );
  XNOR U899 ( .A(n726), .B(n722), .Z(n775) );
  AND U900 ( .A(n793), .B(n794), .Z(n792) );
  OR U901 ( .A(n795), .B(n796), .Z(n794) );
  AND U902 ( .A(n797), .B(n798), .Z(n793) );
  NANDN U903 ( .B(n201), .A(n799), .Z(n798) );
  NANDN U904 ( .B(n800), .A(n801), .Z(n797) );
  XNOR U905 ( .A(n805), .B(n744), .Z(n734) );
  XNOR U906 ( .A(n731), .B(n732), .Z(n744) );
  NAND U907 ( .A(n327), .B(n555), .Z(n732) );
  XNOR U908 ( .A(n730), .B(n806), .Z(n731) );
  AND U909 ( .A(n490), .B(n368), .Z(n806) );
  XNOR U910 ( .A(n743), .B(n733), .Z(n805) );
  XNOR U911 ( .A(n738), .B(n814), .Z(n739) );
  AND U912 ( .A(n389), .B(n475), .Z(n814) );
  XOR U913 ( .A(n818), .B(n740), .Z(n813) );
  NAND U914 ( .A(n421), .B(n438), .Z(n740) );
  IV U915 ( .A(n742), .Z(n818) );
  XNOR U916 ( .A(n747), .B(n823), .Z(n750) );
  AND U917 ( .A(n620), .B(n295), .Z(n823) );
  XOR U918 ( .A(n824), .B(n825), .Z(n747) );
  ANDN U919 ( .A(n826), .B(n827), .Z(n825) );
  XNOR U920 ( .A(n828), .B(n824), .Z(n826) );
  XOR U921 ( .A(n829), .B(n751), .Z(n822) );
  NAND U922 ( .A(n257), .B(n688), .Z(n751) );
  IV U923 ( .A(n753), .Z(n829) );
  XNOR U924 ( .A(n760), .B(n761), .Z(n755) );
  OR U925 ( .A(n833), .B(n202), .Z(n761) );
  XNOR U926 ( .A(n759), .B(n834), .Z(n760) );
  ANDN U927 ( .A(n226), .B(n756), .Z(n834) );
  ANDN U928 ( .A(n835), .B(n836), .Z(n759) );
  NANDN U929 ( .B(n837), .A(n838), .Z(n835) );
  NAND U930 ( .A(n841), .B(n842), .Z(\_MxM/n217 ) );
  NANDN U931 ( .B(n117), .A(o[0]), .Z(n842) );
  AND U932 ( .A(n843), .B(n844), .Z(n841) );
  NANDN U933 ( .B(n164), .A(o[0]), .Z(n844) );
  IV U934 ( .A(n845), .Z(n164) );
  OR U935 ( .A(n169), .B(n115), .Z(n843) );
  IV U936 ( .A(\_MxM/Y0[1] ), .Z(n121) );
  XOR U937 ( .A(n846), .B(n847), .Z(n840) );
  XNOR U938 ( .A(n848), .B(n839), .Z(n846) );
  NAND U939 ( .A(\_MxM/Y0[0] ), .B(n773), .Z(n839) );
  NAND U940 ( .A(n849), .B(n180), .Z(n848) );
  XOR U941 ( .A(e_input[15]), .B(g_input[15]), .Z(n180) );
  XNOR U942 ( .A(n774), .B(n847), .Z(n849) );
  XNOR U943 ( .A(n773), .B(n847), .Z(n774) );
  XNOR U944 ( .A(n791), .B(n790), .Z(n847) );
  XNOR U945 ( .A(n850), .B(n804), .Z(n790) );
  XNOR U946 ( .A(n778), .B(n852), .Z(n779) );
  AND U947 ( .A(n714), .B(n262), .Z(n852) );
  XOR U948 ( .A(n856), .B(n780), .Z(n851) );
  NAND U949 ( .A(n299), .B(n643), .Z(n780) );
  IV U950 ( .A(n782), .Z(n856) );
  XNOR U951 ( .A(n787), .B(n788), .Z(n784) );
  NAND U952 ( .A(n389), .B(n513), .Z(n788) );
  XNOR U953 ( .A(n786), .B(n860), .Z(n787) );
  AND U954 ( .A(n580), .B(n344), .Z(n860) );
  XNOR U955 ( .A(n803), .B(n789), .Z(n850) );
  XNOR U956 ( .A(n867), .B(n800), .Z(n803) );
  XOR U957 ( .A(n868), .B(n795), .Z(n800) );
  NAND U958 ( .A(n227), .B(n799), .Z(n795) );
  NANDN U959 ( .B(n201), .A(n870), .Z(n869) );
  XNOR U960 ( .A(n801), .B(n802), .Z(n867) );
  XNOR U961 ( .A(n880), .B(n821), .Z(n811) );
  XNOR U962 ( .A(n808), .B(n809), .Z(n821) );
  NAND U963 ( .A(n327), .B(n620), .Z(n809) );
  XNOR U964 ( .A(n807), .B(n881), .Z(n808) );
  AND U965 ( .A(n555), .B(n368), .Z(n881) );
  XNOR U966 ( .A(n820), .B(n810), .Z(n880) );
  XNOR U967 ( .A(n815), .B(n889), .Z(n816) );
  AND U968 ( .A(n438), .B(n475), .Z(n889) );
  XOR U969 ( .A(n893), .B(n817), .Z(n888) );
  NAND U970 ( .A(n421), .B(n490), .Z(n817) );
  IV U971 ( .A(n819), .Z(n893) );
  XNOR U972 ( .A(n824), .B(n898), .Z(n827) );
  AND U973 ( .A(n688), .B(n295), .Z(n898) );
  XOR U974 ( .A(n902), .B(n828), .Z(n897) );
  NANDN U975 ( .B(n756), .A(n257), .Z(n828) );
  IV U976 ( .A(n830), .Z(n902) );
  XNOR U977 ( .A(n837), .B(n838), .Z(n832) );
  NANDN U978 ( .B(n202), .A(n906), .Z(n838) );
  ANDN U979 ( .A(n226), .B(n833), .Z(n907) );
  NAND U980 ( .A(n908), .B(n909), .Z(n836) );
  NANDN U981 ( .B(n910), .A(n911), .Z(n908) );
  XNOR U982 ( .A(n866), .B(n865), .Z(n773) );
  XNOR U983 ( .A(n912), .B(n876), .Z(n865) );
  XNOR U984 ( .A(n853), .B(n914), .Z(n854) );
  AND U985 ( .A(n714), .B(n299), .Z(n914) );
  XOR U986 ( .A(n918), .B(n855), .Z(n913) );
  NAND U987 ( .A(n344), .B(n643), .Z(n855) );
  IV U988 ( .A(n857), .Z(n918) );
  XNOR U989 ( .A(n862), .B(n863), .Z(n859) );
  NAND U990 ( .A(n438), .B(n513), .Z(n863) );
  XNOR U991 ( .A(n861), .B(n922), .Z(n862) );
  AND U992 ( .A(n580), .B(n389), .Z(n922) );
  XNOR U993 ( .A(n875), .B(n864), .Z(n912) );
  XOR U994 ( .A(n926), .B(n927), .Z(n864) );
  XNOR U995 ( .A(n928), .B(n879), .Z(n875) );
  NAND U996 ( .A(n262), .B(n799), .Z(n873) );
  XNOR U997 ( .A(n871), .B(n929), .Z(n872) );
  AND U998 ( .A(n870), .B(n227), .Z(n929) );
  XNOR U999 ( .A(n878), .B(n874), .Z(n928) );
  XOR U1000 ( .A(n933), .B(n934), .Z(n874) );
  AND U1001 ( .A(n935), .B(n936), .Z(n934) );
  XOR U1002 ( .A(n937), .B(n938), .Z(n936) );
  XOR U1003 ( .A(n933), .B(n939), .Z(n938) );
  XOR U1004 ( .A(n920), .B(n940), .Z(n935) );
  XOR U1005 ( .A(n933), .B(n921), .Z(n940) );
  NAND U1006 ( .A(n513), .B(n490), .Z(n925) );
  XNOR U1007 ( .A(n923), .B(n941), .Z(n924) );
  AND U1008 ( .A(n580), .B(n438), .Z(n941) );
  XNOR U1009 ( .A(n915), .B(n946), .Z(n916) );
  AND U1010 ( .A(n714), .B(n344), .Z(n946) );
  XOR U1011 ( .A(n947), .B(n948), .Z(n915) );
  ANDN U1012 ( .A(n949), .B(n950), .Z(n948) );
  XNOR U1013 ( .A(n951), .B(n947), .Z(n949) );
  XOR U1014 ( .A(n952), .B(n917), .Z(n945) );
  NAND U1015 ( .A(n389), .B(n643), .Z(n917) );
  IV U1016 ( .A(n919), .Z(n952) );
  XOR U1017 ( .A(n956), .B(n957), .Z(n933) );
  AND U1018 ( .A(n958), .B(n959), .Z(n957) );
  XOR U1019 ( .A(n960), .B(n961), .Z(n959) );
  XOR U1020 ( .A(n956), .B(n962), .Z(n961) );
  XOR U1021 ( .A(n954), .B(n963), .Z(n958) );
  XOR U1022 ( .A(n956), .B(n955), .Z(n963) );
  NAND U1023 ( .A(n513), .B(n555), .Z(n944) );
  XNOR U1024 ( .A(n942), .B(n964), .Z(n943) );
  AND U1025 ( .A(n490), .B(n580), .Z(n964) );
  XNOR U1026 ( .A(n947), .B(n969), .Z(n950) );
  AND U1027 ( .A(n714), .B(n389), .Z(n969) );
  XOR U1028 ( .A(n970), .B(n971), .Z(n947) );
  ANDN U1029 ( .A(n972), .B(n973), .Z(n971) );
  XNOR U1030 ( .A(n974), .B(n970), .Z(n972) );
  XOR U1031 ( .A(n975), .B(n951), .Z(n968) );
  NAND U1032 ( .A(n438), .B(n643), .Z(n951) );
  IV U1033 ( .A(n953), .Z(n975) );
  XOR U1034 ( .A(n979), .B(n980), .Z(n956) );
  AND U1035 ( .A(n981), .B(n982), .Z(n980) );
  XOR U1036 ( .A(n983), .B(n984), .Z(n982) );
  XOR U1037 ( .A(n979), .B(n985), .Z(n984) );
  XOR U1038 ( .A(n977), .B(n986), .Z(n981) );
  XOR U1039 ( .A(n979), .B(n978), .Z(n986) );
  NAND U1040 ( .A(n513), .B(n620), .Z(n967) );
  XNOR U1041 ( .A(n965), .B(n987), .Z(n966) );
  AND U1042 ( .A(n555), .B(n580), .Z(n987) );
  XNOR U1043 ( .A(n970), .B(n992), .Z(n973) );
  AND U1044 ( .A(n714), .B(n438), .Z(n992) );
  XOR U1045 ( .A(n993), .B(n994), .Z(n970) );
  ANDN U1046 ( .A(n995), .B(n996), .Z(n994) );
  XNOR U1047 ( .A(n997), .B(n993), .Z(n995) );
  XOR U1048 ( .A(n998), .B(n974), .Z(n991) );
  NAND U1049 ( .A(n643), .B(n490), .Z(n974) );
  IV U1050 ( .A(n976), .Z(n998) );
  XOR U1051 ( .A(n1002), .B(n1003), .Z(n979) );
  AND U1052 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U1053 ( .A(n1006), .B(n1007), .Z(n1005) );
  XOR U1054 ( .A(n1002), .B(n1008), .Z(n1007) );
  XOR U1055 ( .A(n1000), .B(n1009), .Z(n1004) );
  XOR U1056 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U1057 ( .A(n1010), .B(n990), .Z(n1001) );
  NAND U1058 ( .A(n513), .B(n688), .Z(n990) );
  IV U1059 ( .A(n989), .Z(n1010) );
  XNOR U1060 ( .A(n988), .B(n1011), .Z(n989) );
  AND U1061 ( .A(n620), .B(n580), .Z(n1011) );
  XOR U1062 ( .A(n1012), .B(n1013), .Z(n988) );
  ANDN U1063 ( .A(n1014), .B(n1015), .Z(n1013) );
  XNOR U1064 ( .A(n1016), .B(n1012), .Z(n1014) );
  XNOR U1065 ( .A(n1017), .B(n1018), .Z(n1000) );
  IV U1066 ( .A(n996), .Z(n1018) );
  XNOR U1067 ( .A(n993), .B(n1019), .Z(n996) );
  AND U1068 ( .A(n490), .B(n714), .Z(n1019) );
  XOR U1069 ( .A(n1020), .B(n1021), .Z(n993) );
  ANDN U1070 ( .A(n1022), .B(n1023), .Z(n1021) );
  XNOR U1071 ( .A(n1024), .B(n1020), .Z(n1022) );
  XOR U1072 ( .A(n1025), .B(n997), .Z(n1017) );
  NAND U1073 ( .A(n643), .B(n555), .Z(n997) );
  IV U1074 ( .A(n999), .Z(n1025) );
  XOR U1075 ( .A(n1029), .B(n1030), .Z(n1002) );
  AND U1076 ( .A(n1031), .B(n1032), .Z(n1030) );
  XOR U1077 ( .A(n1033), .B(n1034), .Z(n1032) );
  XOR U1078 ( .A(n1029), .B(n1035), .Z(n1034) );
  XOR U1079 ( .A(n1027), .B(n1036), .Z(n1031) );
  XOR U1080 ( .A(n1029), .B(n1028), .Z(n1036) );
  XNOR U1081 ( .A(n1037), .B(n1016), .Z(n1028) );
  NANDN U1082 ( .B(n756), .A(n513), .Z(n1016) );
  IV U1083 ( .A(n1015), .Z(n1037) );
  XNOR U1084 ( .A(n1012), .B(n1038), .Z(n1015) );
  AND U1085 ( .A(n688), .B(n580), .Z(n1038) );
  XOR U1086 ( .A(n1039), .B(n1040), .Z(n1012) );
  ANDN U1087 ( .A(n1041), .B(n1042), .Z(n1040) );
  XNOR U1088 ( .A(n1043), .B(n1039), .Z(n1041) );
  XNOR U1089 ( .A(n1044), .B(n1045), .Z(n1027) );
  IV U1090 ( .A(n1023), .Z(n1045) );
  XNOR U1091 ( .A(n1020), .B(n1046), .Z(n1023) );
  AND U1092 ( .A(n555), .B(n714), .Z(n1046) );
  XOR U1093 ( .A(n1047), .B(n1048), .Z(n1020) );
  ANDN U1094 ( .A(n1049), .B(n1050), .Z(n1048) );
  XNOR U1095 ( .A(n1051), .B(n1047), .Z(n1049) );
  XOR U1096 ( .A(n1052), .B(n1024), .Z(n1044) );
  NAND U1097 ( .A(n643), .B(n620), .Z(n1024) );
  IV U1098 ( .A(n1026), .Z(n1052) );
  XOR U1099 ( .A(n1056), .B(n1057), .Z(n1029) );
  AND U1100 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR U1101 ( .A(n1060), .B(n1061), .Z(n1059) );
  XOR U1102 ( .A(n1056), .B(n1062), .Z(n1061) );
  XOR U1103 ( .A(n1054), .B(n1063), .Z(n1058) );
  XOR U1104 ( .A(n1056), .B(n1055), .Z(n1063) );
  XNOR U1105 ( .A(n1064), .B(n1043), .Z(n1055) );
  NANDN U1106 ( .B(n833), .A(n513), .Z(n1043) );
  IV U1107 ( .A(n1042), .Z(n1064) );
  XNOR U1108 ( .A(n1039), .B(n1065), .Z(n1042) );
  ANDN U1109 ( .A(n580), .B(n756), .Z(n1065) );
  XOR U1110 ( .A(n1066), .B(n1067), .Z(n1039) );
  ANDN U1111 ( .A(n1068), .B(n1069), .Z(n1067) );
  XNOR U1112 ( .A(n1070), .B(n1066), .Z(n1068) );
  XNOR U1113 ( .A(n1071), .B(n1072), .Z(n1054) );
  IV U1114 ( .A(n1050), .Z(n1072) );
  XNOR U1115 ( .A(n1047), .B(n1073), .Z(n1050) );
  AND U1116 ( .A(n620), .B(n714), .Z(n1073) );
  XOR U1117 ( .A(n1074), .B(n1075), .Z(n1047) );
  ANDN U1118 ( .A(n1076), .B(n1077), .Z(n1075) );
  XNOR U1119 ( .A(n1078), .B(n1074), .Z(n1076) );
  XOR U1120 ( .A(n1079), .B(n1051), .Z(n1071) );
  NAND U1121 ( .A(n643), .B(n688), .Z(n1051) );
  IV U1122 ( .A(n1053), .Z(n1079) );
  XOR U1123 ( .A(n1083), .B(n1084), .Z(n1056) );
  AND U1124 ( .A(n1085), .B(n1086), .Z(n1084) );
  XOR U1125 ( .A(n1087), .B(n1088), .Z(n1086) );
  XOR U1126 ( .A(n1083), .B(n1089), .Z(n1088) );
  XOR U1127 ( .A(n1081), .B(n1090), .Z(n1085) );
  XOR U1128 ( .A(n1083), .B(n1082), .Z(n1090) );
  XNOR U1129 ( .A(n1091), .B(n1070), .Z(n1082) );
  NAND U1130 ( .A(n513), .B(n906), .Z(n1070) );
  IV U1131 ( .A(n1069), .Z(n1091) );
  XNOR U1132 ( .A(n1066), .B(n1092), .Z(n1069) );
  ANDN U1133 ( .A(n580), .B(n833), .Z(n1092) );
  XOR U1134 ( .A(n1093), .B(n1094), .Z(n1066) );
  ANDN U1135 ( .A(n1095), .B(n1096), .Z(n1094) );
  XNOR U1136 ( .A(n1097), .B(n1093), .Z(n1095) );
  XNOR U1137 ( .A(n1098), .B(n1099), .Z(n1081) );
  IV U1138 ( .A(n1077), .Z(n1099) );
  XNOR U1139 ( .A(n1074), .B(n1100), .Z(n1077) );
  AND U1140 ( .A(n688), .B(n714), .Z(n1100) );
  XOR U1141 ( .A(n1101), .B(n1102), .Z(n1074) );
  ANDN U1142 ( .A(n1103), .B(n1104), .Z(n1102) );
  XNOR U1143 ( .A(n1105), .B(n1101), .Z(n1103) );
  XOR U1144 ( .A(n1106), .B(n1078), .Z(n1098) );
  NANDN U1145 ( .B(n756), .A(n643), .Z(n1078) );
  IV U1146 ( .A(n1080), .Z(n1106) );
  XOR U1147 ( .A(n1111), .B(n1112), .Z(n927) );
  XNOR U1148 ( .A(n1113), .B(n1110), .Z(n1111) );
  XNOR U1149 ( .A(n1101), .B(n1115), .Z(n1104) );
  ANDN U1150 ( .A(n714), .B(n756), .Z(n1115) );
  XOR U1151 ( .A(n1118), .B(n1116), .Z(n1117) );
  ANDN U1152 ( .A(n714), .B(n833), .Z(n1118) );
  AND U1153 ( .A(n906), .B(n643), .Z(n1119) );
  XOR U1154 ( .A(n1120), .B(n1121), .Z(n1116) );
  ANDN U1155 ( .A(n1122), .B(n1123), .Z(n1121) );
  XNOR U1156 ( .A(n1124), .B(n1120), .Z(n1122) );
  XOR U1157 ( .A(n1125), .B(n1105), .Z(n1114) );
  NANDN U1158 ( .B(n833), .A(n643), .Z(n1105) );
  IV U1159 ( .A(n1107), .Z(n1125) );
  NAND U1160 ( .A(n643), .B(n1126), .Z(n1124) );
  XNOR U1161 ( .A(n1120), .B(n1127), .Z(n1123) );
  AND U1162 ( .A(n906), .B(n714), .Z(n1127) );
  AND U1163 ( .A(n1128), .B(g_input[0]), .Z(n1120) );
  NANDN U1164 ( .B(n643), .A(n1129), .Z(n1128) );
  NAND U1165 ( .A(n1126), .B(n714), .Z(n1129) );
  XNOR U1166 ( .A(n1096), .B(n1097), .Z(n1109) );
  NAND U1167 ( .A(n513), .B(n1126), .Z(n1097) );
  XNOR U1168 ( .A(n1093), .B(n1132), .Z(n1096) );
  AND U1169 ( .A(n906), .B(n580), .Z(n1132) );
  AND U1170 ( .A(n1133), .B(g_input[0]), .Z(n1093) );
  NANDN U1171 ( .B(n513), .A(n1134), .Z(n1133) );
  NAND U1172 ( .A(n1126), .B(n580), .Z(n1134) );
  XOR U1173 ( .A(n1137), .B(n1138), .Z(n1110) );
  XOR U1174 ( .A(n1139), .B(n1140), .Z(n878) );
  AND U1175 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1176 ( .B(n201), .A(n1143), .Z(n1142) );
  NANDN U1177 ( .B(n1144), .A(n1145), .Z(n201) );
  AND U1178 ( .A(n1146), .B(g_input[15]), .Z(n1145) );
  OR U1179 ( .A(n1147), .B(n1148), .Z(n1141) );
  IV U1180 ( .A(n877), .Z(n1139) );
  NAND U1181 ( .A(n299), .B(n799), .Z(n932) );
  XNOR U1182 ( .A(n930), .B(n1150), .Z(n931) );
  AND U1183 ( .A(n870), .B(n262), .Z(n1150) );
  XOR U1184 ( .A(n1158), .B(n1147), .Z(n1154) );
  NAND U1185 ( .A(n227), .B(n1143), .Z(n1147) );
  IV U1186 ( .A(n1149), .Z(n1158) );
  NAND U1187 ( .A(n344), .B(n799), .Z(n1153) );
  XNOR U1188 ( .A(n1151), .B(n1160), .Z(n1152) );
  AND U1189 ( .A(n870), .B(n299), .Z(n1160) );
  XNOR U1190 ( .A(n1155), .B(n1165), .Z(n1156) );
  AND U1191 ( .A(n227), .B(e_input[0]), .Z(n1165) );
  XNOR U1192 ( .A(n1146), .B(g_input[14]), .Z(n1144) );
  NOR U1193 ( .A(n1166), .B(n1167), .Z(n1146) );
  XOR U1194 ( .A(n1171), .B(n1157), .Z(n1164) );
  NAND U1195 ( .A(n262), .B(n1143), .Z(n1157) );
  IV U1196 ( .A(n1159), .Z(n1171) );
  NAND U1197 ( .A(n389), .B(n799), .Z(n1163) );
  XNOR U1198 ( .A(n1161), .B(n1173), .Z(n1162) );
  AND U1199 ( .A(n870), .B(n344), .Z(n1173) );
  XOR U1200 ( .A(n1174), .B(n1175), .Z(n1161) );
  ANDN U1201 ( .A(n1176), .B(n1177), .Z(n1175) );
  XNOR U1202 ( .A(n1178), .B(n1174), .Z(n1176) );
  XNOR U1203 ( .A(n1168), .B(n1180), .Z(n1169) );
  AND U1204 ( .A(n262), .B(e_input[0]), .Z(n1180) );
  XOR U1205 ( .A(n1166), .B(g_input[13]), .Z(n1167) );
  NANDN U1206 ( .B(n1181), .A(n1182), .Z(n1166) );
  XOR U1207 ( .A(n1186), .B(n1170), .Z(n1179) );
  NAND U1208 ( .A(n299), .B(n1143), .Z(n1170) );
  IV U1209 ( .A(n1172), .Z(n1186) );
  XNOR U1210 ( .A(n1188), .B(n1178), .Z(n1006) );
  NAND U1211 ( .A(n438), .B(n799), .Z(n1178) );
  IV U1212 ( .A(n1177), .Z(n1188) );
  XNOR U1213 ( .A(n1174), .B(n1189), .Z(n1177) );
  AND U1214 ( .A(n870), .B(n389), .Z(n1189) );
  XOR U1215 ( .A(n1190), .B(n1191), .Z(n1174) );
  ANDN U1216 ( .A(n1192), .B(n1193), .Z(n1191) );
  XNOR U1217 ( .A(n1194), .B(n1190), .Z(n1192) );
  XNOR U1218 ( .A(n1195), .B(n1196), .Z(n1008) );
  IV U1219 ( .A(n1184), .Z(n1196) );
  XNOR U1220 ( .A(n1183), .B(n1197), .Z(n1184) );
  AND U1221 ( .A(n299), .B(e_input[0]), .Z(n1197) );
  XNOR U1222 ( .A(n1182), .B(g_input[12]), .Z(n1181) );
  NOR U1223 ( .A(n1198), .B(n1199), .Z(n1182) );
  XOR U1224 ( .A(n1200), .B(n1201), .Z(n1183) );
  ANDN U1225 ( .A(n1202), .B(n1203), .Z(n1201) );
  XNOR U1226 ( .A(n1204), .B(n1200), .Z(n1202) );
  XOR U1227 ( .A(n1205), .B(n1185), .Z(n1195) );
  NAND U1228 ( .A(n344), .B(n1143), .Z(n1185) );
  IV U1229 ( .A(n1187), .Z(n1205) );
  XNOR U1230 ( .A(n1207), .B(n1194), .Z(n1033) );
  NAND U1231 ( .A(n490), .B(n799), .Z(n1194) );
  IV U1232 ( .A(n1193), .Z(n1207) );
  XNOR U1233 ( .A(n1190), .B(n1208), .Z(n1193) );
  AND U1234 ( .A(n870), .B(n438), .Z(n1208) );
  XOR U1235 ( .A(n1209), .B(n1210), .Z(n1190) );
  ANDN U1236 ( .A(n1211), .B(n1212), .Z(n1210) );
  XNOR U1237 ( .A(n1213), .B(n1209), .Z(n1211) );
  XNOR U1238 ( .A(n1214), .B(n1215), .Z(n1035) );
  IV U1239 ( .A(n1203), .Z(n1215) );
  XNOR U1240 ( .A(n1200), .B(n1216), .Z(n1203) );
  AND U1241 ( .A(n344), .B(e_input[0]), .Z(n1216) );
  XOR U1242 ( .A(n1198), .B(g_input[11]), .Z(n1199) );
  NANDN U1243 ( .B(n1217), .A(n1218), .Z(n1198) );
  XOR U1244 ( .A(n1219), .B(n1220), .Z(n1200) );
  ANDN U1245 ( .A(n1221), .B(n1222), .Z(n1220) );
  XNOR U1246 ( .A(n1223), .B(n1219), .Z(n1221) );
  XOR U1247 ( .A(n1224), .B(n1204), .Z(n1214) );
  NAND U1248 ( .A(n389), .B(n1143), .Z(n1204) );
  IV U1249 ( .A(n1206), .Z(n1224) );
  XNOR U1250 ( .A(n1226), .B(n1213), .Z(n1060) );
  NAND U1251 ( .A(n555), .B(n799), .Z(n1213) );
  IV U1252 ( .A(n1212), .Z(n1226) );
  XNOR U1253 ( .A(n1209), .B(n1227), .Z(n1212) );
  AND U1254 ( .A(n870), .B(n490), .Z(n1227) );
  XOR U1255 ( .A(n1228), .B(n1229), .Z(n1209) );
  ANDN U1256 ( .A(n1230), .B(n1231), .Z(n1229) );
  XNOR U1257 ( .A(n1232), .B(n1228), .Z(n1230) );
  XNOR U1258 ( .A(n1233), .B(n1234), .Z(n1062) );
  IV U1259 ( .A(n1222), .Z(n1234) );
  XNOR U1260 ( .A(n1219), .B(n1235), .Z(n1222) );
  AND U1261 ( .A(n389), .B(e_input[0]), .Z(n1235) );
  XNOR U1262 ( .A(n1218), .B(g_input[10]), .Z(n1217) );
  NOR U1263 ( .A(n1236), .B(n1237), .Z(n1218) );
  XOR U1264 ( .A(n1238), .B(n1239), .Z(n1219) );
  ANDN U1265 ( .A(n1240), .B(n1241), .Z(n1239) );
  XNOR U1266 ( .A(n1242), .B(n1238), .Z(n1240) );
  XOR U1267 ( .A(n1243), .B(n1223), .Z(n1233) );
  NAND U1268 ( .A(n438), .B(n1143), .Z(n1223) );
  IV U1269 ( .A(n1225), .Z(n1243) );
  XNOR U1270 ( .A(n1245), .B(n1232), .Z(n1087) );
  NAND U1271 ( .A(n620), .B(n799), .Z(n1232) );
  IV U1272 ( .A(n1231), .Z(n1245) );
  XNOR U1273 ( .A(n1228), .B(n1246), .Z(n1231) );
  AND U1274 ( .A(n870), .B(n555), .Z(n1246) );
  XOR U1275 ( .A(n1247), .B(n1248), .Z(n1228) );
  ANDN U1276 ( .A(n1249), .B(n1250), .Z(n1248) );
  XNOR U1277 ( .A(n1251), .B(n1247), .Z(n1249) );
  XNOR U1278 ( .A(n1252), .B(n1253), .Z(n1089) );
  IV U1279 ( .A(n1241), .Z(n1253) );
  XNOR U1280 ( .A(n1238), .B(n1254), .Z(n1241) );
  AND U1281 ( .A(n438), .B(e_input[0]), .Z(n1254) );
  XOR U1282 ( .A(n1236), .B(g_input[9]), .Z(n1237) );
  NANDN U1283 ( .B(n1255), .A(n1256), .Z(n1236) );
  XOR U1284 ( .A(n1257), .B(n1258), .Z(n1238) );
  ANDN U1285 ( .A(n1259), .B(n1260), .Z(n1258) );
  XNOR U1286 ( .A(n1261), .B(n1257), .Z(n1259) );
  XOR U1287 ( .A(n1262), .B(n1242), .Z(n1252) );
  NAND U1288 ( .A(n490), .B(n1143), .Z(n1242) );
  IV U1289 ( .A(n1244), .Z(n1262) );
  NAND U1290 ( .A(n688), .B(n799), .Z(n1251) );
  XNOR U1291 ( .A(n1247), .B(n1264), .Z(n1250) );
  AND U1292 ( .A(n870), .B(n620), .Z(n1264) );
  XNOR U1293 ( .A(n1268), .B(n1265), .Z(n1267) );
  XNOR U1294 ( .A(n1257), .B(n1270), .Z(n1260) );
  AND U1295 ( .A(n490), .B(e_input[0]), .Z(n1270) );
  XNOR U1296 ( .A(n1274), .B(n1271), .Z(n1273) );
  XOR U1297 ( .A(n1275), .B(n1261), .Z(n1269) );
  NAND U1298 ( .A(n555), .B(n1143), .Z(n1261) );
  IV U1299 ( .A(n1263), .Z(n1275) );
  XNOR U1300 ( .A(n1276), .B(n1277), .Z(n1263) );
  AND U1301 ( .A(n1278), .B(n1279), .Z(n1277) );
  XOR U1302 ( .A(n1272), .B(n1280), .Z(n1279) );
  XNOR U1303 ( .A(n1274), .B(n1276), .Z(n1280) );
  NAND U1304 ( .A(n620), .B(n1143), .Z(n1274) );
  XOR U1305 ( .A(n1271), .B(n1281), .Z(n1272) );
  AND U1306 ( .A(n555), .B(e_input[0]), .Z(n1281) );
  XNOR U1307 ( .A(n1285), .B(n1282), .Z(n1284) );
  XOR U1308 ( .A(n1266), .B(n1286), .Z(n1278) );
  XNOR U1309 ( .A(n1268), .B(n1276), .Z(n1286) );
  NANDN U1310 ( .B(n756), .A(n799), .Z(n1268) );
  XOR U1311 ( .A(n1265), .B(n1287), .Z(n1266) );
  AND U1312 ( .A(n870), .B(n688), .Z(n1287) );
  XOR U1313 ( .A(n1288), .B(n1289), .Z(n1265) );
  AND U1314 ( .A(n1290), .B(n1291), .Z(n1289) );
  XNOR U1315 ( .A(n1292), .B(n1288), .Z(n1291) );
  XOR U1316 ( .A(n1293), .B(n1294), .Z(n1276) );
  AND U1317 ( .A(n1295), .B(n1296), .Z(n1294) );
  XOR U1318 ( .A(n1283), .B(n1297), .Z(n1296) );
  XNOR U1319 ( .A(n1285), .B(n1293), .Z(n1297) );
  NAND U1320 ( .A(n688), .B(n1143), .Z(n1285) );
  XOR U1321 ( .A(n1282), .B(n1298), .Z(n1283) );
  AND U1322 ( .A(n620), .B(e_input[0]), .Z(n1298) );
  XNOR U1323 ( .A(n1302), .B(n1299), .Z(n1301) );
  XOR U1324 ( .A(n1290), .B(n1303), .Z(n1295) );
  XNOR U1325 ( .A(n1292), .B(n1293), .Z(n1303) );
  NANDN U1326 ( .B(n833), .A(n799), .Z(n1292) );
  XOR U1327 ( .A(n1288), .B(n1304), .Z(n1290) );
  ANDN U1328 ( .A(n870), .B(n756), .Z(n1304) );
  XOR U1329 ( .A(n1305), .B(n1306), .Z(n1288) );
  AND U1330 ( .A(n1307), .B(n1308), .Z(n1306) );
  XNOR U1331 ( .A(n1309), .B(n1305), .Z(n1308) );
  XOR U1332 ( .A(n1310), .B(n1311), .Z(n1293) );
  AND U1333 ( .A(n1312), .B(n1313), .Z(n1311) );
  XOR U1334 ( .A(n1300), .B(n1314), .Z(n1313) );
  XNOR U1335 ( .A(n1302), .B(n1310), .Z(n1314) );
  NANDN U1336 ( .B(n756), .A(n1143), .Z(n1302) );
  XOR U1337 ( .A(n1299), .B(n1315), .Z(n1300) );
  AND U1338 ( .A(n688), .B(e_input[0]), .Z(n1315) );
  XOR U1339 ( .A(n1307), .B(n1319), .Z(n1312) );
  XNOR U1340 ( .A(n1309), .B(n1310), .Z(n1319) );
  NAND U1341 ( .A(n799), .B(n906), .Z(n1309) );
  XOR U1342 ( .A(n1305), .B(n1320), .Z(n1307) );
  ANDN U1343 ( .A(n870), .B(n833), .Z(n1320) );
  NAND U1344 ( .A(n799), .B(n1126), .Z(n1323) );
  XNOR U1345 ( .A(n1321), .B(n1325), .Z(n1322) );
  AND U1346 ( .A(n906), .B(n870), .Z(n1325) );
  AND U1347 ( .A(n1326), .B(g_input[0]), .Z(n1321) );
  NANDN U1348 ( .B(n799), .A(n1327), .Z(n1326) );
  NAND U1349 ( .A(n1126), .B(n870), .Z(n1327) );
  XNOR U1350 ( .A(n1316), .B(n1331), .Z(n1317) );
  ANDN U1351 ( .A(e_input[0]), .B(n756), .Z(n1331) );
  XOR U1352 ( .A(n1334), .B(n1332), .Z(n1333) );
  ANDN U1353 ( .A(e_input[0]), .B(n833), .Z(n1334) );
  AND U1354 ( .A(n1143), .B(n906), .Z(n1335) );
  XOR U1355 ( .A(n1339), .B(n1318), .Z(n1330) );
  NANDN U1356 ( .B(n833), .A(n1143), .Z(n1318) );
  IV U1357 ( .A(n1324), .Z(n1339) );
  NAND U1358 ( .A(n1143), .B(n1126), .Z(n1338) );
  XNOR U1359 ( .A(n1336), .B(n1340), .Z(n1337) );
  AND U1360 ( .A(n906), .B(e_input[0]), .Z(n1340) );
  AND U1361 ( .A(n1341), .B(g_input[0]), .Z(n1336) );
  NANDN U1362 ( .B(n1143), .A(n1342), .Z(n1341) );
  NAND U1363 ( .A(n1126), .B(e_input[0]), .Z(n1342) );
  XNOR U1364 ( .A(n1344), .B(n896), .Z(n886) );
  XNOR U1365 ( .A(n883), .B(n884), .Z(n896) );
  NAND U1366 ( .A(n327), .B(n688), .Z(n884) );
  XNOR U1367 ( .A(n882), .B(n1345), .Z(n883) );
  AND U1368 ( .A(n620), .B(n368), .Z(n1345) );
  XNOR U1369 ( .A(n1349), .B(n1346), .Z(n1348) );
  XNOR U1370 ( .A(n895), .B(n885), .Z(n1344) );
  XOR U1371 ( .A(n1350), .B(n1351), .Z(n885) );
  XNOR U1372 ( .A(n890), .B(n1353), .Z(n891) );
  AND U1373 ( .A(n490), .B(n475), .Z(n1353) );
  XNOR U1374 ( .A(n1256), .B(g_input[8]), .Z(n1255) );
  NOR U1375 ( .A(n1354), .B(n1355), .Z(n1256) );
  XOR U1376 ( .A(n1356), .B(n1357), .Z(n890) );
  AND U1377 ( .A(n1358), .B(n1359), .Z(n1357) );
  XNOR U1378 ( .A(n1360), .B(n1356), .Z(n1359) );
  XOR U1379 ( .A(n1361), .B(n892), .Z(n1352) );
  NAND U1380 ( .A(n421), .B(n555), .Z(n892) );
  IV U1381 ( .A(n894), .Z(n1361) );
  XNOR U1382 ( .A(n1362), .B(n1363), .Z(n894) );
  AND U1383 ( .A(n1364), .B(n1365), .Z(n1363) );
  XOR U1384 ( .A(n1358), .B(n1366), .Z(n1365) );
  XNOR U1385 ( .A(n1360), .B(n1362), .Z(n1366) );
  NAND U1386 ( .A(n421), .B(n620), .Z(n1360) );
  XOR U1387 ( .A(n1356), .B(n1367), .Z(n1358) );
  AND U1388 ( .A(n555), .B(n475), .Z(n1367) );
  XOR U1389 ( .A(n1354), .B(g_input[7]), .Z(n1355) );
  NANDN U1390 ( .B(n1368), .A(n1369), .Z(n1354) );
  XOR U1391 ( .A(n1370), .B(n1371), .Z(n1356) );
  AND U1392 ( .A(n1372), .B(n1373), .Z(n1371) );
  XNOR U1393 ( .A(n1374), .B(n1370), .Z(n1373) );
  XOR U1394 ( .A(n1347), .B(n1375), .Z(n1364) );
  XNOR U1395 ( .A(n1349), .B(n1362), .Z(n1375) );
  NANDN U1396 ( .B(n756), .A(n327), .Z(n1349) );
  XOR U1397 ( .A(n1346), .B(n1376), .Z(n1347) );
  AND U1398 ( .A(n688), .B(n368), .Z(n1376) );
  XNOR U1399 ( .A(n1380), .B(n1377), .Z(n1379) );
  XOR U1400 ( .A(n1381), .B(n1382), .Z(n1362) );
  AND U1401 ( .A(n1383), .B(n1384), .Z(n1382) );
  XOR U1402 ( .A(n1372), .B(n1385), .Z(n1384) );
  XNOR U1403 ( .A(n1374), .B(n1381), .Z(n1385) );
  NAND U1404 ( .A(n421), .B(n688), .Z(n1374) );
  XOR U1405 ( .A(n1370), .B(n1386), .Z(n1372) );
  AND U1406 ( .A(n620), .B(n475), .Z(n1386) );
  XNOR U1407 ( .A(n1369), .B(g_input[6]), .Z(n1368) );
  NOR U1408 ( .A(n1387), .B(n1388), .Z(n1369) );
  XOR U1409 ( .A(n1389), .B(n1390), .Z(n1370) );
  AND U1410 ( .A(n1391), .B(n1392), .Z(n1390) );
  XNOR U1411 ( .A(n1393), .B(n1389), .Z(n1392) );
  XOR U1412 ( .A(n1378), .B(n1394), .Z(n1383) );
  XNOR U1413 ( .A(n1380), .B(n1381), .Z(n1394) );
  NANDN U1414 ( .B(n833), .A(n327), .Z(n1380) );
  XOR U1415 ( .A(n1377), .B(n1395), .Z(n1378) );
  ANDN U1416 ( .A(n368), .B(n756), .Z(n1395) );
  XNOR U1417 ( .A(n1399), .B(n1396), .Z(n1398) );
  XOR U1418 ( .A(n1400), .B(n1401), .Z(n1381) );
  AND U1419 ( .A(n1402), .B(n1403), .Z(n1401) );
  XOR U1420 ( .A(n1391), .B(n1404), .Z(n1403) );
  XNOR U1421 ( .A(n1393), .B(n1400), .Z(n1404) );
  NANDN U1422 ( .B(n756), .A(n421), .Z(n1393) );
  XOR U1423 ( .A(n1389), .B(n1405), .Z(n1391) );
  AND U1424 ( .A(n688), .B(n475), .Z(n1405) );
  XOR U1425 ( .A(n1387), .B(g_input[5]), .Z(n1388) );
  NANDN U1426 ( .B(n1406), .A(n1407), .Z(n1387) );
  XOR U1427 ( .A(n1408), .B(n1409), .Z(n1389) );
  ANDN U1428 ( .A(n1410), .B(n1411), .Z(n1409) );
  XNOR U1429 ( .A(n1412), .B(n1408), .Z(n1410) );
  XOR U1430 ( .A(n1397), .B(n1413), .Z(n1402) );
  XNOR U1431 ( .A(n1399), .B(n1400), .Z(n1413) );
  NAND U1432 ( .A(n327), .B(n906), .Z(n1399) );
  XOR U1433 ( .A(n1396), .B(n1414), .Z(n1397) );
  ANDN U1434 ( .A(n368), .B(n833), .Z(n1414) );
  XOR U1435 ( .A(n1415), .B(n1416), .Z(n1396) );
  ANDN U1436 ( .A(n1417), .B(n1418), .Z(n1416) );
  XNOR U1437 ( .A(n1419), .B(n1415), .Z(n1417) );
  NAND U1438 ( .A(n327), .B(n1126), .Z(n1419) );
  XNOR U1439 ( .A(n1415), .B(n1421), .Z(n1418) );
  AND U1440 ( .A(n906), .B(n368), .Z(n1421) );
  AND U1441 ( .A(n1422), .B(g_input[0]), .Z(n1415) );
  NANDN U1442 ( .B(n327), .A(n1423), .Z(n1422) );
  NAND U1443 ( .A(n1126), .B(n368), .Z(n1423) );
  XNOR U1444 ( .A(n1408), .B(n1427), .Z(n1411) );
  ANDN U1445 ( .A(n475), .B(n756), .Z(n1427) );
  XOR U1446 ( .A(n1428), .B(n1429), .Z(n1408) );
  AND U1447 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U1448 ( .A(n1432), .B(n1428), .Z(n1431) );
  ANDN U1449 ( .A(n475), .B(n833), .Z(n1432) );
  XOR U1450 ( .A(n1433), .B(n1428), .Z(n1430) );
  AND U1451 ( .A(n906), .B(n421), .Z(n1433) );
  XOR U1452 ( .A(n1434), .B(n1435), .Z(n1428) );
  ANDN U1453 ( .A(n1436), .B(n1437), .Z(n1435) );
  XNOR U1454 ( .A(n1438), .B(n1434), .Z(n1436) );
  XOR U1455 ( .A(n1439), .B(n1412), .Z(n1426) );
  NANDN U1456 ( .B(n833), .A(n421), .Z(n1412) );
  IV U1457 ( .A(n1420), .Z(n1439) );
  XOR U1458 ( .A(n1440), .B(n1438), .Z(n1420) );
  NAND U1459 ( .A(n421), .B(n1126), .Z(n1438) );
  IV U1460 ( .A(n1437), .Z(n1440) );
  XNOR U1461 ( .A(n1434), .B(n1441), .Z(n1437) );
  AND U1462 ( .A(n906), .B(n475), .Z(n1441) );
  AND U1463 ( .A(n1442), .B(g_input[0]), .Z(n1434) );
  NANDN U1464 ( .B(n421), .A(n1443), .Z(n1442) );
  NAND U1465 ( .A(n1126), .B(n475), .Z(n1443) );
  XNOR U1466 ( .A(n899), .B(n1447), .Z(n900) );
  ANDN U1467 ( .A(n295), .B(n756), .Z(n1447) );
  XNOR U1468 ( .A(n1407), .B(g_input[4]), .Z(n1406) );
  NOR U1469 ( .A(n1448), .B(n1449), .Z(n1407) );
  XOR U1470 ( .A(n1450), .B(n1451), .Z(n899) );
  AND U1471 ( .A(n1452), .B(n1453), .Z(n1451) );
  XOR U1472 ( .A(n1454), .B(n1450), .Z(n1453) );
  ANDN U1473 ( .A(n295), .B(n833), .Z(n1454) );
  XOR U1474 ( .A(n1455), .B(n1450), .Z(n1452) );
  AND U1475 ( .A(n906), .B(n257), .Z(n1455) );
  XOR U1476 ( .A(n1456), .B(n1457), .Z(n1450) );
  ANDN U1477 ( .A(n1458), .B(n1459), .Z(n1457) );
  XNOR U1478 ( .A(n1460), .B(n1456), .Z(n1458) );
  XOR U1479 ( .A(n1461), .B(n901), .Z(n1446) );
  NANDN U1480 ( .B(n833), .A(n257), .Z(n901) );
  NANDN U1481 ( .B(n1462), .A(n1463), .Z(n1448) );
  IV U1482 ( .A(n903), .Z(n1461) );
  NAND U1483 ( .A(n257), .B(n1126), .Z(n1460) );
  XNOR U1484 ( .A(n1456), .B(n1464), .Z(n1459) );
  AND U1485 ( .A(n906), .B(n295), .Z(n1464) );
  AND U1486 ( .A(n1465), .B(g_input[0]), .Z(n1456) );
  NANDN U1487 ( .B(n257), .A(n1466), .Z(n1465) );
  NAND U1488 ( .A(n1126), .B(n295), .Z(n1466) );
  XNOR U1489 ( .A(n1467), .B(e_input[12]), .Z(n295) );
  NAND U1490 ( .A(n1468), .B(e_input[15]), .Z(n1467) );
  XOR U1491 ( .A(n1469), .B(e_input[12]), .Z(n1468) );
  XNOR U1492 ( .A(n910), .B(n911), .Z(n905) );
  NANDN U1493 ( .B(n202), .A(n1126), .Z(n911) );
  XNOR U1494 ( .A(n909), .B(n1471), .Z(n910) );
  AND U1495 ( .A(n906), .B(n226), .Z(n1471) );
  XNOR U1496 ( .A(n1463), .B(g_input[2]), .Z(n1462) );
  AND U1497 ( .A(n1473), .B(g_input[0]), .Z(n909) );
  NAND U1498 ( .A(n1474), .B(n202), .Z(n1473) );
  NANDN U1499 ( .B(n1475), .A(n1476), .Z(n202) );
  ANDN U1500 ( .A(e_input[15]), .B(n1477), .Z(n1476) );
  NAND U1501 ( .A(n1126), .B(n226), .Z(n1474) );
  XOR U1502 ( .A(n1477), .B(e_input[14]), .Z(n1475) );
  OR U1503 ( .A(n1470), .B(n1478), .Z(n1477) );
  XOR U1504 ( .A(n1478), .B(e_input[13]), .Z(n1470) );
  OR U1505 ( .A(n1469), .B(n1479), .Z(n1478) );
  XOR U1506 ( .A(n1479), .B(e_input[12]), .Z(n1469) );
  OR U1507 ( .A(n1425), .B(n1480), .Z(n1479) );
  XOR U1508 ( .A(n1480), .B(e_input[11]), .Z(n1425) );
  OR U1509 ( .A(n1424), .B(n1481), .Z(n1480) );
  XOR U1510 ( .A(n1481), .B(e_input[10]), .Z(n1424) );
  OR U1511 ( .A(n1445), .B(n1482), .Z(n1481) );
  XOR U1512 ( .A(n1482), .B(e_input[9]), .Z(n1445) );
  OR U1513 ( .A(n1444), .B(n1483), .Z(n1482) );
  XOR U1514 ( .A(n1483), .B(e_input[8]), .Z(n1444) );
  OR U1515 ( .A(n1136), .B(n1484), .Z(n1483) );
  XOR U1516 ( .A(n1484), .B(e_input[7]), .Z(n1136) );
  OR U1517 ( .A(n1135), .B(n1485), .Z(n1484) );
  XOR U1518 ( .A(n1485), .B(e_input[6]), .Z(n1135) );
  OR U1519 ( .A(n1131), .B(n1486), .Z(n1485) );
  XOR U1520 ( .A(n1486), .B(e_input[5]), .Z(n1131) );
  OR U1521 ( .A(n1130), .B(n1487), .Z(n1486) );
  XOR U1522 ( .A(n1487), .B(e_input[4]), .Z(n1130) );
  OR U1523 ( .A(n1329), .B(n1488), .Z(n1487) );
  XOR U1524 ( .A(n1488), .B(e_input[3]), .Z(n1329) );
  OR U1525 ( .A(n1328), .B(n1489), .Z(n1488) );
  XOR U1526 ( .A(n1489), .B(e_input[2]), .Z(n1328) );
  NANDN U1527 ( .B(e_input[0]), .A(n1343), .Z(n1489) );
  XNOR U1528 ( .A(e_input[0]), .B(e_input[1]), .Z(n1343) );
  XOR U1529 ( .A(g_input[0]), .B(g_input[1]), .Z(n1472) );
  NANDN U1530 ( .B(n845), .A(n117), .Z(n169) );
  IV U1531 ( .A(rst), .Z(n117) );
  NAND U1532 ( .A(n1490), .B(n1491), .Z(n845) );
  AND U1533 ( .A(n1492), .B(n1493), .Z(n1491) );
  ANDN U1534 ( .A(n1494), .B(\_MxM/n[3] ), .Z(n1493) );
  NOR U1535 ( .A(\_MxM/n[8] ), .B(\_MxM/n[9] ), .Z(n1494) );
  ANDN U1536 ( .A(n1495), .B(\_MxM/n[13] ), .Z(n1492) );
  NOR U1537 ( .A(\_MxM/n[1] ), .B(\_MxM/n[2] ), .Z(n1495) );
  AND U1538 ( .A(n1496), .B(n1497), .Z(n1490) );
  ANDN U1539 ( .A(n1498), .B(n108), .Z(n1497) );
  OR U1540 ( .A(\_MxM/n[6] ), .B(\_MxM/n[7] ), .Z(n108) );
  NOR U1541 ( .A(\_MxM/n[0] ), .B(\_MxM/n[10] ), .Z(n1498) );
  NOR U1542 ( .A(n106), .B(n107), .Z(n1496) );
  OR U1543 ( .A(\_MxM/n[4] ), .B(\_MxM/n[5] ), .Z(n107) );
  OR U1544 ( .A(\_MxM/n[12] ), .B(\_MxM/n[11] ), .Z(n106) );
endmodule

