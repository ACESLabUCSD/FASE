
module MxM_TG_W32_N100 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \_MxM/n171 , \_MxM/n168 , \_MxM/n165 , \_MxM/n162 , \_MxM/n159 ,
         \_MxM/n156 , \_MxM/n153 , \_MxM/n150 , \_MxM/n147 , \_MxM/n144 ,
         \_MxM/n141 , \_MxM/n138 , \_MxM/n135 , \_MxM/n132 , \_MxM/n129 ,
         \_MxM/n126 , \_MxM/n123 , \_MxM/n120 , \_MxM/n117 , \_MxM/n114 ,
         \_MxM/n111 , \_MxM/n108 , \_MxM/n105 , \_MxM/n102 , \_MxM/n99 ,
         \_MxM/n96 , \_MxM/n93 , \_MxM/n90 , \_MxM/n87 , \_MxM/n84 ,
         \_MxM/n81 , \_MxM/n78 , \_MxM/N17 , \_MxM/N16 , \_MxM/N15 ,
         \_MxM/N14 , \_MxM/N13 , \_MxM/N12 , \_MxM/N11 , \_MxM/N9 , \_MxM/N8 ,
         \_MxM/N7 , \_MxM/N6 , \_MxM/N5 , \_MxM/n[0] , \_MxM/n[1] ,
         \_MxM/n[2] , \_MxM/n[3] , \_MxM/n[4] , \_MxM/n[5] , \_MxM/n[6] ,
         \_MxM/Y1[0] , \_MxM/Y1[1] , \_MxM/Y1[2] , \_MxM/Y1[3] , \_MxM/Y1[4] ,
         \_MxM/Y1[5] , \_MxM/Y1[6] , \_MxM/Y1[7] , \_MxM/Y1[8] , \_MxM/Y1[9] ,
         \_MxM/Y1[10] , \_MxM/Y1[11] , \_MxM/Y1[12] , \_MxM/Y1[13] ,
         \_MxM/Y1[14] , \_MxM/Y1[15] , \_MxM/Y1[16] , \_MxM/Y1[17] ,
         \_MxM/Y1[18] , \_MxM/Y1[19] , \_MxM/Y1[20] , \_MxM/Y1[21] ,
         \_MxM/Y1[22] , \_MxM/Y1[23] , \_MxM/Y1[24] , \_MxM/Y1[25] ,
         \_MxM/Y1[26] , \_MxM/Y1[27] , \_MxM/Y1[28] , \_MxM/Y1[29] ,
         \_MxM/Y1[30] , \_MxM/Y1[31] , \_MxM/Y0[31] , \_MxM/Y0[30] ,
         \_MxM/Y0[29] , \_MxM/Y0[28] , \_MxM/Y0[27] , \_MxM/Y0[26] ,
         \_MxM/Y0[25] , \_MxM/Y0[24] , \_MxM/Y0[23] , \_MxM/Y0[22] ,
         \_MxM/Y0[21] , \_MxM/Y0[20] , \_MxM/Y0[19] , \_MxM/Y0[18] ,
         \_MxM/Y0[17] , \_MxM/Y0[16] , \_MxM/Y0[15] , \_MxM/Y0[14] ,
         \_MxM/Y0[13] , \_MxM/Y0[12] , \_MxM/Y0[11] , \_MxM/Y0[10] ,
         \_MxM/Y0[9] , \_MxM/Y0[8] , \_MxM/Y0[7] , \_MxM/Y0[6] , \_MxM/Y0[5] ,
         \_MxM/Y0[4] , \_MxM/Y0[3] , \_MxM/Y0[2] , \_MxM/Y0[1] , \_MxM/Y0[0] ,
         \_MxM/add_43/carry[6] , \_MxM/add_43/carry[5] ,
         \_MxM/add_43/carry[4] , \_MxM/add_43/carry[3] ,
         \_MxM/add_43/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216;

  DFF \_MxM/Y_reg[31]  ( .D(\_MxM/n78 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[31]) );
  DFF \_MxM/Y0_reg[31]  ( .D(\_MxM/Y1[31] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[31] ) );
  DFF \_MxM/Y_reg[30]  ( .D(\_MxM/n81 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[30]) );
  DFF \_MxM/Y0_reg[30]  ( .D(\_MxM/Y1[30] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[30] ) );
  DFF \_MxM/Y_reg[29]  ( .D(\_MxM/n84 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[29]) );
  DFF \_MxM/Y0_reg[29]  ( .D(\_MxM/Y1[29] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[29] ) );
  DFF \_MxM/Y_reg[28]  ( .D(\_MxM/n87 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[28]) );
  DFF \_MxM/Y0_reg[28]  ( .D(\_MxM/Y1[28] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[28] ) );
  DFF \_MxM/Y_reg[27]  ( .D(\_MxM/n90 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[27]) );
  DFF \_MxM/Y0_reg[27]  ( .D(\_MxM/Y1[27] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[27] ) );
  DFF \_MxM/Y_reg[26]  ( .D(\_MxM/n93 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[26]) );
  DFF \_MxM/Y0_reg[26]  ( .D(\_MxM/Y1[26] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[26] ) );
  DFF \_MxM/Y_reg[25]  ( .D(\_MxM/n96 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[25]) );
  DFF \_MxM/Y0_reg[25]  ( .D(\_MxM/Y1[25] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[25] ) );
  DFF \_MxM/Y_reg[24]  ( .D(\_MxM/n99 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[24]) );
  DFF \_MxM/Y0_reg[24]  ( .D(\_MxM/Y1[24] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[24] ) );
  DFF \_MxM/Y_reg[23]  ( .D(\_MxM/n102 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[23]) );
  DFF \_MxM/Y0_reg[23]  ( .D(\_MxM/Y1[23] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[23] ) );
  DFF \_MxM/Y_reg[22]  ( .D(\_MxM/n105 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[22]) );
  DFF \_MxM/Y0_reg[22]  ( .D(\_MxM/Y1[22] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[22] ) );
  DFF \_MxM/Y_reg[21]  ( .D(\_MxM/n108 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[21]) );
  DFF \_MxM/Y0_reg[21]  ( .D(\_MxM/Y1[21] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[21] ) );
  DFF \_MxM/Y_reg[20]  ( .D(\_MxM/n111 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[20]) );
  DFF \_MxM/Y0_reg[20]  ( .D(\_MxM/Y1[20] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[20] ) );
  DFF \_MxM/Y_reg[19]  ( .D(\_MxM/n114 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[19]) );
  DFF \_MxM/Y0_reg[19]  ( .D(\_MxM/Y1[19] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[19] ) );
  DFF \_MxM/Y_reg[18]  ( .D(\_MxM/n117 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[18]) );
  DFF \_MxM/Y0_reg[18]  ( .D(\_MxM/Y1[18] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[18] ) );
  DFF \_MxM/Y_reg[17]  ( .D(\_MxM/n120 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[17]) );
  DFF \_MxM/Y0_reg[17]  ( .D(\_MxM/Y1[17] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[17] ) );
  DFF \_MxM/Y_reg[16]  ( .D(\_MxM/n123 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[16]) );
  DFF \_MxM/Y0_reg[16]  ( .D(\_MxM/Y1[16] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[16] ) );
  DFF \_MxM/Y_reg[15]  ( .D(\_MxM/n126 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[15]) );
  DFF \_MxM/Y0_reg[15]  ( .D(\_MxM/Y1[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[15] ) );
  DFF \_MxM/Y_reg[14]  ( .D(\_MxM/n129 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[14]) );
  DFF \_MxM/Y0_reg[14]  ( .D(\_MxM/Y1[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[14] ) );
  DFF \_MxM/Y_reg[13]  ( .D(\_MxM/n132 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[13]) );
  DFF \_MxM/Y0_reg[13]  ( .D(\_MxM/Y1[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[13] ) );
  DFF \_MxM/Y_reg[12]  ( .D(\_MxM/n135 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[12]) );
  DFF \_MxM/Y0_reg[12]  ( .D(\_MxM/Y1[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[12] ) );
  DFF \_MxM/Y_reg[11]  ( .D(\_MxM/n138 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[11]) );
  DFF \_MxM/Y0_reg[11]  ( .D(\_MxM/Y1[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[11] ) );
  DFF \_MxM/Y_reg[10]  ( .D(\_MxM/n141 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[10]) );
  DFF \_MxM/Y0_reg[10]  ( .D(\_MxM/Y1[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\_MxM/Y0[10] ) );
  DFF \_MxM/Y_reg[9]  ( .D(\_MxM/n144 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[9]) );
  DFF \_MxM/Y0_reg[9]  ( .D(\_MxM/Y1[9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[9] ) );
  DFF \_MxM/Y_reg[8]  ( .D(\_MxM/n147 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[8]) );
  DFF \_MxM/Y0_reg[8]  ( .D(\_MxM/Y1[8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[8] ) );
  DFF \_MxM/Y_reg[7]  ( .D(\_MxM/n150 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[7]) );
  DFF \_MxM/Y0_reg[7]  ( .D(\_MxM/Y1[7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[7] ) );
  DFF \_MxM/Y_reg[6]  ( .D(\_MxM/n153 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[6]) );
  DFF \_MxM/Y0_reg[6]  ( .D(\_MxM/Y1[6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[6] ) );
  DFF \_MxM/Y_reg[5]  ( .D(\_MxM/n156 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[5]) );
  DFF \_MxM/Y0_reg[5]  ( .D(\_MxM/Y1[5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[5] ) );
  DFF \_MxM/Y_reg[4]  ( .D(\_MxM/n159 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[4]) );
  DFF \_MxM/Y0_reg[4]  ( .D(\_MxM/Y1[4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[4] ) );
  DFF \_MxM/Y_reg[3]  ( .D(\_MxM/n162 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[3]) );
  DFF \_MxM/Y0_reg[3]  ( .D(\_MxM/Y1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[3] ) );
  DFF \_MxM/Y_reg[2]  ( .D(\_MxM/n165 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[2]) );
  DFF \_MxM/Y0_reg[2]  ( .D(\_MxM/Y1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[2] ) );
  DFF \_MxM/Y_reg[1]  ( .D(\_MxM/n168 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[1]) );
  DFF \_MxM/Y0_reg[1]  ( .D(\_MxM/Y1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[1] ) );
  DFF \_MxM/Y_reg[0]  ( .D(\_MxM/n171 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o[0]) );
  DFF \_MxM/Y0_reg[0]  ( .D(\_MxM/Y1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/Y0[0] ) );
  DFF \_MxM/n_reg[6]  ( .D(\_MxM/N17 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[6] ) );
  DFF \_MxM/n_reg[5]  ( .D(\_MxM/N16 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[5] ) );
  DFF \_MxM/n_reg[4]  ( .D(\_MxM/N15 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[4] ) );
  DFF \_MxM/n_reg[3]  ( .D(\_MxM/N14 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[3] ) );
  DFF \_MxM/n_reg[2]  ( .D(\_MxM/N13 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[2] ) );
  DFF \_MxM/n_reg[1]  ( .D(\_MxM/N12 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[1] ) );
  DFF \_MxM/n_reg[0]  ( .D(\_MxM/N11 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \_MxM/n[0] ) );
  HADDER \_MxM/add_43/U1_1_1  ( .IN0(\_MxM/n[1] ), .IN1(\_MxM/n[0] ), .COUT(
        \_MxM/add_43/carry[2] ), .SUM(\_MxM/N5 ) );
  HADDER \_MxM/add_43/U1_1_2  ( .IN0(\_MxM/n[2] ), .IN1(\_MxM/add_43/carry[2] ), .COUT(\_MxM/add_43/carry[3] ), .SUM(\_MxM/N6 ) );
  HADDER \_MxM/add_43/U1_1_3  ( .IN0(\_MxM/n[3] ), .IN1(\_MxM/add_43/carry[3] ), .COUT(\_MxM/add_43/carry[4] ), .SUM(\_MxM/N7 ) );
  HADDER \_MxM/add_43/U1_1_4  ( .IN0(\_MxM/n[4] ), .IN1(\_MxM/add_43/carry[4] ), .COUT(\_MxM/add_43/carry[5] ), .SUM(\_MxM/N8 ) );
  HADDER \_MxM/add_43/U1_1_5  ( .IN0(\_MxM/n[5] ), .IN1(\_MxM/add_43/carry[5] ), .COUT(\_MxM/add_43/carry[6] ), .SUM(\_MxM/N9 ) );
  MUX U1 ( .IN0(n3740), .IN1(n3738), .SEL(n3739), .F(n3700) );
  XOR U2 ( .A(n4517), .B(n4507), .Z(n4117) );
  XOR U3 ( .A(n4487), .B(n4488), .Z(n4099) );
  MUX U4 ( .IN0(n4092), .IN1(n4090), .SEL(n4091), .F(n4073) );
  MUX U5 ( .IN0(n4861), .IN1(n4859), .SEL(n4860), .F(n4838) );
  XOR U6 ( .A(n4398), .B(n4390), .Z(n3964) );
  MUX U7 ( .IN0(n1), .IN1(n2817), .SEL(n2818), .F(n2685) );
  IV U8 ( .A(n2819), .Z(n1) );
  MUX U9 ( .IN0(n2), .IN1(n1376), .SEL(n1377), .F(n1305) );
  IV U10 ( .A(n1378), .Z(n2) );
  MUX U11 ( .IN0(n2733), .IN1(n2731), .SEL(n2732), .F(n2604) );
  MUX U12 ( .IN0(n2401), .IN1(n2399), .SEL(n2400), .F(n2284) );
  MUX U13 ( .IN0(n2432), .IN1(n2430), .SEL(n2431), .F(n2309) );
  MUX U14 ( .IN0(n2029), .IN1(n2027), .SEL(n2028), .F(n1922) );
  MUX U15 ( .IN0(n1637), .IN1(n1635), .SEL(n1636), .F(n1543) );
  MUX U16 ( .IN0(n1494), .IN1(n1492), .SEL(n1493), .F(n1407) );
  MUX U17 ( .IN0(n1351), .IN1(n3), .SEL(n1350), .F(n1282) );
  IV U18 ( .A(n1349), .Z(n3) );
  MUX U19 ( .IN0(n1139), .IN1(n1137), .SEL(n1138), .F(n1073) );
  MUX U20 ( .IN0(n853), .IN1(n851), .SEL(n852), .F(n811) );
  XOR U21 ( .A(n103), .B(n1425), .Z(n1355) );
  MUX U22 ( .IN0(n4), .IN1(n977), .SEL(n978), .F(n921) );
  IV U23 ( .A(n979), .Z(n4) );
  MUX U24 ( .IN0(n2546), .IN1(n2544), .SEL(n2545), .F(n2420) );
  MUX U25 ( .IN0(n5), .IN1(n1083), .SEL(n1084), .F(n1024) );
  IV U26 ( .A(n1085), .Z(n5) );
  MUX U27 ( .IN0(n6), .IN1(n1021), .SEL(n1022), .F(n966) );
  IV U28 ( .A(n1023), .Z(n6) );
  XNOR U29 ( .A(n708), .B(n707), .Z(n705) );
  MUX U30 ( .IN0(n2070), .IN1(n7), .SEL(n2071), .F(n1965) );
  IV U31 ( .A(n2072), .Z(n7) );
  OR U32 ( .A(n790), .B(n791), .Z(n757) );
  XNOR U33 ( .A(n732), .B(n729), .Z(n728) );
  MUX U34 ( .IN0(n8), .IN1(n3734), .SEL(n3735), .F(n3696) );
  IV U35 ( .A(n3736), .Z(n8) );
  MUX U36 ( .IN0(n9), .IN1(n4128), .SEL(n4129), .F(n4111) );
  IV U37 ( .A(n4130), .Z(n9) );
  MUX U38 ( .IN0(n10), .IN1(n4120), .SEL(n4121), .F(n4103) );
  IV U39 ( .A(n4122), .Z(n10) );
  MUX U40 ( .IN0(n3759), .IN1(n3761), .SEL(n3760), .F(n3721) );
  XOR U41 ( .A(n4502), .B(n4494), .Z(n4100) );
  MUX U42 ( .IN0(n3664), .IN1(n3662), .SEL(n3663), .F(n3624) );
  XNOR U43 ( .A(n4084), .B(n4070), .Z(n4074) );
  XOR U44 ( .A(n4450), .B(n4442), .Z(n4032) );
  MUX U45 ( .IN0(n3512), .IN1(n3510), .SEL(n3511), .F(n3472) );
  MUX U46 ( .IN0(n11), .IN1(n4600), .SEL(n4601), .F(n4589) );
  IV U47 ( .A(n4602), .Z(n11) );
  MUX U48 ( .IN0(n4987), .IN1(n12), .SEL(n4865), .F(n4974) );
  IV U49 ( .A(n4864), .Z(n12) );
  MUX U50 ( .IN0(n4271), .IN1(n13), .SEL(n4272), .F(n4250) );
  IV U51 ( .A(n4273), .Z(n13) );
  MUX U52 ( .IN0(n4817), .IN1(n14), .SEL(n4818), .F(n4796) );
  IV U53 ( .A(n4819), .Z(n14) );
  MUX U54 ( .IN0(n4582), .IN1(n15), .SEL(n4238), .F(n4571) );
  IV U55 ( .A(n4236), .Z(n15) );
  MUX U56 ( .IN0(n16), .IN1(n4204), .SEL(n4205), .F(n4183) );
  IV U57 ( .A(n4206), .Z(n16) );
  MUX U58 ( .IN0(n4393), .IN1(n17), .SEL(n3964), .F(n4380) );
  IV U59 ( .A(n3963), .Z(n17) );
  MUX U60 ( .IN0(n3284), .IN1(n3282), .SEL(n3283), .F(n3244) );
  MUX U61 ( .IN0(n3905), .IN1(n3903), .SEL(n3904), .F(n3883) );
  XOR U62 ( .A(n4346), .B(n4335), .Z(n3896) );
  XOR U63 ( .A(n4901), .B(n4893), .Z(n4721) );
  MUX U64 ( .IN0(n18), .IN1(n3053), .SEL(n3054), .F(n2917) );
  IV U65 ( .A(n3055), .Z(n18) );
  MUX U66 ( .IN0(n19), .IN1(n2329), .SEL(n2330), .F(n2213) );
  IV U67 ( .A(n2331), .Z(n19) );
  MUX U68 ( .IN0(n20), .IN1(n2239), .SEL(n2240), .F(n2128) );
  IV U69 ( .A(n2241), .Z(n20) );
  MUX U70 ( .IN0(n21), .IN1(n2086), .SEL(n2087), .F(n1981) );
  IV U71 ( .A(n2088), .Z(n21) );
  MUX U72 ( .IN0(n22), .IN1(n2078), .SEL(n2079), .F(n1973) );
  IV U73 ( .A(n2080), .Z(n22) );
  MUX U74 ( .IN0(n23), .IN1(n1792), .SEL(n1793), .F(n1696) );
  IV U75 ( .A(n1794), .Z(n23) );
  MUX U76 ( .IN0(n24), .IN1(n1672), .SEL(n1673), .F(n1581) );
  IV U77 ( .A(n1674), .Z(n24) );
  MUX U78 ( .IN0(n25), .IN1(n1331), .SEL(n1332), .F(n1261) );
  IV U79 ( .A(n1333), .Z(n25) );
  MUX U80 ( .IN0(n26), .IN1(n1226), .SEL(n1227), .F(n1160) );
  IV U81 ( .A(n1228), .Z(n26) );
  MUX U82 ( .IN0(n27), .IN1(n992), .SEL(n993), .F(n934) );
  IV U83 ( .A(n994), .Z(n27) );
  MUX U84 ( .IN0(n3042), .IN1(n3040), .SEL(n3041), .F(n2904) );
  MUX U85 ( .IN0(n2953), .IN1(n2951), .SEL(n2952), .F(n2813) );
  MUX U86 ( .IN0(n2511), .IN1(n2513), .SEL(n2512), .F(n2390) );
  MUX U87 ( .IN0(n2482), .IN1(n2480), .SEL(n2481), .F(n2359) );
  MUX U88 ( .IN0(n2286), .IN1(n2284), .SEL(n2285), .F(n2172) );
  MUX U89 ( .IN0(n2311), .IN1(n2309), .SEL(n2310), .F(n2193) );
  MUX U90 ( .IN0(n1824), .IN1(n1822), .SEL(n1823), .F(n1726) );
  MUX U91 ( .IN0(n1813), .IN1(n1815), .SEL(n1814), .F(n1717) );
  MUX U92 ( .IN0(n1459), .IN1(n1457), .SEL(n1458), .F(n1380) );
  MUX U93 ( .IN0(n1175), .IN1(n1173), .SEL(n1174), .F(n1111) );
  MUX U94 ( .IN0(n1102), .IN1(n1104), .SEL(n1103), .F(n1043) );
  MUX U95 ( .IN0(n28), .IN1(n2983), .SEL(n2984), .F(n2845) );
  IV U96 ( .A(n2985), .Z(n28) );
  MUX U97 ( .IN0(n29), .IN1(n2754), .SEL(n2755), .F(n2628) );
  IV U98 ( .A(n2756), .Z(n29) );
  MUX U99 ( .IN0(n30), .IN1(n2009), .SEL(n2010), .F(n1904) );
  IV U100 ( .A(n2011), .Z(n30) );
  MUX U101 ( .IN0(n31), .IN1(n1617), .SEL(n1618), .F(n1525) );
  IV U102 ( .A(n1619), .Z(n31) );
  MUX U103 ( .IN0(n32), .IN1(n1422), .SEL(n1423), .F(n1352) );
  IV U104 ( .A(n1424), .Z(n32) );
  MUX U105 ( .IN0(n1356), .IN1(n103), .SEL(n1355), .F(n33) );
  IV U106 ( .A(n33), .Z(n1276) );
  MUX U107 ( .IN0(n813), .IN1(n811), .SEL(n812), .F(n771) );
  MUX U108 ( .IN0(n2422), .IN1(n2420), .SEL(n2421), .F(n2295) );
  MUX U109 ( .IN0(n34), .IN1(n2316), .SEL(n2317), .F(n2200) );
  IV U110 ( .A(n2318), .Z(n34) );
  MUX U111 ( .IN0(n35), .IN1(n1342), .SEL(n1343), .F(n1272) );
  IV U112 ( .A(n1344), .Z(n35) );
  MUX U113 ( .IN0(n1147), .IN1(n1149), .SEL(n1148), .F(n1086) );
  MUX U114 ( .IN0(n36), .IN1(n1024), .SEL(n1025), .F(n969) );
  IV U115 ( .A(n1026), .Z(n36) );
  NANDN U116 ( .B(n1968), .A(n1969), .Z(n1863) );
  MUX U117 ( .IN0(n37), .IN1(n1577), .SEL(n1576), .F(n1482) );
  IV U118 ( .A(n1575), .Z(n37) );
  AND U119 ( .A(n1004), .B(n1005), .Z(n946) );
  OR U120 ( .A(n704), .B(n705), .Z(n682) );
  OR U121 ( .A(n727), .B(n728), .Z(n702) );
  OR U122 ( .A(n1189), .B(n1190), .Z(n1128) );
  XNOR U123 ( .A(n871), .B(n870), .Z(n869) );
  MUX U124 ( .IN0(n4126), .IN1(n4124), .SEL(n4125), .F(n4107) );
  MUX U125 ( .IN0(n38), .IN1(n4103), .SEL(n4104), .F(n4086) );
  IV U126 ( .A(n4105), .Z(n38) );
  MUX U127 ( .IN0(n39), .IN1(n3717), .SEL(n3718), .F(n3679) );
  IV U128 ( .A(n3719), .Z(n39) );
  XNOR U129 ( .A(n3694), .B(n3659), .Z(n3663) );
  MUX U130 ( .IN0(n4497), .IN1(n40), .SEL(n4100), .F(n4484) );
  IV U131 ( .A(n4099), .Z(n40) );
  XNOR U132 ( .A(n3580), .B(n3545), .Z(n3549) );
  XOR U133 ( .A(n3601), .B(n3566), .Z(n3570) );
  MUX U134 ( .IN0(n4041), .IN1(n4039), .SEL(n4040), .F(n4022) );
  MUX U135 ( .IN0(n4445), .IN1(n41), .SEL(n4032), .F(n4432) );
  IV U136 ( .A(n4031), .Z(n41) );
  MUX U137 ( .IN0(n42), .IN1(n4976), .SEL(n4977), .F(n4963) );
  IV U138 ( .A(n4978), .Z(n42) );
  MUX U139 ( .IN0(n43), .IN1(n4983), .SEL(n4984), .F(n4970) );
  IV U140 ( .A(n4985), .Z(n43) );
  MUX U141 ( .IN0(n4615), .IN1(n44), .SEL(n4298), .F(n4604) );
  IV U142 ( .A(n4297), .Z(n44) );
  MUX U143 ( .IN0(n4294), .IN1(n4292), .SEL(n4293), .F(n4271) );
  MUX U144 ( .IN0(n45), .IN1(n4834), .SEL(n4835), .F(n4813) );
  IV U145 ( .A(n4836), .Z(n45) );
  MUX U146 ( .IN0(n3436), .IN1(n3434), .SEL(n3435), .F(n3396) );
  MUX U147 ( .IN0(n46), .IN1(n4589), .SEL(n4590), .F(n4578) );
  IV U148 ( .A(n4591), .Z(n46) );
  MUX U149 ( .IN0(n3973), .IN1(n3971), .SEL(n3972), .F(n3954) );
  MUX U150 ( .IN0(n4948), .IN1(n47), .SEL(n4805), .F(n4935) );
  IV U151 ( .A(n4803), .Z(n47) );
  XOR U152 ( .A(n3373), .B(n3338), .Z(n3342) );
  MUX U153 ( .IN0(n4571), .IN1(n48), .SEL(n4217), .F(n4560) );
  IV U154 ( .A(n4215), .Z(n48) );
  MUX U155 ( .IN0(n4208), .IN1(n49), .SEL(n4209), .F(n4187) );
  IV U156 ( .A(n4210), .Z(n49) );
  XOR U157 ( .A(n4372), .B(n4364), .Z(n3930) );
  MUX U158 ( .IN0(n50), .IN1(n3240), .SEL(n3241), .F(n3202) );
  IV U159 ( .A(n3242), .Z(n50) );
  MUX U160 ( .IN0(n4754), .IN1(n51), .SEL(n4755), .F(n4733) );
  IV U161 ( .A(n4756), .Z(n51) );
  XNOR U162 ( .A(n3914), .B(n3900), .Z(n3904) );
  XOR U163 ( .A(n4339), .B(n4340), .Z(n3895) );
  MUX U164 ( .IN0(n3227), .IN1(n3229), .SEL(n3228), .F(n3160) );
  MUX U165 ( .IN0(n52), .IN1(n3082), .SEL(n3083), .F(n2947) );
  IV U166 ( .A(n3084), .Z(n52) );
  MUX U167 ( .IN0(n53), .IN1(n3027), .SEL(n3028), .F(n2891) );
  IV U168 ( .A(n3029), .Z(n53) );
  XOR U169 ( .A(n4713), .B(n4714), .Z(n4719) );
  MUX U170 ( .IN0(n54), .IN1(n2727), .SEL(n2728), .F(n2600) );
  IV U171 ( .A(n2729), .Z(n54) );
  MUX U172 ( .IN0(n55), .IN1(n2516), .SEL(n2517), .F(n2395) );
  IV U173 ( .A(n2518), .Z(n55) );
  MUX U174 ( .IN0(n56), .IN1(n2507), .SEL(n2508), .F(n2386) );
  IV U175 ( .A(n2509), .Z(n56) );
  MUX U176 ( .IN0(n57), .IN1(n2550), .SEL(n2551), .F(n2426) );
  IV U177 ( .A(n2552), .Z(n57) );
  MUX U178 ( .IN0(n58), .IN1(n2102), .SEL(n2103), .F(n1997) );
  IV U179 ( .A(n2104), .Z(n58) );
  MUX U180 ( .IN0(n59), .IN1(n2128), .SEL(n2129), .F(n2023) );
  IV U181 ( .A(n2130), .Z(n59) );
  MUX U182 ( .IN0(n60), .IN1(n2014), .SEL(n2015), .F(n1909) );
  IV U183 ( .A(n2016), .Z(n60) );
  MUX U184 ( .IN0(n61), .IN1(n1868), .SEL(n1869), .F(n1768) );
  IV U185 ( .A(n1870), .Z(n61) );
  MUX U186 ( .IN0(n3059), .IN1(n3057), .SEL(n3058), .F(n2921) );
  XOR U187 ( .A(n476), .B(n4321), .Z(n3077) );
  MUX U188 ( .IN0(n3003), .IN1(n3001), .SEL(n3002), .F(n2863) );
  MUX U189 ( .IN0(n2906), .IN1(n2904), .SEL(n2905), .F(n2772) );
  MUX U190 ( .IN0(n2763), .IN1(n2765), .SEL(n2764), .F(n2637) );
  MUX U191 ( .IN0(n2815), .IN1(n2813), .SEL(n2814), .F(n2681) );
  MUX U192 ( .IN0(n2854), .IN1(n2856), .SEL(n2855), .F(n2722) );
  MUX U193 ( .IN0(n2269), .IN1(n2271), .SEL(n2270), .F(n62) );
  IV U194 ( .A(n62), .Z(n2163) );
  MUX U195 ( .IN0(n2245), .IN1(n2243), .SEL(n2244), .F(n2132) );
  MUX U196 ( .IN0(n2065), .IN1(n2063), .SEL(n2064), .F(n1958) );
  MUX U197 ( .IN0(n2084), .IN1(n2082), .SEL(n2083), .F(n1977) );
  MUX U198 ( .IN0(n1896), .IN1(n1898), .SEL(n1897), .F(n1796) );
  MUX U199 ( .IN0(n1717), .IN1(n1719), .SEL(n1718), .F(n1626) );
  MUX U200 ( .IN0(n1678), .IN1(n1676), .SEL(n1677), .F(n1585) );
  MUX U201 ( .IN0(n1511), .IN1(n1513), .SEL(n1512), .F(n63) );
  IV U202 ( .A(n63), .Z(n1431) );
  MUX U203 ( .IN0(n1337), .IN1(n1335), .SEL(n1336), .F(n1265) );
  MUX U204 ( .IN0(n1382), .IN1(n1380), .SEL(n1381), .F(n1309) );
  MUX U205 ( .IN0(n1300), .IN1(n1302), .SEL(n1301), .F(n1230) );
  MUX U206 ( .IN0(n1054), .IN1(n1052), .SEL(n1053), .F(n996) );
  MUX U207 ( .IN0(n987), .IN1(n989), .SEL(n988), .F(n929) );
  MUX U208 ( .IN0(n64), .IN1(n2628), .SEL(n2629), .F(n2502) );
  IV U209 ( .A(n2630), .Z(n64) );
  MUX U210 ( .IN0(n65), .IN1(n2713), .SEL(n2714), .F(n2586) );
  IV U211 ( .A(n2715), .Z(n65) );
  XNOR U212 ( .A(n1916), .B(n1819), .Z(n1823) );
  MUX U213 ( .IN0(n66), .IN1(n1525), .SEL(n1526), .F(n1439) );
  IV U214 ( .A(n1527), .Z(n66) );
  XOR U215 ( .A(n1350), .B(n1351), .Z(n1356) );
  MUX U216 ( .IN0(n1213), .IN1(n1211), .SEL(n1212), .F(n1147) );
  XNOR U217 ( .A(n1131), .B(n1076), .Z(n1074) );
  MUX U218 ( .IN0(n67), .IN1(n878), .SEL(n879), .F(n839) );
  IV U219 ( .A(n880), .Z(n67) );
  AND U220 ( .A(n798), .B(n794), .Z(n797) );
  XNOR U221 ( .A(n804), .B(n767), .Z(n772) );
  MUX U222 ( .IN0(n2297), .IN1(n2295), .SEL(n2296), .F(n2182) );
  MUX U223 ( .IN0(n68), .IN1(n2089), .SEL(n2090), .F(n1984) );
  IV U224 ( .A(n2091), .Z(n68) );
  MUX U225 ( .IN0(n69), .IN1(n1144), .SEL(n1145), .F(n1083) );
  IV U226 ( .A(n1146), .Z(n69) );
  ANDN U227 ( .A(n960), .B(n961), .Z(n959) );
  MUX U228 ( .IN0(n1860), .IN1(n70), .SEL(n1861), .F(n1760) );
  IV U229 ( .A(n1862), .Z(n70) );
  MUX U230 ( .IN0(n1482), .IN1(n1484), .SEL(n1483), .F(n1397) );
  AND U231 ( .A(n1119), .B(n1120), .Z(n1060) );
  OR U232 ( .A(n1012), .B(n1013), .Z(n954) );
  OR U233 ( .A(n828), .B(n829), .Z(n788) );
  XNOR U234 ( .A(n728), .B(n727), .Z(n726) );
  ANDN U235 ( .A(n681), .B(n680), .Z(n679) );
  XNOR U236 ( .A(n3732), .B(n3697), .Z(n3701) );
  MUX U237 ( .IN0(n71), .IN1(n4514), .SEL(n4515), .F(n4499) );
  IV U238 ( .A(n4516), .Z(n71) );
  MUX U239 ( .IN0(n4109), .IN1(n4107), .SEL(n4108), .F(n4090) );
  MUX U240 ( .IN0(n72), .IN1(n3762), .SEL(n3177), .F(n3724) );
  IV U241 ( .A(n3176), .Z(n72) );
  XOR U242 ( .A(n3715), .B(n3680), .Z(n3684) );
  XOR U243 ( .A(n4489), .B(n4481), .Z(n4083) );
  XOR U244 ( .A(n4461), .B(n4462), .Z(n4065) );
  MUX U245 ( .IN0(n3588), .IN1(n3586), .SEL(n3587), .F(n3548) );
  MUX U246 ( .IN0(n73), .IN1(n3506), .SEL(n3507), .F(n3468) );
  IV U247 ( .A(n3508), .Z(n73) );
  XNOR U248 ( .A(n4050), .B(n4036), .Z(n4040) );
  XOR U249 ( .A(n3563), .B(n3528), .Z(n3532) );
  XOR U250 ( .A(n4437), .B(n4429), .Z(n4015) );
  MUX U251 ( .IN0(n74), .IN1(n4595), .SEL(n4596), .F(n4584) );
  IV U252 ( .A(n4597), .Z(n74) );
  MUX U253 ( .IN0(n75), .IN1(n4963), .SEL(n4964), .F(n4950) );
  IV U254 ( .A(n4965), .Z(n75) );
  XOR U255 ( .A(n4979), .B(n4971), .Z(n4847) );
  XNOR U256 ( .A(n3999), .B(n3985), .Z(n3989) );
  XNOR U257 ( .A(n3428), .B(n3393), .Z(n3397) );
  XOR U258 ( .A(n4598), .B(n4590), .Z(n4259) );
  XOR U259 ( .A(n4853), .B(n4835), .Z(n4839) );
  XOR U260 ( .A(n3449), .B(n3414), .Z(n3418) );
  XOR U261 ( .A(n4265), .B(n4247), .Z(n4251) );
  MUX U262 ( .IN0(n76), .IN1(n4395), .SEL(n4396), .F(n4382) );
  IV U263 ( .A(n4397), .Z(n76) );
  MUX U264 ( .IN0(n77), .IN1(n3324), .SEL(n3325), .F(n3286) );
  IV U265 ( .A(n3326), .Z(n77) );
  MUX U266 ( .IN0(n78), .IN1(n3941), .SEL(n3942), .F(n3924) );
  IV U267 ( .A(n3943), .Z(n78) );
  XOR U268 ( .A(n4385), .B(n4377), .Z(n3947) );
  XOR U269 ( .A(n4940), .B(n4932), .Z(n4784) );
  XNOR U270 ( .A(n3948), .B(n3934), .Z(n3938) );
  MUX U271 ( .IN0(n4775), .IN1(n79), .SEL(n4776), .F(n4754) );
  IV U272 ( .A(n4777), .Z(n79) );
  XOR U273 ( .A(n3335), .B(n3300), .Z(n3304) );
  MUX U274 ( .IN0(n4560), .IN1(n80), .SEL(n4196), .F(n4549) );
  IV U275 ( .A(n4194), .Z(n80) );
  MUX U276 ( .IN0(n4187), .IN1(n81), .SEL(n4188), .F(n4166) );
  IV U277 ( .A(n4189), .Z(n81) );
  XOR U278 ( .A(n4725), .B(n4726), .Z(n4735) );
  MUX U279 ( .IN0(n3246), .IN1(n3244), .SEL(n3245), .F(n3206) );
  XOR U280 ( .A(n4706), .B(n4707), .Z(n4703) );
  MUX U281 ( .IN0(n82), .IN1(n3165), .SEL(n3166), .F(n3036) );
  IV U282 ( .A(n3167), .Z(n82) );
  MUX U283 ( .IN0(n3885), .IN1(n3883), .SEL(n3884), .F(n3185) );
  MUX U284 ( .IN0(n83), .IN1(n3895), .SEL(n3896), .F(n4327) );
  IV U285 ( .A(n4341), .Z(n83) );
  MUX U286 ( .IN0(n4896), .IN1(n84), .SEL(n4721), .F(n3110) );
  IV U287 ( .A(n4719), .Z(n84) );
  MUX U288 ( .IN0(n3160), .IN1(n3162), .SEL(n3161), .F(n3031) );
  MUX U289 ( .IN0(n85), .IN1(n2971), .SEL(n2972), .F(n2833) );
  IV U290 ( .A(n2973), .Z(n85) );
  MUX U291 ( .IN0(n86), .IN1(n2947), .SEL(n2948), .F(n2809) );
  IV U292 ( .A(n2949), .Z(n86) );
  MUX U293 ( .IN0(n87), .IN1(n2759), .SEL(n2760), .F(n2633) );
  IV U294 ( .A(n2761), .Z(n87) );
  MUX U295 ( .IN0(n88), .IN1(n2850), .SEL(n2851), .F(n2718) );
  IV U296 ( .A(n2852), .Z(n88) );
  MUX U297 ( .IN0(n89), .IN1(n2917), .SEL(n2918), .F(n2793) );
  IV U298 ( .A(n2919), .Z(n89) );
  MUX U299 ( .IN0(n90), .IN1(n2426), .SEL(n2427), .F(n2305) );
  IV U300 ( .A(n2428), .Z(n90) );
  MUX U301 ( .IN0(n91), .IN1(n2450), .SEL(n2451), .F(n2329) );
  IV U302 ( .A(n2452), .Z(n91) );
  MUX U303 ( .IN0(n92), .IN1(n2338), .SEL(n2339), .F(n2222) );
  IV U304 ( .A(n2340), .Z(n92) );
  MUX U305 ( .IN0(n93), .IN1(n2346), .SEL(n2347), .F(n2230) );
  IV U306 ( .A(n2348), .Z(n93) );
  MUX U307 ( .IN0(n94), .IN1(n2168), .SEL(n2169), .F(n2059) );
  IV U308 ( .A(n2170), .Z(n94) );
  MUX U309 ( .IN0(n95), .IN1(n1818), .SEL(n1819), .F(n1722) );
  IV U310 ( .A(n1820), .Z(n95) );
  MUX U311 ( .IN0(n96), .IN1(n1809), .SEL(n1810), .F(n1713) );
  IV U312 ( .A(n1811), .Z(n96) );
  MUX U313 ( .IN0(n97), .IN1(n1581), .SEL(n1582), .F(n1488) );
  IV U314 ( .A(n1583), .Z(n97) );
  MUX U315 ( .IN0(n98), .IN1(n1444), .SEL(n1445), .F(n1367) );
  IV U316 ( .A(n1446), .Z(n98) );
  MUX U317 ( .IN0(n99), .IN1(n1261), .SEL(n1262), .F(n1195) );
  IV U318 ( .A(n1263), .Z(n99) );
  MUX U319 ( .IN0(n100), .IN1(n1235), .SEL(n1236), .F(n1169) );
  IV U320 ( .A(n1237), .Z(n100) );
  MUX U321 ( .IN0(n101), .IN1(n1039), .SEL(n1040), .F(n983) );
  IV U322 ( .A(n1041), .Z(n101) );
  MUX U323 ( .IN0(n102), .IN1(n891), .SEL(n892), .F(n847) );
  IV U324 ( .A(n893), .Z(n102) );
  XOR U325 ( .A(n3072), .B(n3073), .Z(n3078) );
  MUX U326 ( .IN0(n2774), .IN1(n2772), .SEL(n2773), .F(n2646) );
  XNOR U327 ( .A(n2785), .B(n2786), .Z(n2784) );
  MUX U328 ( .IN0(n2683), .IN1(n2681), .SEL(n2682), .F(n2554) );
  MUX U329 ( .IN0(n2705), .IN1(n2707), .SEL(n2706), .F(n2578) );
  MUX U330 ( .IN0(n2595), .IN1(n2597), .SEL(n2596), .F(n2471) );
  MUX U331 ( .IN0(n2390), .IN1(n2392), .SEL(n2391), .F(n2269) );
  MUX U332 ( .IN0(n2195), .IN1(n2193), .SEL(n2194), .F(n2082) );
  MUX U333 ( .IN0(n2217), .IN1(n2219), .SEL(n2218), .F(n2106) );
  MUX U334 ( .IN0(n2134), .IN1(n2132), .SEL(n2133), .F(n2027) );
  MUX U335 ( .IN0(n2123), .IN1(n2125), .SEL(n2124), .F(n2018) );
  MUX U336 ( .IN0(n1960), .IN1(n1958), .SEL(n1959), .F(n1845) );
  MUX U337 ( .IN0(n1796), .IN1(n1798), .SEL(n1797), .F(n1700) );
  MUX U338 ( .IN0(n1774), .IN1(n1772), .SEL(n1773), .F(n1676) );
  MUX U339 ( .IN0(n1626), .IN1(n1628), .SEL(n1627), .F(n1534) );
  MUX U340 ( .IN0(n1545), .IN1(n1543), .SEL(n1544), .F(n1457) );
  MUX U341 ( .IN0(n1409), .IN1(n1407), .SEL(n1408), .F(n1335) );
  MUX U342 ( .IN0(n1433), .IN1(n1431), .SEL(n1432), .F(n103) );
  MUX U343 ( .IN0(n929), .IN1(n931), .SEL(n930), .F(n883) );
  MUX U344 ( .IN0(n104), .IN1(n3118), .SEL(n3119), .F(n2983) );
  IV U345 ( .A(n3120), .Z(n104) );
  MUX U346 ( .IN0(n2966), .IN1(n105), .SEL(n2967), .F(n2828) );
  IV U347 ( .A(n2968), .Z(n105) );
  XNOR U348 ( .A(n2725), .B(n2601), .Z(n2605) );
  MUX U349 ( .IN0(n106), .IN1(n2502), .SEL(n2503), .F(n2381) );
  IV U350 ( .A(n2504), .Z(n106) );
  MUX U351 ( .IN0(n107), .IN1(n2462), .SEL(n2463), .F(n2341) );
  IV U352 ( .A(n2464), .Z(n107) );
  MUX U353 ( .IN0(n2051), .IN1(n108), .SEL(n2052), .F(n1949) );
  IV U354 ( .A(n2053), .Z(n108) );
  MUX U355 ( .IN0(n109), .IN1(n1904), .SEL(n1905), .F(n1804) );
  IV U356 ( .A(n1906), .Z(n109) );
  MUX U357 ( .IN0(n110), .IN1(n1362), .SEL(n1363), .F(n1291) );
  IV U358 ( .A(n1364), .Z(n110) );
  MUX U359 ( .IN0(n1285), .IN1(n111), .SEL(n1284), .F(n1211) );
  IV U360 ( .A(n1283), .Z(n111) );
  MUX U361 ( .IN0(n112), .IN1(n1093), .SEL(n1094), .F(n1034) );
  IV U362 ( .A(n1095), .Z(n112) );
  MUX U363 ( .IN0(n1075), .IN1(n1073), .SEL(n1074), .F(n1015) );
  MUX U364 ( .IN0(n113), .IN1(n839), .SEL(n840), .F(n801) );
  IV U365 ( .A(n841), .Z(n113) );
  AND U366 ( .A(n800), .B(n799), .Z(n796) );
  MUX U367 ( .IN0(n114), .IN1(n2928), .SEL(n2929), .F(n2800) );
  IV U368 ( .A(n2930), .Z(n114) );
  MUX U369 ( .IN0(n115), .IN1(n2820), .SEL(n2821), .F(n2688) );
  IV U370 ( .A(n2822), .Z(n115) );
  MUX U371 ( .IN0(n116), .IN1(n2200), .SEL(n2201), .F(n2089) );
  IV U372 ( .A(n2202), .Z(n116) );
  MUX U373 ( .IN0(n117), .IN1(n1683), .SEL(n1684), .F(n1592) );
  IV U374 ( .A(n1685), .Z(n117) );
  MUX U375 ( .IN0(n118), .IN1(n1206), .SEL(n1207), .F(n1144) );
  IV U376 ( .A(n1208), .Z(n118) );
  MUX U377 ( .IN0(n773), .IN1(n771), .SEL(n772), .F(n735) );
  MUX U378 ( .IN0(n2529), .IN1(n119), .SEL(n2530), .F(n2406) );
  IV U379 ( .A(n2531), .Z(n119) );
  XNOR U380 ( .A(n2267), .B(n2266), .Z(n2297) );
  MUX U381 ( .IN0(n1965), .IN1(n120), .SEL(n1966), .F(n1860) );
  IV U382 ( .A(n1967), .Z(n120) );
  ANDN U383 ( .A(n2036), .B(n2037), .Z(n1931) );
  NANDN U384 ( .B(n1763), .A(n1764), .Z(n1667) );
  ANDN U385 ( .A(n1552), .B(n1553), .Z(n1466) );
  ANDN U386 ( .A(n1248), .B(n1249), .Z(n1181) );
  OR U387 ( .A(n870), .B(n871), .Z(n830) );
  XNOR U388 ( .A(n1397), .B(n1479), .Z(n1474) );
  OR U389 ( .A(n1068), .B(n1069), .Z(n1012) );
  XNOR U390 ( .A(n971), .B(n970), .Z(n955) );
  MUX U391 ( .IN0(n121), .IN1(n905), .SEL(n906), .F(n861) );
  IV U392 ( .A(\_MxM/Y0[24] ), .Z(n121) );
  AND U393 ( .A(n859), .B(n860), .Z(n819) );
  OR U394 ( .A(n755), .B(n756), .Z(n725) );
  OR U395 ( .A(n702), .B(n703), .Z(n680) );
  MUX U396 ( .IN0(n122), .IN1(n2615), .SEL(n657), .F(n2491) );
  IV U397 ( .A(\_MxM/Y0[4] ), .Z(n122) );
  MUX U398 ( .IN0(n2143), .IN1(n123), .SEL(n653), .F(n2038) );
  IV U399 ( .A(\_MxM/Y0[8] ), .Z(n123) );
  MUX U400 ( .IN0(n1739), .IN1(n124), .SEL(n1740), .F(n1646) );
  IV U401 ( .A(\_MxM/Y0[12] ), .Z(n124) );
  MUX U402 ( .IN0(n1391), .IN1(n125), .SEL(n1392), .F(n1320) );
  IV U403 ( .A(\_MxM/Y0[16] ), .Z(n125) );
  MUX U404 ( .IN0(n126), .IN1(n1121), .SEL(n1122), .F(n1062) );
  IV U405 ( .A(\_MxM/Y0[20] ), .Z(n126) );
  MUX U406 ( .IN0(n127), .IN1(n3666), .SEL(n3667), .F(n3628) );
  IV U407 ( .A(n3668), .Z(n127) );
  MUX U408 ( .IN0(n128), .IN1(n3658), .SEL(n3659), .F(n3620) );
  IV U409 ( .A(n3660), .Z(n128) );
  MUX U410 ( .IN0(n129), .IN1(n4521), .SEL(n4522), .F(n4506) );
  IV U411 ( .A(n4523), .Z(n129) );
  MUX U412 ( .IN0(n130), .IN1(n4131), .SEL(n3765), .F(n4114) );
  IV U413 ( .A(n3764), .Z(n130) );
  XNOR U414 ( .A(n4118), .B(n4104), .Z(n4108) );
  MUX U415 ( .IN0(n131), .IN1(n4094), .SEL(n4095), .F(n4077) );
  IV U416 ( .A(n4096), .Z(n131) );
  MUX U417 ( .IN0(n132), .IN1(n4499), .SEL(n4500), .F(n4486) );
  IV U418 ( .A(n4501), .Z(n132) );
  MUX U419 ( .IN0(n3712), .IN1(n133), .SEL(n3713), .F(n3674) );
  IV U420 ( .A(n3714), .Z(n133) );
  XOR U421 ( .A(n3677), .B(n3642), .Z(n3646) );
  XOR U422 ( .A(n4476), .B(n4468), .Z(n4066) );
  XNOR U423 ( .A(n4067), .B(n4053), .Z(n4057) );
  XOR U424 ( .A(n4448), .B(n4449), .Z(n4048) );
  MUX U425 ( .IN0(n134), .IN1(n3514), .SEL(n3515), .F(n3476) );
  IV U426 ( .A(n3516), .Z(n134) );
  XNOR U427 ( .A(n3542), .B(n3507), .Z(n3511) );
  XOR U428 ( .A(n4435), .B(n4436), .Z(n4031) );
  MUX U429 ( .IN0(n135), .IN1(n4288), .SEL(n4289), .F(n4267) );
  IV U430 ( .A(n4290), .Z(n135) );
  XOR U431 ( .A(n4422), .B(n4423), .Z(n4014) );
  XNOR U432 ( .A(n4016), .B(n4002), .Z(n4006) );
  XOR U433 ( .A(n3525), .B(n3490), .Z(n3494) );
  XOR U434 ( .A(n4409), .B(n4410), .Z(n3997) );
  MUX U435 ( .IN0(n136), .IN1(n4970), .SEL(n4971), .F(n4957) );
  IV U436 ( .A(n4972), .Z(n136) );
  MUX U437 ( .IN0(n137), .IN1(n4428), .SEL(n4429), .F(n4415) );
  IV U438 ( .A(n4430), .Z(n137) );
  MUX U439 ( .IN0(n4604), .IN1(n138), .SEL(n4280), .F(n4593) );
  IV U440 ( .A(n4278), .Z(n138) );
  MUX U441 ( .IN0(n139), .IN1(n4584), .SEL(n4585), .F(n4573) );
  IV U442 ( .A(n4586), .Z(n139) );
  MUX U443 ( .IN0(n4974), .IN1(n140), .SEL(n4847), .F(n4961) );
  IV U444 ( .A(n4845), .Z(n140) );
  MUX U445 ( .IN0(n4838), .IN1(n141), .SEL(n4839), .F(n4817) );
  IV U446 ( .A(n4840), .Z(n141) );
  MUX U447 ( .IN0(n3398), .IN1(n3396), .SEL(n3397), .F(n3358) );
  MUX U448 ( .IN0(n142), .IN1(n3354), .SEL(n3355), .F(n3316) );
  IV U449 ( .A(n3356), .Z(n142) );
  MUX U450 ( .IN0(n143), .IN1(n4671), .SEL(n4672), .F(n4656) );
  IV U451 ( .A(n4673), .Z(n143) );
  MUX U452 ( .IN0(n144), .IN1(n4666), .SEL(n4667), .F(n4650) );
  IV U453 ( .A(n4668), .Z(n144) );
  MUX U454 ( .IN0(n145), .IN1(n4578), .SEL(n4579), .F(n4567) );
  IV U455 ( .A(n4580), .Z(n145) );
  MUX U456 ( .IN0(n4250), .IN1(n146), .SEL(n4251), .F(n4229) );
  IV U457 ( .A(n4252), .Z(n146) );
  MUX U458 ( .IN0(n147), .IN1(n5043), .SEL(n5044), .F(n5028) );
  IV U459 ( .A(n5045), .Z(n147) );
  MUX U460 ( .IN0(n148), .IN1(n5038), .SEL(n5039), .F(n5022) );
  IV U461 ( .A(n5040), .Z(n148) );
  MUX U462 ( .IN0(n149), .IN1(n4787), .SEL(n4788), .F(n4766) );
  IV U463 ( .A(n4789), .Z(n149) );
  MUX U464 ( .IN0(n150), .IN1(n4792), .SEL(n4793), .F(n4771) );
  IV U465 ( .A(n4794), .Z(n150) );
  XNOR U466 ( .A(n3965), .B(n3951), .Z(n3955) );
  XOR U467 ( .A(n3411), .B(n3376), .Z(n3380) );
  MUX U468 ( .IN0(n151), .IN1(n3819), .SEL(n3820), .F(n3803) );
  IV U469 ( .A(n3821), .Z(n151) );
  XOR U470 ( .A(n4200), .B(n4201), .Z(n4210) );
  MUX U471 ( .IN0(n152), .IN1(n5128), .SEL(n5129), .F(n5110) );
  IV U472 ( .A(n5130), .Z(n152) );
  MUX U473 ( .IN0(n153), .IN1(n4924), .SEL(n4925), .F(n4911) );
  IV U474 ( .A(n4926), .Z(n153) );
  MUX U475 ( .IN0(n154), .IN1(n3924), .SEL(n3925), .F(n3907) );
  IV U476 ( .A(n3926), .Z(n154) );
  XOR U477 ( .A(n4179), .B(n4180), .Z(n4189) );
  MUX U478 ( .IN0(n155), .IN1(n4369), .SEL(n4370), .F(n4356) );
  IV U479 ( .A(n4371), .Z(n155) );
  XOR U480 ( .A(n4927), .B(n4919), .Z(n4763) );
  MUX U481 ( .IN0(n156), .IN1(n3944), .SEL(n3350), .F(n3927) );
  IV U482 ( .A(n3348), .Z(n156) );
  XNOR U483 ( .A(n3276), .B(n3241), .Z(n3245) );
  XOR U484 ( .A(n4554), .B(n4546), .Z(n4175) );
  XOR U485 ( .A(n4158), .B(n4159), .Z(n4168) );
  MUX U486 ( .IN0(n157), .IN1(n4162), .SEL(n4163), .F(n4137) );
  IV U487 ( .A(n4164), .Z(n157) );
  MUX U488 ( .IN0(n158), .IN1(n5165), .SEL(n5166), .F(n5161) );
  IV U489 ( .A(n5167), .Z(n158) );
  MUX U490 ( .IN0(n159), .IN1(n3210), .SEL(n3211), .F(n3173) );
  IV U491 ( .A(n3212), .Z(n159) );
  XOR U492 ( .A(n3297), .B(n3262), .Z(n3266) );
  MUX U493 ( .IN0(n4354), .IN1(n160), .SEL(n3913), .F(n4341) );
  IV U494 ( .A(n3912), .Z(n160) );
  XOR U495 ( .A(n4748), .B(n4730), .Z(n4734) );
  XNOR U496 ( .A(n3897), .B(n3880), .Z(n3884) );
  MUX U497 ( .IN0(n161), .IN1(n2833), .SEL(n2834), .F(n2701) );
  IV U498 ( .A(n2835), .Z(n161) );
  MUX U499 ( .IN0(n162), .IN1(n2718), .SEL(n2719), .F(n2591) );
  IV U500 ( .A(n2720), .Z(n162) );
  MUX U501 ( .IN0(n163), .IN1(n2685), .SEL(n2686), .F(n2558) );
  IV U502 ( .A(n2687), .Z(n163) );
  MUX U503 ( .IN0(n164), .IN1(n2386), .SEL(n2387), .F(n2275) );
  IV U504 ( .A(n2388), .Z(n164) );
  MUX U505 ( .IN0(n165), .IN1(n2230), .SEL(n2231), .F(n2119) );
  IV U506 ( .A(n2232), .Z(n165) );
  MUX U507 ( .IN0(n166), .IN1(n1981), .SEL(n1982), .F(n1876) );
  IV U508 ( .A(n1983), .Z(n166) );
  MUX U509 ( .IN0(n167), .IN1(n1997), .SEL(n1998), .F(n1892) );
  IV U510 ( .A(n1999), .Z(n167) );
  MUX U511 ( .IN0(n168), .IN1(n1713), .SEL(n1714), .F(n1622) );
  IV U512 ( .A(n1715), .Z(n168) );
  MUX U513 ( .IN0(n169), .IN1(n1589), .SEL(n1590), .F(n1496) );
  IV U514 ( .A(n1591), .Z(n169) );
  MUX U515 ( .IN0(n170), .IN1(n1962), .SEL(n1963), .F(n1857) );
  IV U516 ( .A(n1964), .Z(n170) );
  MUX U517 ( .IN0(n171), .IN1(n1954), .SEL(n1955), .F(n1853) );
  IV U518 ( .A(n1956), .Z(n171) );
  MUX U519 ( .IN0(n172), .IN1(n1367), .SEL(n1368), .F(n1296) );
  IV U520 ( .A(n1369), .Z(n172) );
  MUX U521 ( .IN0(n173), .IN1(n1098), .SEL(n1099), .F(n1039) );
  IV U522 ( .A(n1100), .Z(n173) );
  MUX U523 ( .IN0(n174), .IN1(n1107), .SEL(n1108), .F(n1048) );
  IV U524 ( .A(n1109), .Z(n174) );
  MUX U525 ( .IN0(n175), .IN1(n1195), .SEL(n1196), .F(n1132) );
  IV U526 ( .A(n1197), .Z(n175) );
  MUX U527 ( .IN0(n176), .IN1(n1203), .SEL(n1204), .F(n1141) );
  IV U528 ( .A(n1205), .Z(n176) );
  MUX U529 ( .IN0(n3110), .IN1(n3112), .SEL(n3111), .F(n2975) );
  XNOR U530 ( .A(n3163), .B(n3037), .Z(n3041) );
  XOR U531 ( .A(n3154), .B(n3028), .Z(n3032) );
  MUX U532 ( .IN0(n3876), .IN1(n177), .SEL(n3198), .F(n3074) );
  IV U533 ( .A(n3197), .Z(n177) );
  MUX U534 ( .IN0(n2992), .IN1(n2994), .SEL(n2993), .F(n2854) );
  MUX U535 ( .IN0(n2923), .IN1(n2921), .SEL(n2922), .F(n2785) );
  MUX U536 ( .IN0(n2637), .IN1(n2639), .SEL(n2638), .F(n2511) );
  MUX U537 ( .IN0(n2648), .IN1(n2646), .SEL(n2647), .F(n2520) );
  MUX U538 ( .IN0(n2578), .IN1(n2580), .SEL(n2579), .F(n2454) );
  MUX U539 ( .IN0(n2471), .IN1(n2473), .SEL(n2472), .F(n2350) );
  MUX U540 ( .IN0(n2174), .IN1(n2172), .SEL(n2173), .F(n2063) );
  MUX U541 ( .IN0(n2165), .IN1(n178), .SEL(n2164), .F(n2054) );
  IV U542 ( .A(n2163), .Z(n178) );
  MUX U543 ( .IN0(n2106), .IN1(n2108), .SEL(n2107), .F(n2001) );
  MUX U544 ( .IN0(n2018), .IN1(n2020), .SEL(n2019), .F(n1913) );
  XNOR U545 ( .A(n1845), .B(n1846), .Z(n1844) );
  MUX U546 ( .IN0(n1534), .IN1(n1536), .SEL(n1535), .F(n1448) );
  MUX U547 ( .IN0(n1311), .IN1(n1309), .SEL(n1310), .F(n1239) );
  MUX U548 ( .IN0(n1230), .IN1(n1232), .SEL(n1231), .F(n1164) );
  MUX U549 ( .IN0(n940), .IN1(n938), .SEL(n939), .F(n895) );
  XNOR U550 ( .A(n3130), .B(n2998), .Z(n3002) );
  XNOR U551 ( .A(n3080), .B(n2948), .Z(n2952) );
  MUX U552 ( .IN0(n3078), .IN1(n476), .SEL(n3077), .F(n2940) );
  MUX U553 ( .IN0(n179), .IN1(n2845), .SEL(n2846), .F(n2713) );
  IV U554 ( .A(n2847), .Z(n179) );
  MUX U555 ( .IN0(n2696), .IN1(n180), .SEL(n2697), .F(n2569) );
  IV U556 ( .A(n2698), .Z(n180) );
  XNOR U557 ( .A(n2548), .B(n2427), .Z(n2431) );
  XNOR U558 ( .A(n2598), .B(n2477), .Z(n2481) );
  MUX U559 ( .IN0(n181), .IN1(n2381), .SEL(n2382), .F(n2265) );
  IV U560 ( .A(n2383), .Z(n181) );
  MUX U561 ( .IN0(n2535), .IN1(n2533), .SEL(n2534), .F(n2419) );
  MUX U562 ( .IN0(n182), .IN1(n2341), .SEL(n2342), .F(n2225) );
  IV U563 ( .A(n2343), .Z(n182) );
  XNOR U564 ( .A(n2237), .B(n2129), .Z(n2133) );
  MUX U565 ( .IN0(n2208), .IN1(n183), .SEL(n2209), .F(n2097) );
  IV U566 ( .A(n2210), .Z(n183) );
  XNOR U567 ( .A(n1971), .B(n1869), .Z(n1873) );
  MUX U568 ( .IN0(n1949), .IN1(n184), .SEL(n1950), .F(n1840) );
  IV U569 ( .A(n1951), .Z(n184) );
  XNOR U570 ( .A(n1816), .B(n1723), .Z(n1729) );
  MUX U571 ( .IN0(n185), .IN1(n1804), .SEL(n1805), .F(n1708) );
  IV U572 ( .A(n1806), .Z(n185) );
  MUX U573 ( .IN0(n1787), .IN1(n186), .SEL(n1788), .F(n1691) );
  IV U574 ( .A(n1789), .Z(n186) );
  XOR U575 ( .A(n1694), .B(n1606), .Z(n1610) );
  XNOR U576 ( .A(n1579), .B(n1489), .Z(n1493) );
  XOR U577 ( .A(n1420), .B(n1421), .Z(n1433) );
  MUX U578 ( .IN0(n187), .IN1(n1439), .SEL(n1440), .F(n1362) );
  IV U579 ( .A(n1441), .Z(n187) );
  MUX U580 ( .IN0(n188), .IN1(n1352), .SEL(n1353), .F(n1283) );
  IV U581 ( .A(n1354), .Z(n188) );
  MUX U582 ( .IN0(n189), .IN1(n1155), .SEL(n1156), .F(n1093) );
  IV U583 ( .A(n1157), .Z(n189) );
  XOR U584 ( .A(n980), .B(n926), .Z(n930) );
  MUX U585 ( .IN0(n803), .IN1(n190), .SEL(n802), .F(n761) );
  IV U586 ( .A(n801), .Z(n190) );
  MUX U587 ( .IN0(n191), .IN1(n816), .SEL(n817), .F(n776) );
  IV U588 ( .A(n818), .Z(n191) );
  MUX U589 ( .IN0(n192), .IN1(n3093), .SEL(n3094), .F(n2958) );
  IV U590 ( .A(n3095), .Z(n192) );
  MUX U591 ( .IN0(n193), .IN1(n2800), .SEL(n2801), .F(n2671) );
  IV U592 ( .A(n2802), .Z(n193) );
  MUX U593 ( .IN0(n194), .IN1(n2561), .SEL(n2562), .F(n2437) );
  IV U594 ( .A(n2563), .Z(n194) );
  MUX U595 ( .IN0(n195), .IN1(n1984), .SEL(n1985), .F(n1879) );
  IV U596 ( .A(n1986), .Z(n195) );
  MUX U597 ( .IN0(n196), .IN1(n1592), .SEL(n1593), .F(n1499) );
  IV U598 ( .A(n1594), .Z(n196) );
  MUX U599 ( .IN0(n197), .IN1(n1272), .SEL(n1273), .F(n1206) );
  IV U600 ( .A(n1274), .Z(n197) );
  OR U601 ( .A(n1086), .B(n1087), .Z(n1027) );
  XNOR U602 ( .A(n765), .B(n738), .Z(n736) );
  ANDN U603 ( .A(n2614), .B(n2613), .Z(n2489) );
  MUX U604 ( .IN0(n2291), .IN1(n198), .SEL(n2292), .F(n2179) );
  IV U605 ( .A(n2293), .Z(n198) );
  MUX U606 ( .IN0(n2182), .IN1(n2294), .SEL(n2184), .F(n2073) );
  ANDN U607 ( .A(n2141), .B(n2142), .Z(n2036) );
  MUX U608 ( .IN0(n1760), .IN1(n199), .SEL(n1761), .F(n1664) );
  IV U609 ( .A(n1762), .Z(n199) );
  NANDN U610 ( .B(n1667), .A(n1668), .Z(n1561) );
  ANDN U611 ( .A(n1466), .B(n1467), .Z(n1389) );
  AND U612 ( .A(n1181), .B(n1182), .Z(n1119) );
  XNOR U613 ( .A(n1036), .B(n1035), .Z(n1026) );
  AND U614 ( .A(n946), .B(n947), .Z(n903) );
  MUX U615 ( .IN0(n1399), .IN1(n1397), .SEL(n1398), .F(n1326) );
  OR U616 ( .A(n1128), .B(n1129), .Z(n1068) );
  OR U617 ( .A(n911), .B(n912), .Z(n868) );
  XNOR U618 ( .A(n833), .B(n830), .Z(n829) );
  AND U619 ( .A(n779), .B(n780), .Z(n746) );
  OR U620 ( .A(n725), .B(n726), .Z(n700) );
  MUX U621 ( .IN0(n2491), .IN1(n200), .SEL(n656), .F(n2370) );
  IV U622 ( .A(\_MxM/Y0[5] ), .Z(n200) );
  MUX U623 ( .IN0(n2038), .IN1(n201), .SEL(n652), .F(n1933) );
  IV U624 ( .A(\_MxM/Y0[9] ), .Z(n201) );
  MUX U625 ( .IN0(n1646), .IN1(n202), .SEL(n1647), .F(n1554) );
  IV U626 ( .A(\_MxM/Y0[13] ), .Z(n202) );
  MUX U627 ( .IN0(n1320), .IN1(n203), .SEL(n1321), .F(n1250) );
  IV U628 ( .A(\_MxM/Y0[17] ), .Z(n203) );
  MUX U629 ( .IN0(n204), .IN1(n1062), .SEL(n1063), .F(n1006) );
  IV U630 ( .A(\_MxM/Y0[21] ), .Z(n204) );
  AND U631 ( .A(n688), .B(n689), .Z(n684) );
  MUX U632 ( .IN0(n205), .IN1(n3747), .SEL(n3748), .F(n3709) );
  IV U633 ( .A(n3749), .Z(n205) );
  MUX U634 ( .IN0(n3702), .IN1(n3700), .SEL(n3701), .F(n3662) );
  MUX U635 ( .IN0(n206), .IN1(n3679), .SEL(n3680), .F(n3641) );
  IV U636 ( .A(n3681), .Z(n206) );
  MUX U637 ( .IN0(n207), .IN1(n3620), .SEL(n3621), .F(n3582) );
  IV U638 ( .A(n3622), .Z(n207) );
  MUX U639 ( .IN0(n208), .IN1(n4506), .SEL(n4507), .F(n4493) );
  IV U640 ( .A(n4508), .Z(n208) );
  XNOR U641 ( .A(n4101), .B(n4087), .Z(n4091) );
  MUX U642 ( .IN0(n209), .IN1(n4077), .SEL(n4078), .F(n4060) );
  IV U643 ( .A(n4079), .Z(n209) );
  MUX U644 ( .IN0(n3683), .IN1(n3685), .SEL(n3684), .F(n3645) );
  MUX U645 ( .IN0(n210), .IN1(n4486), .SEL(n4487), .F(n4473) );
  IV U646 ( .A(n4488), .Z(n210) );
  MUX U647 ( .IN0(n211), .IN1(n4080), .SEL(n3654), .F(n4063) );
  IV U648 ( .A(n3652), .Z(n211) );
  MUX U649 ( .IN0(n3636), .IN1(n212), .SEL(n3637), .F(n3598) );
  IV U650 ( .A(n3638), .Z(n212) );
  XOR U651 ( .A(n4463), .B(n4455), .Z(n4049) );
  MUX U652 ( .IN0(n3550), .IN1(n3548), .SEL(n3549), .F(n3510) );
  MUX U653 ( .IN0(n213), .IN1(n3527), .SEL(n3528), .F(n3489) );
  IV U654 ( .A(n3529), .Z(n213) );
  MUX U655 ( .IN0(n214), .IN1(n3476), .SEL(n3477), .F(n3438) );
  IV U656 ( .A(n3478), .Z(n214) );
  MUX U657 ( .IN0(n215), .IN1(n3468), .SEL(n3469), .F(n3430) );
  IV U658 ( .A(n3470), .Z(n215) );
  XNOR U659 ( .A(n4033), .B(n4019), .Z(n4023) );
  MUX U660 ( .IN0(n216), .IN1(n4009), .SEL(n4010), .F(n3992) );
  IV U661 ( .A(n4011), .Z(n216) );
  MUX U662 ( .IN0(n3531), .IN1(n3533), .SEL(n3532), .F(n3493) );
  MUX U663 ( .IN0(n217), .IN1(n4606), .SEL(n4607), .F(n4595) );
  IV U664 ( .A(n4608), .Z(n217) );
  XOR U665 ( .A(n4830), .B(n4831), .Z(n4840) );
  MUX U666 ( .IN0(n218), .IN1(n4012), .SEL(n3502), .F(n3995) );
  IV U667 ( .A(n3500), .Z(n218) );
  MUX U668 ( .IN0(n3484), .IN1(n219), .SEL(n3485), .F(n3446) );
  IV U669 ( .A(n3486), .Z(n219) );
  XOR U670 ( .A(n4286), .B(n4268), .Z(n4272) );
  XOR U671 ( .A(n4242), .B(n4243), .Z(n4252) );
  XOR U672 ( .A(n4411), .B(n4403), .Z(n3981) );
  MUX U673 ( .IN0(n220), .IN1(n4950), .SEL(n4951), .F(n4937) );
  IV U674 ( .A(n4952), .Z(n220) );
  XOR U675 ( .A(n4966), .B(n4958), .Z(n4826) );
  XOR U676 ( .A(n4809), .B(n4810), .Z(n4819) );
  MUX U677 ( .IN0(n221), .IN1(n4813), .SEL(n4814), .F(n4792) );
  IV U678 ( .A(n4815), .Z(n221) );
  XNOR U679 ( .A(n3982), .B(n3968), .Z(n3972) );
  XNOR U680 ( .A(n3390), .B(n3355), .Z(n3359) );
  XOR U681 ( .A(n4587), .B(n4579), .Z(n4238) );
  XOR U682 ( .A(n4221), .B(n4222), .Z(n4231) );
  MUX U683 ( .IN0(n222), .IN1(n4225), .SEL(n4226), .F(n4204) );
  IV U684 ( .A(n4227), .Z(n222) );
  XOR U685 ( .A(n4788), .B(n4789), .Z(n4798) );
  MUX U686 ( .IN0(n3379), .IN1(n3381), .SEL(n3380), .F(n3341) );
  MUX U687 ( .IN0(n223), .IN1(n4319), .SEL(n4320), .F(n4660) );
  IV U688 ( .A(n4674), .Z(n223) );
  MUX U689 ( .IN0(n4650), .IN1(n4665), .SEL(n4652), .F(n4634) );
  MUX U690 ( .IN0(n224), .IN1(n4562), .SEL(n4563), .F(n4551) );
  IV U691 ( .A(n4564), .Z(n224) );
  XOR U692 ( .A(n4370), .B(n4371), .Z(n3946) );
  MUX U693 ( .IN0(n225), .IN1(n4886), .SEL(n4887), .F(n5032) );
  IV U694 ( .A(n5046), .Z(n225) );
  MUX U695 ( .IN0(n5022), .IN1(n5037), .SEL(n5024), .F(n5006) );
  MUX U696 ( .IN0(n226), .IN1(n4931), .SEL(n4932), .F(n4918) );
  IV U697 ( .A(n4933), .Z(n226) );
  MUX U698 ( .IN0(n227), .IN1(n3772), .SEL(n3773), .F(n3813) );
  IV U699 ( .A(n3827), .Z(n227) );
  MUX U700 ( .IN0(n3803), .IN1(n3818), .SEL(n3805), .F(n3787) );
  MUX U701 ( .IN0(n228), .IN1(n5073), .SEL(n5074), .F(n5120) );
  IV U702 ( .A(n5136), .Z(n228) );
  MUX U703 ( .IN0(n229), .IN1(n3248), .SEL(n3249), .F(n3210) );
  IV U704 ( .A(n3250), .Z(n229) );
  MUX U705 ( .IN0(n230), .IN1(n4376), .SEL(n4377), .F(n4363) );
  IV U706 ( .A(n4378), .Z(n230) );
  XNOR U707 ( .A(n3931), .B(n3917), .Z(n3921) );
  MUX U708 ( .IN0(n231), .IN1(n3907), .SEL(n3908), .F(n3887) );
  IV U709 ( .A(n3909), .Z(n231) );
  MUX U710 ( .IN0(n232), .IN1(n3253), .SEL(n3254), .F(n3215) );
  IV U711 ( .A(n3255), .Z(n232) );
  MUX U712 ( .IN0(n3332), .IN1(n233), .SEL(n3333), .F(n3294) );
  IV U713 ( .A(n3334), .Z(n233) );
  MUX U714 ( .IN0(n4922), .IN1(n234), .SEL(n4763), .F(n4909) );
  IV U715 ( .A(n4761), .Z(n234) );
  MUX U716 ( .IN0(n235), .IN1(n4729), .SEL(n4730), .F(n4697) );
  IV U717 ( .A(n4731), .Z(n235) );
  MUX U718 ( .IN0(n236), .IN1(n3223), .SEL(n3224), .F(n3156) );
  IV U719 ( .A(n3225), .Z(n236) );
  XNOR U720 ( .A(n3238), .B(n3203), .Z(n3207) );
  MUX U721 ( .IN0(n4549), .IN1(n237), .SEL(n4175), .F(n4538) );
  IV U722 ( .A(n4173), .Z(n237) );
  XOR U723 ( .A(n4181), .B(n4163), .Z(n4167) );
  XOR U724 ( .A(n4146), .B(n4147), .Z(n4143) );
  MUX U725 ( .IN0(n5069), .IN1(n5097), .SEL(n5071), .F(n3115) );
  MUX U726 ( .IN0(n4733), .IN1(n238), .SEL(n4734), .F(n4701) );
  IV U727 ( .A(n4735), .Z(n238) );
  MUX U728 ( .IN0(n239), .IN1(n4338), .SEL(n4339), .F(n3873) );
  IV U729 ( .A(n4340), .Z(n239) );
  MUX U730 ( .IN0(n240), .IN1(n3123), .SEL(n3124), .F(n2988) );
  IV U731 ( .A(n3125), .Z(n240) );
  MUX U732 ( .IN0(n241), .IN1(n3132), .SEL(n3133), .F(n2997) );
  IV U733 ( .A(n3134), .Z(n241) );
  MUX U734 ( .IN0(n242), .IN1(n3098), .SEL(n3099), .F(n2963) );
  IV U735 ( .A(n3100), .Z(n242) );
  MUX U736 ( .IN0(n243), .IN1(n3106), .SEL(n3107), .F(n2971) );
  IV U737 ( .A(n3108), .Z(n243) );
  NAND U738 ( .A(n4326), .B(n4330), .Z(n4329) );
  MUX U739 ( .IN0(n3187), .IN1(n3185), .SEL(n3186), .F(n3057) );
  MUX U740 ( .IN0(n244), .IN1(n2908), .SEL(n2909), .F(n2776) );
  IV U741 ( .A(n2910), .Z(n244) );
  MUX U742 ( .IN0(n245), .IN1(n2925), .SEL(n2926), .F(n2797) );
  IV U743 ( .A(n2927), .Z(n245) );
  MUX U744 ( .IN0(n246), .IN1(n2642), .SEL(n2643), .F(n2516) );
  IV U745 ( .A(n2644), .Z(n246) );
  MUX U746 ( .IN0(n247), .IN1(n2566), .SEL(n2567), .F(n2442) );
  IV U747 ( .A(n2568), .Z(n247) );
  MUX U748 ( .IN0(n248), .IN1(n2574), .SEL(n2575), .F(n2450) );
  IV U749 ( .A(n2576), .Z(n248) );
  MUX U750 ( .IN0(n249), .IN1(n2558), .SEL(n2559), .F(n2434) );
  IV U751 ( .A(n2560), .Z(n249) );
  MUX U752 ( .IN0(n250), .IN1(n2403), .SEL(n2404), .F(n2288) );
  IV U753 ( .A(n2405), .Z(n250) );
  MUX U754 ( .IN0(n251), .IN1(n2467), .SEL(n2468), .F(n2346) );
  IV U755 ( .A(n2469), .Z(n251) );
  MUX U756 ( .IN0(n252), .IN1(n2059), .SEL(n2060), .F(n1954) );
  IV U757 ( .A(n2061), .Z(n252) );
  MUX U758 ( .IN0(n253), .IN1(n2094), .SEL(n2095), .F(n1989) );
  IV U759 ( .A(n2096), .Z(n253) );
  MUX U760 ( .IN0(n254), .IN1(n1901), .SEL(n1902), .F(n1801) );
  IV U761 ( .A(n1903), .Z(n254) );
  MUX U762 ( .IN0(n255), .IN1(n1688), .SEL(n1689), .F(n1597) );
  IV U763 ( .A(n1690), .Z(n255) );
  MUX U764 ( .IN0(n256), .IN1(n1696), .SEL(n1697), .F(n1605) );
  IV U765 ( .A(n1698), .Z(n256) );
  MUX U766 ( .IN0(n257), .IN1(n1522), .SEL(n1523), .F(n1436) );
  IV U767 ( .A(n1524), .Z(n257) );
  MUX U768 ( .IN0(n258), .IN1(n1530), .SEL(n1531), .F(n1444) );
  IV U769 ( .A(n1532), .Z(n258) );
  MUX U770 ( .IN0(n259), .IN1(n1453), .SEL(n1454), .F(n1376) );
  IV U771 ( .A(n1455), .Z(n259) );
  MUX U772 ( .IN0(n260), .IN1(n1218), .SEL(n1219), .F(n1152) );
  IV U773 ( .A(n1220), .Z(n260) );
  MUX U774 ( .IN0(n261), .IN1(n1169), .SEL(n1170), .F(n1107) );
  IV U775 ( .A(n1171), .Z(n261) );
  MUX U776 ( .IN0(n262), .IN1(n1116), .SEL(n1117), .F(n1057) );
  IV U777 ( .A(n1118), .Z(n262) );
  MUX U778 ( .IN0(n263), .IN1(n934), .SEL(n935), .F(n891) );
  IV U779 ( .A(n936), .Z(n263) );
  MUX U780 ( .IN0(n264), .IN1(n918), .SEL(n919), .F(n875) );
  IV U781 ( .A(n920), .Z(n264) );
  MUX U782 ( .IN0(n265), .IN1(n900), .SEL(n901), .F(n856) );
  IV U783 ( .A(n902), .Z(n265) );
  MUX U784 ( .IN0(n3151), .IN1(n266), .SEL(n3152), .F(n3022) );
  IV U785 ( .A(n3153), .Z(n266) );
  MUX U786 ( .IN0(n2895), .IN1(n2897), .SEL(n2896), .F(n2763) );
  MUX U787 ( .IN0(n2837), .IN1(n2839), .SEL(n2838), .F(n2705) );
  MUX U788 ( .IN0(n2865), .IN1(n2863), .SEL(n2864), .F(n2731) );
  MUX U789 ( .IN0(n2795), .IN1(n267), .SEL(n2794), .F(n2662) );
  IV U790 ( .A(n2793), .Z(n267) );
  MUX U791 ( .IN0(n2722), .IN1(n2724), .SEL(n2723), .F(n2595) );
  MUX U792 ( .IN0(n2333), .IN1(n2335), .SEL(n2334), .F(n2217) );
  MUX U793 ( .IN0(n2234), .IN1(n2236), .SEL(n2235), .F(n2123) );
  MUX U794 ( .IN0(n1979), .IN1(n1977), .SEL(n1978), .F(n1872) );
  MUX U795 ( .IN0(n1587), .IN1(n1585), .SEL(n1586), .F(n1492) );
  MUX U796 ( .IN0(n268), .IN1(n1857), .SEL(n1858), .F(n1757) );
  IV U797 ( .A(n1859), .Z(n268) );
  MUX U798 ( .IN0(n1371), .IN1(n1373), .SEL(n1372), .F(n1300) );
  MUX U799 ( .IN0(n1267), .IN1(n1265), .SEL(n1266), .F(n1199) );
  MUX U800 ( .IN0(n1241), .IN1(n1239), .SEL(n1240), .F(n1173) );
  MUX U801 ( .IN0(n269), .IN1(n1141), .SEL(n1142), .F(n1080) );
  IV U802 ( .A(n1143), .Z(n269) );
  MUX U803 ( .IN0(n998), .IN1(n996), .SEL(n997), .F(n938) );
  MUX U804 ( .IN0(n3101), .IN1(n270), .SEL(n3102), .F(n2966) );
  IV U805 ( .A(n3103), .Z(n270) );
  XNOR U806 ( .A(n3034), .B(n2901), .Z(n2905) );
  XNOR U807 ( .A(n2945), .B(n2810), .Z(n2814) );
  MUX U808 ( .IN0(n2943), .IN1(n271), .SEL(n2942), .F(n2803) );
  IV U809 ( .A(n2941), .Z(n271) );
  MUX U810 ( .IN0(n2569), .IN1(n272), .SEL(n2570), .F(n2445) );
  IV U811 ( .A(n2571), .Z(n272) );
  MUX U812 ( .IN0(n273), .IN1(n2586), .SEL(n2587), .F(n2462) );
  IV U813 ( .A(n2588), .Z(n273) );
  XOR U814 ( .A(n2384), .B(n2276), .Z(n2270) );
  XNOR U815 ( .A(n2393), .B(n2281), .Z(n2285) );
  XNOR U816 ( .A(n2424), .B(n2306), .Z(n2310) );
  NAND U817 ( .A(n2416), .B(n2537), .Z(n2536) );
  XNOR U818 ( .A(n2353), .B(n2240), .Z(n2244) );
  MUX U819 ( .IN0(n2097), .IN1(n274), .SEL(n2098), .F(n1992) );
  IV U820 ( .A(n2099), .Z(n274) );
  MUX U821 ( .IN0(n275), .IN1(n2114), .SEL(n2115), .F(n2009) );
  IV U822 ( .A(n2116), .Z(n275) );
  XOR U823 ( .A(n1995), .B(n1893), .Z(n1897) );
  NAND U824 ( .A(n1753), .B(n1851), .Z(n1850) );
  XOR U825 ( .A(n1907), .B(n1810), .Z(n1814) );
  MUX U826 ( .IN0(n276), .IN1(n1708), .SEL(n1709), .F(n1617) );
  IV U827 ( .A(n1710), .Z(n276) );
  XNOR U828 ( .A(n1720), .B(n1632), .Z(n1636) );
  MUX U829 ( .IN0(n1691), .IN1(n277), .SEL(n1692), .F(n1600) );
  IV U830 ( .A(n1693), .Z(n277) );
  NAND U831 ( .A(n1282), .B(n1347), .Z(n1346) );
  MUX U832 ( .IN0(n278), .IN1(n1291), .SEL(n1292), .F(n1221) );
  IV U833 ( .A(n1293), .Z(n278) );
  XOR U834 ( .A(n1158), .B(n1099), .Z(n1103) );
  MUX U835 ( .IN0(n279), .IN1(n1034), .SEL(n1035), .F(n977) );
  IV U836 ( .A(n1036), .Z(n279) );
  OR U837 ( .A(n1076), .B(n1077), .Z(n1071) );
  XNOR U838 ( .A(n845), .B(n808), .Z(n812) );
  MUX U839 ( .IN0(n842), .IN1(n844), .SEL(n843), .F(n280) );
  IV U840 ( .A(n280), .Z(n794) );
  XNOR U841 ( .A(n3003), .B(n3002), .Z(n2985) );
  MUX U842 ( .IN0(n281), .IN1(n2688), .SEL(n2689), .F(n2561) );
  IV U843 ( .A(n2690), .Z(n281) );
  MUX U844 ( .IN0(n1840), .IN1(n282), .SEL(n1841), .F(n1747) );
  IV U845 ( .A(n1842), .Z(n282) );
  MUX U846 ( .IN0(n283), .IN1(n1879), .SEL(n1880), .F(n1779) );
  IV U847 ( .A(n1881), .Z(n283) );
  MUX U848 ( .IN0(n284), .IN1(n1499), .SEL(n1500), .F(n1414) );
  IV U849 ( .A(n1501), .Z(n284) );
  XNOR U850 ( .A(n773), .B(n772), .Z(n763) );
  MUX U851 ( .IN0(n3047), .IN1(n285), .SEL(n3048), .F(n2911) );
  IV U852 ( .A(n3049), .Z(n285) );
  XNOR U853 ( .A(n2756), .B(n2755), .Z(n2802) );
  XNOR U854 ( .A(n2504), .B(n2503), .Z(n2546) );
  MUX U855 ( .IN0(n2406), .IN1(n286), .SEL(n2407), .F(n2291) );
  IV U856 ( .A(n2408), .Z(n286) );
  ANDN U857 ( .A(n2252), .B(n2253), .Z(n2141) );
  ANDN U858 ( .A(n1831), .B(n1832), .Z(n1737) );
  MUX U859 ( .IN0(n1664), .IN1(n287), .SEL(n1665), .F(n1575) );
  IV U860 ( .A(n1666), .Z(n287) );
  NANDN U861 ( .B(n1561), .A(n1562), .Z(n1479) );
  ANDN U862 ( .A(n1389), .B(n1390), .Z(n1318) );
  XOR U863 ( .A(n1086), .B(n1083), .Z(n1130) );
  AND U864 ( .A(n1060), .B(n1061), .Z(n1004) );
  MUX U865 ( .IN0(n915), .IN1(n288), .SEL(n914), .F(n870) );
  IV U866 ( .A(n913), .Z(n288) );
  XNOR U867 ( .A(n687), .B(n686), .Z(n683) );
  XOR U868 ( .A(n1968), .B(n1965), .Z(n2043) );
  OR U869 ( .A(n1326), .B(n1327), .Z(n1256) );
  XNOR U870 ( .A(n1146), .B(n1145), .Z(n1129) );
  OR U871 ( .A(n954), .B(n955), .Z(n911) );
  OR U872 ( .A(n788), .B(n789), .Z(n755) );
  AND U873 ( .A(n819), .B(n820), .Z(n779) );
  MUX U874 ( .IN0(n289), .IN1(n748), .SEL(n749), .F(n716) );
  IV U875 ( .A(\_MxM/Y0[28] ), .Z(n289) );
  XNOR U876 ( .A(n703), .B(n702), .Z(n701) );
  MUX U877 ( .IN0(n290), .IN1(n2872), .SEL(n1123), .F(n2740) );
  IV U878 ( .A(\_MxM/Y0[2] ), .Z(n290) );
  MUX U879 ( .IN0(n2370), .IN1(n291), .SEL(n655), .F(n2254) );
  IV U880 ( .A(\_MxM/Y0[6] ), .Z(n291) );
  MUX U881 ( .IN0(n1933), .IN1(n292), .SEL(n651), .F(n1833) );
  IV U882 ( .A(\_MxM/Y0[10] ), .Z(n292) );
  MUX U883 ( .IN0(n1554), .IN1(n293), .SEL(n1555), .F(n1468) );
  IV U884 ( .A(\_MxM/Y0[14] ), .Z(n293) );
  MUX U885 ( .IN0(n1250), .IN1(n294), .SEL(n1251), .F(n1183) );
  IV U886 ( .A(\_MxM/Y0[18] ), .Z(n294) );
  MUX U887 ( .IN0(n295), .IN1(n1006), .SEL(n1007), .F(n948) );
  IV U888 ( .A(\_MxM/Y0[22] ), .Z(n295) );
  NAND U889 ( .A(n669), .B(n670), .Z(n668) );
  MUX U890 ( .IN0(n296), .IN1(n3755), .SEL(n3756), .F(n3717) );
  IV U891 ( .A(n3757), .Z(n296) );
  MUX U892 ( .IN0(n297), .IN1(n4111), .SEL(n4112), .F(n4094) );
  IV U893 ( .A(n4113), .Z(n297) );
  MUX U894 ( .IN0(n298), .IN1(n3709), .SEL(n3710), .F(n3671) );
  IV U895 ( .A(n3711), .Z(n298) );
  MUX U896 ( .IN0(n299), .IN1(n3750), .SEL(n3751), .F(n3712) );
  IV U897 ( .A(n3752), .Z(n299) );
  MUX U898 ( .IN0(n300), .IN1(n3628), .SEL(n3629), .F(n3590) );
  IV U899 ( .A(n3630), .Z(n300) );
  MUX U900 ( .IN0(n301), .IN1(n4114), .SEL(n3730), .F(n4097) );
  IV U901 ( .A(n3728), .Z(n301) );
  XNOR U902 ( .A(n3656), .B(n3621), .Z(n3625) );
  XOR U903 ( .A(n4474), .B(n4475), .Z(n4082) );
  MUX U904 ( .IN0(n302), .IN1(n4493), .SEL(n4494), .F(n4480) );
  IV U905 ( .A(n4495), .Z(n302) );
  MUX U906 ( .IN0(n4075), .IN1(n4073), .SEL(n4074), .F(n4056) );
  MUX U907 ( .IN0(n3645), .IN1(n3647), .SEL(n3646), .F(n3607) );
  MUX U908 ( .IN0(n303), .IN1(n3603), .SEL(n3604), .F(n3565) );
  IV U909 ( .A(n3605), .Z(n303) );
  MUX U910 ( .IN0(n304), .IN1(n4043), .SEL(n4044), .F(n4026) );
  IV U911 ( .A(n4045), .Z(n304) );
  MUX U912 ( .IN0(n305), .IN1(n4035), .SEL(n4036), .F(n4018) );
  IV U913 ( .A(n4037), .Z(n305) );
  MUX U914 ( .IN0(n306), .IN1(n3557), .SEL(n3558), .F(n3519) );
  IV U915 ( .A(n3559), .Z(n306) );
  MUX U916 ( .IN0(n3598), .IN1(n307), .SEL(n3599), .F(n3560) );
  IV U917 ( .A(n3600), .Z(n307) );
  MUX U918 ( .IN0(n308), .IN1(n4447), .SEL(n4448), .F(n4434) );
  IV U919 ( .A(n4449), .Z(n308) );
  MUX U920 ( .IN0(n309), .IN1(n4046), .SEL(n3578), .F(n4029) );
  IV U921 ( .A(n3576), .Z(n309) );
  XNOR U922 ( .A(n3504), .B(n3469), .Z(n3473) );
  MUX U923 ( .IN0(n310), .IN1(n4283), .SEL(n4284), .F(n4262) );
  IV U924 ( .A(n4285), .Z(n310) );
  MUX U925 ( .IN0(n311), .IN1(n4611), .SEL(n4612), .F(n4600) );
  IV U926 ( .A(n4613), .Z(n311) );
  MUX U927 ( .IN0(n312), .IN1(n3438), .SEL(n3439), .F(n3400) );
  IV U928 ( .A(n3440), .Z(n312) );
  MUX U929 ( .IN0(n313), .IN1(n4441), .SEL(n4442), .F(n4428) );
  IV U930 ( .A(n4443), .Z(n313) );
  MUX U931 ( .IN0(n4007), .IN1(n4005), .SEL(n4006), .F(n3988) );
  MUX U932 ( .IN0(n3493), .IN1(n3495), .SEL(n3494), .F(n3455) );
  MUX U933 ( .IN0(n314), .IN1(n3451), .SEL(n3452), .F(n3413) );
  IV U934 ( .A(n3453), .Z(n314) );
  MUX U935 ( .IN0(n315), .IN1(n3975), .SEL(n3976), .F(n3958) );
  IV U936 ( .A(n3977), .Z(n315) );
  MUX U937 ( .IN0(n316), .IN1(n3967), .SEL(n3968), .F(n3950) );
  IV U938 ( .A(n3969), .Z(n316) );
  MUX U939 ( .IN0(n317), .IN1(n3405), .SEL(n3406), .F(n3367) );
  IV U940 ( .A(n3407), .Z(n317) );
  MUX U941 ( .IN0(n318), .IN1(n4295), .SEL(n3870), .F(n4274) );
  IV U942 ( .A(n3869), .Z(n318) );
  MUX U943 ( .IN0(n4419), .IN1(n319), .SEL(n3998), .F(n4406) );
  IV U944 ( .A(n3997), .Z(n319) );
  MUX U945 ( .IN0(n320), .IN1(n4862), .SEL(n4709), .F(n4841) );
  IV U946 ( .A(n4708), .Z(n320) );
  MUX U947 ( .IN0(n321), .IN1(n4957), .SEL(n4958), .F(n4944) );
  IV U948 ( .A(n4959), .Z(n321) );
  MUX U949 ( .IN0(n3446), .IN1(n322), .SEL(n3447), .F(n3408) );
  IV U950 ( .A(n3448), .Z(n322) );
  MUX U951 ( .IN0(n4593), .IN1(n323), .SEL(n4259), .F(n4582) );
  IV U952 ( .A(n4257), .Z(n323) );
  MUX U953 ( .IN0(n4961), .IN1(n324), .SEL(n4826), .F(n4948) );
  IV U954 ( .A(n4824), .Z(n324) );
  MUX U955 ( .IN0(n3360), .IN1(n3358), .SEL(n3359), .F(n3320) );
  MUX U956 ( .IN0(n325), .IN1(n3316), .SEL(n3317), .F(n3278) );
  IV U957 ( .A(n3318), .Z(n325) );
  MUX U958 ( .IN0(n326), .IN1(n3978), .SEL(n3426), .F(n3961) );
  IV U959 ( .A(n3424), .Z(n326) );
  MUX U960 ( .IN0(n327), .IN1(n3824), .SEL(n3825), .F(n3809) );
  IV U961 ( .A(n3826), .Z(n327) );
  MUX U962 ( .IN0(n328), .IN1(n4199), .SEL(n4200), .F(n4178) );
  IV U963 ( .A(n4201), .Z(n328) );
  MUX U964 ( .IN0(n4656), .IN1(n4670), .SEL(n4658), .F(n4640) );
  MUX U965 ( .IN0(n329), .IN1(n4686), .SEL(n4687), .F(n4682) );
  IV U966 ( .A(n4688), .Z(n329) );
  MUX U967 ( .IN0(n330), .IN1(n4567), .SEL(n4568), .F(n4556) );
  IV U968 ( .A(n4569), .Z(n330) );
  XOR U969 ( .A(n4244), .B(n4226), .Z(n4230) );
  MUX U970 ( .IN0(n331), .IN1(n4382), .SEL(n4383), .F(n4369) );
  IV U971 ( .A(n4384), .Z(n331) );
  MUX U972 ( .IN0(n332), .IN1(n5133), .SEL(n5134), .F(n5116) );
  IV U973 ( .A(n5135), .Z(n332) );
  MUX U974 ( .IN0(n5028), .IN1(n5042), .SEL(n5030), .F(n5012) );
  MUX U975 ( .IN0(n333), .IN1(n5058), .SEL(n5059), .F(n5054) );
  IV U976 ( .A(n5060), .Z(n333) );
  MUX U977 ( .IN0(n334), .IN1(n4766), .SEL(n4767), .F(n4745) );
  IV U978 ( .A(n4768), .Z(n334) );
  MUX U979 ( .IN0(n4796), .IN1(n335), .SEL(n4797), .F(n4775) );
  IV U980 ( .A(n4798), .Z(n335) );
  MUX U981 ( .IN0(n336), .IN1(n4771), .SEL(n4772), .F(n4750) );
  IV U982 ( .A(n4773), .Z(n336) );
  MUX U983 ( .IN0(n3939), .IN1(n3937), .SEL(n3938), .F(n3920) );
  MUX U984 ( .IN0(n3341), .IN1(n3343), .SEL(n3342), .F(n3303) );
  MUX U985 ( .IN0(n337), .IN1(n3299), .SEL(n3300), .F(n3261) );
  IV U986 ( .A(n3301), .Z(n337) );
  MUX U987 ( .IN0(n338), .IN1(n3840), .SEL(n3841), .F(n3836) );
  IV U988 ( .A(n3842), .Z(n338) );
  MUX U989 ( .IN0(n339), .IN1(n4305), .SEL(n4306), .F(n4301) );
  IV U990 ( .A(n4307), .Z(n339) );
  XOR U991 ( .A(n4563), .B(n4564), .Z(n4215) );
  MUX U992 ( .IN0(n340), .IN1(n4872), .SEL(n4873), .F(n4868) );
  IV U993 ( .A(n4874), .Z(n340) );
  MUX U994 ( .IN0(n341), .IN1(n3899), .SEL(n3900), .F(n3879) );
  IV U995 ( .A(n3901), .Z(n341) );
  MUX U996 ( .IN0(n342), .IN1(n3855), .SEL(n3856), .F(n3851) );
  IV U997 ( .A(n3857), .Z(n342) );
  MUX U998 ( .IN0(n343), .IN1(n4540), .SEL(n4541), .F(n4529) );
  IV U999 ( .A(n4542), .Z(n343) );
  MUX U1000 ( .IN0(n4367), .IN1(n344), .SEL(n3930), .F(n4354) );
  IV U1001 ( .A(n3929), .Z(n344) );
  MUX U1002 ( .IN0(n5144), .IN1(n5147), .SEL(n5145), .F(n5128) );
  MUX U1003 ( .IN0(n345), .IN1(n4898), .SEL(n4899), .F(n4712) );
  IV U1004 ( .A(n4900), .Z(n345) );
  XOR U1005 ( .A(n4914), .B(n4906), .Z(n4742) );
  MUX U1006 ( .IN0(n346), .IN1(n3887), .SEL(n3888), .F(n3189) );
  IV U1007 ( .A(n3889), .Z(n346) );
  MUX U1008 ( .IN0(n3294), .IN1(n347), .SEL(n3295), .F(n3256) );
  IV U1009 ( .A(n3296), .Z(n347) );
  MUX U1010 ( .IN0(n348), .IN1(n4137), .SEL(n4138), .F(n4120) );
  IV U1011 ( .A(n4139), .Z(n348) );
  XOR U1012 ( .A(n4543), .B(n4535), .Z(n4154) );
  MUX U1013 ( .IN0(n4166), .IN1(n349), .SEL(n4167), .F(n4141) );
  IV U1014 ( .A(n4168), .Z(n349) );
  MUX U1015 ( .IN0(n5079), .IN1(n5089), .SEL(n5081), .F(n3123) );
  MUX U1016 ( .IN0(n3208), .IN1(n3206), .SEL(n3207), .F(n3169) );
  MUX U1017 ( .IN0(n350), .IN1(n3148), .SEL(n3149), .F(n3019) );
  IV U1018 ( .A(n3150), .Z(n350) );
  MUX U1019 ( .IN0(n351), .IN1(n3910), .SEL(n3274), .F(n3893) );
  IV U1020 ( .A(n3272), .Z(n351) );
  MUX U1021 ( .IN0(n352), .IN1(n3090), .SEL(n3091), .F(n2955) );
  IV U1022 ( .A(n3092), .Z(n352) );
  MUX U1023 ( .IN0(n353), .IN1(n3036), .SEL(n3037), .F(n2900) );
  IV U1024 ( .A(n3038), .Z(n353) );
  XOR U1025 ( .A(n3874), .B(n3875), .Z(n3891) );
  MUX U1026 ( .IN0(n4701), .IN1(n354), .SEL(n4702), .F(n3086) );
  IV U1027 ( .A(n4703), .Z(n354) );
  MUX U1028 ( .IN0(n4336), .IN1(n355), .SEL(n4335), .F(n4326) );
  IV U1029 ( .A(n4334), .Z(n355) );
  XOR U1030 ( .A(n3221), .B(n3157), .Z(n3161) );
  MUX U1031 ( .IN0(n356), .IN1(n2776), .SEL(n2777), .F(n2650) );
  IV U1032 ( .A(n2778), .Z(n356) );
  MUX U1033 ( .IN0(n357), .IN1(n2842), .SEL(n2843), .F(n2710) );
  IV U1034 ( .A(n2844), .Z(n357) );
  MUX U1035 ( .IN0(n358), .IN1(n2625), .SEL(n2626), .F(n2499) );
  IV U1036 ( .A(n2627), .Z(n358) );
  MUX U1037 ( .IN0(n359), .IN1(n2701), .SEL(n2702), .F(n2574) );
  IV U1038 ( .A(n2703), .Z(n359) );
  MUX U1039 ( .IN0(n360), .IN1(n2591), .SEL(n2592), .F(n2467) );
  IV U1040 ( .A(n2593), .Z(n360) );
  MUX U1041 ( .IN0(n361), .IN1(n2395), .SEL(n2396), .F(n2280) );
  IV U1042 ( .A(n2397), .Z(n361) );
  MUX U1043 ( .IN0(n362), .IN1(n2434), .SEL(n2435), .F(n2313) );
  IV U1044 ( .A(n2436), .Z(n362) );
  MUX U1045 ( .IN0(n363), .IN1(n2288), .SEL(n2289), .F(n2176) );
  IV U1046 ( .A(n2290), .Z(n363) );
  MUX U1047 ( .IN0(n364), .IN1(n2213), .SEL(n2214), .F(n2102) );
  IV U1048 ( .A(n2215), .Z(n364) );
  MUX U1049 ( .IN0(n365), .IN1(n2119), .SEL(n2120), .F(n2014) );
  IV U1050 ( .A(n2121), .Z(n365) );
  MUX U1051 ( .IN0(n366), .IN1(n1973), .SEL(n1974), .F(n1868) );
  IV U1052 ( .A(n1975), .Z(n366) );
  MUX U1053 ( .IN0(n367), .IN1(n1776), .SEL(n1777), .F(n1680) );
  IV U1054 ( .A(n1778), .Z(n367) );
  MUX U1055 ( .IN0(n368), .IN1(n1488), .SEL(n1489), .F(n1403) );
  IV U1056 ( .A(n1490), .Z(n368) );
  MUX U1057 ( .IN0(n369), .IN1(n1605), .SEL(n1606), .F(n1517) );
  IV U1058 ( .A(n1607), .Z(n369) );
  MUX U1059 ( .IN0(n370), .IN1(n1411), .SEL(n1412), .F(n1339) );
  IV U1060 ( .A(n1413), .Z(n370) );
  MUX U1061 ( .IN0(n371), .IN1(n1436), .SEL(n1437), .F(n1359) );
  IV U1062 ( .A(n1438), .Z(n371) );
  MUX U1063 ( .IN0(n372), .IN1(n1305), .SEL(n1306), .F(n1235) );
  IV U1064 ( .A(n1307), .Z(n372) );
  MUX U1065 ( .IN0(n373), .IN1(n1152), .SEL(n1153), .F(n1090) );
  IV U1066 ( .A(n1154), .Z(n373) );
  MUX U1067 ( .IN0(n374), .IN1(n1160), .SEL(n1161), .F(n1098) );
  IV U1068 ( .A(n1162), .Z(n374) );
  MUX U1069 ( .IN0(n375), .IN1(n1048), .SEL(n1049), .F(n992) );
  IV U1070 ( .A(n1050), .Z(n375) );
  MUX U1071 ( .IN0(n376), .IN1(n1001), .SEL(n1002), .F(n943) );
  IV U1072 ( .A(n1003), .Z(n376) );
  XNOR U1073 ( .A(n5157), .B(n3133), .Z(n3137) );
  XNOR U1074 ( .A(n3179), .B(n3054), .Z(n3058) );
  MUX U1075 ( .IN0(n2975), .IN1(n2977), .SEL(n2976), .F(n2837) );
  XOR U1076 ( .A(n2486), .B(n2608), .Z(n2487) );
  MUX U1077 ( .IN0(n2454), .IN1(n2456), .SEL(n2455), .F(n2333) );
  MUX U1078 ( .IN0(n377), .IN1(n2666), .SEL(n2667), .F(n2539) );
  IV U1079 ( .A(n2668), .Z(n377) );
  MUX U1080 ( .IN0(n2350), .IN1(n2352), .SEL(n2351), .F(n2234) );
  MUX U1081 ( .IN0(n2277), .IN1(n378), .SEL(n2276), .F(n2162) );
  IV U1082 ( .A(n2275), .Z(n378) );
  MUX U1083 ( .IN0(n379), .IN1(n2151), .SEL(n2152), .F(n2048) );
  IV U1084 ( .A(n2153), .Z(n379) );
  MUX U1085 ( .IN0(n2001), .IN1(n2003), .SEL(n2002), .F(n1896) );
  MUX U1086 ( .IN0(n1913), .IN1(n1915), .SEL(n1914), .F(n1813) );
  XOR U1087 ( .A(n1641), .B(n1732), .Z(n1642) );
  MUX U1088 ( .IN0(n1609), .IN1(n1611), .SEL(n1610), .F(n1511) );
  MUX U1089 ( .IN0(n1113), .IN1(n1111), .SEL(n1112), .F(n1052) );
  MUX U1090 ( .IN0(n1043), .IN1(n1045), .SEL(n1044), .F(n987) );
  MUX U1091 ( .IN0(n1134), .IN1(n380), .SEL(n1133), .F(n1076) );
  IV U1092 ( .A(n1132), .Z(n380) );
  MUX U1093 ( .IN0(n927), .IN1(n381), .SEL(n926), .F(n887) );
  IV U1094 ( .A(n925), .Z(n381) );
  MUX U1095 ( .IN0(n897), .IN1(n895), .SEL(n896), .F(n851) );
  MUX U1096 ( .IN0(n382), .IN1(n847), .SEL(n848), .F(n807) );
  IV U1097 ( .A(n849), .Z(n382) );
  MUX U1098 ( .IN0(n383), .IN1(n3022), .SEL(n3023), .F(n2886) );
  IV U1099 ( .A(n3024), .Z(n383) );
  XOR U1100 ( .A(n2986), .B(n2851), .Z(n2855) );
  XNOR U1101 ( .A(n2766), .B(n2643), .Z(n2647) );
  XOR U1102 ( .A(n2757), .B(n2634), .Z(n2638) );
  NAND U1103 ( .A(n2662), .B(n2791), .Z(n2790) );
  MUX U1104 ( .IN0(n2828), .IN1(n384), .SEL(n2829), .F(n2696) );
  IV U1105 ( .A(n2830), .Z(n384) );
  XNOR U1106 ( .A(n2807), .B(n2678), .Z(n2682) );
  XNOR U1107 ( .A(n2857), .B(n2728), .Z(n2732) );
  XNOR U1108 ( .A(n2474), .B(n2356), .Z(n2360) );
  MUX U1109 ( .IN0(n385), .IN1(n2265), .SEL(n2266), .F(n2154) );
  IV U1110 ( .A(n2267), .Z(n385) );
  MUX U1111 ( .IN0(n2324), .IN1(n386), .SEL(n2325), .F(n2208) );
  IV U1112 ( .A(n2326), .Z(n386) );
  XNOR U1113 ( .A(n2303), .B(n2190), .Z(n2194) );
  MUX U1114 ( .IN0(n387), .IN1(n2225), .SEL(n2226), .F(n2114) );
  IV U1115 ( .A(n2227), .Z(n387) );
  XNOR U1116 ( .A(n2057), .B(n1955), .Z(n1959) );
  XNOR U1117 ( .A(n2021), .B(n1919), .Z(n1923) );
  MUX U1118 ( .IN0(n1887), .IN1(n388), .SEL(n1888), .F(n1787) );
  IV U1119 ( .A(n1889), .Z(n388) );
  XNOR U1120 ( .A(n1766), .B(n1673), .Z(n1677) );
  XOR U1121 ( .A(n1620), .B(n1531), .Z(n1535) );
  XNOR U1122 ( .A(n1629), .B(n1540), .Z(n1544) );
  MUX U1123 ( .IN0(n1507), .IN1(n389), .SEL(n1508), .F(n1422) );
  IV U1124 ( .A(n1509), .Z(n389) );
  XNOR U1125 ( .A(n1329), .B(n1262), .Z(n1266) );
  XOR U1126 ( .A(n1365), .B(n1297), .Z(n1301) );
  MUX U1127 ( .IN0(n390), .IN1(n1221), .SEL(n1222), .F(n1155) );
  IV U1128 ( .A(n1223), .Z(n390) );
  MUX U1129 ( .IN0(n391), .IN1(n1080), .SEL(n1081), .F(n1021) );
  IV U1130 ( .A(n1082), .Z(n391) );
  MUX U1131 ( .IN0(n392), .IN1(n921), .SEL(n922), .F(n878) );
  IV U1132 ( .A(n923), .Z(n392) );
  MUX U1133 ( .IN0(n393), .IN1(n2958), .SEL(n2959), .F(n2820) );
  IV U1134 ( .A(n2960), .Z(n393) );
  XNOR U1135 ( .A(n2865), .B(n2864), .Z(n2847) );
  XNOR U1136 ( .A(n2803), .B(n2931), .Z(n2804) );
  MUX U1137 ( .IN0(n394), .IN1(n2437), .SEL(n2438), .F(n2316) );
  IV U1138 ( .A(n2439), .Z(n394) );
  XNOR U1139 ( .A(n1849), .B(n1848), .Z(n1842) );
  MUX U1140 ( .IN0(n395), .IN1(n1779), .SEL(n1780), .F(n1683) );
  IV U1141 ( .A(n1781), .Z(n395) );
  MUX U1142 ( .IN0(n1657), .IN1(n1655), .SEL(n1656), .F(n1572) );
  MUX U1143 ( .IN0(n396), .IN1(n1414), .SEL(n1415), .F(n1342) );
  IV U1144 ( .A(n1416), .Z(n396) );
  NANDN U1145 ( .B(n1214), .A(n1215), .Z(n1209) );
  MUX U1146 ( .IN0(n397), .IN1(n969), .SEL(n970), .F(n913) );
  IV U1147 ( .A(n971), .Z(n397) );
  XOR U1148 ( .A(n761), .B(n799), .Z(n792) );
  MUX U1149 ( .IN0(n2653), .IN1(n398), .SEL(n2654), .F(n2529) );
  IV U1150 ( .A(n2655), .Z(n398) );
  XNOR U1151 ( .A(n2420), .B(n2414), .Z(n2532) );
  ANDN U1152 ( .A(n2368), .B(n2369), .Z(n2252) );
  MUX U1153 ( .IN0(n2179), .IN1(n399), .SEL(n2180), .F(n2070) );
  IV U1154 ( .A(n2181), .Z(n399) );
  NANDN U1155 ( .B(n2073), .A(n2074), .Z(n1968) );
  ANDN U1156 ( .A(n1931), .B(n1932), .Z(n1831) );
  ANDN U1157 ( .A(n1318), .B(n1319), .Z(n1248) );
  OR U1158 ( .A(n738), .B(n739), .Z(n733) );
  MUX U1159 ( .IN0(n400), .IN1(n743), .SEL(n744), .F(n711) );
  IV U1160 ( .A(n745), .Z(n400) );
  XNOR U1161 ( .A(n1986), .B(n1985), .Z(n1967) );
  XOR U1162 ( .A(n1667), .B(n1664), .Z(n1745) );
  XNOR U1163 ( .A(n1594), .B(n1593), .Z(n1577) );
  OR U1164 ( .A(n1256), .B(n1257), .Z(n1189) );
  XNOR U1165 ( .A(n1085), .B(n1084), .Z(n1069) );
  XNOR U1166 ( .A(n1026), .B(n1025), .Z(n1013) );
  OR U1167 ( .A(n868), .B(n869), .Z(n828) );
  AND U1168 ( .A(n903), .B(n904), .Z(n859) );
  XNOR U1169 ( .A(n791), .B(n790), .Z(n789) );
  AND U1170 ( .A(n746), .B(n747), .Z(n714) );
  ANDN U1171 ( .A(n683), .B(n682), .Z(n678) );
  MUX U1172 ( .IN0(n401), .IN1(n2740), .SEL(n695), .F(n2615) );
  IV U1173 ( .A(\_MxM/Y0[3] ), .Z(n401) );
  MUX U1174 ( .IN0(n2254), .IN1(n402), .SEL(n654), .F(n2143) );
  IV U1175 ( .A(\_MxM/Y0[7] ), .Z(n402) );
  MUX U1176 ( .IN0(n1833), .IN1(n403), .SEL(n1834), .F(n1739) );
  IV U1177 ( .A(\_MxM/Y0[11] ), .Z(n403) );
  MUX U1178 ( .IN0(n1468), .IN1(n404), .SEL(n1469), .F(n1391) );
  IV U1179 ( .A(\_MxM/Y0[15] ), .Z(n404) );
  MUX U1180 ( .IN0(n405), .IN1(n1183), .SEL(n1184), .F(n1121) );
  IV U1181 ( .A(\_MxM/Y0[19] ), .Z(n405) );
  MUX U1182 ( .IN0(n406), .IN1(n948), .SEL(n949), .F(n905) );
  IV U1183 ( .A(\_MxM/Y0[23] ), .Z(n406) );
  XNOR U1184 ( .A(n716), .B(n717), .Z(n694) );
  OR U1185 ( .A(n700), .B(n701), .Z(n671) );
  MUX U1186 ( .IN0(n407), .IN1(n3742), .SEL(n3743), .F(n3704) );
  IV U1187 ( .A(n3744), .Z(n407) );
  XOR U1188 ( .A(n3753), .B(n3718), .Z(n3722) );
  MUX U1189 ( .IN0(n408), .IN1(n3590), .SEL(n3591), .F(n3552) );
  IV U1190 ( .A(n3592), .Z(n408) );
  MUX U1191 ( .IN0(n3626), .IN1(n3624), .SEL(n3625), .F(n3586) );
  MUX U1192 ( .IN0(n409), .IN1(n3582), .SEL(n3583), .F(n3544) );
  IV U1193 ( .A(n3584), .Z(n409) );
  MUX U1194 ( .IN0(n410), .IN1(n4060), .SEL(n4061), .F(n4043) );
  IV U1195 ( .A(n4062), .Z(n410) );
  MUX U1196 ( .IN0(n411), .IN1(n4052), .SEL(n4053), .F(n4035) );
  IV U1197 ( .A(n4054), .Z(n411) );
  MUX U1198 ( .IN0(n412), .IN1(n3595), .SEL(n3596), .F(n3557) );
  IV U1199 ( .A(n3597), .Z(n412) );
  MUX U1200 ( .IN0(n3674), .IN1(n413), .SEL(n3675), .F(n3636) );
  IV U1201 ( .A(n3676), .Z(n413) );
  MUX U1202 ( .IN0(n4484), .IN1(n414), .SEL(n4083), .F(n4471) );
  IV U1203 ( .A(n4082), .Z(n414) );
  MUX U1204 ( .IN0(n415), .IN1(n4480), .SEL(n4481), .F(n4467) );
  IV U1205 ( .A(n4482), .Z(n415) );
  XOR U1206 ( .A(n3639), .B(n3604), .Z(n3608) );
  MUX U1207 ( .IN0(n416), .IN1(n4460), .SEL(n4461), .F(n4447) );
  IV U1208 ( .A(n4462), .Z(n416) );
  MUX U1209 ( .IN0(n417), .IN1(n4063), .SEL(n3616), .F(n4046) );
  IV U1210 ( .A(n3614), .Z(n417) );
  MUX U1211 ( .IN0(n4024), .IN1(n4022), .SEL(n4023), .F(n4005) );
  MUX U1212 ( .IN0(n418), .IN1(n4850), .SEL(n4851), .F(n4829) );
  IV U1213 ( .A(n4852), .Z(n418) );
  MUX U1214 ( .IN0(n419), .IN1(n4855), .SEL(n4856), .F(n4834) );
  IV U1215 ( .A(n4857), .Z(n419) );
  MUX U1216 ( .IN0(n3474), .IN1(n3472), .SEL(n3473), .F(n3434) );
  MUX U1217 ( .IN0(n420), .IN1(n3430), .SEL(n3431), .F(n3392) );
  IV U1218 ( .A(n3432), .Z(n420) );
  MUX U1219 ( .IN0(n421), .IN1(n3992), .SEL(n3993), .F(n3975) );
  IV U1220 ( .A(n3994), .Z(n421) );
  MUX U1221 ( .IN0(n422), .IN1(n3984), .SEL(n3985), .F(n3967) );
  IV U1222 ( .A(n3986), .Z(n422) );
  MUX U1223 ( .IN0(n423), .IN1(n3443), .SEL(n3444), .F(n3405) );
  IV U1224 ( .A(n3445), .Z(n423) );
  MUX U1225 ( .IN0(n3522), .IN1(n424), .SEL(n3523), .F(n3484) );
  IV U1226 ( .A(n3524), .Z(n424) );
  MUX U1227 ( .IN0(n425), .IN1(n4262), .SEL(n4263), .F(n4241) );
  IV U1228 ( .A(n4264), .Z(n425) );
  XOR U1229 ( .A(n4609), .B(n4601), .Z(n4280) );
  MUX U1230 ( .IN0(n426), .IN1(n4267), .SEL(n4268), .F(n4246) );
  IV U1231 ( .A(n4269), .Z(n426) );
  MUX U1232 ( .IN0(n4432), .IN1(n427), .SEL(n4015), .F(n4419) );
  IV U1233 ( .A(n4014), .Z(n427) );
  XOR U1234 ( .A(n3487), .B(n3452), .Z(n3456) );
  MUX U1235 ( .IN0(n428), .IN1(n4408), .SEL(n4409), .F(n4395) );
  IV U1236 ( .A(n4410), .Z(n428) );
  MUX U1237 ( .IN0(n429), .IN1(n3362), .SEL(n3363), .F(n3324) );
  IV U1238 ( .A(n3364), .Z(n429) );
  MUX U1239 ( .IN0(n430), .IN1(n4415), .SEL(n4416), .F(n4402) );
  IV U1240 ( .A(n4417), .Z(n430) );
  MUX U1241 ( .IN0(n431), .IN1(n3995), .SEL(n3464), .F(n3978) );
  IV U1242 ( .A(n3462), .Z(n431) );
  MUX U1243 ( .IN0(n432), .IN1(n3375), .SEL(n3376), .F(n3337) );
  IV U1244 ( .A(n3377), .Z(n432) );
  XOR U1245 ( .A(n4953), .B(n4945), .Z(n4805) );
  MUX U1246 ( .IN0(n3956), .IN1(n3954), .SEL(n3955), .F(n3937) );
  XNOR U1247 ( .A(n3352), .B(n3317), .Z(n3321) );
  XOR U1248 ( .A(n4576), .B(n4568), .Z(n4217) );
  MUX U1249 ( .IN0(n4229), .IN1(n433), .SEL(n4230), .F(n4208) );
  IV U1250 ( .A(n4231), .Z(n433) );
  XOR U1251 ( .A(n4811), .B(n4793), .Z(n4797) );
  XOR U1252 ( .A(n4767), .B(n4768), .Z(n4777) );
  MUX U1253 ( .IN0(n434), .IN1(n3916), .SEL(n3917), .F(n3899) );
  IV U1254 ( .A(n3918), .Z(n434) );
  MUX U1255 ( .IN0(n435), .IN1(n3291), .SEL(n3292), .F(n3253) );
  IV U1256 ( .A(n3293), .Z(n435) );
  MUX U1257 ( .IN0(n3370), .IN1(n436), .SEL(n3371), .F(n3332) );
  IV U1258 ( .A(n3372), .Z(n436) );
  MUX U1259 ( .IN0(n3809), .IN1(n3823), .SEL(n3811), .F(n3793) );
  MUX U1260 ( .IN0(n437), .IN1(n4178), .SEL(n4179), .F(n4157) );
  IV U1261 ( .A(n4180), .Z(n437) );
  MUX U1262 ( .IN0(n4640), .IN1(n4655), .SEL(n4642), .F(n4617) );
  MUX U1263 ( .IN0(n4634), .IN1(n4649), .SEL(n4636), .F(n4623) );
  MUX U1264 ( .IN0(n438), .IN1(n4551), .SEL(n4552), .F(n4540) );
  IV U1265 ( .A(n4553), .Z(n438) );
  MUX U1266 ( .IN0(n439), .IN1(n4183), .SEL(n4184), .F(n4162) );
  IV U1267 ( .A(n4185), .Z(n439) );
  MUX U1268 ( .IN0(n4380), .IN1(n440), .SEL(n3947), .F(n4367) );
  IV U1269 ( .A(n3946), .Z(n440) );
  MUX U1270 ( .IN0(n5110), .IN1(n5125), .SEL(n5112), .F(n5092) );
  MUX U1271 ( .IN0(n5012), .IN1(n5027), .SEL(n5014), .F(n4989) );
  MUX U1272 ( .IN0(n5006), .IN1(n5021), .SEL(n5008), .F(n4995) );
  XOR U1273 ( .A(n4925), .B(n4926), .Z(n4782) );
  XOR U1274 ( .A(n4746), .B(n4747), .Z(n4756) );
  MUX U1275 ( .IN0(n441), .IN1(n4750), .SEL(n4751), .F(n4729) );
  IV U1276 ( .A(n4752), .Z(n441) );
  XNOR U1277 ( .A(n3284), .B(n3283), .Z(n3296) );
  MUX U1278 ( .IN0(n3787), .IN1(n3802), .SEL(n3789), .F(n3776) );
  XNOR U1279 ( .A(n4687), .B(n4688), .Z(n4674) );
  MUX U1280 ( .IN0(n442), .IN1(n4545), .SEL(n4546), .F(n4534) );
  IV U1281 ( .A(n4547), .Z(n442) );
  MUX U1282 ( .IN0(n443), .IN1(n4356), .SEL(n4357), .F(n4343) );
  IV U1283 ( .A(n4358), .Z(n443) );
  NOR U1284 ( .A(g_input[0]), .B(n5177), .Z(n5170) );
  MUX U1285 ( .IN0(n5098), .IN1(n5115), .SEL(n5100), .F(n5069) );
  XNOR U1286 ( .A(n5059), .B(n5060), .Z(n5046) );
  XOR U1287 ( .A(n4912), .B(n4913), .Z(n4761) );
  MUX U1288 ( .IN0(n444), .IN1(n4905), .SEL(n4906), .F(n4892) );
  IV U1289 ( .A(n4907), .Z(n444) );
  MUX U1290 ( .IN0(n445), .IN1(n4363), .SEL(n4364), .F(n4350) );
  IV U1291 ( .A(n4365), .Z(n445) );
  MUX U1292 ( .IN0(n446), .IN1(n3927), .SEL(n3312), .F(n3910) );
  IV U1293 ( .A(n3310), .Z(n446) );
  XNOR U1294 ( .A(n3246), .B(n3245), .Z(n3258) );
  XNOR U1295 ( .A(n3841), .B(n3842), .Z(n3827) );
  XNOR U1296 ( .A(n4306), .B(n4307), .Z(n4292) );
  MUX U1297 ( .IN0(n5161), .IN1(n5164), .SEL(n5162), .F(n3132) );
  XNOR U1298 ( .A(n5149), .B(n5150), .Z(n5136) );
  XNOR U1299 ( .A(n4873), .B(n4874), .Z(n4859) );
  XOR U1300 ( .A(n4899), .B(n4900), .Z(n4740) );
  MUX U1301 ( .IN0(n447), .IN1(n4705), .SEL(n4706), .F(n3090) );
  IV U1302 ( .A(n4707), .Z(n447) );
  MUX U1303 ( .IN0(n448), .IN1(n3189), .SEL(n3190), .F(n3061) );
  IV U1304 ( .A(n3191), .Z(n448) );
  XOR U1305 ( .A(n3259), .B(n3224), .Z(n3228) );
  XNOR U1306 ( .A(n3208), .B(n3207), .Z(n3220) );
  MUX U1307 ( .IN0(n4141), .IN1(n449), .SEL(n4142), .F(n4124) );
  IV U1308 ( .A(n4143), .Z(n449) );
  MUX U1309 ( .IN0(n4538), .IN1(n450), .SEL(n4154), .F(n4525) );
  IV U1310 ( .A(n4152), .Z(n450) );
  MUX U1311 ( .IN0(n451), .IN1(n3019), .SEL(n3020), .F(n2883) );
  IV U1312 ( .A(n3021), .Z(n451) );
  XNOR U1313 ( .A(n3877), .B(n3182), .Z(n3186) );
  XNOR U1314 ( .A(n3171), .B(n3170), .Z(n3153) );
  XNOR U1315 ( .A(n3849), .B(n3735), .Z(n3739) );
  MUX U1316 ( .IN0(n452), .IN1(n2963), .SEL(n2964), .F(n2825) );
  IV U1317 ( .A(n2965), .Z(n452) );
  MUX U1318 ( .IN0(n453), .IN1(n2988), .SEL(n2989), .F(n2850) );
  IV U1319 ( .A(n2990), .Z(n453) );
  MUX U1320 ( .IN0(n454), .IN1(n2900), .SEL(n2901), .F(n2768) );
  IV U1321 ( .A(n2902), .Z(n454) );
  MUX U1322 ( .IN0(n455), .IN1(n2633), .SEL(n2634), .F(n2507) );
  IV U1323 ( .A(n2635), .Z(n455) );
  MUX U1324 ( .IN0(n456), .IN1(n2650), .SEL(n2651), .F(n2526) );
  IV U1325 ( .A(n2652), .Z(n456) );
  MUX U1326 ( .IN0(n457), .IN1(n2710), .SEL(n2711), .F(n2583) );
  IV U1327 ( .A(n2712), .Z(n457) );
  MUX U1328 ( .IN0(n458), .IN1(n2499), .SEL(n2500), .F(n2378) );
  IV U1329 ( .A(n2501), .Z(n458) );
  MUX U1330 ( .IN0(n459), .IN1(n2600), .SEL(n2601), .F(n2476) );
  IV U1331 ( .A(n2602), .Z(n459) );
  MUX U1332 ( .IN0(n460), .IN1(n2442), .SEL(n2443), .F(n2321) );
  IV U1333 ( .A(n2444), .Z(n460) );
  MUX U1334 ( .IN0(n461), .IN1(n2313), .SEL(n2314), .F(n2197) );
  IV U1335 ( .A(n2315), .Z(n461) );
  MUX U1336 ( .IN0(n462), .IN1(n2176), .SEL(n2177), .F(n2067) );
  IV U1337 ( .A(n2178), .Z(n462) );
  MUX U1338 ( .IN0(n463), .IN1(n2222), .SEL(n2223), .F(n2111) );
  IV U1339 ( .A(n2224), .Z(n463) );
  MUX U1340 ( .IN0(n464), .IN1(n1989), .SEL(n1990), .F(n1884) );
  IV U1341 ( .A(n1991), .Z(n464) );
  MUX U1342 ( .IN0(n465), .IN1(n1892), .SEL(n1893), .F(n1792) );
  IV U1343 ( .A(n1894), .Z(n465) );
  MUX U1344 ( .IN0(n466), .IN1(n1876), .SEL(n1877), .F(n1776) );
  IV U1345 ( .A(n1878), .Z(n466) );
  MUX U1346 ( .IN0(n467), .IN1(n1801), .SEL(n1802), .F(n1705) );
  IV U1347 ( .A(n1803), .Z(n467) );
  MUX U1348 ( .IN0(n468), .IN1(n1722), .SEL(n1723), .F(n1631) );
  IV U1349 ( .A(n1724), .Z(n468) );
  MUX U1350 ( .IN0(n469), .IN1(n1597), .SEL(n1598), .F(n1504) );
  IV U1351 ( .A(n1599), .Z(n469) );
  MUX U1352 ( .IN0(n470), .IN1(n1622), .SEL(n1623), .F(n1530) );
  IV U1353 ( .A(n1624), .Z(n470) );
  MUX U1354 ( .IN0(n471), .IN1(n1496), .SEL(n1497), .F(n1411) );
  IV U1355 ( .A(n1498), .Z(n471) );
  MUX U1356 ( .IN0(n472), .IN1(n1296), .SEL(n1297), .F(n1226) );
  IV U1357 ( .A(n1298), .Z(n472) );
  MUX U1358 ( .IN0(n473), .IN1(n974), .SEL(n975), .F(n918) );
  IV U1359 ( .A(n976), .Z(n473) );
  MUX U1360 ( .IN0(n474), .IN1(n943), .SEL(n944), .F(n900) );
  IV U1361 ( .A(n945), .Z(n474) );
  MUX U1362 ( .IN0(n475), .IN1(n983), .SEL(n984), .F(n925) );
  IV U1363 ( .A(n985), .Z(n475) );
  MUX U1364 ( .IN0(n3127), .IN1(n3129), .SEL(n3128), .F(n2992) );
  MUX U1365 ( .IN0(n3891), .IN1(n4327), .SEL(n3892), .F(n476) );
  XNOR U1366 ( .A(n4695), .B(n3083), .Z(n3087) );
  MUX U1367 ( .IN0(n3073), .IN1(n477), .SEL(n3072), .F(n2935) );
  IV U1368 ( .A(n3071), .Z(n477) );
  MUX U1369 ( .IN0(n2664), .IN1(n2784), .SEL(n2663), .F(n2533) );
  XOR U1370 ( .A(n2033), .B(n2136), .Z(n2034) );
  MUX U1371 ( .IN0(n1700), .IN1(n1702), .SEL(n1701), .F(n1609) );
  XOR U1372 ( .A(n1463), .B(n1547), .Z(n1464) );
  MUX U1373 ( .IN0(n1519), .IN1(n478), .SEL(n1518), .F(n1430) );
  IV U1374 ( .A(n1517), .Z(n478) );
  MUX U1375 ( .IN0(n1448), .IN1(n1450), .SEL(n1449), .F(n1371) );
  MUX U1376 ( .IN0(n1201), .IN1(n1199), .SEL(n1200), .F(n1137) );
  MUX U1377 ( .IN0(n1164), .IN1(n1166), .SEL(n1165), .F(n1102) );
  MUX U1378 ( .IN0(n883), .IN1(n885), .SEL(n884), .F(n842) );
  XOR U1379 ( .A(n3104), .B(n2972), .Z(n2976) );
  XOR U1380 ( .A(n3025), .B(n2892), .Z(n2896) );
  MUX U1381 ( .IN0(n479), .IN1(n3074), .SEL(n3075), .F(n2941) );
  IV U1382 ( .A(n3076), .Z(n479) );
  XNOR U1383 ( .A(n3138), .B(n3137), .Z(n3120) );
  XNOR U1384 ( .A(n3042), .B(n3041), .Z(n3024) );
  XNOR U1385 ( .A(n2995), .B(n2860), .Z(n2864) );
  XNOR U1386 ( .A(n2640), .B(n2517), .Z(n2523) );
  XOR U1387 ( .A(n2716), .B(n2592), .Z(n2596) );
  XNOR U1388 ( .A(n2675), .B(n2551), .Z(n2555) );
  XOR U1389 ( .A(n2699), .B(n2575), .Z(n2579) );
  MUX U1390 ( .IN0(n2445), .IN1(n480), .SEL(n2446), .F(n2324) );
  IV U1391 ( .A(n2447), .Z(n480) );
  MUX U1392 ( .IN0(n2541), .IN1(n481), .SEL(n2540), .F(n2416) );
  IV U1393 ( .A(n2539), .Z(n481) );
  NAND U1394 ( .A(n2162), .B(n2273), .Z(n2272) );
  XNOR U1395 ( .A(n2278), .B(n2169), .Z(n2173) );
  XOR U1396 ( .A(n2327), .B(n2214), .Z(n2218) );
  XOR U1397 ( .A(n2344), .B(n2231), .Z(n2235) );
  XNOR U1398 ( .A(n2187), .B(n2079), .Z(n2083) );
  XNOR U1399 ( .A(n2126), .B(n2024), .Z(n2028) );
  MUX U1400 ( .IN0(n2050), .IN1(n482), .SEL(n2049), .F(n1943) );
  IV U1401 ( .A(n2048), .Z(n482) );
  XNOR U1402 ( .A(n1952), .B(n1854), .Z(n1848) );
  XOR U1403 ( .A(n2012), .B(n1910), .Z(n1914) );
  MUX U1404 ( .IN0(n1992), .IN1(n483), .SEL(n1993), .F(n1887) );
  IV U1405 ( .A(n1994), .Z(n483) );
  XNOR U1406 ( .A(n1866), .B(n1769), .Z(n1773) );
  MUX U1407 ( .IN0(n1600), .IN1(n484), .SEL(n1601), .F(n1507) );
  IV U1408 ( .A(n1602), .Z(n484) );
  MUX U1409 ( .IN0(n485), .IN1(n1757), .SEL(n1758), .F(n1661) );
  IV U1410 ( .A(n1759), .Z(n485) );
  XNOR U1411 ( .A(n1486), .B(n1404), .Z(n1408) );
  XNOR U1412 ( .A(n1537), .B(n1454), .Z(n1458) );
  XNOR U1413 ( .A(n1303), .B(n1236), .Z(n1240) );
  OR U1414 ( .A(n1276), .B(n1277), .Z(n1214) );
  XNOR U1415 ( .A(n1105), .B(n1049), .Z(n1053) );
  XNOR U1416 ( .A(n932), .B(n892), .Z(n896) );
  XNOR U1417 ( .A(n2953), .B(n2952), .Z(n2968) );
  XNOR U1418 ( .A(n2906), .B(n2905), .Z(n2888) );
  XNOR U1419 ( .A(n2789), .B(n2788), .Z(n2805) );
  MUX U1420 ( .IN0(n2673), .IN1(n486), .SEL(n2672), .F(n2544) );
  IV U1421 ( .A(n2671), .Z(n486) );
  XNOR U1422 ( .A(n2606), .B(n2605), .Z(n2588) );
  XNOR U1423 ( .A(n2245), .B(n2244), .Z(n2227) );
  XNOR U1424 ( .A(n1924), .B(n1923), .Z(n1906) );
  XNOR U1425 ( .A(n1337), .B(n1336), .Z(n1354) );
  XNOR U1426 ( .A(n1382), .B(n1381), .Z(n1364) );
  XNOR U1427 ( .A(n1267), .B(n1266), .Z(n1285) );
  XNOR U1428 ( .A(n1175), .B(n1174), .Z(n1157) );
  NOR U1429 ( .A(n1027), .B(n1028), .Z(n960) );
  XNOR U1430 ( .A(n998), .B(n997), .Z(n979) );
  ANDN U1431 ( .A(n965), .B(n964), .Z(n963) );
  XNOR U1432 ( .A(n853), .B(n852), .Z(n841) );
  XNOR U1433 ( .A(n813), .B(n812), .Z(n803) );
  XNOR U1434 ( .A(n2985), .B(n2984), .Z(n2960) );
  MUX U1435 ( .IN0(n2779), .IN1(n487), .SEL(n2780), .F(n2653) );
  IV U1436 ( .A(n2781), .Z(n487) );
  XNOR U1437 ( .A(n2715), .B(n2714), .Z(n2690) );
  XNOR U1438 ( .A(n2383), .B(n2382), .Z(n2422) );
  XNOR U1439 ( .A(n2464), .B(n2463), .Z(n2439) );
  XNOR U1440 ( .A(n2343), .B(n2342), .Z(n2318) );
  ANDN U1441 ( .A(n2489), .B(n2490), .Z(n2368) );
  XNOR U1442 ( .A(n2116), .B(n2115), .Z(n2091) );
  XNOR U1443 ( .A(n1806), .B(n1805), .Z(n1781) );
  ANDN U1444 ( .A(n1480), .B(n1481), .Z(n1478) );
  XNOR U1445 ( .A(n1293), .B(n1292), .Z(n1274) );
  XNOR U1446 ( .A(n1095), .B(n1094), .Z(n1085) );
  XNOR U1447 ( .A(n923), .B(n922), .Z(n915) );
  XOR U1448 ( .A(n2073), .B(n2070), .Z(n2148) );
  XOR U1449 ( .A(n1763), .B(n1760), .Z(n1839) );
  XNOR U1450 ( .A(n1685), .B(n1684), .Z(n1666) );
  XNOR U1451 ( .A(n1501), .B(n1500), .Z(n1484) );
  MUX U1452 ( .IN0(n488), .IN1(n861), .SEL(n862), .F(n821) );
  IV U1453 ( .A(\_MxM/Y0[25] ), .Z(n488) );
  XNOR U1454 ( .A(n760), .B(n757), .Z(n756) );
  MUX U1455 ( .IN0(n708), .IN1(n706), .SEL(n707), .F(n686) );
  AND U1456 ( .A(n714), .B(n715), .Z(n669) );
  XOR U1457 ( .A(n1190), .B(n1189), .Z(n1253) );
  XNOR U1458 ( .A(n1013), .B(n1012), .Z(n1065) );
  XNOR U1459 ( .A(n869), .B(n868), .Z(n908) );
  ANDN U1460 ( .A(n672), .B(n671), .Z(n665) );
  MUX U1461 ( .IN0(\_MxM/Y0[30] ), .IN1(n694), .SEL(n693), .F(n661) );
  XOR U1462 ( .A(n2615), .B(n2618), .Z(n2616) );
  XOR U1463 ( .A(n2254), .B(n2257), .Z(n2255) );
  XOR U1464 ( .A(n1933), .B(n1936), .Z(n1934) );
  XOR U1465 ( .A(n1646), .B(n1650), .Z(n1648) );
  XOR U1466 ( .A(n1391), .B(n1395), .Z(n1393) );
  XOR U1467 ( .A(n1183), .B(n1187), .Z(n1185) );
  XOR U1468 ( .A(n1006), .B(n1010), .Z(n1008) );
  MUX U1469 ( .IN0(n489), .IN1(n3704), .SEL(n3705), .F(n3666) );
  IV U1470 ( .A(n3706), .Z(n489) );
  XOR U1471 ( .A(n4500), .B(n4501), .Z(n4116) );
  MUX U1472 ( .IN0(n490), .IN1(n4086), .SEL(n4087), .F(n4069) );
  IV U1473 ( .A(n4088), .Z(n490) );
  MUX U1474 ( .IN0(n491), .IN1(n3671), .SEL(n3672), .F(n3633) );
  IV U1475 ( .A(n3673), .Z(n491) );
  MUX U1476 ( .IN0(n492), .IN1(n4097), .SEL(n3692), .F(n4080) );
  IV U1477 ( .A(n3690), .Z(n492) );
  XNOR U1478 ( .A(n3618), .B(n3583), .Z(n3587) );
  MUX U1479 ( .IN0(n493), .IN1(n4473), .SEL(n4474), .F(n4460) );
  IV U1480 ( .A(n4475), .Z(n493) );
  MUX U1481 ( .IN0(n494), .IN1(n3552), .SEL(n3553), .F(n3514) );
  IV U1482 ( .A(n3554), .Z(n494) );
  MUX U1483 ( .IN0(n4058), .IN1(n4056), .SEL(n4057), .F(n4039) );
  MUX U1484 ( .IN0(n3607), .IN1(n3609), .SEL(n3608), .F(n3569) );
  MUX U1485 ( .IN0(n495), .IN1(n3565), .SEL(n3566), .F(n3527) );
  IV U1486 ( .A(n3567), .Z(n495) );
  MUX U1487 ( .IN0(n496), .IN1(n4467), .SEL(n4468), .F(n4454) );
  IV U1488 ( .A(n4469), .Z(n496) );
  MUX U1489 ( .IN0(n497), .IN1(n4026), .SEL(n4027), .F(n4009) );
  IV U1490 ( .A(n4028), .Z(n497) );
  MUX U1491 ( .IN0(n498), .IN1(n4018), .SEL(n4019), .F(n4001) );
  IV U1492 ( .A(n4020), .Z(n498) );
  MUX U1493 ( .IN0(n499), .IN1(n3519), .SEL(n3520), .F(n3481) );
  IV U1494 ( .A(n3521), .Z(n499) );
  MUX U1495 ( .IN0(n4458), .IN1(n500), .SEL(n4049), .F(n4445) );
  IV U1496 ( .A(n4048), .Z(n500) );
  MUX U1497 ( .IN0(n3560), .IN1(n501), .SEL(n3561), .F(n3522) );
  IV U1498 ( .A(n3562), .Z(n501) );
  MUX U1499 ( .IN0(n502), .IN1(n4029), .SEL(n3540), .F(n4012) );
  IV U1500 ( .A(n3538), .Z(n502) );
  XNOR U1501 ( .A(n3466), .B(n3431), .Z(n3435) );
  XOR U1502 ( .A(n4263), .B(n4264), .Z(n4273) );
  MUX U1503 ( .IN0(n503), .IN1(n4421), .SEL(n4422), .F(n4408) );
  IV U1504 ( .A(n4423), .Z(n503) );
  MUX U1505 ( .IN0(n504), .IN1(n3400), .SEL(n3401), .F(n3362) );
  IV U1506 ( .A(n3402), .Z(n504) );
  MUX U1507 ( .IN0(n3990), .IN1(n3988), .SEL(n3989), .F(n3971) );
  MUX U1508 ( .IN0(n3455), .IN1(n3457), .SEL(n3456), .F(n3417) );
  MUX U1509 ( .IN0(n505), .IN1(n3413), .SEL(n3414), .F(n3375) );
  IV U1510 ( .A(n3415), .Z(n505) );
  XOR U1511 ( .A(n4596), .B(n4597), .Z(n4278) );
  MUX U1512 ( .IN0(n506), .IN1(n4246), .SEL(n4247), .F(n4225) );
  IV U1513 ( .A(n4248), .Z(n506) );
  XOR U1514 ( .A(n4964), .B(n4965), .Z(n4845) );
  MUX U1515 ( .IN0(n507), .IN1(n4808), .SEL(n4809), .F(n4787) );
  IV U1516 ( .A(n4810), .Z(n507) );
  MUX U1517 ( .IN0(n508), .IN1(n3958), .SEL(n3959), .F(n3941) );
  IV U1518 ( .A(n3960), .Z(n508) );
  MUX U1519 ( .IN0(n509), .IN1(n3950), .SEL(n3951), .F(n3933) );
  IV U1520 ( .A(n3952), .Z(n509) );
  MUX U1521 ( .IN0(n510), .IN1(n3367), .SEL(n3368), .F(n3329) );
  IV U1522 ( .A(n3369), .Z(n510) );
  MUX U1523 ( .IN0(n511), .IN1(n4220), .SEL(n4221), .F(n4199) );
  IV U1524 ( .A(n4222), .Z(n511) );
  MUX U1525 ( .IN0(n512), .IN1(n4573), .SEL(n4574), .F(n4562) );
  IV U1526 ( .A(n4575), .Z(n512) );
  MUX U1527 ( .IN0(n4406), .IN1(n513), .SEL(n3981), .F(n4393) );
  IV U1528 ( .A(n3980), .Z(n513) );
  XOR U1529 ( .A(n4951), .B(n4952), .Z(n4824) );
  MUX U1530 ( .IN0(n514), .IN1(n4944), .SEL(n4945), .F(n4931) );
  IV U1531 ( .A(n4946), .Z(n514) );
  MUX U1532 ( .IN0(n515), .IN1(n4402), .SEL(n4403), .F(n4389) );
  IV U1533 ( .A(n4404), .Z(n515) );
  MUX U1534 ( .IN0(n3408), .IN1(n516), .SEL(n3409), .F(n3370) );
  IV U1535 ( .A(n3410), .Z(n516) );
  XOR U1536 ( .A(n4938), .B(n4939), .Z(n4803) );
  MUX U1537 ( .IN0(n3322), .IN1(n3320), .SEL(n3321), .F(n3282) );
  MUX U1538 ( .IN0(n517), .IN1(n3278), .SEL(n3279), .F(n3240) );
  IV U1539 ( .A(n3280), .Z(n517) );
  MUX U1540 ( .IN0(n518), .IN1(n3961), .SEL(n3388), .F(n3944) );
  IV U1541 ( .A(n3386), .Z(n518) );
  MUX U1542 ( .IN0(n4682), .IN1(n4685), .SEL(n4683), .F(n4666) );
  XOR U1543 ( .A(n4565), .B(n4557), .Z(n4196) );
  XOR U1544 ( .A(n4357), .B(n4358), .Z(n3929) );
  MUX U1545 ( .IN0(n519), .IN1(n5148), .SEL(n5149), .F(n5144) );
  IV U1546 ( .A(n5150), .Z(n519) );
  MUX U1547 ( .IN0(n5054), .IN1(n5057), .SEL(n5055), .F(n5038) );
  XOR U1548 ( .A(n4790), .B(n4772), .Z(n4776) );
  MUX U1549 ( .IN0(n520), .IN1(n4911), .SEL(n4912), .F(n4898) );
  IV U1550 ( .A(n4913), .Z(n520) );
  MUX U1551 ( .IN0(n3922), .IN1(n3920), .SEL(n3921), .F(n3903) );
  MUX U1552 ( .IN0(n3303), .IN1(n3305), .SEL(n3304), .F(n3265) );
  MUX U1553 ( .IN0(n521), .IN1(n3261), .SEL(n3262), .F(n3223) );
  IV U1554 ( .A(n3263), .Z(n521) );
  MUX U1555 ( .IN0(n3793), .IN1(n3808), .SEL(n3795), .F(n3768) );
  MUX U1556 ( .IN0(n3836), .IN1(n3839), .SEL(n3837), .F(n3819) );
  MUX U1557 ( .IN0(n4623), .IN1(n4633), .SEL(n4625), .F(n4611) );
  XOR U1558 ( .A(n4202), .B(n4184), .Z(n4188) );
  XOR U1559 ( .A(n4344), .B(n4345), .Z(n3912) );
  MUX U1560 ( .IN0(n5092), .IN1(n5107), .SEL(n5094), .F(n5079) );
  MUX U1561 ( .IN0(n4995), .IN1(n5005), .SEL(n4997), .F(n4983) );
  MUX U1562 ( .IN0(n522), .IN1(n4724), .SEL(n4725), .F(n4705) );
  IV U1563 ( .A(n4726), .Z(n522) );
  MUX U1564 ( .IN0(n523), .IN1(n3879), .SEL(n3880), .F(n3181) );
  IV U1565 ( .A(n3881), .Z(n523) );
  MUX U1566 ( .IN0(n524), .IN1(n3215), .SEL(n3216), .F(n3148) );
  IV U1567 ( .A(n3217), .Z(n524) );
  MUX U1568 ( .IN0(n3851), .IN1(n3854), .SEL(n3852), .F(n3734) );
  MUX U1569 ( .IN0(n525), .IN1(n4145), .SEL(n4146), .F(n4128) );
  IV U1570 ( .A(n4147), .Z(n525) );
  XOR U1571 ( .A(n4672), .B(n4673), .Z(n4319) );
  MUX U1572 ( .IN0(n526), .IN1(n4534), .SEL(n4535), .F(n4521) );
  IV U1573 ( .A(n4536), .Z(n526) );
  XOR U1574 ( .A(n4541), .B(n4542), .Z(n4173) );
  XOR U1575 ( .A(n5044), .B(n5045), .Z(n4886) );
  MUX U1576 ( .IN0(n4909), .IN1(n527), .SEL(n4742), .F(n4896) );
  IV U1577 ( .A(n4740), .Z(n527) );
  MUX U1578 ( .IN0(n528), .IN1(n4892), .SEL(n4893), .F(n3106) );
  IV U1579 ( .A(n4894), .Z(n528) );
  MUX U1580 ( .IN0(n529), .IN1(n3173), .SEL(n3174), .F(n3044) );
  IV U1581 ( .A(n3175), .Z(n529) );
  MUX U1582 ( .IN0(n530), .IN1(n4350), .SEL(n4351), .F(n4334) );
  IV U1583 ( .A(n4352), .Z(n530) );
  XNOR U1584 ( .A(n3200), .B(n3166), .Z(n3170) );
  MUX U1585 ( .IN0(n3256), .IN1(n531), .SEL(n3257), .F(n3218) );
  IV U1586 ( .A(n3258), .Z(n531) );
  XOR U1587 ( .A(n3825), .B(n3826), .Z(n3772) );
  XNOR U1588 ( .A(n4299), .B(n4289), .Z(n4293) );
  XOR U1589 ( .A(n4607), .B(n4608), .Z(n4297) );
  XOR U1590 ( .A(n4530), .B(n4531), .Z(n4152) );
  XOR U1591 ( .A(n5159), .B(g_input[3]), .Z(n5160) );
  MUX U1592 ( .IN0(n532), .IN1(n3115), .SEL(n3116), .F(n2980) );
  IV U1593 ( .A(n3117), .Z(n532) );
  MUX U1594 ( .IN0(n533), .IN1(n3061), .SEL(n3062), .F(n2925) );
  IV U1595 ( .A(n3063), .Z(n533) );
  XNOR U1596 ( .A(n5166), .B(n5167), .Z(n3136) );
  XOR U1597 ( .A(n5134), .B(n5135), .Z(n5073) );
  XNOR U1598 ( .A(n4866), .B(n4856), .Z(n4860) );
  XOR U1599 ( .A(n4977), .B(n4978), .Z(n4864) );
  XOR U1600 ( .A(n4727), .B(n4698), .Z(n4702) );
  MUX U1601 ( .IN0(n534), .IN1(n3893), .SEL(n3236), .F(n3876) );
  IV U1602 ( .A(n3234), .Z(n534) );
  XOR U1603 ( .A(n3774), .B(n3756), .Z(n3760) );
  XNOR U1604 ( .A(n4135), .B(n4121), .Z(n4125) );
  XOR U1605 ( .A(n4515), .B(n4516), .Z(n4133) );
  MUX U1606 ( .IN0(n535), .IN1(n2997), .SEL(n2998), .F(n2859) );
  IV U1607 ( .A(n2999), .Z(n535) );
  MUX U1608 ( .IN0(n536), .IN1(n2891), .SEL(n2892), .F(n2759) );
  IV U1609 ( .A(n2893), .Z(n536) );
  MUX U1610 ( .IN0(n537), .IN1(n3873), .SEL(n3874), .F(n3071) );
  IV U1611 ( .A(n3875), .Z(n537) );
  MUX U1612 ( .IN0(n538), .IN1(n2751), .SEL(n2752), .F(n2625) );
  IV U1613 ( .A(n2753), .Z(n538) );
  MUX U1614 ( .IN0(n539), .IN1(n2825), .SEL(n2826), .F(n2693) );
  IV U1615 ( .A(n2827), .Z(n539) );
  MUX U1616 ( .IN0(n540), .IN1(n2809), .SEL(n2810), .F(n2677) );
  IV U1617 ( .A(n2811), .Z(n540) );
  MUX U1618 ( .IN0(n541), .IN1(n2526), .SEL(n2527), .F(n2403) );
  IV U1619 ( .A(n2528), .Z(n541) );
  MUX U1620 ( .IN0(n542), .IN1(n2583), .SEL(n2584), .F(n2459) );
  IV U1621 ( .A(n2585), .Z(n542) );
  MUX U1622 ( .IN0(n543), .IN1(n2476), .SEL(n2477), .F(n2355) );
  IV U1623 ( .A(n2478), .Z(n543) );
  MUX U1624 ( .IN0(n544), .IN1(n2321), .SEL(n2322), .F(n2205) );
  IV U1625 ( .A(n2323), .Z(n544) );
  MUX U1626 ( .IN0(n545), .IN1(n2305), .SEL(n2306), .F(n2189) );
  IV U1627 ( .A(n2307), .Z(n545) );
  MUX U1628 ( .IN0(n546), .IN1(n2067), .SEL(n2068), .F(n1962) );
  IV U1629 ( .A(n2069), .Z(n546) );
  MUX U1630 ( .IN0(n547), .IN1(n2111), .SEL(n2112), .F(n2006) );
  IV U1631 ( .A(n2113), .Z(n547) );
  MUX U1632 ( .IN0(n548), .IN1(n2262), .SEL(n2263), .F(n2151) );
  IV U1633 ( .A(n2264), .Z(n548) );
  MUX U1634 ( .IN0(n549), .IN1(n2023), .SEL(n2024), .F(n1918) );
  IV U1635 ( .A(n2025), .Z(n549) );
  MUX U1636 ( .IN0(n550), .IN1(n1884), .SEL(n1885), .F(n1784) );
  IV U1637 ( .A(n1886), .Z(n550) );
  MUX U1638 ( .IN0(n551), .IN1(n1909), .SEL(n1910), .F(n1809) );
  IV U1639 ( .A(n1911), .Z(n551) );
  MUX U1640 ( .IN0(n552), .IN1(n1705), .SEL(n1706), .F(n1614) );
  IV U1641 ( .A(n1707), .Z(n552) );
  MUX U1642 ( .IN0(n553), .IN1(n1680), .SEL(n1681), .F(n1589) );
  IV U1643 ( .A(n1682), .Z(n553) );
  MUX U1644 ( .IN0(n554), .IN1(n1631), .SEL(n1632), .F(n1539) );
  IV U1645 ( .A(n1633), .Z(n554) );
  MUX U1646 ( .IN0(n555), .IN1(n1504), .SEL(n1505), .F(n1419) );
  IV U1647 ( .A(n1506), .Z(n555) );
  MUX U1648 ( .IN0(n556), .IN1(n1339), .SEL(n1340), .F(n1269) );
  IV U1649 ( .A(n1341), .Z(n556) );
  MUX U1650 ( .IN0(n557), .IN1(n1359), .SEL(n1360), .F(n1288) );
  IV U1651 ( .A(n1361), .Z(n557) );
  MUX U1652 ( .IN0(n558), .IN1(n1090), .SEL(n1091), .F(n1031) );
  IV U1653 ( .A(n1092), .Z(n558) );
  MUX U1654 ( .IN0(n559), .IN1(n1057), .SEL(n1058), .F(n1001) );
  IV U1655 ( .A(n1059), .Z(n559) );
  MUX U1656 ( .IN0(n3031), .IN1(n3033), .SEL(n3032), .F(n2895) );
  XNOR U1657 ( .A(n3740), .B(n3739), .Z(n3752) );
  XOR U1658 ( .A(n2737), .B(n2867), .Z(n2738) );
  MUX U1659 ( .IN0(n2361), .IN1(n2359), .SEL(n2360), .F(n2243) );
  MUX U1660 ( .IN0(n560), .IN1(n875), .SEL(n876), .F(n836) );
  IV U1661 ( .A(n877), .Z(n560) );
  XOR U1662 ( .A(n3121), .B(n2989), .Z(n2993) );
  XNOR U1663 ( .A(n3051), .B(n2918), .Z(n2922) );
  XNOR U1664 ( .A(n3088), .B(n3087), .Z(n3103) );
  XOR U1665 ( .A(n2969), .B(n2834), .Z(n2838) );
  XNOR U1666 ( .A(n2898), .B(n2769), .Z(n2773) );
  MUX U1667 ( .IN0(n561), .IN1(n2886), .SEL(n2887), .F(n2754) );
  IV U1668 ( .A(n2888), .Z(n561) );
  XOR U1669 ( .A(n2667), .B(n2668), .Z(n2664) );
  XOR U1670 ( .A(n2631), .B(n2508), .Z(n2512) );
  XOR U1671 ( .A(n2540), .B(n2541), .Z(n2535) );
  XNOR U1672 ( .A(n2514), .B(n2396), .Z(n2400) );
  XOR U1673 ( .A(n2572), .B(n2451), .Z(n2455) );
  XOR U1674 ( .A(n2589), .B(n2468), .Z(n2472) );
  MUX U1675 ( .IN0(n2154), .IN1(n562), .SEL(n2155), .F(n2051) );
  IV U1676 ( .A(n2156), .Z(n562) );
  XNOR U1677 ( .A(n2166), .B(n2060), .Z(n2064) );
  XOR U1678 ( .A(n2228), .B(n2120), .Z(n2124) );
  XOR U1679 ( .A(n2211), .B(n2103), .Z(n2107) );
  MUX U1680 ( .IN0(n2056), .IN1(n2054), .SEL(n2055), .F(n563) );
  IV U1681 ( .A(n563), .Z(n1948) );
  XNOR U1682 ( .A(n2076), .B(n1974), .Z(n1978) );
  XOR U1683 ( .A(n1890), .B(n1793), .Z(n1797) );
  XOR U1684 ( .A(n1711), .B(n1623), .Z(n1627) );
  XNOR U1685 ( .A(n1670), .B(n1582), .Z(n1586) );
  XOR U1686 ( .A(n1603), .B(n1518), .Z(n1512) );
  MUX U1687 ( .IN0(n1755), .IN1(n1844), .SEL(n1754), .F(n1655) );
  XNOR U1688 ( .A(n1401), .B(n1332), .Z(n1336) );
  XNOR U1689 ( .A(n1451), .B(n1377), .Z(n1381) );
  XOR U1690 ( .A(n1442), .B(n1368), .Z(n1372) );
  XOR U1691 ( .A(n1224), .B(n1161), .Z(n1165) );
  XNOR U1692 ( .A(n1233), .B(n1170), .Z(n1174) );
  XNOR U1693 ( .A(n1192), .B(n1133), .Z(n1138) );
  XOR U1694 ( .A(n1037), .B(n984), .Z(n988) );
  XNOR U1695 ( .A(n1046), .B(n993), .Z(n997) );
  OR U1696 ( .A(n887), .B(n888), .Z(n881) );
  XNOR U1697 ( .A(n889), .B(n848), .Z(n852) );
  MUX U1698 ( .IN0(n564), .IN1(n3064), .SEL(n3065), .F(n2928) );
  IV U1699 ( .A(n3066), .Z(n564) );
  XNOR U1700 ( .A(n3120), .B(n3119), .Z(n3095) );
  XNOR U1701 ( .A(n2815), .B(n2814), .Z(n2830) );
  MUX U1702 ( .IN0(n2805), .IN1(n2803), .SEL(n2804), .F(n565) );
  IV U1703 ( .A(n565), .Z(n2670) );
  XNOR U1704 ( .A(n2556), .B(n2555), .Z(n2571) );
  XNOR U1705 ( .A(n2432), .B(n2431), .Z(n2447) );
  XNOR U1706 ( .A(n2482), .B(n2481), .Z(n2464) );
  XNOR U1707 ( .A(n2195), .B(n2194), .Z(n2210) );
  XNOR U1708 ( .A(n2134), .B(n2133), .Z(n2116) );
  XNOR U1709 ( .A(n2084), .B(n2083), .Z(n2099) );
  XNOR U1710 ( .A(n1874), .B(n1873), .Z(n1889) );
  XNOR U1711 ( .A(n1774), .B(n1773), .Z(n1789) );
  XNOR U1712 ( .A(n1824), .B(n1823), .Z(n1806) );
  XNOR U1713 ( .A(n1637), .B(n1636), .Z(n1619) );
  XNOR U1714 ( .A(n1545), .B(n1544), .Z(n1527) );
  MUX U1715 ( .IN0(n566), .IN1(n1661), .SEL(n1662), .F(n1574) );
  IV U1716 ( .A(n1663), .Z(n566) );
  XOR U1717 ( .A(n1276), .B(n1283), .Z(n1345) );
  XNOR U1718 ( .A(n1311), .B(n1310), .Z(n1293) );
  XNOR U1719 ( .A(n1201), .B(n1200), .Z(n1213) );
  XNOR U1720 ( .A(n1113), .B(n1112), .Z(n1095) );
  AND U1721 ( .A(n966), .B(n967), .Z(n962) );
  XNOR U1722 ( .A(n940), .B(n939), .Z(n923) );
  MUX U1723 ( .IN0(n763), .IN1(n761), .SEL(n762), .F(n729) );
  MUX U1724 ( .IN0(n768), .IN1(n567), .SEL(n767), .F(n738) );
  IV U1725 ( .A(n766), .Z(n567) );
  MUX U1726 ( .IN0(n568), .IN1(n776), .SEL(n777), .F(n743) );
  IV U1727 ( .A(n778), .Z(n568) );
  XNOR U1728 ( .A(n2847), .B(n2846), .Z(n2822) );
  MUX U1729 ( .IN0(n2911), .IN1(n569), .SEL(n2912), .F(n2779) );
  IV U1730 ( .A(n2913), .Z(n569) );
  XNOR U1731 ( .A(n2630), .B(n2629), .Z(n2673) );
  XNOR U1732 ( .A(n2588), .B(n2587), .Z(n2563) );
  XNOR U1733 ( .A(n2295), .B(n2409), .Z(n2296) );
  XNOR U1734 ( .A(n2227), .B(n2226), .Z(n2202) );
  XNOR U1735 ( .A(n2011), .B(n2010), .Z(n1986) );
  XNOR U1736 ( .A(n1906), .B(n1905), .Z(n1881) );
  XNOR U1737 ( .A(n1710), .B(n1709), .Z(n1685) );
  ANDN U1738 ( .A(n1737), .B(n1738), .Z(n1644) );
  XNOR U1739 ( .A(n1441), .B(n1440), .Z(n1416) );
  XNOR U1740 ( .A(n1223), .B(n1222), .Z(n1208) );
  XOR U1741 ( .A(n1027), .B(n1024), .Z(n1070) );
  XNOR U1742 ( .A(n880), .B(n879), .Z(n871) );
  XNOR U1743 ( .A(n803), .B(n802), .Z(n791) );
  XNOR U1744 ( .A(n2690), .B(n2689), .Z(n2655) );
  XNOR U1745 ( .A(n2318), .B(n2317), .Z(n2293) );
  XOR U1746 ( .A(n1863), .B(n1860), .Z(n1938) );
  XOR U1747 ( .A(n1561), .B(n1575), .Z(n1652) );
  MUX U1748 ( .IN0(n570), .IN1(n821), .SEL(n822), .F(n781) );
  IV U1749 ( .A(\_MxM/Y0[26] ), .Z(n570) );
  ANDN U1750 ( .A(n687), .B(n686), .Z(n685) );
  XNOR U1751 ( .A(n681), .B(n680), .Z(n672) );
  MUX U1752 ( .IN0(n3010), .IN1(n571), .SEL(n3011), .F(n2872) );
  IV U1753 ( .A(\_MxM/Y0[1] ), .Z(n571) );
  XOR U1754 ( .A(n1327), .B(n1326), .Z(n1394) );
  XNOR U1755 ( .A(n1129), .B(n1128), .Z(n1186) );
  XNOR U1756 ( .A(n955), .B(n954), .Z(n1009) );
  XNOR U1757 ( .A(n829), .B(n828), .Z(n865) );
  XNOR U1758 ( .A(n756), .B(n755), .Z(n785) );
  XNOR U1759 ( .A(n701), .B(n700), .Z(n722) );
  XOR U1760 ( .A(n2491), .B(n2494), .Z(n2492) );
  XOR U1761 ( .A(n2143), .B(n2146), .Z(n2144) );
  XOR U1762 ( .A(n1833), .B(n1837), .Z(n1835) );
  XOR U1763 ( .A(n1554), .B(n1558), .Z(n1556) );
  XOR U1764 ( .A(n1320), .B(n1324), .Z(n1322) );
  XOR U1765 ( .A(n1121), .B(n1126), .Z(n1124) );
  XOR U1766 ( .A(n948), .B(n952), .Z(n950) );
  MUX U1767 ( .IN0(\_MxM/Y0[31] ), .IN1(n661), .SEL(n662), .F(n658) );
  MUX U1768 ( .IN0(n572), .IN1(n3696), .SEL(n3697), .F(n3658) );
  IV U1769 ( .A(n3698), .Z(n572) );
  MUX U1770 ( .IN0(n3721), .IN1(n3723), .SEL(n3722), .F(n3683) );
  XNOR U1771 ( .A(n3702), .B(n3701), .Z(n3714) );
  XNOR U1772 ( .A(n4109), .B(n4108), .Z(n3728) );
  MUX U1773 ( .IN0(n573), .IN1(n4069), .SEL(n4070), .F(n4052) );
  IV U1774 ( .A(n4071), .Z(n573) );
  MUX U1775 ( .IN0(n574), .IN1(n3633), .SEL(n3634), .F(n3595) );
  IV U1776 ( .A(n3635), .Z(n574) );
  MUX U1777 ( .IN0(n575), .IN1(n3641), .SEL(n3642), .F(n3603) );
  IV U1778 ( .A(n3643), .Z(n575) );
  XNOR U1779 ( .A(n3664), .B(n3663), .Z(n3676) );
  XNOR U1780 ( .A(n4092), .B(n4091), .Z(n3690) );
  XNOR U1781 ( .A(n3626), .B(n3625), .Z(n3638) );
  MUX U1782 ( .IN0(n576), .IN1(n3544), .SEL(n3545), .F(n3506) );
  IV U1783 ( .A(n3546), .Z(n576) );
  XNOR U1784 ( .A(n4075), .B(n4074), .Z(n3652) );
  XNOR U1785 ( .A(n3588), .B(n3587), .Z(n3600) );
  MUX U1786 ( .IN0(n4471), .IN1(n577), .SEL(n4066), .F(n4458) );
  IV U1787 ( .A(n4065), .Z(n577) );
  XNOR U1788 ( .A(n4058), .B(n4057), .Z(n3614) );
  MUX U1789 ( .IN0(n3569), .IN1(n3571), .SEL(n3570), .F(n3531) );
  XNOR U1790 ( .A(n3550), .B(n3549), .Z(n3562) );
  MUX U1791 ( .IN0(n578), .IN1(n4454), .SEL(n4455), .F(n4441) );
  IV U1792 ( .A(n4456), .Z(n578) );
  XNOR U1793 ( .A(n4041), .B(n4040), .Z(n3576) );
  MUX U1794 ( .IN0(n579), .IN1(n4001), .SEL(n4002), .F(n3984) );
  IV U1795 ( .A(n4003), .Z(n579) );
  MUX U1796 ( .IN0(n580), .IN1(n3481), .SEL(n3482), .F(n3443) );
  IV U1797 ( .A(n3483), .Z(n580) );
  MUX U1798 ( .IN0(n581), .IN1(n3489), .SEL(n3490), .F(n3451) );
  IV U1799 ( .A(n3491), .Z(n581) );
  XNOR U1800 ( .A(n3512), .B(n3511), .Z(n3524) );
  MUX U1801 ( .IN0(n582), .IN1(n4434), .SEL(n4435), .F(n4421) );
  IV U1802 ( .A(n4436), .Z(n582) );
  XNOR U1803 ( .A(n4024), .B(n4023), .Z(n3538) );
  XNOR U1804 ( .A(n3474), .B(n3473), .Z(n3486) );
  XOR U1805 ( .A(n4424), .B(n4416), .Z(n3998) );
  MUX U1806 ( .IN0(n583), .IN1(n4829), .SEL(n4830), .F(n4808) );
  IV U1807 ( .A(n4831), .Z(n583) );
  MUX U1808 ( .IN0(n584), .IN1(n3392), .SEL(n3393), .F(n3354) );
  IV U1809 ( .A(n3394), .Z(n584) );
  XNOR U1810 ( .A(n4007), .B(n4006), .Z(n3500) );
  XNOR U1811 ( .A(n3436), .B(n3435), .Z(n3448) );
  MUX U1812 ( .IN0(n585), .IN1(n4241), .SEL(n4242), .F(n4220) );
  IV U1813 ( .A(n4243), .Z(n585) );
  XOR U1814 ( .A(n4396), .B(n4397), .Z(n3980) );
  XNOR U1815 ( .A(n3990), .B(n3989), .Z(n3462) );
  MUX U1816 ( .IN0(n3417), .IN1(n3419), .SEL(n3418), .F(n3379) );
  XNOR U1817 ( .A(n3398), .B(n3397), .Z(n3410) );
  XOR U1818 ( .A(n4585), .B(n4586), .Z(n4257) );
  XOR U1819 ( .A(n4383), .B(n4384), .Z(n3963) );
  XOR U1820 ( .A(n4832), .B(n4814), .Z(n4818) );
  MUX U1821 ( .IN0(n586), .IN1(n4937), .SEL(n4938), .F(n4924) );
  IV U1822 ( .A(n4939), .Z(n586) );
  XNOR U1823 ( .A(n3973), .B(n3972), .Z(n3424) );
  MUX U1824 ( .IN0(n587), .IN1(n3933), .SEL(n3934), .F(n3916) );
  IV U1825 ( .A(n3935), .Z(n587) );
  MUX U1826 ( .IN0(n588), .IN1(n3329), .SEL(n3330), .F(n3291) );
  IV U1827 ( .A(n3331), .Z(n588) );
  MUX U1828 ( .IN0(n589), .IN1(n3337), .SEL(n3338), .F(n3299) );
  IV U1829 ( .A(n3339), .Z(n589) );
  XNOR U1830 ( .A(n3360), .B(n3359), .Z(n3372) );
  XOR U1831 ( .A(n4574), .B(n4575), .Z(n4236) );
  MUX U1832 ( .IN0(n590), .IN1(n3286), .SEL(n3287), .F(n3248) );
  IV U1833 ( .A(n3288), .Z(n590) );
  MUX U1834 ( .IN0(n591), .IN1(n4389), .SEL(n4390), .F(n4376) );
  IV U1835 ( .A(n4391), .Z(n591) );
  XNOR U1836 ( .A(n3956), .B(n3955), .Z(n3386) );
  XNOR U1837 ( .A(n3322), .B(n3321), .Z(n3334) );
  XNOR U1838 ( .A(n3314), .B(n3279), .Z(n3283) );
  MUX U1839 ( .IN0(n592), .IN1(n4556), .SEL(n4557), .F(n4545) );
  IV U1840 ( .A(n4558), .Z(n592) );
  XOR U1841 ( .A(n4223), .B(n4205), .Z(n4209) );
  MUX U1842 ( .IN0(n5116), .IN1(n5132), .SEL(n5118), .F(n5098) );
  MUX U1843 ( .IN0(n4935), .IN1(n593), .SEL(n4784), .F(n4922) );
  IV U1844 ( .A(n4782), .Z(n593) );
  MUX U1845 ( .IN0(n594), .IN1(n4918), .SEL(n4919), .F(n4905) );
  IV U1846 ( .A(n4920), .Z(n594) );
  MUX U1847 ( .IN0(n595), .IN1(n4745), .SEL(n4746), .F(n4724) );
  IV U1848 ( .A(n4747), .Z(n595) );
  XNOR U1849 ( .A(n3939), .B(n3938), .Z(n3348) );
  MUX U1850 ( .IN0(n596), .IN1(n4157), .SEL(n4158), .F(n4145) );
  IV U1851 ( .A(n4159), .Z(n596) );
  MUX U1852 ( .IN0(n4301), .IN1(n4304), .SEL(n4302), .F(n4288) );
  MUX U1853 ( .IN0(n4617), .IN1(n4639), .SEL(n4619), .F(n4606) );
  XOR U1854 ( .A(n4552), .B(n4553), .Z(n4194) );
  XOR U1855 ( .A(n4359), .B(n4351), .Z(n3913) );
  MUX U1856 ( .IN0(n4868), .IN1(n4871), .SEL(n4869), .F(n4855) );
  MUX U1857 ( .IN0(n4989), .IN1(n5011), .SEL(n4991), .F(n4976) );
  XOR U1858 ( .A(n4769), .B(n4751), .Z(n4755) );
  MUX U1859 ( .IN0(n597), .IN1(n3202), .SEL(n3203), .F(n3165) );
  IV U1860 ( .A(n3204), .Z(n597) );
  XNOR U1861 ( .A(n3922), .B(n3921), .Z(n3310) );
  MUX U1862 ( .IN0(n3265), .IN1(n3267), .SEL(n3266), .F(n3227) );
  MUX U1863 ( .IN0(n3768), .IN1(n3792), .SEL(n3770), .F(n3747) );
  MUX U1864 ( .IN0(n3776), .IN1(n3786), .SEL(n3778), .F(n3755) );
  XOR U1865 ( .A(n4680), .B(n4667), .Z(n4320) );
  MUX U1866 ( .IN0(n598), .IN1(n4529), .SEL(n4530), .F(n4514) );
  IV U1867 ( .A(n4531), .Z(n598) );
  MUX U1868 ( .IN0(n599), .IN1(n4343), .SEL(n4344), .F(n4338) );
  IV U1869 ( .A(n4345), .Z(n599) );
  MUX U1870 ( .IN0(g_input[1]), .IN1(n5177), .SEL(g_input[31]), .F(n3828) );
  XOR U1871 ( .A(n5052), .B(n5039), .Z(n4887) );
  MUX U1872 ( .IN0(n600), .IN1(n4712), .SEL(n4713), .F(n3098) );
  IV U1873 ( .A(n4714), .Z(n600) );
  MUX U1874 ( .IN0(n601), .IN1(n4697), .SEL(n4698), .F(n3082) );
  IV U1875 ( .A(n4699), .Z(n601) );
  MUX U1876 ( .IN0(n602), .IN1(n3156), .SEL(n3157), .F(n3027) );
  IV U1877 ( .A(n3158), .Z(n602) );
  MUX U1878 ( .IN0(n603), .IN1(n3181), .SEL(n3182), .F(n3053) );
  IV U1879 ( .A(n3183), .Z(n603) );
  MUX U1880 ( .IN0(e_input[1]), .IN1(n604), .SEL(e_input[31]), .F(n4324) );
  IV U1881 ( .A(n4693), .Z(n604) );
  XNOR U1882 ( .A(n3905), .B(n3904), .Z(n3272) );
  XOR U1883 ( .A(n3834), .B(n3820), .Z(n3773) );
  XNOR U1884 ( .A(n3856), .B(n3857), .Z(n3738) );
  XOR U1885 ( .A(n4621), .B(n4612), .Z(n4298) );
  XOR U1886 ( .A(n4160), .B(n4138), .Z(n4142) );
  MUX U1887 ( .IN0(g_input[2]), .IN1(n5169), .SEL(g_input[31]), .F(n3139) );
  MUX U1888 ( .IN0(n605), .IN1(n3044), .SEL(n3045), .F(n2908) );
  IV U1889 ( .A(n3046), .Z(n605) );
  XOR U1890 ( .A(n5142), .B(n5129), .Z(n5074) );
  XOR U1891 ( .A(n4993), .B(n4984), .Z(n4865) );
  MUX U1892 ( .IN0(n3171), .IN1(n3169), .SEL(n3170), .F(n3040) );
  XNOR U1893 ( .A(n3885), .B(n3884), .Z(n3234) );
  MUX U1894 ( .IN0(n3218), .IN1(n606), .SEL(n3219), .F(n3151) );
  IV U1895 ( .A(n3220), .Z(n606) );
  XNOR U1896 ( .A(n4294), .B(n4293), .Z(n3869) );
  XOR U1897 ( .A(n4532), .B(n4522), .Z(n4134) );
  MUX U1898 ( .IN0(n607), .IN1(n2955), .SEL(n2956), .F(n2817) );
  IV U1899 ( .A(n2957), .Z(n607) );
  MUX U1900 ( .IN0(n608), .IN1(n2980), .SEL(n2981), .F(n2842) );
  IV U1901 ( .A(n2982), .Z(n608) );
  MUX U1902 ( .IN0(g_input[3]), .IN1(n5160), .SEL(g_input[31]), .F(n609) );
  IV U1903 ( .A(n609), .Z(n3004) );
  MUX U1904 ( .IN0(n610), .IN1(n2883), .SEL(n2884), .F(n2751) );
  IV U1905 ( .A(n2885), .Z(n610) );
  MUX U1906 ( .IN0(n611), .IN1(n2768), .SEL(n2769), .F(n2642) );
  IV U1907 ( .A(n2770), .Z(n611) );
  MUX U1908 ( .IN0(e_input[4]), .IN1(n4312), .SEL(e_input[31]), .F(n2792) );
  MUX U1909 ( .IN0(g_input[4]), .IN1(n5126), .SEL(g_input[31]), .F(n612) );
  IV U1910 ( .A(n612), .Z(n2866) );
  MUX U1911 ( .IN0(n613), .IN1(n2859), .SEL(n2860), .F(n2727) );
  IV U1912 ( .A(n2861), .Z(n613) );
  MUX U1913 ( .IN0(g_input[5]), .IN1(n5109), .SEL(g_input[31]), .F(n2734) );
  MUX U1914 ( .IN0(n614), .IN1(n2677), .SEL(n2678), .F(n2550) );
  IV U1915 ( .A(n2679), .Z(n614) );
  MUX U1916 ( .IN0(n615), .IN1(n2693), .SEL(n2694), .F(n2566) );
  IV U1917 ( .A(n2695), .Z(n615) );
  MUX U1918 ( .IN0(g_input[6]), .IN1(n5090), .SEL(g_input[31]), .F(n2607) );
  MUX U1919 ( .IN0(n616), .IN1(n2378), .SEL(n2379), .F(n2262) );
  IV U1920 ( .A(n2380), .Z(n616) );
  MUX U1921 ( .IN0(n617), .IN1(n2459), .SEL(n2460), .F(n2338) );
  IV U1922 ( .A(n2461), .Z(n617) );
  MUX U1923 ( .IN0(g_input[7]), .IN1(n5078), .SEL(g_input[31]), .F(n2483) );
  MUX U1924 ( .IN0(n618), .IN1(n2797), .SEL(n2798), .F(n2666) );
  IV U1925 ( .A(n2799), .Z(n618) );
  MUX U1926 ( .IN0(e_input[8]), .IN1(n3847), .SEL(e_input[31]), .F(n2274) );
  MUX U1927 ( .IN0(n619), .IN1(n2280), .SEL(n2281), .F(n2168) );
  IV U1928 ( .A(n2282), .Z(n619) );
  MUX U1929 ( .IN0(g_input[8]), .IN1(n4981), .SEL(g_input[31]), .F(n2362) );
  MUX U1930 ( .IN0(n620), .IN1(n2355), .SEL(n2356), .F(n2239) );
  IV U1931 ( .A(n2357), .Z(n620) );
  MUX U1932 ( .IN0(e_input[9]), .IN1(n3848), .SEL(e_input[31]), .F(n2160) );
  MUX U1933 ( .IN0(g_input[9]), .IN1(n4969), .SEL(g_input[31]), .F(n2246) );
  MUX U1934 ( .IN0(n621), .IN1(n2197), .SEL(n2198), .F(n2086) );
  IV U1935 ( .A(n2199), .Z(n621) );
  MUX U1936 ( .IN0(n622), .IN1(n2189), .SEL(n2190), .F(n2078) );
  IV U1937 ( .A(n2191), .Z(n622) );
  MUX U1938 ( .IN0(n623), .IN1(n2205), .SEL(n2206), .F(n2094) );
  IV U1939 ( .A(n2207), .Z(n623) );
  MUX U1940 ( .IN0(g_input[10]), .IN1(n4955), .SEL(g_input[31]), .F(n2135) );
  MUX U1941 ( .IN0(n624), .IN1(n2006), .SEL(n2007), .F(n1901) );
  IV U1942 ( .A(n2008), .Z(n624) );
  MUX U1943 ( .IN0(g_input[11]), .IN1(n4943), .SEL(g_input[31]), .F(n2030) );
  MUX U1944 ( .IN0(e_input[12]), .IN1(n3862), .SEL(e_input[31]), .F(n1852) );
  MUX U1945 ( .IN0(g_input[12]), .IN1(n4929), .SEL(g_input[31]), .F(n1925) );
  MUX U1946 ( .IN0(n625), .IN1(n1918), .SEL(n1919), .F(n1818) );
  IV U1947 ( .A(n1920), .Z(n625) );
  MUX U1948 ( .IN0(g_input[13]), .IN1(n4917), .SEL(g_input[31]), .F(n1825) );
  MUX U1949 ( .IN0(n626), .IN1(n1784), .SEL(n1785), .F(n1688) );
  IV U1950 ( .A(n1786), .Z(n626) );
  MUX U1951 ( .IN0(n627), .IN1(n1768), .SEL(n1769), .F(n1672) );
  IV U1952 ( .A(n1770), .Z(n627) );
  MUX U1953 ( .IN0(g_input[14]), .IN1(n4903), .SEL(g_input[31]), .F(n1731) );
  MUX U1954 ( .IN0(n628), .IN1(n1614), .SEL(n1615), .F(n1522) );
  IV U1955 ( .A(n1616), .Z(n628) );
  MUX U1956 ( .IN0(g_input[15]), .IN1(n4891), .SEL(g_input[31]), .F(n1638) );
  MUX U1957 ( .IN0(e_input[16]), .IN1(n5065), .SEL(e_input[31]), .F(n1516) );
  MUX U1958 ( .IN0(g_input[16]), .IN1(n4519), .SEL(g_input[31]), .F(n1546) );
  MUX U1959 ( .IN0(n629), .IN1(n1539), .SEL(n1540), .F(n1453) );
  IV U1960 ( .A(n1541), .Z(n629) );
  MUX U1961 ( .IN0(e_input[17]), .IN1(n5066), .SEL(e_input[31]), .F(n1428) );
  MUX U1962 ( .IN0(n630), .IN1(n1403), .SEL(n1404), .F(n1331) );
  IV U1963 ( .A(n1405), .Z(n630) );
  MUX U1964 ( .IN0(g_input[17]), .IN1(n4505), .SEL(g_input[31]), .F(n1460) );
  MUX U1965 ( .IN0(g_input[18]), .IN1(n4491), .SEL(g_input[31]), .F(n1383) );
  MUX U1966 ( .IN0(n631), .IN1(n1269), .SEL(n1270), .F(n1203) );
  IV U1967 ( .A(n1271), .Z(n631) );
  MUX U1968 ( .IN0(n632), .IN1(n1419), .SEL(n1420), .F(n1349) );
  IV U1969 ( .A(n1421), .Z(n632) );
  MUX U1970 ( .IN0(g_input[19]), .IN1(n4479), .SEL(g_input[31]), .F(n1312) );
  MUX U1971 ( .IN0(n633), .IN1(n1288), .SEL(n1289), .F(n1218) );
  IV U1972 ( .A(n1290), .Z(n633) );
  MUX U1973 ( .IN0(g_input[20]), .IN1(n4465), .SEL(g_input[31]), .F(n1242) );
  MUX U1974 ( .IN0(e_input[20]), .IN1(n4879), .SEL(e_input[31]), .F(n1194) );
  MUX U1975 ( .IN0(e_input[21]), .IN1(n4880), .SEL(e_input[31]), .F(n1136) );
  MUX U1976 ( .IN0(g_input[21]), .IN1(n4453), .SEL(g_input[31]), .F(n1176) );
  MUX U1977 ( .IN0(n634), .IN1(n1178), .SEL(n1179), .F(n1116) );
  IV U1978 ( .A(n1180), .Z(n634) );
  MUX U1979 ( .IN0(g_input[22]), .IN1(n4439), .SEL(g_input[31]), .F(n1114) );
  MUX U1980 ( .IN0(n635), .IN1(n1031), .SEL(n1032), .F(n974) );
  IV U1981 ( .A(n1033), .Z(n635) );
  MUX U1982 ( .IN0(g_input[23]), .IN1(n4427), .SEL(g_input[31]), .F(n1055) );
  MUX U1983 ( .IN0(g_input[24]), .IN1(n4413), .SEL(g_input[31]), .F(n999) );
  MUX U1984 ( .IN0(e_input[24]), .IN1(n5155), .SEL(e_input[31]), .F(n982) );
  MUX U1985 ( .IN0(e_input[25]), .IN1(n5156), .SEL(e_input[31]), .F(n928) );
  MUX U1986 ( .IN0(g_input[25]), .IN1(n4401), .SEL(g_input[31]), .F(n941) );
  MUX U1987 ( .IN0(g_input[26]), .IN1(n4387), .SEL(g_input[31]), .F(n898) );
  MUX U1988 ( .IN0(e_input[27]), .IN1(n5140), .SEL(e_input[31]), .F(n636) );
  IV U1989 ( .A(n636), .Z(n835) );
  MUX U1990 ( .IN0(e_input[26]), .IN1(n5141), .SEL(e_input[31]), .F(n874) );
  MUX U1991 ( .IN0(g_input[27]), .IN1(n4375), .SEL(g_input[31]), .F(n854) );
  XOR U1992 ( .A(n3007), .B(n3140), .Z(n3008) );
  MUX U1993 ( .IN0(n3138), .IN1(n3136), .SEL(n3137), .F(n3001) );
  MUX U1994 ( .IN0(n3088), .IN1(n3086), .SEL(n3087), .F(n2951) );
  MUX U1995 ( .IN0(e_input[2]), .IN1(n4678), .SEL(e_input[31]), .F(n3070) );
  XOR U1996 ( .A(n5075), .B(n3124), .Z(n3128) );
  XNOR U1997 ( .A(n4861), .B(n4860), .Z(n4708) );
  XOR U1998 ( .A(n4888), .B(n3107), .Z(n3111) );
  XNOR U1999 ( .A(n3187), .B(n3186), .Z(n3197) );
  XNOR U2000 ( .A(n4126), .B(n4125), .Z(n3764) );
  MUX U2001 ( .IN0(e_input[3]), .IN1(n4679), .SEL(e_input[31]), .F(n2938) );
  MUX U2002 ( .IN0(e_input[5]), .IN1(n4313), .SEL(e_input[31]), .F(n2660) );
  MUX U2003 ( .IN0(n2556), .IN1(n2554), .SEL(n2555), .F(n2430) );
  MUX U2004 ( .IN0(n2606), .IN1(n2604), .SEL(n2605), .F(n2480) );
  MUX U2005 ( .IN0(e_input[6]), .IN1(n4317), .SEL(e_input[31]), .F(n2538) );
  XOR U2006 ( .A(n2249), .B(n2363), .Z(n2250) );
  MUX U2007 ( .IN0(e_input[10]), .IN1(n3832), .SEL(e_input[31]), .F(n2047) );
  MUX U2008 ( .IN0(e_input[11]), .IN1(n3833), .SEL(e_input[31]), .F(n1946) );
  MUX U2009 ( .IN0(n1874), .IN1(n1872), .SEL(n1873), .F(n1772) );
  XOR U2010 ( .A(n1828), .B(n1926), .Z(n1829) );
  MUX U2011 ( .IN0(n1924), .IN1(n1922), .SEL(n1923), .F(n1822) );
  MUX U2012 ( .IN0(e_input[13]), .IN1(n3863), .SEL(e_input[31]), .F(n1751) );
  MUX U2013 ( .IN0(n1855), .IN1(n637), .SEL(n1854), .F(n1753) );
  IV U2014 ( .A(n1853), .Z(n637) );
  MUX U2015 ( .IN0(e_input[18]), .IN1(n5050), .SEL(e_input[31]), .F(n1348) );
  MUX U2016 ( .IN0(e_input[19]), .IN1(n5051), .SEL(e_input[31]), .F(n1280) );
  MUX U2017 ( .IN0(e_input[22]), .IN1(n4885), .SEL(e_input[31]), .F(n1079) );
  MUX U2018 ( .IN0(e_input[23]), .IN1(n4884), .SEL(e_input[31]), .F(n638) );
  IV U2019 ( .A(n638), .Z(n1020) );
  MUX U2020 ( .IN0(e_input[28]), .IN1(n5174), .SEL(e_input[31]), .F(n806) );
  MUX U2021 ( .IN0(e_input[29]), .IN1(n5175), .SEL(e_input[31]), .F(n770) );
  MUX U2022 ( .IN0(n639), .IN1(n856), .SEL(n857), .F(n816) );
  IV U2023 ( .A(n858), .Z(n639) );
  MUX U2024 ( .IN0(g_input[28]), .IN1(n4361), .SEL(g_input[31]), .F(n814) );
  NAND U2025 ( .A(n2935), .B(n3069), .Z(n3068) );
  XNOR U2026 ( .A(n3059), .B(n3058), .Z(n3076) );
  XNOR U2027 ( .A(n3752), .B(n3751), .Z(n3176) );
  XOR U2028 ( .A(n2889), .B(n2760), .Z(n2764) );
  XNOR U2029 ( .A(n2915), .B(n2794), .Z(n2788) );
  XOR U2030 ( .A(n2831), .B(n2702), .Z(n2706) );
  XOR U2031 ( .A(n2848), .B(n2719), .Z(n2723) );
  XOR U2032 ( .A(n2505), .B(n2387), .Z(n2391) );
  MUX U2033 ( .IN0(e_input[7]), .IN1(n4318), .SEL(e_input[31]), .F(n2413) );
  XOR U2034 ( .A(n2465), .B(n2347), .Z(n2351) );
  XOR U2035 ( .A(n2448), .B(n2330), .Z(n2334) );
  XNOR U2036 ( .A(n2054), .B(n2157), .Z(n2055) );
  NAND U2037 ( .A(n1943), .B(n2046), .Z(n2045) );
  XOR U2038 ( .A(n2100), .B(n1998), .Z(n2002) );
  XOR U2039 ( .A(n2117), .B(n2015), .Z(n2019) );
  XOR U2040 ( .A(n1758), .B(n1759), .Z(n1755) );
  XOR U2041 ( .A(n1807), .B(n1714), .Z(n1718) );
  XOR U2042 ( .A(n1790), .B(n1697), .Z(n1701) );
  XOR U2043 ( .A(n1662), .B(n1663), .Z(n1657) );
  MUX U2044 ( .IN0(e_input[14]), .IN1(n3867), .SEL(e_input[31]), .F(n1660) );
  NAND U2045 ( .A(n1430), .B(n1515), .Z(n1514) );
  XOR U2046 ( .A(n1528), .B(n1445), .Z(n1449) );
  XNOR U2047 ( .A(n1374), .B(n1306), .Z(n1310) );
  XNOR U2048 ( .A(n1259), .B(n1196), .Z(n1200) );
  XOR U2049 ( .A(n1294), .B(n1227), .Z(n1231) );
  XNOR U2050 ( .A(n1167), .B(n1108), .Z(n1112) );
  XOR U2051 ( .A(n1096), .B(n1040), .Z(n1044) );
  XNOR U2052 ( .A(n990), .B(n935), .Z(n939) );
  XNOR U2053 ( .A(n883), .B(n888), .Z(n924) );
  MUX U2054 ( .IN0(n640), .IN1(n836), .SEL(n837), .F(n799) );
  IV U2055 ( .A(n838), .Z(n640) );
  MUX U2056 ( .IN0(n641), .IN1(n807), .SEL(n808), .F(n766) );
  IV U2057 ( .A(n809), .Z(n641) );
  MUX U2058 ( .IN0(g_input[29]), .IN1(n4349), .SEL(g_input[31]), .F(n774) );
  XNOR U2059 ( .A(n2923), .B(n2922), .Z(n2943) );
  XNOR U2060 ( .A(n3024), .B(n3023), .Z(n3066) );
  XNOR U2061 ( .A(n2774), .B(n2773), .Z(n2756) );
  XNOR U2062 ( .A(n2648), .B(n2647), .Z(n2630) );
  XNOR U2063 ( .A(n2683), .B(n2682), .Z(n2698) );
  XNOR U2064 ( .A(n2733), .B(n2732), .Z(n2715) );
  XNOR U2065 ( .A(n2524), .B(n2523), .Z(n2504) );
  XNOR U2066 ( .A(n2401), .B(n2400), .Z(n2383) );
  XNOR U2067 ( .A(n2286), .B(n2285), .Z(n2267) );
  XNOR U2068 ( .A(n2361), .B(n2360), .Z(n2343) );
  XNOR U2069 ( .A(n2311), .B(n2310), .Z(n2326) );
  XNOR U2070 ( .A(n2174), .B(n2173), .Z(n2156) );
  XNOR U2071 ( .A(n2065), .B(n2064), .Z(n2053) );
  XNOR U2072 ( .A(n1960), .B(n1959), .Z(n1951) );
  XNOR U2073 ( .A(n1979), .B(n1978), .Z(n1994) );
  XNOR U2074 ( .A(n2029), .B(n2028), .Z(n2011) );
  XNOR U2075 ( .A(n1730), .B(n1729), .Z(n1710) );
  XNOR U2076 ( .A(n1678), .B(n1677), .Z(n1693) );
  XNOR U2077 ( .A(n1587), .B(n1586), .Z(n1602) );
  XNOR U2078 ( .A(n1494), .B(n1493), .Z(n1509) );
  MUX U2079 ( .IN0(e_input[15]), .IN1(n3868), .SEL(e_input[31]), .F(n1566) );
  XNOR U2080 ( .A(n1409), .B(n1408), .Z(n1424) );
  XNOR U2081 ( .A(n1459), .B(n1458), .Z(n1441) );
  XNOR U2082 ( .A(n1211), .B(n1215), .Z(n1275) );
  XNOR U2083 ( .A(n1241), .B(n1240), .Z(n1223) );
  XNOR U2084 ( .A(n1139), .B(n1138), .Z(n1149) );
  XNOR U2085 ( .A(n1075), .B(n1074), .Z(n1087) );
  XNOR U2086 ( .A(n1054), .B(n1053), .Z(n1036) );
  XNOR U2087 ( .A(n1019), .B(n1018), .Z(n1028) );
  XNOR U2088 ( .A(n965), .B(n964), .Z(n961) );
  XNOR U2089 ( .A(n897), .B(n896), .Z(n880) );
  MUX U2090 ( .IN0(g_input[30]), .IN1(n4331), .SEL(g_input[31]), .F(n740) );
  MUX U2091 ( .IN0(e_input[30]), .IN1(n5180), .SEL(e_input[31]), .F(n742) );
  XNOR U2092 ( .A(n2888), .B(n2887), .Z(n2930) );
  XNOR U2093 ( .A(n3095), .B(n3094), .Z(n3049) );
  XNOR U2094 ( .A(n2544), .B(n2543), .Z(n2656) );
  XOR U2095 ( .A(n2294), .B(n2182), .Z(n2183) );
  NANDN U2096 ( .B(n1863), .A(n1864), .Z(n1763) );
  XNOR U2097 ( .A(n1619), .B(n1618), .Z(n1594) );
  XNOR U2098 ( .A(n1527), .B(n1526), .Z(n1501) );
  ANDN U2099 ( .A(n1644), .B(n1645), .Z(n1552) );
  XNOR U2100 ( .A(n1364), .B(n1363), .Z(n1344) );
  XNOR U2101 ( .A(n1157), .B(n1156), .Z(n1146) );
  XNOR U2102 ( .A(n979), .B(n978), .Z(n971) );
  XNOR U2103 ( .A(n841), .B(n840), .Z(n833) );
  MUX U2104 ( .IN0(n737), .IN1(n735), .SEL(n736), .F(n706) );
  XNOR U2105 ( .A(n705), .B(n704), .Z(n703) );
  XNOR U2106 ( .A(n2960), .B(n2959), .Z(n2913) );
  XNOR U2107 ( .A(n2822), .B(n2821), .Z(n2781) );
  XNOR U2108 ( .A(n2563), .B(n2562), .Z(n2531) );
  XNOR U2109 ( .A(n2439), .B(n2438), .Z(n2408) );
  XNOR U2110 ( .A(n2202), .B(n2201), .Z(n2181) );
  XNOR U2111 ( .A(n2091), .B(n2090), .Z(n2072) );
  XNOR U2112 ( .A(n1881), .B(n1880), .Z(n1862) );
  XNOR U2113 ( .A(n1781), .B(n1780), .Z(n1762) );
  XNOR U2114 ( .A(n1482), .B(n1481), .Z(n1560) );
  MUX U2115 ( .IN0(n642), .IN1(n781), .SEL(n782), .F(n748) );
  IV U2116 ( .A(\_MxM/Y0[27] ), .Z(n642) );
  MUX U2117 ( .IN0(n643), .IN1(n711), .SEL(n712), .F(n688) );
  IV U2118 ( .A(n713), .Z(n643) );
  XOR U2119 ( .A(n1257), .B(n1256), .Z(n1323) );
  XNOR U2120 ( .A(n1069), .B(n1068), .Z(n1125) );
  XNOR U2121 ( .A(n912), .B(n911), .Z(n951) );
  XNOR U2122 ( .A(n789), .B(n788), .Z(n825) );
  XNOR U2123 ( .A(n726), .B(n725), .Z(n752) );
  XNOR U2124 ( .A(n672), .B(n671), .Z(n697) );
  XOR U2125 ( .A(n2740), .B(n2743), .Z(n2741) );
  XOR U2126 ( .A(n2370), .B(n2373), .Z(n2371) );
  XOR U2127 ( .A(n2038), .B(n2041), .Z(n2039) );
  XOR U2128 ( .A(n1739), .B(n1743), .Z(n1741) );
  XOR U2129 ( .A(n1468), .B(n1472), .Z(n1470) );
  XOR U2130 ( .A(n1250), .B(n1254), .Z(n1252) );
  XOR U2131 ( .A(n1062), .B(n1066), .Z(n1064) );
  XOR U2132 ( .A(n905), .B(n909), .Z(n907) );
  MUX U2133 ( .IN0(n658), .IN1(\_MxM/Y1[30] ), .SEL(n659), .F(\_MxM/Y1[31] )
         );
  MUX U2134 ( .IN0(\_MxM/Y1[24] ), .IN1(o[24]), .SEL(n644), .F(\_MxM/n99 ) );
  MUX U2135 ( .IN0(\_MxM/Y1[25] ), .IN1(o[25]), .SEL(n644), .F(\_MxM/n96 ) );
  MUX U2136 ( .IN0(\_MxM/Y1[26] ), .IN1(o[26]), .SEL(n644), .F(\_MxM/n93 ) );
  MUX U2137 ( .IN0(\_MxM/Y1[27] ), .IN1(o[27]), .SEL(n644), .F(\_MxM/n90 ) );
  MUX U2138 ( .IN0(\_MxM/Y1[28] ), .IN1(o[28]), .SEL(n644), .F(\_MxM/n87 ) );
  MUX U2139 ( .IN0(\_MxM/Y1[29] ), .IN1(o[29]), .SEL(n644), .F(\_MxM/n84 ) );
  MUX U2140 ( .IN0(\_MxM/Y1[30] ), .IN1(o[30]), .SEL(n644), .F(\_MxM/n81 ) );
  MUX U2141 ( .IN0(\_MxM/Y1[31] ), .IN1(o[31]), .SEL(n644), .F(\_MxM/n78 ) );
  MUX U2142 ( .IN0(\_MxM/Y1[0] ), .IN1(o[0]), .SEL(n644), .F(\_MxM/n171 ) );
  MUX U2143 ( .IN0(\_MxM/Y1[1] ), .IN1(o[1]), .SEL(n644), .F(\_MxM/n168 ) );
  MUX U2144 ( .IN0(\_MxM/Y1[2] ), .IN1(o[2]), .SEL(n644), .F(\_MxM/n165 ) );
  MUX U2145 ( .IN0(\_MxM/Y1[3] ), .IN1(o[3]), .SEL(n644), .F(\_MxM/n162 ) );
  MUX U2146 ( .IN0(\_MxM/Y1[4] ), .IN1(o[4]), .SEL(n644), .F(\_MxM/n159 ) );
  MUX U2147 ( .IN0(\_MxM/Y1[5] ), .IN1(o[5]), .SEL(n644), .F(\_MxM/n156 ) );
  MUX U2148 ( .IN0(\_MxM/Y1[6] ), .IN1(o[6]), .SEL(n644), .F(\_MxM/n153 ) );
  MUX U2149 ( .IN0(\_MxM/Y1[7] ), .IN1(o[7]), .SEL(n644), .F(\_MxM/n150 ) );
  MUX U2150 ( .IN0(\_MxM/Y1[8] ), .IN1(o[8]), .SEL(n644), .F(\_MxM/n147 ) );
  MUX U2151 ( .IN0(\_MxM/Y1[9] ), .IN1(o[9]), .SEL(n644), .F(\_MxM/n144 ) );
  MUX U2152 ( .IN0(\_MxM/Y1[10] ), .IN1(o[10]), .SEL(n644), .F(\_MxM/n141 ) );
  MUX U2153 ( .IN0(\_MxM/Y1[11] ), .IN1(o[11]), .SEL(n644), .F(\_MxM/n138 ) );
  MUX U2154 ( .IN0(\_MxM/Y1[12] ), .IN1(o[12]), .SEL(n644), .F(\_MxM/n135 ) );
  MUX U2155 ( .IN0(\_MxM/Y1[13] ), .IN1(o[13]), .SEL(n644), .F(\_MxM/n132 ) );
  MUX U2156 ( .IN0(\_MxM/Y1[14] ), .IN1(o[14]), .SEL(n644), .F(\_MxM/n129 ) );
  MUX U2157 ( .IN0(\_MxM/Y1[15] ), .IN1(o[15]), .SEL(n644), .F(\_MxM/n126 ) );
  MUX U2158 ( .IN0(\_MxM/Y1[16] ), .IN1(o[16]), .SEL(n644), .F(\_MxM/n123 ) );
  MUX U2159 ( .IN0(\_MxM/Y1[17] ), .IN1(o[17]), .SEL(n644), .F(\_MxM/n120 ) );
  MUX U2160 ( .IN0(\_MxM/Y1[18] ), .IN1(o[18]), .SEL(n644), .F(\_MxM/n117 ) );
  MUX U2161 ( .IN0(\_MxM/Y1[19] ), .IN1(o[19]), .SEL(n644), .F(\_MxM/n114 ) );
  MUX U2162 ( .IN0(\_MxM/Y1[20] ), .IN1(o[20]), .SEL(n644), .F(\_MxM/n111 ) );
  MUX U2163 ( .IN0(\_MxM/Y1[21] ), .IN1(o[21]), .SEL(n644), .F(\_MxM/n108 ) );
  IV U2164 ( .A(n645), .Z(n644) );
  MUX U2165 ( .IN0(o[22]), .IN1(\_MxM/Y1[22] ), .SEL(n645), .F(\_MxM/n105 ) );
  MUX U2166 ( .IN0(o[23]), .IN1(\_MxM/Y1[23] ), .SEL(n645), .F(\_MxM/n102 ) );
  AND U2167 ( .A(n646), .B(n647), .Z(n645) );
  ANDN U2168 ( .A(n648), .B(\_MxM/n[2] ), .Z(n647) );
  NOR U2169 ( .A(\_MxM/n[6] ), .B(\_MxM/n[5] ), .Z(n648) );
  ANDN U2170 ( .A(n649), .B(n650), .Z(n646) );
  ANDN U2171 ( .A(\_MxM/N11 ), .B(\_MxM/n[1] ), .Z(n649) );
  XOR U2172 ( .A(n651), .B(\_MxM/Y0[10] ), .Z(\_MxM/Y1[9] ) );
  XOR U2173 ( .A(n652), .B(\_MxM/Y0[9] ), .Z(\_MxM/Y1[8] ) );
  XOR U2174 ( .A(n653), .B(\_MxM/Y0[8] ), .Z(\_MxM/Y1[7] ) );
  XOR U2175 ( .A(n654), .B(\_MxM/Y0[7] ), .Z(\_MxM/Y1[6] ) );
  XOR U2176 ( .A(n655), .B(\_MxM/Y0[6] ), .Z(\_MxM/Y1[5] ) );
  XOR U2177 ( .A(n656), .B(\_MxM/Y0[5] ), .Z(\_MxM/Y1[4] ) );
  XNOR U2178 ( .A(n657), .B(\_MxM/Y0[4] ), .Z(\_MxM/Y1[3] ) );
  XNOR U2179 ( .A(\_MxM/Y0[31] ), .B(n660), .Z(n659) );
  XNOR U2180 ( .A(n662), .B(\_MxM/Y0[31] ), .Z(\_MxM/Y1[30] ) );
  XOR U2181 ( .A(n661), .B(n660), .Z(n662) );
  XOR U2182 ( .A(n663), .B(n664), .Z(n660) );
  XOR U2183 ( .A(n665), .B(n666), .Z(n664) );
  AND U2184 ( .A(n667), .B(n668), .Z(n666) );
  XNOR U2185 ( .A(n673), .B(n671), .Z(n663) );
  XOR U2186 ( .A(n674), .B(n675), .Z(n673) );
  XOR U2187 ( .A(n676), .B(n677), .Z(n675) );
  XOR U2188 ( .A(n678), .B(n679), .Z(n677) );
  XOR U2189 ( .A(n684), .B(n685), .Z(n676) );
  XOR U2190 ( .A(n690), .B(n691), .Z(n674) );
  XNOR U2191 ( .A(n680), .B(n692), .Z(n691) );
  XOR U2192 ( .A(n688), .B(n686), .Z(n690) );
  XNOR U2193 ( .A(n695), .B(\_MxM/Y0[3] ), .Z(\_MxM/Y1[2] ) );
  XNOR U2194 ( .A(n693), .B(\_MxM/Y0[30] ), .Z(\_MxM/Y1[29] ) );
  XNOR U2195 ( .A(n696), .B(n697), .Z(n693) );
  XNOR U2196 ( .A(n694), .B(n698), .Z(n696) );
  AND U2197 ( .A(n667), .B(n699), .Z(n698) );
  XOR U2198 ( .A(n670), .B(n697), .Z(n699) );
  XNOR U2199 ( .A(n669), .B(n697), .Z(n670) );
  XOR U2200 ( .A(n683), .B(n692), .Z(n681) );
  IV U2201 ( .A(n682), .Z(n692) );
  XOR U2202 ( .A(n688), .B(n689), .Z(n687) );
  OR U2203 ( .A(n709), .B(n710), .Z(n689) );
  ANDN U2204 ( .A(n718), .B(n719), .Z(n717) );
  XOR U2205 ( .A(\_MxM/Y0[29] ), .B(n720), .Z(n718) );
  XNOR U2206 ( .A(n719), .B(\_MxM/Y0[29] ), .Z(\_MxM/Y1[28] ) );
  XNOR U2207 ( .A(n721), .B(n722), .Z(n719) );
  XNOR U2208 ( .A(n720), .B(n723), .Z(n721) );
  AND U2209 ( .A(n667), .B(n724), .Z(n723) );
  XOR U2210 ( .A(n715), .B(n722), .Z(n724) );
  XNOR U2211 ( .A(n714), .B(n722), .Z(n715) );
  XOR U2212 ( .A(n729), .B(n730), .Z(n704) );
  ANDN U2213 ( .A(n731), .B(n729), .Z(n730) );
  XOR U2214 ( .A(n729), .B(n732), .Z(n731) );
  XOR U2215 ( .A(n733), .B(n734), .Z(n707) );
  IV U2216 ( .A(n706), .Z(n734) );
  XNOR U2217 ( .A(n712), .B(n713), .Z(n708) );
  NANDN U2218 ( .B(n709), .A(n740), .Z(n713) );
  XNOR U2219 ( .A(n711), .B(n741), .Z(n712) );
  ANDN U2220 ( .A(n742), .B(n710), .Z(n741) );
  IV U2221 ( .A(n716), .Z(n720) );
  XNOR U2222 ( .A(n749), .B(\_MxM/Y0[28] ), .Z(\_MxM/Y1[27] ) );
  XNOR U2223 ( .A(n751), .B(n752), .Z(n749) );
  XNOR U2224 ( .A(n750), .B(n753), .Z(n751) );
  AND U2225 ( .A(n667), .B(n754), .Z(n753) );
  XOR U2226 ( .A(n747), .B(n752), .Z(n754) );
  XNOR U2227 ( .A(n746), .B(n752), .Z(n747) );
  XOR U2228 ( .A(n757), .B(n758), .Z(n727) );
  ANDN U2229 ( .A(n759), .B(n757), .Z(n758) );
  XOR U2230 ( .A(n757), .B(n760), .Z(n759) );
  XOR U2231 ( .A(n737), .B(n764), .Z(n732) );
  IV U2232 ( .A(n736), .Z(n764) );
  XOR U2233 ( .A(n769), .B(n739), .Z(n765) );
  NANDN U2234 ( .B(n710), .A(n770), .Z(n739) );
  IV U2235 ( .A(n735), .Z(n769) );
  XNOR U2236 ( .A(n744), .B(n745), .Z(n737) );
  NANDN U2237 ( .B(n709), .A(n774), .Z(n745) );
  XNOR U2238 ( .A(n743), .B(n775), .Z(n744) );
  AND U2239 ( .A(n740), .B(n742), .Z(n775) );
  IV U2240 ( .A(n748), .Z(n750) );
  XNOR U2241 ( .A(n782), .B(\_MxM/Y0[27] ), .Z(\_MxM/Y1[26] ) );
  XNOR U2242 ( .A(n784), .B(n785), .Z(n782) );
  XNOR U2243 ( .A(n783), .B(n786), .Z(n784) );
  AND U2244 ( .A(n667), .B(n787), .Z(n786) );
  XOR U2245 ( .A(n780), .B(n785), .Z(n787) );
  XNOR U2246 ( .A(n779), .B(n785), .Z(n780) );
  XNOR U2247 ( .A(n763), .B(n762), .Z(n760) );
  XOR U2248 ( .A(n792), .B(n793), .Z(n762) );
  XOR U2249 ( .A(n794), .B(n795), .Z(n793) );
  XOR U2250 ( .A(n796), .B(n797), .Z(n795) );
  XNOR U2251 ( .A(n766), .B(n805), .Z(n767) );
  ANDN U2252 ( .A(n806), .B(n710), .Z(n805) );
  XOR U2253 ( .A(n810), .B(n768), .Z(n804) );
  NAND U2254 ( .A(n770), .B(n740), .Z(n768) );
  IV U2255 ( .A(n771), .Z(n810) );
  XNOR U2256 ( .A(n777), .B(n778), .Z(n773) );
  NANDN U2257 ( .B(n709), .A(n814), .Z(n778) );
  XNOR U2258 ( .A(n776), .B(n815), .Z(n777) );
  AND U2259 ( .A(n774), .B(n742), .Z(n815) );
  IV U2260 ( .A(n781), .Z(n783) );
  XNOR U2261 ( .A(n822), .B(\_MxM/Y0[26] ), .Z(\_MxM/Y1[25] ) );
  XNOR U2262 ( .A(n824), .B(n825), .Z(n822) );
  XNOR U2263 ( .A(n823), .B(n826), .Z(n824) );
  AND U2264 ( .A(n667), .B(n827), .Z(n826) );
  XOR U2265 ( .A(n820), .B(n825), .Z(n827) );
  XNOR U2266 ( .A(n819), .B(n825), .Z(n820) );
  XOR U2267 ( .A(n830), .B(n831), .Z(n790) );
  ANDN U2268 ( .A(n832), .B(n830), .Z(n831) );
  XOR U2269 ( .A(n830), .B(n833), .Z(n832) );
  XNOR U2270 ( .A(n834), .B(n798), .Z(n802) );
  XOR U2271 ( .A(n799), .B(n800), .Z(n798) );
  OR U2272 ( .A(n710), .B(n835), .Z(n800) );
  XNOR U2273 ( .A(n794), .B(n801), .Z(n834) );
  XNOR U2274 ( .A(n807), .B(n846), .Z(n808) );
  AND U2275 ( .A(n740), .B(n806), .Z(n846) );
  XOR U2276 ( .A(n850), .B(n809), .Z(n845) );
  NAND U2277 ( .A(n770), .B(n774), .Z(n809) );
  IV U2278 ( .A(n811), .Z(n850) );
  XNOR U2279 ( .A(n817), .B(n818), .Z(n813) );
  NANDN U2280 ( .B(n709), .A(n854), .Z(n818) );
  XNOR U2281 ( .A(n816), .B(n855), .Z(n817) );
  AND U2282 ( .A(n814), .B(n742), .Z(n855) );
  IV U2283 ( .A(n821), .Z(n823) );
  XNOR U2284 ( .A(n862), .B(\_MxM/Y0[25] ), .Z(\_MxM/Y1[24] ) );
  XNOR U2285 ( .A(n864), .B(n865), .Z(n862) );
  XNOR U2286 ( .A(n863), .B(n866), .Z(n864) );
  AND U2287 ( .A(n667), .B(n867), .Z(n866) );
  XOR U2288 ( .A(n860), .B(n865), .Z(n867) );
  XNOR U2289 ( .A(n859), .B(n865), .Z(n860) );
  XNOR U2290 ( .A(n872), .B(n844), .Z(n840) );
  XNOR U2291 ( .A(n837), .B(n838), .Z(n844) );
  NANDN U2292 ( .B(n835), .A(n740), .Z(n838) );
  XNOR U2293 ( .A(n836), .B(n873), .Z(n837) );
  ANDN U2294 ( .A(n874), .B(n710), .Z(n873) );
  XNOR U2295 ( .A(n843), .B(n839), .Z(n872) );
  XNOR U2296 ( .A(n881), .B(n882), .Z(n843) );
  IV U2297 ( .A(n842), .Z(n882) );
  XNOR U2298 ( .A(n847), .B(n890), .Z(n848) );
  AND U2299 ( .A(n774), .B(n806), .Z(n890) );
  XOR U2300 ( .A(n894), .B(n849), .Z(n889) );
  NAND U2301 ( .A(n770), .B(n814), .Z(n849) );
  IV U2302 ( .A(n851), .Z(n894) );
  XNOR U2303 ( .A(n857), .B(n858), .Z(n853) );
  NANDN U2304 ( .B(n709), .A(n898), .Z(n858) );
  XNOR U2305 ( .A(n856), .B(n899), .Z(n857) );
  AND U2306 ( .A(n854), .B(n742), .Z(n899) );
  IV U2307 ( .A(n861), .Z(n863) );
  XNOR U2308 ( .A(n906), .B(\_MxM/Y0[24] ), .Z(\_MxM/Y1[23] ) );
  XNOR U2309 ( .A(n907), .B(n908), .Z(n906) );
  AND U2310 ( .A(n667), .B(n910), .Z(n909) );
  XOR U2311 ( .A(n904), .B(n908), .Z(n910) );
  XNOR U2312 ( .A(n903), .B(n908), .Z(n904) );
  XNOR U2313 ( .A(n916), .B(n885), .Z(n879) );
  XNOR U2314 ( .A(n876), .B(n877), .Z(n885) );
  NANDN U2315 ( .B(n835), .A(n774), .Z(n877) );
  XNOR U2316 ( .A(n875), .B(n917), .Z(n876) );
  AND U2317 ( .A(n740), .B(n874), .Z(n917) );
  XNOR U2318 ( .A(n884), .B(n878), .Z(n916) );
  XNOR U2319 ( .A(n924), .B(n886), .Z(n884) );
  IV U2320 ( .A(n887), .Z(n886) );
  NANDN U2321 ( .B(n710), .A(n928), .Z(n888) );
  XNOR U2322 ( .A(n891), .B(n933), .Z(n892) );
  AND U2323 ( .A(n814), .B(n806), .Z(n933) );
  XOR U2324 ( .A(n937), .B(n893), .Z(n932) );
  NAND U2325 ( .A(n770), .B(n854), .Z(n893) );
  IV U2326 ( .A(n895), .Z(n937) );
  XNOR U2327 ( .A(n901), .B(n902), .Z(n897) );
  NANDN U2328 ( .B(n709), .A(n941), .Z(n902) );
  XNOR U2329 ( .A(n900), .B(n942), .Z(n901) );
  AND U2330 ( .A(n898), .B(n742), .Z(n942) );
  XNOR U2331 ( .A(n949), .B(\_MxM/Y0[23] ), .Z(\_MxM/Y1[22] ) );
  XNOR U2332 ( .A(n950), .B(n951), .Z(n949) );
  AND U2333 ( .A(n667), .B(n953), .Z(n952) );
  XOR U2334 ( .A(n947), .B(n951), .Z(n953) );
  XNOR U2335 ( .A(n946), .B(n951), .Z(n947) );
  XNOR U2336 ( .A(n915), .B(n914), .Z(n912) );
  XOR U2337 ( .A(n956), .B(n957), .Z(n914) );
  XOR U2338 ( .A(n958), .B(n959), .Z(n957) );
  XOR U2339 ( .A(n962), .B(n963), .Z(n958) );
  XOR U2340 ( .A(n968), .B(n913), .Z(n956) );
  XOR U2341 ( .A(n966), .B(n964), .Z(n968) );
  XNOR U2342 ( .A(n972), .B(n931), .Z(n922) );
  XNOR U2343 ( .A(n919), .B(n920), .Z(n931) );
  NANDN U2344 ( .B(n835), .A(n814), .Z(n920) );
  XNOR U2345 ( .A(n918), .B(n973), .Z(n919) );
  AND U2346 ( .A(n774), .B(n874), .Z(n973) );
  XNOR U2347 ( .A(n930), .B(n921), .Z(n972) );
  XNOR U2348 ( .A(n925), .B(n981), .Z(n926) );
  ANDN U2349 ( .A(n982), .B(n710), .Z(n981) );
  XOR U2350 ( .A(n986), .B(n927), .Z(n980) );
  NAND U2351 ( .A(n928), .B(n740), .Z(n927) );
  IV U2352 ( .A(n929), .Z(n986) );
  XNOR U2353 ( .A(n934), .B(n991), .Z(n935) );
  AND U2354 ( .A(n854), .B(n806), .Z(n991) );
  XOR U2355 ( .A(n995), .B(n936), .Z(n990) );
  NAND U2356 ( .A(n770), .B(n898), .Z(n936) );
  IV U2357 ( .A(n938), .Z(n995) );
  XNOR U2358 ( .A(n944), .B(n945), .Z(n940) );
  NANDN U2359 ( .B(n709), .A(n999), .Z(n945) );
  XNOR U2360 ( .A(n943), .B(n1000), .Z(n944) );
  AND U2361 ( .A(n941), .B(n742), .Z(n1000) );
  XNOR U2362 ( .A(n1007), .B(\_MxM/Y0[22] ), .Z(\_MxM/Y1[21] ) );
  XNOR U2363 ( .A(n1008), .B(n1009), .Z(n1007) );
  AND U2364 ( .A(n667), .B(n1011), .Z(n1010) );
  XOR U2365 ( .A(n1005), .B(n1009), .Z(n1011) );
  XNOR U2366 ( .A(n1004), .B(n1009), .Z(n1005) );
  XNOR U2367 ( .A(n1014), .B(n961), .Z(n970) );
  XOR U2368 ( .A(n1015), .B(n1016), .Z(n964) );
  ANDN U2369 ( .A(n1017), .B(n1018), .Z(n1016) );
  XOR U2370 ( .A(n1015), .B(n1019), .Z(n1017) );
  XOR U2371 ( .A(n966), .B(n967), .Z(n965) );
  OR U2372 ( .A(n710), .B(n1020), .Z(n967) );
  XNOR U2373 ( .A(n960), .B(n969), .Z(n1014) );
  XNOR U2374 ( .A(n1029), .B(n989), .Z(n978) );
  XNOR U2375 ( .A(n975), .B(n976), .Z(n989) );
  NANDN U2376 ( .B(n835), .A(n854), .Z(n976) );
  XNOR U2377 ( .A(n974), .B(n1030), .Z(n975) );
  AND U2378 ( .A(n814), .B(n874), .Z(n1030) );
  XNOR U2379 ( .A(n988), .B(n977), .Z(n1029) );
  XNOR U2380 ( .A(n983), .B(n1038), .Z(n984) );
  AND U2381 ( .A(n740), .B(n982), .Z(n1038) );
  XOR U2382 ( .A(n1042), .B(n985), .Z(n1037) );
  NAND U2383 ( .A(n928), .B(n774), .Z(n985) );
  IV U2384 ( .A(n987), .Z(n1042) );
  XNOR U2385 ( .A(n992), .B(n1047), .Z(n993) );
  AND U2386 ( .A(n898), .B(n806), .Z(n1047) );
  XOR U2387 ( .A(n1051), .B(n994), .Z(n1046) );
  NAND U2388 ( .A(n770), .B(n941), .Z(n994) );
  IV U2389 ( .A(n996), .Z(n1051) );
  XNOR U2390 ( .A(n1002), .B(n1003), .Z(n998) );
  NANDN U2391 ( .B(n709), .A(n1055), .Z(n1003) );
  XNOR U2392 ( .A(n1001), .B(n1056), .Z(n1002) );
  AND U2393 ( .A(n999), .B(n742), .Z(n1056) );
  XNOR U2394 ( .A(n1063), .B(\_MxM/Y0[21] ), .Z(\_MxM/Y1[20] ) );
  XNOR U2395 ( .A(n1064), .B(n1065), .Z(n1063) );
  AND U2396 ( .A(n667), .B(n1067), .Z(n1066) );
  XOR U2397 ( .A(n1061), .B(n1065), .Z(n1067) );
  XNOR U2398 ( .A(n1060), .B(n1065), .Z(n1061) );
  XNOR U2399 ( .A(n1070), .B(n1028), .Z(n1025) );
  XOR U2400 ( .A(n1071), .B(n1072), .Z(n1018) );
  IV U2401 ( .A(n1015), .Z(n1072) );
  XNOR U2402 ( .A(n1022), .B(n1023), .Z(n1019) );
  NANDN U2403 ( .B(n1020), .A(n740), .Z(n1023) );
  XNOR U2404 ( .A(n1021), .B(n1078), .Z(n1022) );
  ANDN U2405 ( .A(n1079), .B(n710), .Z(n1078) );
  XNOR U2406 ( .A(n1088), .B(n1045), .Z(n1035) );
  XNOR U2407 ( .A(n1032), .B(n1033), .Z(n1045) );
  NANDN U2408 ( .B(n835), .A(n898), .Z(n1033) );
  XNOR U2409 ( .A(n1031), .B(n1089), .Z(n1032) );
  AND U2410 ( .A(n854), .B(n874), .Z(n1089) );
  XNOR U2411 ( .A(n1044), .B(n1034), .Z(n1088) );
  XNOR U2412 ( .A(n1039), .B(n1097), .Z(n1040) );
  AND U2413 ( .A(n774), .B(n982), .Z(n1097) );
  XOR U2414 ( .A(n1101), .B(n1041), .Z(n1096) );
  NAND U2415 ( .A(n928), .B(n814), .Z(n1041) );
  IV U2416 ( .A(n1043), .Z(n1101) );
  XNOR U2417 ( .A(n1048), .B(n1106), .Z(n1049) );
  AND U2418 ( .A(n941), .B(n806), .Z(n1106) );
  XOR U2419 ( .A(n1110), .B(n1050), .Z(n1105) );
  NAND U2420 ( .A(n770), .B(n999), .Z(n1050) );
  IV U2421 ( .A(n1052), .Z(n1110) );
  XNOR U2422 ( .A(n1058), .B(n1059), .Z(n1054) );
  NANDN U2423 ( .B(n709), .A(n1114), .Z(n1059) );
  XNOR U2424 ( .A(n1057), .B(n1115), .Z(n1058) );
  AND U2425 ( .A(n1055), .B(n742), .Z(n1115) );
  XNOR U2426 ( .A(n1123), .B(\_MxM/Y0[2] ), .Z(\_MxM/Y1[1] ) );
  XNOR U2427 ( .A(n1122), .B(\_MxM/Y0[20] ), .Z(\_MxM/Y1[19] ) );
  XNOR U2428 ( .A(n1124), .B(n1125), .Z(n1122) );
  AND U2429 ( .A(n667), .B(n1127), .Z(n1126) );
  XOR U2430 ( .A(n1120), .B(n1125), .Z(n1127) );
  XNOR U2431 ( .A(n1119), .B(n1125), .Z(n1120) );
  XNOR U2432 ( .A(n1130), .B(n1087), .Z(n1084) );
  XOR U2433 ( .A(n1135), .B(n1077), .Z(n1131) );
  NANDN U2434 ( .B(n710), .A(n1136), .Z(n1077) );
  IV U2435 ( .A(n1073), .Z(n1135) );
  XNOR U2436 ( .A(n1081), .B(n1082), .Z(n1075) );
  NANDN U2437 ( .B(n1020), .A(n774), .Z(n1082) );
  XNOR U2438 ( .A(n1080), .B(n1140), .Z(n1081) );
  AND U2439 ( .A(n740), .B(n1079), .Z(n1140) );
  XNOR U2440 ( .A(n1150), .B(n1104), .Z(n1094) );
  XNOR U2441 ( .A(n1091), .B(n1092), .Z(n1104) );
  NANDN U2442 ( .B(n835), .A(n941), .Z(n1092) );
  XNOR U2443 ( .A(n1090), .B(n1151), .Z(n1091) );
  AND U2444 ( .A(n898), .B(n874), .Z(n1151) );
  XNOR U2445 ( .A(n1103), .B(n1093), .Z(n1150) );
  XNOR U2446 ( .A(n1098), .B(n1159), .Z(n1099) );
  AND U2447 ( .A(n814), .B(n982), .Z(n1159) );
  XOR U2448 ( .A(n1163), .B(n1100), .Z(n1158) );
  NAND U2449 ( .A(n928), .B(n854), .Z(n1100) );
  IV U2450 ( .A(n1102), .Z(n1163) );
  XNOR U2451 ( .A(n1107), .B(n1168), .Z(n1108) );
  AND U2452 ( .A(n999), .B(n806), .Z(n1168) );
  XOR U2453 ( .A(n1172), .B(n1109), .Z(n1167) );
  NAND U2454 ( .A(n770), .B(n1055), .Z(n1109) );
  IV U2455 ( .A(n1111), .Z(n1172) );
  XNOR U2456 ( .A(n1117), .B(n1118), .Z(n1113) );
  NANDN U2457 ( .B(n709), .A(n1176), .Z(n1118) );
  XNOR U2458 ( .A(n1116), .B(n1177), .Z(n1117) );
  AND U2459 ( .A(n1114), .B(n742), .Z(n1177) );
  XNOR U2460 ( .A(n1184), .B(\_MxM/Y0[19] ), .Z(\_MxM/Y1[18] ) );
  XNOR U2461 ( .A(n1185), .B(n1186), .Z(n1184) );
  AND U2462 ( .A(n667), .B(n1188), .Z(n1187) );
  XOR U2463 ( .A(n1182), .B(n1186), .Z(n1188) );
  XNOR U2464 ( .A(n1181), .B(n1186), .Z(n1182) );
  XNOR U2465 ( .A(n1191), .B(n1149), .Z(n1145) );
  XNOR U2466 ( .A(n1132), .B(n1193), .Z(n1133) );
  ANDN U2467 ( .A(n1194), .B(n710), .Z(n1193) );
  XOR U2468 ( .A(n1198), .B(n1134), .Z(n1192) );
  NAND U2469 ( .A(n1136), .B(n740), .Z(n1134) );
  IV U2470 ( .A(n1137), .Z(n1198) );
  XNOR U2471 ( .A(n1142), .B(n1143), .Z(n1139) );
  NANDN U2472 ( .B(n1020), .A(n814), .Z(n1143) );
  XNOR U2473 ( .A(n1141), .B(n1202), .Z(n1142) );
  AND U2474 ( .A(n774), .B(n1079), .Z(n1202) );
  XNOR U2475 ( .A(n1148), .B(n1144), .Z(n1191) );
  XNOR U2476 ( .A(n1209), .B(n1210), .Z(n1148) );
  IV U2477 ( .A(n1147), .Z(n1210) );
  XNOR U2478 ( .A(n1216), .B(n1166), .Z(n1156) );
  XNOR U2479 ( .A(n1153), .B(n1154), .Z(n1166) );
  NANDN U2480 ( .B(n835), .A(n999), .Z(n1154) );
  XNOR U2481 ( .A(n1152), .B(n1217), .Z(n1153) );
  AND U2482 ( .A(n941), .B(n874), .Z(n1217) );
  XNOR U2483 ( .A(n1165), .B(n1155), .Z(n1216) );
  XNOR U2484 ( .A(n1160), .B(n1225), .Z(n1161) );
  AND U2485 ( .A(n854), .B(n982), .Z(n1225) );
  XOR U2486 ( .A(n1229), .B(n1162), .Z(n1224) );
  NAND U2487 ( .A(n928), .B(n898), .Z(n1162) );
  IV U2488 ( .A(n1164), .Z(n1229) );
  XNOR U2489 ( .A(n1169), .B(n1234), .Z(n1170) );
  AND U2490 ( .A(n1055), .B(n806), .Z(n1234) );
  XOR U2491 ( .A(n1238), .B(n1171), .Z(n1233) );
  NAND U2492 ( .A(n770), .B(n1114), .Z(n1171) );
  IV U2493 ( .A(n1173), .Z(n1238) );
  XNOR U2494 ( .A(n1179), .B(n1180), .Z(n1175) );
  NANDN U2495 ( .B(n709), .A(n1242), .Z(n1180) );
  XNOR U2496 ( .A(n1178), .B(n1243), .Z(n1179) );
  AND U2497 ( .A(n1176), .B(n742), .Z(n1243) );
  ANDN U2498 ( .A(n1244), .B(n1245), .Z(n1178) );
  NANDN U2499 ( .B(n1246), .A(n1247), .Z(n1244) );
  XOR U2500 ( .A(n1251), .B(\_MxM/Y0[18] ), .Z(\_MxM/Y1[17] ) );
  XNOR U2501 ( .A(n1252), .B(n1253), .Z(n1251) );
  AND U2502 ( .A(n667), .B(n1255), .Z(n1254) );
  XOR U2503 ( .A(n1249), .B(n1253), .Z(n1255) );
  XNOR U2504 ( .A(n1248), .B(n1253), .Z(n1249) );
  XNOR U2505 ( .A(n1208), .B(n1207), .Z(n1190) );
  XOR U2506 ( .A(n1258), .B(n1213), .Z(n1207) );
  XNOR U2507 ( .A(n1195), .B(n1260), .Z(n1196) );
  AND U2508 ( .A(n740), .B(n1194), .Z(n1260) );
  XOR U2509 ( .A(n1264), .B(n1197), .Z(n1259) );
  NAND U2510 ( .A(n1136), .B(n774), .Z(n1197) );
  IV U2511 ( .A(n1199), .Z(n1264) );
  XNOR U2512 ( .A(n1204), .B(n1205), .Z(n1201) );
  NANDN U2513 ( .B(n1020), .A(n854), .Z(n1205) );
  XNOR U2514 ( .A(n1203), .B(n1268), .Z(n1204) );
  AND U2515 ( .A(n814), .B(n1079), .Z(n1268) );
  XNOR U2516 ( .A(n1212), .B(n1206), .Z(n1258) );
  XOR U2517 ( .A(n1275), .B(n1214), .Z(n1212) );
  NAND U2518 ( .A(n1278), .B(n1279), .Z(n1215) );
  NANDN U2519 ( .B(n710), .A(n1280), .Z(n1279) );
  OR U2520 ( .A(n1281), .B(n1282), .Z(n1278) );
  XNOR U2521 ( .A(n1286), .B(n1232), .Z(n1222) );
  XNOR U2522 ( .A(n1219), .B(n1220), .Z(n1232) );
  NANDN U2523 ( .B(n835), .A(n1055), .Z(n1220) );
  XNOR U2524 ( .A(n1218), .B(n1287), .Z(n1219) );
  AND U2525 ( .A(n999), .B(n874), .Z(n1287) );
  XNOR U2526 ( .A(n1231), .B(n1221), .Z(n1286) );
  XNOR U2527 ( .A(n1226), .B(n1295), .Z(n1227) );
  AND U2528 ( .A(n898), .B(n982), .Z(n1295) );
  XOR U2529 ( .A(n1299), .B(n1228), .Z(n1294) );
  NAND U2530 ( .A(n928), .B(n941), .Z(n1228) );
  IV U2531 ( .A(n1230), .Z(n1299) );
  XNOR U2532 ( .A(n1235), .B(n1304), .Z(n1236) );
  AND U2533 ( .A(n1114), .B(n806), .Z(n1304) );
  XOR U2534 ( .A(n1308), .B(n1237), .Z(n1303) );
  NAND U2535 ( .A(n770), .B(n1176), .Z(n1237) );
  IV U2536 ( .A(n1239), .Z(n1308) );
  XNOR U2537 ( .A(n1246), .B(n1247), .Z(n1241) );
  NANDN U2538 ( .B(n709), .A(n1312), .Z(n1247) );
  XOR U2539 ( .A(n1245), .B(n1313), .Z(n1246) );
  AND U2540 ( .A(n1242), .B(n742), .Z(n1313) );
  NAND U2541 ( .A(n1314), .B(n1315), .Z(n1245) );
  NANDN U2542 ( .B(n1316), .A(n1317), .Z(n1314) );
  XOR U2543 ( .A(n1321), .B(\_MxM/Y0[17] ), .Z(\_MxM/Y1[16] ) );
  XNOR U2544 ( .A(n1322), .B(n1323), .Z(n1321) );
  AND U2545 ( .A(n667), .B(n1325), .Z(n1324) );
  XOR U2546 ( .A(n1319), .B(n1323), .Z(n1325) );
  XNOR U2547 ( .A(n1318), .B(n1323), .Z(n1319) );
  XNOR U2548 ( .A(n1274), .B(n1273), .Z(n1257) );
  XOR U2549 ( .A(n1328), .B(n1285), .Z(n1273) );
  XNOR U2550 ( .A(n1261), .B(n1330), .Z(n1262) );
  AND U2551 ( .A(n774), .B(n1194), .Z(n1330) );
  XOR U2552 ( .A(n1334), .B(n1263), .Z(n1329) );
  NAND U2553 ( .A(n1136), .B(n814), .Z(n1263) );
  IV U2554 ( .A(n1265), .Z(n1334) );
  XNOR U2555 ( .A(n1270), .B(n1271), .Z(n1267) );
  NANDN U2556 ( .B(n1020), .A(n898), .Z(n1271) );
  XNOR U2557 ( .A(n1269), .B(n1338), .Z(n1270) );
  AND U2558 ( .A(n854), .B(n1079), .Z(n1338) );
  XNOR U2559 ( .A(n1284), .B(n1272), .Z(n1328) );
  XNOR U2560 ( .A(n1345), .B(n1277), .Z(n1284) );
  XOR U2561 ( .A(n1346), .B(n1281), .Z(n1277) );
  NAND U2562 ( .A(n1280), .B(n740), .Z(n1281) );
  NANDN U2563 ( .B(n710), .A(n1348), .Z(n1347) );
  XNOR U2564 ( .A(n1357), .B(n1302), .Z(n1292) );
  XNOR U2565 ( .A(n1289), .B(n1290), .Z(n1302) );
  NANDN U2566 ( .B(n835), .A(n1114), .Z(n1290) );
  XNOR U2567 ( .A(n1288), .B(n1358), .Z(n1289) );
  AND U2568 ( .A(n1055), .B(n874), .Z(n1358) );
  XNOR U2569 ( .A(n1301), .B(n1291), .Z(n1357) );
  XNOR U2570 ( .A(n1296), .B(n1366), .Z(n1297) );
  AND U2571 ( .A(n941), .B(n982), .Z(n1366) );
  XOR U2572 ( .A(n1370), .B(n1298), .Z(n1365) );
  NAND U2573 ( .A(n928), .B(n999), .Z(n1298) );
  IV U2574 ( .A(n1300), .Z(n1370) );
  XNOR U2575 ( .A(n1305), .B(n1375), .Z(n1306) );
  AND U2576 ( .A(n1176), .B(n806), .Z(n1375) );
  XOR U2577 ( .A(n1379), .B(n1307), .Z(n1374) );
  NAND U2578 ( .A(n770), .B(n1242), .Z(n1307) );
  IV U2579 ( .A(n1309), .Z(n1379) );
  XNOR U2580 ( .A(n1316), .B(n1317), .Z(n1311) );
  NANDN U2581 ( .B(n709), .A(n1383), .Z(n1317) );
  XNOR U2582 ( .A(n1315), .B(n1384), .Z(n1316) );
  AND U2583 ( .A(n1312), .B(n742), .Z(n1384) );
  AND U2584 ( .A(n1385), .B(n1386), .Z(n1315) );
  NANDN U2585 ( .B(n1387), .A(n1388), .Z(n1385) );
  XOR U2586 ( .A(n1392), .B(\_MxM/Y0[16] ), .Z(\_MxM/Y1[15] ) );
  XNOR U2587 ( .A(n1393), .B(n1394), .Z(n1392) );
  AND U2588 ( .A(n667), .B(n1396), .Z(n1395) );
  XOR U2589 ( .A(n1390), .B(n1394), .Z(n1396) );
  XNOR U2590 ( .A(n1389), .B(n1394), .Z(n1390) );
  XNOR U2591 ( .A(n1344), .B(n1343), .Z(n1327) );
  XOR U2592 ( .A(n1400), .B(n1354), .Z(n1343) );
  XNOR U2593 ( .A(n1331), .B(n1402), .Z(n1332) );
  AND U2594 ( .A(n814), .B(n1194), .Z(n1402) );
  XOR U2595 ( .A(n1406), .B(n1333), .Z(n1401) );
  NAND U2596 ( .A(n1136), .B(n854), .Z(n1333) );
  IV U2597 ( .A(n1335), .Z(n1406) );
  XNOR U2598 ( .A(n1340), .B(n1341), .Z(n1337) );
  NANDN U2599 ( .B(n1020), .A(n941), .Z(n1341) );
  XNOR U2600 ( .A(n1339), .B(n1410), .Z(n1340) );
  AND U2601 ( .A(n898), .B(n1079), .Z(n1410) );
  XNOR U2602 ( .A(n1353), .B(n1342), .Z(n1400) );
  XNOR U2603 ( .A(n1417), .B(n1356), .Z(n1353) );
  NAND U2604 ( .A(n1280), .B(n774), .Z(n1351) );
  XNOR U2605 ( .A(n1349), .B(n1418), .Z(n1350) );
  AND U2606 ( .A(n740), .B(n1348), .Z(n1418) );
  XNOR U2607 ( .A(n1355), .B(n1352), .Z(n1417) );
  AND U2608 ( .A(n1426), .B(n1427), .Z(n1425) );
  NANDN U2609 ( .B(n710), .A(n1428), .Z(n1427) );
  OR U2610 ( .A(n1429), .B(n1430), .Z(n1426) );
  XNOR U2611 ( .A(n1434), .B(n1373), .Z(n1363) );
  XNOR U2612 ( .A(n1360), .B(n1361), .Z(n1373) );
  NANDN U2613 ( .B(n835), .A(n1176), .Z(n1361) );
  XNOR U2614 ( .A(n1359), .B(n1435), .Z(n1360) );
  AND U2615 ( .A(n1114), .B(n874), .Z(n1435) );
  XNOR U2616 ( .A(n1372), .B(n1362), .Z(n1434) );
  XNOR U2617 ( .A(n1367), .B(n1443), .Z(n1368) );
  AND U2618 ( .A(n999), .B(n982), .Z(n1443) );
  XOR U2619 ( .A(n1447), .B(n1369), .Z(n1442) );
  NAND U2620 ( .A(n928), .B(n1055), .Z(n1369) );
  IV U2621 ( .A(n1371), .Z(n1447) );
  XNOR U2622 ( .A(n1376), .B(n1452), .Z(n1377) );
  AND U2623 ( .A(n1242), .B(n806), .Z(n1452) );
  XOR U2624 ( .A(n1456), .B(n1378), .Z(n1451) );
  NAND U2625 ( .A(n770), .B(n1312), .Z(n1378) );
  IV U2626 ( .A(n1380), .Z(n1456) );
  XNOR U2627 ( .A(n1387), .B(n1388), .Z(n1382) );
  NANDN U2628 ( .B(n709), .A(n1460), .Z(n1388) );
  XNOR U2629 ( .A(n1386), .B(n1461), .Z(n1387) );
  AND U2630 ( .A(n1383), .B(n742), .Z(n1461) );
  ANDN U2631 ( .A(n1462), .B(n1463), .Z(n1386) );
  NANDN U2632 ( .B(n1464), .A(n1465), .Z(n1462) );
  XOR U2633 ( .A(n1469), .B(\_MxM/Y0[15] ), .Z(\_MxM/Y1[14] ) );
  XNOR U2634 ( .A(n1470), .B(n1471), .Z(n1469) );
  AND U2635 ( .A(n667), .B(n1473), .Z(n1472) );
  XOR U2636 ( .A(n1467), .B(n1471), .Z(n1473) );
  XNOR U2637 ( .A(n1466), .B(n1471), .Z(n1467) );
  XOR U2638 ( .A(n1399), .B(n1398), .Z(n1471) );
  XOR U2639 ( .A(n1474), .B(n1475), .Z(n1398) );
  XOR U2640 ( .A(n1476), .B(n1477), .Z(n1475) );
  XOR U2641 ( .A(n1478), .B(n1476), .Z(n1477) );
  IV U2642 ( .A(n1479), .Z(n1480) );
  XNOR U2643 ( .A(n1416), .B(n1415), .Z(n1399) );
  XOR U2644 ( .A(n1485), .B(n1424), .Z(n1415) );
  XNOR U2645 ( .A(n1403), .B(n1487), .Z(n1404) );
  AND U2646 ( .A(n854), .B(n1194), .Z(n1487) );
  XOR U2647 ( .A(n1491), .B(n1405), .Z(n1486) );
  NAND U2648 ( .A(n1136), .B(n898), .Z(n1405) );
  IV U2649 ( .A(n1407), .Z(n1491) );
  XNOR U2650 ( .A(n1412), .B(n1413), .Z(n1409) );
  NANDN U2651 ( .B(n1020), .A(n999), .Z(n1413) );
  XNOR U2652 ( .A(n1411), .B(n1495), .Z(n1412) );
  AND U2653 ( .A(n941), .B(n1079), .Z(n1495) );
  XNOR U2654 ( .A(n1423), .B(n1414), .Z(n1485) );
  XNOR U2655 ( .A(n1502), .B(n1433), .Z(n1423) );
  NAND U2656 ( .A(n1280), .B(n814), .Z(n1421) );
  XNOR U2657 ( .A(n1419), .B(n1503), .Z(n1420) );
  AND U2658 ( .A(n774), .B(n1348), .Z(n1503) );
  XNOR U2659 ( .A(n1432), .B(n1422), .Z(n1502) );
  XNOR U2660 ( .A(n1510), .B(n1431), .Z(n1432) );
  XNOR U2661 ( .A(n1514), .B(n1429), .Z(n1510) );
  NAND U2662 ( .A(n1428), .B(n740), .Z(n1429) );
  NANDN U2663 ( .B(n710), .A(n1516), .Z(n1515) );
  XNOR U2664 ( .A(n1520), .B(n1450), .Z(n1440) );
  XNOR U2665 ( .A(n1437), .B(n1438), .Z(n1450) );
  NANDN U2666 ( .B(n835), .A(n1242), .Z(n1438) );
  XNOR U2667 ( .A(n1436), .B(n1521), .Z(n1437) );
  AND U2668 ( .A(n1176), .B(n874), .Z(n1521) );
  XNOR U2669 ( .A(n1449), .B(n1439), .Z(n1520) );
  XNOR U2670 ( .A(n1444), .B(n1529), .Z(n1445) );
  AND U2671 ( .A(n1055), .B(n982), .Z(n1529) );
  XOR U2672 ( .A(n1533), .B(n1446), .Z(n1528) );
  NAND U2673 ( .A(n928), .B(n1114), .Z(n1446) );
  IV U2674 ( .A(n1448), .Z(n1533) );
  XNOR U2675 ( .A(n1453), .B(n1538), .Z(n1454) );
  AND U2676 ( .A(n1312), .B(n806), .Z(n1538) );
  XOR U2677 ( .A(n1542), .B(n1455), .Z(n1537) );
  NAND U2678 ( .A(n770), .B(n1383), .Z(n1455) );
  IV U2679 ( .A(n1457), .Z(n1542) );
  XNOR U2680 ( .A(n1464), .B(n1465), .Z(n1459) );
  NANDN U2681 ( .B(n709), .A(n1546), .Z(n1465) );
  AND U2682 ( .A(n1460), .B(n742), .Z(n1547) );
  NAND U2683 ( .A(n1548), .B(n1549), .Z(n1463) );
  NANDN U2684 ( .B(n1550), .A(n1551), .Z(n1548) );
  XOR U2685 ( .A(n1555), .B(\_MxM/Y0[14] ), .Z(\_MxM/Y1[13] ) );
  XNOR U2686 ( .A(n1556), .B(n1557), .Z(n1555) );
  AND U2687 ( .A(n667), .B(n1559), .Z(n1558) );
  XOR U2688 ( .A(n1553), .B(n1557), .Z(n1559) );
  XNOR U2689 ( .A(n1552), .B(n1557), .Z(n1553) );
  XNOR U2690 ( .A(n1484), .B(n1483), .Z(n1557) );
  XNOR U2691 ( .A(n1560), .B(n1479), .Z(n1483) );
  NAND U2692 ( .A(n1476), .B(n1563), .Z(n1481) );
  AND U2693 ( .A(n1564), .B(n1565), .Z(n1563) );
  NANDN U2694 ( .B(n710), .A(n1566), .Z(n1565) );
  NANDN U2695 ( .B(n1567), .A(n1568), .Z(n1564) );
  AND U2696 ( .A(n1569), .B(n1570), .Z(n1476) );
  NANDN U2697 ( .B(n1571), .A(n1572), .Z(n1570) );
  NANDN U2698 ( .B(n1573), .A(n1574), .Z(n1569) );
  XNOR U2699 ( .A(n1578), .B(n1509), .Z(n1500) );
  XNOR U2700 ( .A(n1488), .B(n1580), .Z(n1489) );
  AND U2701 ( .A(n898), .B(n1194), .Z(n1580) );
  XOR U2702 ( .A(n1584), .B(n1490), .Z(n1579) );
  NAND U2703 ( .A(n1136), .B(n941), .Z(n1490) );
  IV U2704 ( .A(n1492), .Z(n1584) );
  XNOR U2705 ( .A(n1497), .B(n1498), .Z(n1494) );
  NANDN U2706 ( .B(n1020), .A(n1055), .Z(n1498) );
  XNOR U2707 ( .A(n1496), .B(n1588), .Z(n1497) );
  AND U2708 ( .A(n999), .B(n1079), .Z(n1588) );
  XNOR U2709 ( .A(n1508), .B(n1499), .Z(n1578) );
  XOR U2710 ( .A(n1595), .B(n1513), .Z(n1508) );
  XNOR U2711 ( .A(n1505), .B(n1506), .Z(n1513) );
  NAND U2712 ( .A(n1280), .B(n854), .Z(n1506) );
  XNOR U2713 ( .A(n1504), .B(n1596), .Z(n1505) );
  AND U2714 ( .A(n814), .B(n1348), .Z(n1596) );
  XNOR U2715 ( .A(n1512), .B(n1507), .Z(n1595) );
  XNOR U2716 ( .A(n1517), .B(n1604), .Z(n1518) );
  AND U2717 ( .A(n740), .B(n1516), .Z(n1604) );
  XOR U2718 ( .A(n1608), .B(n1519), .Z(n1603) );
  NAND U2719 ( .A(n1428), .B(n774), .Z(n1519) );
  IV U2720 ( .A(n1511), .Z(n1608) );
  XNOR U2721 ( .A(n1612), .B(n1536), .Z(n1526) );
  XNOR U2722 ( .A(n1523), .B(n1524), .Z(n1536) );
  NANDN U2723 ( .B(n835), .A(n1312), .Z(n1524) );
  XNOR U2724 ( .A(n1522), .B(n1613), .Z(n1523) );
  AND U2725 ( .A(n1242), .B(n874), .Z(n1613) );
  XNOR U2726 ( .A(n1535), .B(n1525), .Z(n1612) );
  XNOR U2727 ( .A(n1530), .B(n1621), .Z(n1531) );
  AND U2728 ( .A(n1114), .B(n982), .Z(n1621) );
  XOR U2729 ( .A(n1625), .B(n1532), .Z(n1620) );
  NAND U2730 ( .A(n928), .B(n1176), .Z(n1532) );
  IV U2731 ( .A(n1534), .Z(n1625) );
  XNOR U2732 ( .A(n1539), .B(n1630), .Z(n1540) );
  AND U2733 ( .A(n1383), .B(n806), .Z(n1630) );
  XOR U2734 ( .A(n1634), .B(n1541), .Z(n1629) );
  NAND U2735 ( .A(n770), .B(n1460), .Z(n1541) );
  IV U2736 ( .A(n1543), .Z(n1634) );
  XNOR U2737 ( .A(n1550), .B(n1551), .Z(n1545) );
  NANDN U2738 ( .B(n709), .A(n1638), .Z(n1551) );
  XNOR U2739 ( .A(n1549), .B(n1639), .Z(n1550) );
  AND U2740 ( .A(n1546), .B(n742), .Z(n1639) );
  ANDN U2741 ( .A(n1640), .B(n1641), .Z(n1549) );
  NANDN U2742 ( .B(n1642), .A(n1643), .Z(n1640) );
  XOR U2743 ( .A(n1647), .B(\_MxM/Y0[13] ), .Z(\_MxM/Y1[12] ) );
  XNOR U2744 ( .A(n1648), .B(n1649), .Z(n1647) );
  AND U2745 ( .A(n667), .B(n1651), .Z(n1650) );
  XOR U2746 ( .A(n1645), .B(n1649), .Z(n1651) );
  XNOR U2747 ( .A(n1644), .B(n1649), .Z(n1645) );
  XNOR U2748 ( .A(n1577), .B(n1576), .Z(n1649) );
  XNOR U2749 ( .A(n1652), .B(n1562), .Z(n1576) );
  XNOR U2750 ( .A(n1568), .B(n1567), .Z(n1562) );
  OR U2751 ( .A(n1653), .B(n1654), .Z(n1567) );
  XNOR U2752 ( .A(n1571), .B(n1572), .Z(n1568) );
  XOR U2753 ( .A(n1658), .B(n1573), .Z(n1571) );
  NAND U2754 ( .A(n740), .B(n1566), .Z(n1573) );
  NANDN U2755 ( .B(n1574), .A(n1659), .Z(n1658) );
  NANDN U2756 ( .B(n710), .A(n1660), .Z(n1659) );
  XNOR U2757 ( .A(n1669), .B(n1602), .Z(n1593) );
  XNOR U2758 ( .A(n1581), .B(n1671), .Z(n1582) );
  AND U2759 ( .A(n941), .B(n1194), .Z(n1671) );
  XOR U2760 ( .A(n1675), .B(n1583), .Z(n1670) );
  NAND U2761 ( .A(n1136), .B(n999), .Z(n1583) );
  IV U2762 ( .A(n1585), .Z(n1675) );
  XNOR U2763 ( .A(n1590), .B(n1591), .Z(n1587) );
  NANDN U2764 ( .B(n1020), .A(n1114), .Z(n1591) );
  XNOR U2765 ( .A(n1589), .B(n1679), .Z(n1590) );
  AND U2766 ( .A(n1055), .B(n1079), .Z(n1679) );
  XNOR U2767 ( .A(n1601), .B(n1592), .Z(n1669) );
  XOR U2768 ( .A(n1686), .B(n1611), .Z(n1601) );
  XNOR U2769 ( .A(n1598), .B(n1599), .Z(n1611) );
  NAND U2770 ( .A(n1280), .B(n898), .Z(n1599) );
  XNOR U2771 ( .A(n1597), .B(n1687), .Z(n1598) );
  AND U2772 ( .A(n854), .B(n1348), .Z(n1687) );
  XNOR U2773 ( .A(n1610), .B(n1600), .Z(n1686) );
  XNOR U2774 ( .A(n1605), .B(n1695), .Z(n1606) );
  AND U2775 ( .A(n774), .B(n1516), .Z(n1695) );
  XOR U2776 ( .A(n1699), .B(n1607), .Z(n1694) );
  NAND U2777 ( .A(n1428), .B(n814), .Z(n1607) );
  IV U2778 ( .A(n1609), .Z(n1699) );
  XNOR U2779 ( .A(n1703), .B(n1628), .Z(n1618) );
  XNOR U2780 ( .A(n1615), .B(n1616), .Z(n1628) );
  NANDN U2781 ( .B(n835), .A(n1383), .Z(n1616) );
  XNOR U2782 ( .A(n1614), .B(n1704), .Z(n1615) );
  AND U2783 ( .A(n1312), .B(n874), .Z(n1704) );
  XNOR U2784 ( .A(n1627), .B(n1617), .Z(n1703) );
  XNOR U2785 ( .A(n1622), .B(n1712), .Z(n1623) );
  AND U2786 ( .A(n1176), .B(n982), .Z(n1712) );
  XOR U2787 ( .A(n1716), .B(n1624), .Z(n1711) );
  NAND U2788 ( .A(n928), .B(n1242), .Z(n1624) );
  IV U2789 ( .A(n1626), .Z(n1716) );
  XNOR U2790 ( .A(n1631), .B(n1721), .Z(n1632) );
  AND U2791 ( .A(n1460), .B(n806), .Z(n1721) );
  XOR U2792 ( .A(n1725), .B(n1633), .Z(n1720) );
  NAND U2793 ( .A(n770), .B(n1546), .Z(n1633) );
  IV U2794 ( .A(n1635), .Z(n1725) );
  XOR U2795 ( .A(n1726), .B(n1727), .Z(n1635) );
  ANDN U2796 ( .A(n1728), .B(n1729), .Z(n1727) );
  XOR U2797 ( .A(n1726), .B(n1730), .Z(n1728) );
  XNOR U2798 ( .A(n1642), .B(n1643), .Z(n1637) );
  NANDN U2799 ( .B(n709), .A(n1731), .Z(n1643) );
  AND U2800 ( .A(n1638), .B(n742), .Z(n1732) );
  NAND U2801 ( .A(n1733), .B(n1734), .Z(n1641) );
  NANDN U2802 ( .B(n1735), .A(n1736), .Z(n1733) );
  XOR U2803 ( .A(n1740), .B(\_MxM/Y0[12] ), .Z(\_MxM/Y1[11] ) );
  XNOR U2804 ( .A(n1741), .B(n1742), .Z(n1740) );
  AND U2805 ( .A(n667), .B(n1744), .Z(n1743) );
  XOR U2806 ( .A(n1738), .B(n1742), .Z(n1744) );
  XNOR U2807 ( .A(n1737), .B(n1742), .Z(n1738) );
  XNOR U2808 ( .A(n1666), .B(n1665), .Z(n1742) );
  XNOR U2809 ( .A(n1745), .B(n1668), .Z(n1665) );
  XOR U2810 ( .A(n1654), .B(n1653), .Z(n1668) );
  NANDN U2811 ( .B(n1746), .A(n1747), .Z(n1653) );
  XOR U2812 ( .A(n1657), .B(n1656), .Z(n1654) );
  XOR U2813 ( .A(n1655), .B(n1748), .Z(n1656) );
  AND U2814 ( .A(n1749), .B(n1750), .Z(n1748) );
  NANDN U2815 ( .B(n710), .A(n1751), .Z(n1750) );
  OR U2816 ( .A(n1752), .B(n1753), .Z(n1749) );
  NAND U2817 ( .A(n774), .B(n1566), .Z(n1663) );
  XNOR U2818 ( .A(n1661), .B(n1756), .Z(n1662) );
  AND U2819 ( .A(n1660), .B(n740), .Z(n1756) );
  XNOR U2820 ( .A(n1765), .B(n1693), .Z(n1684) );
  XNOR U2821 ( .A(n1672), .B(n1767), .Z(n1673) );
  AND U2822 ( .A(n999), .B(n1194), .Z(n1767) );
  XOR U2823 ( .A(n1771), .B(n1674), .Z(n1766) );
  NAND U2824 ( .A(n1136), .B(n1055), .Z(n1674) );
  IV U2825 ( .A(n1676), .Z(n1771) );
  XNOR U2826 ( .A(n1681), .B(n1682), .Z(n1678) );
  NANDN U2827 ( .B(n1020), .A(n1176), .Z(n1682) );
  XNOR U2828 ( .A(n1680), .B(n1775), .Z(n1681) );
  AND U2829 ( .A(n1114), .B(n1079), .Z(n1775) );
  XNOR U2830 ( .A(n1692), .B(n1683), .Z(n1765) );
  XOR U2831 ( .A(n1782), .B(n1702), .Z(n1692) );
  XNOR U2832 ( .A(n1689), .B(n1690), .Z(n1702) );
  NAND U2833 ( .A(n1280), .B(n941), .Z(n1690) );
  XNOR U2834 ( .A(n1688), .B(n1783), .Z(n1689) );
  AND U2835 ( .A(n898), .B(n1348), .Z(n1783) );
  XNOR U2836 ( .A(n1701), .B(n1691), .Z(n1782) );
  XNOR U2837 ( .A(n1696), .B(n1791), .Z(n1697) );
  AND U2838 ( .A(n814), .B(n1516), .Z(n1791) );
  XOR U2839 ( .A(n1795), .B(n1698), .Z(n1790) );
  NAND U2840 ( .A(n1428), .B(n854), .Z(n1698) );
  IV U2841 ( .A(n1700), .Z(n1795) );
  XNOR U2842 ( .A(n1799), .B(n1719), .Z(n1709) );
  XNOR U2843 ( .A(n1706), .B(n1707), .Z(n1719) );
  NANDN U2844 ( .B(n835), .A(n1460), .Z(n1707) );
  XNOR U2845 ( .A(n1705), .B(n1800), .Z(n1706) );
  AND U2846 ( .A(n1383), .B(n874), .Z(n1800) );
  XNOR U2847 ( .A(n1718), .B(n1708), .Z(n1799) );
  XNOR U2848 ( .A(n1713), .B(n1808), .Z(n1714) );
  AND U2849 ( .A(n1242), .B(n982), .Z(n1808) );
  XOR U2850 ( .A(n1812), .B(n1715), .Z(n1807) );
  NAND U2851 ( .A(n928), .B(n1312), .Z(n1715) );
  IV U2852 ( .A(n1717), .Z(n1812) );
  XNOR U2853 ( .A(n1722), .B(n1817), .Z(n1723) );
  AND U2854 ( .A(n1546), .B(n806), .Z(n1817) );
  XOR U2855 ( .A(n1821), .B(n1724), .Z(n1816) );
  NAND U2856 ( .A(n770), .B(n1638), .Z(n1724) );
  IV U2857 ( .A(n1726), .Z(n1821) );
  XNOR U2858 ( .A(n1735), .B(n1736), .Z(n1730) );
  NANDN U2859 ( .B(n709), .A(n1825), .Z(n1736) );
  XNOR U2860 ( .A(n1734), .B(n1826), .Z(n1735) );
  AND U2861 ( .A(n1731), .B(n742), .Z(n1826) );
  ANDN U2862 ( .A(n1827), .B(n1828), .Z(n1734) );
  NANDN U2863 ( .B(n1829), .A(n1830), .Z(n1827) );
  XOR U2864 ( .A(n1834), .B(\_MxM/Y0[11] ), .Z(\_MxM/Y1[10] ) );
  XNOR U2865 ( .A(n1835), .B(n1836), .Z(n1834) );
  AND U2866 ( .A(n667), .B(n1838), .Z(n1837) );
  XOR U2867 ( .A(n1832), .B(n1836), .Z(n1838) );
  XNOR U2868 ( .A(n1831), .B(n1836), .Z(n1832) );
  XNOR U2869 ( .A(n1762), .B(n1761), .Z(n1836) );
  XNOR U2870 ( .A(n1839), .B(n1764), .Z(n1761) );
  XNOR U2871 ( .A(n1746), .B(n1747), .Z(n1764) );
  XOR U2872 ( .A(n1755), .B(n1754), .Z(n1746) );
  XNOR U2873 ( .A(n1843), .B(n1844), .Z(n1754) );
  ANDN U2874 ( .A(n1847), .B(n1848), .Z(n1846) );
  XOR U2875 ( .A(n1845), .B(n1849), .Z(n1847) );
  XNOR U2876 ( .A(n1850), .B(n1752), .Z(n1843) );
  NAND U2877 ( .A(n740), .B(n1751), .Z(n1752) );
  NANDN U2878 ( .B(n710), .A(n1852), .Z(n1851) );
  NAND U2879 ( .A(n814), .B(n1566), .Z(n1759) );
  XNOR U2880 ( .A(n1757), .B(n1856), .Z(n1758) );
  AND U2881 ( .A(n1660), .B(n774), .Z(n1856) );
  XNOR U2882 ( .A(n1865), .B(n1789), .Z(n1780) );
  XNOR U2883 ( .A(n1768), .B(n1867), .Z(n1769) );
  AND U2884 ( .A(n1055), .B(n1194), .Z(n1867) );
  XOR U2885 ( .A(n1871), .B(n1770), .Z(n1866) );
  NAND U2886 ( .A(n1136), .B(n1114), .Z(n1770) );
  IV U2887 ( .A(n1772), .Z(n1871) );
  XNOR U2888 ( .A(n1777), .B(n1778), .Z(n1774) );
  NANDN U2889 ( .B(n1020), .A(n1242), .Z(n1778) );
  XNOR U2890 ( .A(n1776), .B(n1875), .Z(n1777) );
  AND U2891 ( .A(n1176), .B(n1079), .Z(n1875) );
  XNOR U2892 ( .A(n1788), .B(n1779), .Z(n1865) );
  XOR U2893 ( .A(n1882), .B(n1798), .Z(n1788) );
  XNOR U2894 ( .A(n1785), .B(n1786), .Z(n1798) );
  NAND U2895 ( .A(n1280), .B(n999), .Z(n1786) );
  XNOR U2896 ( .A(n1784), .B(n1883), .Z(n1785) );
  AND U2897 ( .A(n941), .B(n1348), .Z(n1883) );
  XNOR U2898 ( .A(n1797), .B(n1787), .Z(n1882) );
  XNOR U2899 ( .A(n1792), .B(n1891), .Z(n1793) );
  AND U2900 ( .A(n854), .B(n1516), .Z(n1891) );
  XOR U2901 ( .A(n1895), .B(n1794), .Z(n1890) );
  NAND U2902 ( .A(n1428), .B(n898), .Z(n1794) );
  IV U2903 ( .A(n1796), .Z(n1895) );
  XNOR U2904 ( .A(n1899), .B(n1815), .Z(n1805) );
  XNOR U2905 ( .A(n1802), .B(n1803), .Z(n1815) );
  NANDN U2906 ( .B(n835), .A(n1546), .Z(n1803) );
  XNOR U2907 ( .A(n1801), .B(n1900), .Z(n1802) );
  AND U2908 ( .A(n1460), .B(n874), .Z(n1900) );
  XNOR U2909 ( .A(n1814), .B(n1804), .Z(n1899) );
  XNOR U2910 ( .A(n1809), .B(n1908), .Z(n1810) );
  AND U2911 ( .A(n1312), .B(n982), .Z(n1908) );
  XOR U2912 ( .A(n1912), .B(n1811), .Z(n1907) );
  NAND U2913 ( .A(n928), .B(n1383), .Z(n1811) );
  IV U2914 ( .A(n1813), .Z(n1912) );
  XNOR U2915 ( .A(n1818), .B(n1917), .Z(n1819) );
  AND U2916 ( .A(n1638), .B(n806), .Z(n1917) );
  XOR U2917 ( .A(n1921), .B(n1820), .Z(n1916) );
  NAND U2918 ( .A(n770), .B(n1731), .Z(n1820) );
  IV U2919 ( .A(n1822), .Z(n1921) );
  XNOR U2920 ( .A(n1829), .B(n1830), .Z(n1824) );
  NANDN U2921 ( .B(n709), .A(n1925), .Z(n1830) );
  AND U2922 ( .A(n1825), .B(n742), .Z(n1926) );
  NAND U2923 ( .A(n1927), .B(n1928), .Z(n1828) );
  NANDN U2924 ( .B(n1929), .A(n1930), .Z(n1927) );
  XNOR U2925 ( .A(n1934), .B(n1935), .Z(n651) );
  AND U2926 ( .A(n667), .B(n1937), .Z(n1936) );
  XOR U2927 ( .A(n1932), .B(n1935), .Z(n1937) );
  XNOR U2928 ( .A(n1931), .B(n1935), .Z(n1932) );
  XNOR U2929 ( .A(n1862), .B(n1861), .Z(n1935) );
  XNOR U2930 ( .A(n1938), .B(n1864), .Z(n1861) );
  XNOR U2931 ( .A(n1842), .B(n1841), .Z(n1864) );
  XNOR U2932 ( .A(n1840), .B(n1939), .Z(n1841) );
  AND U2933 ( .A(n1940), .B(n1941), .Z(n1939) );
  OR U2934 ( .A(n1942), .B(n1943), .Z(n1941) );
  AND U2935 ( .A(n1944), .B(n1945), .Z(n1940) );
  NANDN U2936 ( .B(n710), .A(n1946), .Z(n1945) );
  NAND U2937 ( .A(n1947), .B(n1948), .Z(n1944) );
  XNOR U2938 ( .A(n1853), .B(n1953), .Z(n1854) );
  AND U2939 ( .A(n1852), .B(n740), .Z(n1953) );
  XOR U2940 ( .A(n1957), .B(n1855), .Z(n1952) );
  NAND U2941 ( .A(n774), .B(n1751), .Z(n1855) );
  IV U2942 ( .A(n1845), .Z(n1957) );
  XNOR U2943 ( .A(n1858), .B(n1859), .Z(n1849) );
  NAND U2944 ( .A(n854), .B(n1566), .Z(n1859) );
  XNOR U2945 ( .A(n1857), .B(n1961), .Z(n1858) );
  AND U2946 ( .A(n1660), .B(n814), .Z(n1961) );
  XNOR U2947 ( .A(n1970), .B(n1889), .Z(n1880) );
  XNOR U2948 ( .A(n1868), .B(n1972), .Z(n1869) );
  AND U2949 ( .A(n1114), .B(n1194), .Z(n1972) );
  XOR U2950 ( .A(n1976), .B(n1870), .Z(n1971) );
  NAND U2951 ( .A(n1136), .B(n1176), .Z(n1870) );
  IV U2952 ( .A(n1872), .Z(n1976) );
  XNOR U2953 ( .A(n1877), .B(n1878), .Z(n1874) );
  NANDN U2954 ( .B(n1020), .A(n1312), .Z(n1878) );
  XNOR U2955 ( .A(n1876), .B(n1980), .Z(n1877) );
  AND U2956 ( .A(n1242), .B(n1079), .Z(n1980) );
  XNOR U2957 ( .A(n1888), .B(n1879), .Z(n1970) );
  XOR U2958 ( .A(n1987), .B(n1898), .Z(n1888) );
  XNOR U2959 ( .A(n1885), .B(n1886), .Z(n1898) );
  NAND U2960 ( .A(n1280), .B(n1055), .Z(n1886) );
  XNOR U2961 ( .A(n1884), .B(n1988), .Z(n1885) );
  AND U2962 ( .A(n999), .B(n1348), .Z(n1988) );
  XNOR U2963 ( .A(n1897), .B(n1887), .Z(n1987) );
  XNOR U2964 ( .A(n1892), .B(n1996), .Z(n1893) );
  AND U2965 ( .A(n898), .B(n1516), .Z(n1996) );
  XOR U2966 ( .A(n2000), .B(n1894), .Z(n1995) );
  NAND U2967 ( .A(n1428), .B(n941), .Z(n1894) );
  IV U2968 ( .A(n1896), .Z(n2000) );
  XNOR U2969 ( .A(n2004), .B(n1915), .Z(n1905) );
  XNOR U2970 ( .A(n1902), .B(n1903), .Z(n1915) );
  NANDN U2971 ( .B(n835), .A(n1638), .Z(n1903) );
  XNOR U2972 ( .A(n1901), .B(n2005), .Z(n1902) );
  AND U2973 ( .A(n1546), .B(n874), .Z(n2005) );
  XNOR U2974 ( .A(n1914), .B(n1904), .Z(n2004) );
  XNOR U2975 ( .A(n1909), .B(n2013), .Z(n1910) );
  AND U2976 ( .A(n1383), .B(n982), .Z(n2013) );
  XOR U2977 ( .A(n2017), .B(n1911), .Z(n2012) );
  NAND U2978 ( .A(n928), .B(n1460), .Z(n1911) );
  IV U2979 ( .A(n1913), .Z(n2017) );
  XNOR U2980 ( .A(n1918), .B(n2022), .Z(n1919) );
  AND U2981 ( .A(n1731), .B(n806), .Z(n2022) );
  XOR U2982 ( .A(n2026), .B(n1920), .Z(n2021) );
  NAND U2983 ( .A(n770), .B(n1825), .Z(n1920) );
  IV U2984 ( .A(n1922), .Z(n2026) );
  XNOR U2985 ( .A(n1929), .B(n1930), .Z(n1924) );
  NANDN U2986 ( .B(n709), .A(n2030), .Z(n1930) );
  XNOR U2987 ( .A(n1928), .B(n2031), .Z(n1929) );
  AND U2988 ( .A(n1925), .B(n742), .Z(n2031) );
  ANDN U2989 ( .A(n2032), .B(n2033), .Z(n1928) );
  NANDN U2990 ( .B(n2034), .A(n2035), .Z(n2032) );
  XNOR U2991 ( .A(n2039), .B(n2040), .Z(n652) );
  AND U2992 ( .A(n667), .B(n2042), .Z(n2041) );
  XOR U2993 ( .A(n2037), .B(n2040), .Z(n2042) );
  XNOR U2994 ( .A(n2036), .B(n2040), .Z(n2037) );
  XNOR U2995 ( .A(n1967), .B(n1966), .Z(n2040) );
  XNOR U2996 ( .A(n2043), .B(n1969), .Z(n1966) );
  XNOR U2997 ( .A(n1951), .B(n1950), .Z(n1969) );
  XNOR U2998 ( .A(n2044), .B(n1947), .Z(n1950) );
  XNOR U2999 ( .A(n2045), .B(n1942), .Z(n1947) );
  NAND U3000 ( .A(n740), .B(n1946), .Z(n1942) );
  NANDN U3001 ( .B(n710), .A(n2047), .Z(n2046) );
  XNOR U3002 ( .A(n1948), .B(n1949), .Z(n2044) );
  XNOR U3003 ( .A(n1954), .B(n2058), .Z(n1955) );
  AND U3004 ( .A(n1852), .B(n774), .Z(n2058) );
  XOR U3005 ( .A(n2062), .B(n1956), .Z(n2057) );
  NAND U3006 ( .A(n814), .B(n1751), .Z(n1956) );
  IV U3007 ( .A(n1958), .Z(n2062) );
  XNOR U3008 ( .A(n1963), .B(n1964), .Z(n1960) );
  NAND U3009 ( .A(n898), .B(n1566), .Z(n1964) );
  XNOR U3010 ( .A(n1962), .B(n2066), .Z(n1963) );
  AND U3011 ( .A(n1660), .B(n854), .Z(n2066) );
  XNOR U3012 ( .A(n2075), .B(n1994), .Z(n1985) );
  XNOR U3013 ( .A(n1973), .B(n2077), .Z(n1974) );
  AND U3014 ( .A(n1176), .B(n1194), .Z(n2077) );
  XOR U3015 ( .A(n2081), .B(n1975), .Z(n2076) );
  NAND U3016 ( .A(n1136), .B(n1242), .Z(n1975) );
  IV U3017 ( .A(n1977), .Z(n2081) );
  XNOR U3018 ( .A(n1982), .B(n1983), .Z(n1979) );
  NANDN U3019 ( .B(n1020), .A(n1383), .Z(n1983) );
  XNOR U3020 ( .A(n1981), .B(n2085), .Z(n1982) );
  AND U3021 ( .A(n1312), .B(n1079), .Z(n2085) );
  XNOR U3022 ( .A(n1993), .B(n1984), .Z(n2075) );
  XOR U3023 ( .A(n2092), .B(n2003), .Z(n1993) );
  XNOR U3024 ( .A(n1990), .B(n1991), .Z(n2003) );
  NAND U3025 ( .A(n1280), .B(n1114), .Z(n1991) );
  XNOR U3026 ( .A(n1989), .B(n2093), .Z(n1990) );
  AND U3027 ( .A(n1055), .B(n1348), .Z(n2093) );
  XNOR U3028 ( .A(n2002), .B(n1992), .Z(n2092) );
  XNOR U3029 ( .A(n1997), .B(n2101), .Z(n1998) );
  AND U3030 ( .A(n941), .B(n1516), .Z(n2101) );
  XOR U3031 ( .A(n2105), .B(n1999), .Z(n2100) );
  NAND U3032 ( .A(n1428), .B(n999), .Z(n1999) );
  IV U3033 ( .A(n2001), .Z(n2105) );
  XNOR U3034 ( .A(n2109), .B(n2020), .Z(n2010) );
  XNOR U3035 ( .A(n2007), .B(n2008), .Z(n2020) );
  NANDN U3036 ( .B(n835), .A(n1731), .Z(n2008) );
  XNOR U3037 ( .A(n2006), .B(n2110), .Z(n2007) );
  AND U3038 ( .A(n1638), .B(n874), .Z(n2110) );
  XNOR U3039 ( .A(n2019), .B(n2009), .Z(n2109) );
  XNOR U3040 ( .A(n2014), .B(n2118), .Z(n2015) );
  AND U3041 ( .A(n1460), .B(n982), .Z(n2118) );
  XOR U3042 ( .A(n2122), .B(n2016), .Z(n2117) );
  NAND U3043 ( .A(n928), .B(n1546), .Z(n2016) );
  IV U3044 ( .A(n2018), .Z(n2122) );
  XNOR U3045 ( .A(n2023), .B(n2127), .Z(n2024) );
  AND U3046 ( .A(n1825), .B(n806), .Z(n2127) );
  XOR U3047 ( .A(n2131), .B(n2025), .Z(n2126) );
  NAND U3048 ( .A(n770), .B(n1925), .Z(n2025) );
  IV U3049 ( .A(n2027), .Z(n2131) );
  XNOR U3050 ( .A(n2034), .B(n2035), .Z(n2029) );
  NANDN U3051 ( .B(n709), .A(n2135), .Z(n2035) );
  AND U3052 ( .A(n2030), .B(n742), .Z(n2136) );
  NAND U3053 ( .A(n2137), .B(n2138), .Z(n2033) );
  NANDN U3054 ( .B(n2139), .A(n2140), .Z(n2137) );
  XNOR U3055 ( .A(n2144), .B(n2145), .Z(n653) );
  AND U3056 ( .A(n667), .B(n2147), .Z(n2146) );
  XOR U3057 ( .A(n2142), .B(n2145), .Z(n2147) );
  XNOR U3058 ( .A(n2141), .B(n2145), .Z(n2142) );
  XNOR U3059 ( .A(n2072), .B(n2071), .Z(n2145) );
  XNOR U3060 ( .A(n2148), .B(n2074), .Z(n2071) );
  XNOR U3061 ( .A(n2053), .B(n2052), .Z(n2074) );
  XNOR U3062 ( .A(n2149), .B(n2056), .Z(n2052) );
  XNOR U3063 ( .A(n2049), .B(n2050), .Z(n2056) );
  NAND U3064 ( .A(n774), .B(n1946), .Z(n2050) );
  XNOR U3065 ( .A(n2048), .B(n2150), .Z(n2049) );
  AND U3066 ( .A(n2047), .B(n740), .Z(n2150) );
  XNOR U3067 ( .A(n2055), .B(n2051), .Z(n2149) );
  AND U3068 ( .A(n2158), .B(n2159), .Z(n2157) );
  NANDN U3069 ( .B(n710), .A(n2160), .Z(n2159) );
  OR U3070 ( .A(n2161), .B(n2162), .Z(n2158) );
  XNOR U3071 ( .A(n2059), .B(n2167), .Z(n2060) );
  AND U3072 ( .A(n1852), .B(n814), .Z(n2167) );
  XOR U3073 ( .A(n2171), .B(n2061), .Z(n2166) );
  NAND U3074 ( .A(n854), .B(n1751), .Z(n2061) );
  IV U3075 ( .A(n2063), .Z(n2171) );
  XNOR U3076 ( .A(n2068), .B(n2069), .Z(n2065) );
  NAND U3077 ( .A(n941), .B(n1566), .Z(n2069) );
  XNOR U3078 ( .A(n2067), .B(n2175), .Z(n2068) );
  AND U3079 ( .A(n1660), .B(n898), .Z(n2175) );
  XNOR U3080 ( .A(n2185), .B(n2182), .Z(n2184) );
  XNOR U3081 ( .A(n2186), .B(n2099), .Z(n2090) );
  XNOR U3082 ( .A(n2078), .B(n2188), .Z(n2079) );
  AND U3083 ( .A(n1242), .B(n1194), .Z(n2188) );
  XOR U3084 ( .A(n2192), .B(n2080), .Z(n2187) );
  NAND U3085 ( .A(n1136), .B(n1312), .Z(n2080) );
  IV U3086 ( .A(n2082), .Z(n2192) );
  XNOR U3087 ( .A(n2087), .B(n2088), .Z(n2084) );
  NANDN U3088 ( .B(n1020), .A(n1460), .Z(n2088) );
  XNOR U3089 ( .A(n2086), .B(n2196), .Z(n2087) );
  AND U3090 ( .A(n1383), .B(n1079), .Z(n2196) );
  XNOR U3091 ( .A(n2098), .B(n2089), .Z(n2186) );
  XOR U3092 ( .A(n2203), .B(n2108), .Z(n2098) );
  XNOR U3093 ( .A(n2095), .B(n2096), .Z(n2108) );
  NAND U3094 ( .A(n1280), .B(n1176), .Z(n2096) );
  XNOR U3095 ( .A(n2094), .B(n2204), .Z(n2095) );
  AND U3096 ( .A(n1114), .B(n1348), .Z(n2204) );
  XNOR U3097 ( .A(n2107), .B(n2097), .Z(n2203) );
  XNOR U3098 ( .A(n2102), .B(n2212), .Z(n2103) );
  AND U3099 ( .A(n999), .B(n1516), .Z(n2212) );
  XOR U3100 ( .A(n2216), .B(n2104), .Z(n2211) );
  NAND U3101 ( .A(n1428), .B(n1055), .Z(n2104) );
  IV U3102 ( .A(n2106), .Z(n2216) );
  XNOR U3103 ( .A(n2220), .B(n2125), .Z(n2115) );
  XNOR U3104 ( .A(n2112), .B(n2113), .Z(n2125) );
  NANDN U3105 ( .B(n835), .A(n1825), .Z(n2113) );
  XNOR U3106 ( .A(n2111), .B(n2221), .Z(n2112) );
  AND U3107 ( .A(n1731), .B(n874), .Z(n2221) );
  XNOR U3108 ( .A(n2124), .B(n2114), .Z(n2220) );
  XNOR U3109 ( .A(n2119), .B(n2229), .Z(n2120) );
  AND U3110 ( .A(n1546), .B(n982), .Z(n2229) );
  XOR U3111 ( .A(n2233), .B(n2121), .Z(n2228) );
  NAND U3112 ( .A(n928), .B(n1638), .Z(n2121) );
  IV U3113 ( .A(n2123), .Z(n2233) );
  XNOR U3114 ( .A(n2128), .B(n2238), .Z(n2129) );
  AND U3115 ( .A(n1925), .B(n806), .Z(n2238) );
  XOR U3116 ( .A(n2242), .B(n2130), .Z(n2237) );
  NAND U3117 ( .A(n770), .B(n2030), .Z(n2130) );
  IV U3118 ( .A(n2132), .Z(n2242) );
  XNOR U3119 ( .A(n2139), .B(n2140), .Z(n2134) );
  NANDN U3120 ( .B(n709), .A(n2246), .Z(n2140) );
  XNOR U3121 ( .A(n2138), .B(n2247), .Z(n2139) );
  AND U3122 ( .A(n2135), .B(n742), .Z(n2247) );
  ANDN U3123 ( .A(n2248), .B(n2249), .Z(n2138) );
  NANDN U3124 ( .B(n2250), .A(n2251), .Z(n2248) );
  XNOR U3125 ( .A(n2255), .B(n2256), .Z(n654) );
  AND U3126 ( .A(n667), .B(n2258), .Z(n2257) );
  XOR U3127 ( .A(n2253), .B(n2256), .Z(n2258) );
  XNOR U3128 ( .A(n2252), .B(n2256), .Z(n2253) );
  XNOR U3129 ( .A(n2181), .B(n2180), .Z(n2256) );
  XNOR U3130 ( .A(n2259), .B(n2185), .Z(n2180) );
  XNOR U3131 ( .A(n2156), .B(n2155), .Z(n2185) );
  XNOR U3132 ( .A(n2260), .B(n2165), .Z(n2155) );
  XNOR U3133 ( .A(n2152), .B(n2153), .Z(n2165) );
  NAND U3134 ( .A(n814), .B(n1946), .Z(n2153) );
  XNOR U3135 ( .A(n2151), .B(n2261), .Z(n2152) );
  AND U3136 ( .A(n2047), .B(n774), .Z(n2261) );
  XNOR U3137 ( .A(n2164), .B(n2154), .Z(n2260) );
  XNOR U3138 ( .A(n2268), .B(n2163), .Z(n2164) );
  XNOR U3139 ( .A(n2272), .B(n2161), .Z(n2268) );
  NAND U3140 ( .A(n740), .B(n2160), .Z(n2161) );
  NANDN U3141 ( .B(n710), .A(n2274), .Z(n2273) );
  XNOR U3142 ( .A(n2168), .B(n2279), .Z(n2169) );
  AND U3143 ( .A(n1852), .B(n854), .Z(n2279) );
  XOR U3144 ( .A(n2283), .B(n2170), .Z(n2278) );
  NAND U3145 ( .A(n898), .B(n1751), .Z(n2170) );
  IV U3146 ( .A(n2172), .Z(n2283) );
  XNOR U3147 ( .A(n2177), .B(n2178), .Z(n2174) );
  NAND U3148 ( .A(n999), .B(n1566), .Z(n2178) );
  XNOR U3149 ( .A(n2176), .B(n2287), .Z(n2177) );
  AND U3150 ( .A(n1660), .B(n941), .Z(n2287) );
  XNOR U3151 ( .A(n2183), .B(n2179), .Z(n2259) );
  XOR U3152 ( .A(n2298), .B(n2299), .Z(n2294) );
  NANDN U3153 ( .B(n2300), .A(n2301), .Z(n2298) );
  XNOR U3154 ( .A(n2302), .B(n2210), .Z(n2201) );
  XNOR U3155 ( .A(n2189), .B(n2304), .Z(n2190) );
  AND U3156 ( .A(n1312), .B(n1194), .Z(n2304) );
  XOR U3157 ( .A(n2308), .B(n2191), .Z(n2303) );
  NAND U3158 ( .A(n1136), .B(n1383), .Z(n2191) );
  IV U3159 ( .A(n2193), .Z(n2308) );
  XNOR U3160 ( .A(n2198), .B(n2199), .Z(n2195) );
  NANDN U3161 ( .B(n1020), .A(n1546), .Z(n2199) );
  XNOR U3162 ( .A(n2197), .B(n2312), .Z(n2198) );
  AND U3163 ( .A(n1460), .B(n1079), .Z(n2312) );
  XNOR U3164 ( .A(n2209), .B(n2200), .Z(n2302) );
  XOR U3165 ( .A(n2319), .B(n2219), .Z(n2209) );
  XNOR U3166 ( .A(n2206), .B(n2207), .Z(n2219) );
  NAND U3167 ( .A(n1280), .B(n1242), .Z(n2207) );
  XNOR U3168 ( .A(n2205), .B(n2320), .Z(n2206) );
  AND U3169 ( .A(n1176), .B(n1348), .Z(n2320) );
  XNOR U3170 ( .A(n2218), .B(n2208), .Z(n2319) );
  XNOR U3171 ( .A(n2213), .B(n2328), .Z(n2214) );
  AND U3172 ( .A(n1055), .B(n1516), .Z(n2328) );
  XOR U3173 ( .A(n2332), .B(n2215), .Z(n2327) );
  NAND U3174 ( .A(n1428), .B(n1114), .Z(n2215) );
  IV U3175 ( .A(n2217), .Z(n2332) );
  XNOR U3176 ( .A(n2336), .B(n2236), .Z(n2226) );
  XNOR U3177 ( .A(n2223), .B(n2224), .Z(n2236) );
  NANDN U3178 ( .B(n835), .A(n1925), .Z(n2224) );
  XNOR U3179 ( .A(n2222), .B(n2337), .Z(n2223) );
  AND U3180 ( .A(n1825), .B(n874), .Z(n2337) );
  XNOR U3181 ( .A(n2235), .B(n2225), .Z(n2336) );
  XNOR U3182 ( .A(n2230), .B(n2345), .Z(n2231) );
  AND U3183 ( .A(n1638), .B(n982), .Z(n2345) );
  XOR U3184 ( .A(n2349), .B(n2232), .Z(n2344) );
  NAND U3185 ( .A(n928), .B(n1731), .Z(n2232) );
  IV U3186 ( .A(n2234), .Z(n2349) );
  XNOR U3187 ( .A(n2239), .B(n2354), .Z(n2240) );
  AND U3188 ( .A(n2030), .B(n806), .Z(n2354) );
  XOR U3189 ( .A(n2358), .B(n2241), .Z(n2353) );
  NAND U3190 ( .A(n770), .B(n2135), .Z(n2241) );
  IV U3191 ( .A(n2243), .Z(n2358) );
  XNOR U3192 ( .A(n2250), .B(n2251), .Z(n2245) );
  NANDN U3193 ( .B(n709), .A(n2362), .Z(n2251) );
  AND U3194 ( .A(n2246), .B(n742), .Z(n2363) );
  NAND U3195 ( .A(n2364), .B(n2365), .Z(n2249) );
  NANDN U3196 ( .B(n2366), .A(n2367), .Z(n2364) );
  XNOR U3197 ( .A(n2371), .B(n2372), .Z(n655) );
  AND U3198 ( .A(n667), .B(n2374), .Z(n2373) );
  XOR U3199 ( .A(n2369), .B(n2372), .Z(n2374) );
  XNOR U3200 ( .A(n2368), .B(n2372), .Z(n2369) );
  XNOR U3201 ( .A(n2293), .B(n2292), .Z(n2372) );
  XNOR U3202 ( .A(n2375), .B(n2297), .Z(n2292) );
  XNOR U3203 ( .A(n2376), .B(n2271), .Z(n2266) );
  XNOR U3204 ( .A(n2263), .B(n2264), .Z(n2271) );
  NAND U3205 ( .A(n854), .B(n1946), .Z(n2264) );
  XNOR U3206 ( .A(n2262), .B(n2377), .Z(n2263) );
  AND U3207 ( .A(n2047), .B(n814), .Z(n2377) );
  XNOR U3208 ( .A(n2270), .B(n2265), .Z(n2376) );
  XNOR U3209 ( .A(n2275), .B(n2385), .Z(n2276) );
  AND U3210 ( .A(n2274), .B(n740), .Z(n2385) );
  XOR U3211 ( .A(n2389), .B(n2277), .Z(n2384) );
  NAND U3212 ( .A(n774), .B(n2160), .Z(n2277) );
  IV U3213 ( .A(n2269), .Z(n2389) );
  XNOR U3214 ( .A(n2280), .B(n2394), .Z(n2281) );
  AND U3215 ( .A(n1852), .B(n898), .Z(n2394) );
  XOR U3216 ( .A(n2398), .B(n2282), .Z(n2393) );
  NAND U3217 ( .A(n941), .B(n1751), .Z(n2282) );
  IV U3218 ( .A(n2284), .Z(n2398) );
  XNOR U3219 ( .A(n2289), .B(n2290), .Z(n2286) );
  NAND U3220 ( .A(n1055), .B(n1566), .Z(n2290) );
  XNOR U3221 ( .A(n2288), .B(n2402), .Z(n2289) );
  AND U3222 ( .A(n1660), .B(n999), .Z(n2402) );
  XNOR U3223 ( .A(n2296), .B(n2291), .Z(n2375) );
  AND U3224 ( .A(n2299), .B(n2410), .Z(n2409) );
  AND U3225 ( .A(n2411), .B(n2412), .Z(n2410) );
  NANDN U3226 ( .B(n710), .A(n2413), .Z(n2412) );
  NANDN U3227 ( .B(n2414), .A(n2415), .Z(n2411) );
  ANDN U3228 ( .A(n2301), .B(n2300), .Z(n2299) );
  NOR U3229 ( .A(n2416), .B(n2417), .Z(n2300) );
  NANDN U3230 ( .B(n2418), .A(n2419), .Z(n2301) );
  XNOR U3231 ( .A(n2423), .B(n2326), .Z(n2317) );
  XNOR U3232 ( .A(n2305), .B(n2425), .Z(n2306) );
  AND U3233 ( .A(n1383), .B(n1194), .Z(n2425) );
  XOR U3234 ( .A(n2429), .B(n2307), .Z(n2424) );
  NAND U3235 ( .A(n1136), .B(n1460), .Z(n2307) );
  IV U3236 ( .A(n2309), .Z(n2429) );
  XNOR U3237 ( .A(n2314), .B(n2315), .Z(n2311) );
  NANDN U3238 ( .B(n1020), .A(n1638), .Z(n2315) );
  XNOR U3239 ( .A(n2313), .B(n2433), .Z(n2314) );
  AND U3240 ( .A(n1546), .B(n1079), .Z(n2433) );
  XNOR U3241 ( .A(n2325), .B(n2316), .Z(n2423) );
  XOR U3242 ( .A(n2440), .B(n2335), .Z(n2325) );
  XNOR U3243 ( .A(n2322), .B(n2323), .Z(n2335) );
  NAND U3244 ( .A(n1280), .B(n1312), .Z(n2323) );
  XNOR U3245 ( .A(n2321), .B(n2441), .Z(n2322) );
  AND U3246 ( .A(n1242), .B(n1348), .Z(n2441) );
  XNOR U3247 ( .A(n2334), .B(n2324), .Z(n2440) );
  XNOR U3248 ( .A(n2329), .B(n2449), .Z(n2330) );
  AND U3249 ( .A(n1114), .B(n1516), .Z(n2449) );
  XOR U3250 ( .A(n2453), .B(n2331), .Z(n2448) );
  NAND U3251 ( .A(n1428), .B(n1176), .Z(n2331) );
  IV U3252 ( .A(n2333), .Z(n2453) );
  XNOR U3253 ( .A(n2457), .B(n2352), .Z(n2342) );
  XNOR U3254 ( .A(n2339), .B(n2340), .Z(n2352) );
  NANDN U3255 ( .B(n835), .A(n2030), .Z(n2340) );
  XNOR U3256 ( .A(n2338), .B(n2458), .Z(n2339) );
  AND U3257 ( .A(n1925), .B(n874), .Z(n2458) );
  XNOR U3258 ( .A(n2351), .B(n2341), .Z(n2457) );
  XNOR U3259 ( .A(n2346), .B(n2466), .Z(n2347) );
  AND U3260 ( .A(n1731), .B(n982), .Z(n2466) );
  XOR U3261 ( .A(n2470), .B(n2348), .Z(n2465) );
  NAND U3262 ( .A(n928), .B(n1825), .Z(n2348) );
  IV U3263 ( .A(n2350), .Z(n2470) );
  XNOR U3264 ( .A(n2355), .B(n2475), .Z(n2356) );
  AND U3265 ( .A(n2135), .B(n806), .Z(n2475) );
  XOR U3266 ( .A(n2479), .B(n2357), .Z(n2474) );
  NAND U3267 ( .A(n770), .B(n2246), .Z(n2357) );
  IV U3268 ( .A(n2359), .Z(n2479) );
  XNOR U3269 ( .A(n2366), .B(n2367), .Z(n2361) );
  NANDN U3270 ( .B(n709), .A(n2483), .Z(n2367) );
  XNOR U3271 ( .A(n2365), .B(n2484), .Z(n2366) );
  AND U3272 ( .A(n2362), .B(n742), .Z(n2484) );
  ANDN U3273 ( .A(n2485), .B(n2486), .Z(n2365) );
  NANDN U3274 ( .B(n2487), .A(n2488), .Z(n2485) );
  XNOR U3275 ( .A(n2492), .B(n2493), .Z(n656) );
  AND U3276 ( .A(n667), .B(n2495), .Z(n2494) );
  XOR U3277 ( .A(n2490), .B(n2493), .Z(n2495) );
  XNOR U3278 ( .A(n2489), .B(n2493), .Z(n2490) );
  XNOR U3279 ( .A(n2408), .B(n2407), .Z(n2493) );
  XNOR U3280 ( .A(n2496), .B(n2422), .Z(n2407) );
  XNOR U3281 ( .A(n2497), .B(n2392), .Z(n2382) );
  XNOR U3282 ( .A(n2379), .B(n2380), .Z(n2392) );
  NAND U3283 ( .A(n898), .B(n1946), .Z(n2380) );
  XNOR U3284 ( .A(n2378), .B(n2498), .Z(n2379) );
  AND U3285 ( .A(n2047), .B(n854), .Z(n2498) );
  XNOR U3286 ( .A(n2391), .B(n2381), .Z(n2497) );
  XNOR U3287 ( .A(n2386), .B(n2506), .Z(n2387) );
  AND U3288 ( .A(n2274), .B(n774), .Z(n2506) );
  XOR U3289 ( .A(n2510), .B(n2388), .Z(n2505) );
  NAND U3290 ( .A(n814), .B(n2160), .Z(n2388) );
  IV U3291 ( .A(n2390), .Z(n2510) );
  XNOR U3292 ( .A(n2395), .B(n2515), .Z(n2396) );
  AND U3293 ( .A(n1852), .B(n941), .Z(n2515) );
  XOR U3294 ( .A(n2519), .B(n2397), .Z(n2514) );
  NAND U3295 ( .A(n999), .B(n1751), .Z(n2397) );
  IV U3296 ( .A(n2399), .Z(n2519) );
  XOR U3297 ( .A(n2520), .B(n2521), .Z(n2399) );
  ANDN U3298 ( .A(n2522), .B(n2523), .Z(n2521) );
  XOR U3299 ( .A(n2520), .B(n2524), .Z(n2522) );
  XNOR U3300 ( .A(n2404), .B(n2405), .Z(n2401) );
  NAND U3301 ( .A(n1114), .B(n1566), .Z(n2405) );
  XNOR U3302 ( .A(n2403), .B(n2525), .Z(n2404) );
  AND U3303 ( .A(n1660), .B(n1055), .Z(n2525) );
  XNOR U3304 ( .A(n2421), .B(n2406), .Z(n2496) );
  XOR U3305 ( .A(n2532), .B(n2415), .Z(n2421) );
  XNOR U3306 ( .A(n2418), .B(n2419), .Z(n2415) );
  XOR U3307 ( .A(n2536), .B(n2417), .Z(n2418) );
  NAND U3308 ( .A(n740), .B(n2413), .Z(n2417) );
  NANDN U3309 ( .B(n710), .A(n2538), .Z(n2537) );
  OR U3310 ( .A(n2542), .B(n2543), .Z(n2414) );
  XNOR U3311 ( .A(n2547), .B(n2447), .Z(n2438) );
  XNOR U3312 ( .A(n2426), .B(n2549), .Z(n2427) );
  AND U3313 ( .A(n1460), .B(n1194), .Z(n2549) );
  XOR U3314 ( .A(n2553), .B(n2428), .Z(n2548) );
  NAND U3315 ( .A(n1136), .B(n1546), .Z(n2428) );
  IV U3316 ( .A(n2430), .Z(n2553) );
  XNOR U3317 ( .A(n2435), .B(n2436), .Z(n2432) );
  NANDN U3318 ( .B(n1020), .A(n1731), .Z(n2436) );
  XNOR U3319 ( .A(n2434), .B(n2557), .Z(n2435) );
  AND U3320 ( .A(n1638), .B(n1079), .Z(n2557) );
  XNOR U3321 ( .A(n2446), .B(n2437), .Z(n2547) );
  XOR U3322 ( .A(n2564), .B(n2456), .Z(n2446) );
  XNOR U3323 ( .A(n2443), .B(n2444), .Z(n2456) );
  NAND U3324 ( .A(n1280), .B(n1383), .Z(n2444) );
  XNOR U3325 ( .A(n2442), .B(n2565), .Z(n2443) );
  AND U3326 ( .A(n1312), .B(n1348), .Z(n2565) );
  XNOR U3327 ( .A(n2455), .B(n2445), .Z(n2564) );
  XNOR U3328 ( .A(n2450), .B(n2573), .Z(n2451) );
  AND U3329 ( .A(n1176), .B(n1516), .Z(n2573) );
  XOR U3330 ( .A(n2577), .B(n2452), .Z(n2572) );
  NAND U3331 ( .A(n1428), .B(n1242), .Z(n2452) );
  IV U3332 ( .A(n2454), .Z(n2577) );
  XNOR U3333 ( .A(n2581), .B(n2473), .Z(n2463) );
  XNOR U3334 ( .A(n2460), .B(n2461), .Z(n2473) );
  NANDN U3335 ( .B(n835), .A(n2135), .Z(n2461) );
  XNOR U3336 ( .A(n2459), .B(n2582), .Z(n2460) );
  AND U3337 ( .A(n2030), .B(n874), .Z(n2582) );
  XNOR U3338 ( .A(n2472), .B(n2462), .Z(n2581) );
  XNOR U3339 ( .A(n2467), .B(n2590), .Z(n2468) );
  AND U3340 ( .A(n1825), .B(n982), .Z(n2590) );
  XOR U3341 ( .A(n2594), .B(n2469), .Z(n2589) );
  NAND U3342 ( .A(n928), .B(n1925), .Z(n2469) );
  IV U3343 ( .A(n2471), .Z(n2594) );
  XNOR U3344 ( .A(n2476), .B(n2599), .Z(n2477) );
  AND U3345 ( .A(n2246), .B(n806), .Z(n2599) );
  XOR U3346 ( .A(n2603), .B(n2478), .Z(n2598) );
  NAND U3347 ( .A(n770), .B(n2362), .Z(n2478) );
  IV U3348 ( .A(n2480), .Z(n2603) );
  XNOR U3349 ( .A(n2487), .B(n2488), .Z(n2482) );
  NANDN U3350 ( .B(n709), .A(n2607), .Z(n2488) );
  AND U3351 ( .A(n2483), .B(n742), .Z(n2608) );
  NAND U3352 ( .A(n2609), .B(n2610), .Z(n2486) );
  NANDN U3353 ( .B(n2611), .A(n2612), .Z(n2609) );
  XOR U3354 ( .A(n2616), .B(n2617), .Z(n657) );
  AND U3355 ( .A(n667), .B(n2619), .Z(n2618) );
  XNOR U3356 ( .A(n2614), .B(n2617), .Z(n2619) );
  XNOR U3357 ( .A(n2617), .B(n2613), .Z(n2614) );
  OR U3358 ( .A(n2620), .B(n2621), .Z(n2613) );
  XNOR U3359 ( .A(n2531), .B(n2530), .Z(n2617) );
  XNOR U3360 ( .A(n2622), .B(n2546), .Z(n2530) );
  XNOR U3361 ( .A(n2623), .B(n2513), .Z(n2503) );
  XNOR U3362 ( .A(n2500), .B(n2501), .Z(n2513) );
  NAND U3363 ( .A(n941), .B(n1946), .Z(n2501) );
  XNOR U3364 ( .A(n2499), .B(n2624), .Z(n2500) );
  AND U3365 ( .A(n2047), .B(n898), .Z(n2624) );
  XNOR U3366 ( .A(n2512), .B(n2502), .Z(n2623) );
  XNOR U3367 ( .A(n2507), .B(n2632), .Z(n2508) );
  AND U3368 ( .A(n2274), .B(n814), .Z(n2632) );
  XOR U3369 ( .A(n2636), .B(n2509), .Z(n2631) );
  NAND U3370 ( .A(n854), .B(n2160), .Z(n2509) );
  IV U3371 ( .A(n2511), .Z(n2636) );
  XNOR U3372 ( .A(n2516), .B(n2641), .Z(n2517) );
  AND U3373 ( .A(n1852), .B(n999), .Z(n2641) );
  XOR U3374 ( .A(n2645), .B(n2518), .Z(n2640) );
  NAND U3375 ( .A(n1055), .B(n1751), .Z(n2518) );
  IV U3376 ( .A(n2520), .Z(n2645) );
  XNOR U3377 ( .A(n2527), .B(n2528), .Z(n2524) );
  NAND U3378 ( .A(n1176), .B(n1566), .Z(n2528) );
  XNOR U3379 ( .A(n2526), .B(n2649), .Z(n2527) );
  AND U3380 ( .A(n1660), .B(n1114), .Z(n2649) );
  XNOR U3381 ( .A(n2545), .B(n2529), .Z(n2622) );
  XNOR U3382 ( .A(n2656), .B(n2542), .Z(n2545) );
  XOR U3383 ( .A(n2535), .B(n2534), .Z(n2542) );
  XOR U3384 ( .A(n2533), .B(n2657), .Z(n2534) );
  AND U3385 ( .A(n2658), .B(n2659), .Z(n2657) );
  NANDN U3386 ( .B(n710), .A(n2660), .Z(n2659) );
  OR U3387 ( .A(n2661), .B(n2662), .Z(n2658) );
  NAND U3388 ( .A(n774), .B(n2413), .Z(n2541) );
  XNOR U3389 ( .A(n2539), .B(n2665), .Z(n2540) );
  AND U3390 ( .A(n2538), .B(n740), .Z(n2665) );
  NANDN U3391 ( .B(n2669), .A(n2670), .Z(n2543) );
  XNOR U3392 ( .A(n2674), .B(n2571), .Z(n2562) );
  XNOR U3393 ( .A(n2550), .B(n2676), .Z(n2551) );
  AND U3394 ( .A(n1546), .B(n1194), .Z(n2676) );
  XOR U3395 ( .A(n2680), .B(n2552), .Z(n2675) );
  NAND U3396 ( .A(n1136), .B(n1638), .Z(n2552) );
  IV U3397 ( .A(n2554), .Z(n2680) );
  XNOR U3398 ( .A(n2559), .B(n2560), .Z(n2556) );
  NANDN U3399 ( .B(n1020), .A(n1825), .Z(n2560) );
  XNOR U3400 ( .A(n2558), .B(n2684), .Z(n2559) );
  AND U3401 ( .A(n1731), .B(n1079), .Z(n2684) );
  XNOR U3402 ( .A(n2570), .B(n2561), .Z(n2674) );
  XOR U3403 ( .A(n2691), .B(n2580), .Z(n2570) );
  XNOR U3404 ( .A(n2567), .B(n2568), .Z(n2580) );
  NAND U3405 ( .A(n1280), .B(n1460), .Z(n2568) );
  XNOR U3406 ( .A(n2566), .B(n2692), .Z(n2567) );
  AND U3407 ( .A(n1383), .B(n1348), .Z(n2692) );
  XNOR U3408 ( .A(n2579), .B(n2569), .Z(n2691) );
  XNOR U3409 ( .A(n2574), .B(n2700), .Z(n2575) );
  AND U3410 ( .A(n1242), .B(n1516), .Z(n2700) );
  XOR U3411 ( .A(n2704), .B(n2576), .Z(n2699) );
  NAND U3412 ( .A(n1428), .B(n1312), .Z(n2576) );
  IV U3413 ( .A(n2578), .Z(n2704) );
  XNOR U3414 ( .A(n2708), .B(n2597), .Z(n2587) );
  XNOR U3415 ( .A(n2584), .B(n2585), .Z(n2597) );
  NANDN U3416 ( .B(n835), .A(n2246), .Z(n2585) );
  XNOR U3417 ( .A(n2583), .B(n2709), .Z(n2584) );
  AND U3418 ( .A(n2135), .B(n874), .Z(n2709) );
  XNOR U3419 ( .A(n2596), .B(n2586), .Z(n2708) );
  XNOR U3420 ( .A(n2591), .B(n2717), .Z(n2592) );
  AND U3421 ( .A(n1925), .B(n982), .Z(n2717) );
  XOR U3422 ( .A(n2721), .B(n2593), .Z(n2716) );
  NAND U3423 ( .A(n928), .B(n2030), .Z(n2593) );
  IV U3424 ( .A(n2595), .Z(n2721) );
  XNOR U3425 ( .A(n2600), .B(n2726), .Z(n2601) );
  AND U3426 ( .A(n2362), .B(n806), .Z(n2726) );
  XOR U3427 ( .A(n2730), .B(n2602), .Z(n2725) );
  NAND U3428 ( .A(n770), .B(n2483), .Z(n2602) );
  IV U3429 ( .A(n2604), .Z(n2730) );
  XNOR U3430 ( .A(n2611), .B(n2612), .Z(n2606) );
  NANDN U3431 ( .B(n709), .A(n2734), .Z(n2612) );
  XNOR U3432 ( .A(n2610), .B(n2735), .Z(n2611) );
  AND U3433 ( .A(n2607), .B(n742), .Z(n2735) );
  ANDN U3434 ( .A(n2736), .B(n2737), .Z(n2610) );
  NANDN U3435 ( .B(n2738), .A(n2739), .Z(n2736) );
  XNOR U3436 ( .A(n2741), .B(n2742), .Z(n695) );
  AND U3437 ( .A(n667), .B(n2744), .Z(n2743) );
  XOR U3438 ( .A(n2620), .B(n2745), .Z(n2744) );
  XOR U3439 ( .A(n2745), .B(n2621), .Z(n2620) );
  OR U3440 ( .A(n2746), .B(n2747), .Z(n2621) );
  IV U3441 ( .A(n2742), .Z(n2745) );
  XOR U3442 ( .A(n2655), .B(n2654), .Z(n2742) );
  XNOR U3443 ( .A(n2748), .B(n2673), .Z(n2654) );
  XNOR U3444 ( .A(n2749), .B(n2639), .Z(n2629) );
  XNOR U3445 ( .A(n2626), .B(n2627), .Z(n2639) );
  NAND U3446 ( .A(n999), .B(n1946), .Z(n2627) );
  XNOR U3447 ( .A(n2625), .B(n2750), .Z(n2626) );
  AND U3448 ( .A(n2047), .B(n941), .Z(n2750) );
  XNOR U3449 ( .A(n2638), .B(n2628), .Z(n2749) );
  XNOR U3450 ( .A(n2633), .B(n2758), .Z(n2634) );
  AND U3451 ( .A(n2274), .B(n854), .Z(n2758) );
  XOR U3452 ( .A(n2762), .B(n2635), .Z(n2757) );
  NAND U3453 ( .A(n898), .B(n2160), .Z(n2635) );
  IV U3454 ( .A(n2637), .Z(n2762) );
  XNOR U3455 ( .A(n2642), .B(n2767), .Z(n2643) );
  AND U3456 ( .A(n1852), .B(n1055), .Z(n2767) );
  XOR U3457 ( .A(n2771), .B(n2644), .Z(n2766) );
  NAND U3458 ( .A(n1114), .B(n1751), .Z(n2644) );
  IV U3459 ( .A(n2646), .Z(n2771) );
  XNOR U3460 ( .A(n2651), .B(n2652), .Z(n2648) );
  NAND U3461 ( .A(n1242), .B(n1566), .Z(n2652) );
  XNOR U3462 ( .A(n2650), .B(n2775), .Z(n2651) );
  AND U3463 ( .A(n1660), .B(n1176), .Z(n2775) );
  XNOR U3464 ( .A(n2672), .B(n2653), .Z(n2748) );
  XNOR U3465 ( .A(n2782), .B(n2669), .Z(n2672) );
  XOR U3466 ( .A(n2664), .B(n2663), .Z(n2669) );
  XNOR U3467 ( .A(n2783), .B(n2784), .Z(n2663) );
  ANDN U3468 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR U3469 ( .A(n2785), .B(n2789), .Z(n2787) );
  XNOR U3470 ( .A(n2790), .B(n2661), .Z(n2783) );
  NAND U3471 ( .A(n740), .B(n2660), .Z(n2661) );
  NANDN U3472 ( .B(n710), .A(n2792), .Z(n2791) );
  NAND U3473 ( .A(n814), .B(n2413), .Z(n2668) );
  XNOR U3474 ( .A(n2666), .B(n2796), .Z(n2667) );
  AND U3475 ( .A(n2538), .B(n774), .Z(n2796) );
  XNOR U3476 ( .A(n2670), .B(n2671), .Z(n2782) );
  XNOR U3477 ( .A(n2806), .B(n2698), .Z(n2689) );
  XNOR U3478 ( .A(n2677), .B(n2808), .Z(n2678) );
  AND U3479 ( .A(n1638), .B(n1194), .Z(n2808) );
  XOR U3480 ( .A(n2812), .B(n2679), .Z(n2807) );
  NAND U3481 ( .A(n1136), .B(n1731), .Z(n2679) );
  IV U3482 ( .A(n2681), .Z(n2812) );
  XNOR U3483 ( .A(n2686), .B(n2687), .Z(n2683) );
  NANDN U3484 ( .B(n1020), .A(n1925), .Z(n2687) );
  XNOR U3485 ( .A(n2685), .B(n2816), .Z(n2686) );
  AND U3486 ( .A(n1825), .B(n1079), .Z(n2816) );
  XNOR U3487 ( .A(n2697), .B(n2688), .Z(n2806) );
  XOR U3488 ( .A(n2823), .B(n2707), .Z(n2697) );
  XNOR U3489 ( .A(n2694), .B(n2695), .Z(n2707) );
  NAND U3490 ( .A(n1280), .B(n1546), .Z(n2695) );
  XNOR U3491 ( .A(n2693), .B(n2824), .Z(n2694) );
  AND U3492 ( .A(n1460), .B(n1348), .Z(n2824) );
  XNOR U3493 ( .A(n2706), .B(n2696), .Z(n2823) );
  XNOR U3494 ( .A(n2701), .B(n2832), .Z(n2702) );
  AND U3495 ( .A(n1312), .B(n1516), .Z(n2832) );
  XOR U3496 ( .A(n2836), .B(n2703), .Z(n2831) );
  NAND U3497 ( .A(n1428), .B(n1383), .Z(n2703) );
  IV U3498 ( .A(n2705), .Z(n2836) );
  XNOR U3499 ( .A(n2840), .B(n2724), .Z(n2714) );
  XNOR U3500 ( .A(n2711), .B(n2712), .Z(n2724) );
  NANDN U3501 ( .B(n835), .A(n2362), .Z(n2712) );
  XNOR U3502 ( .A(n2710), .B(n2841), .Z(n2711) );
  AND U3503 ( .A(n2246), .B(n874), .Z(n2841) );
  XNOR U3504 ( .A(n2723), .B(n2713), .Z(n2840) );
  XNOR U3505 ( .A(n2718), .B(n2849), .Z(n2719) );
  AND U3506 ( .A(n2030), .B(n982), .Z(n2849) );
  XOR U3507 ( .A(n2853), .B(n2720), .Z(n2848) );
  NAND U3508 ( .A(n928), .B(n2135), .Z(n2720) );
  IV U3509 ( .A(n2722), .Z(n2853) );
  XNOR U3510 ( .A(n2727), .B(n2858), .Z(n2728) );
  AND U3511 ( .A(n2483), .B(n806), .Z(n2858) );
  XOR U3512 ( .A(n2862), .B(n2729), .Z(n2857) );
  NAND U3513 ( .A(n770), .B(n2607), .Z(n2729) );
  IV U3514 ( .A(n2731), .Z(n2862) );
  XNOR U3515 ( .A(n2738), .B(n2739), .Z(n2733) );
  OR U3516 ( .A(n2866), .B(n709), .Z(n2739) );
  AND U3517 ( .A(n2734), .B(n742), .Z(n2867) );
  NAND U3518 ( .A(n2868), .B(n2869), .Z(n2737) );
  NANDN U3519 ( .B(n2870), .A(n2871), .Z(n2868) );
  XNOR U3520 ( .A(n2873), .B(n2874), .Z(n1123) );
  XOR U3521 ( .A(n2872), .B(n2875), .Z(n2873) );
  AND U3522 ( .A(n667), .B(n2876), .Z(n2875) );
  XOR U3523 ( .A(n2746), .B(n2877), .Z(n2876) );
  XOR U3524 ( .A(n2877), .B(n2747), .Z(n2746) );
  NANDN U3525 ( .B(n2878), .A(n2879), .Z(n2747) );
  IV U3526 ( .A(n2874), .Z(n2877) );
  XOR U3527 ( .A(n2781), .B(n2780), .Z(n2874) );
  XNOR U3528 ( .A(n2880), .B(n2802), .Z(n2780) );
  XNOR U3529 ( .A(n2881), .B(n2765), .Z(n2755) );
  XNOR U3530 ( .A(n2752), .B(n2753), .Z(n2765) );
  NAND U3531 ( .A(n1055), .B(n1946), .Z(n2753) );
  XNOR U3532 ( .A(n2751), .B(n2882), .Z(n2752) );
  AND U3533 ( .A(n2047), .B(n999), .Z(n2882) );
  XNOR U3534 ( .A(n2764), .B(n2754), .Z(n2881) );
  XNOR U3535 ( .A(n2759), .B(n2890), .Z(n2760) );
  AND U3536 ( .A(n2274), .B(n898), .Z(n2890) );
  XOR U3537 ( .A(n2894), .B(n2761), .Z(n2889) );
  NAND U3538 ( .A(n941), .B(n2160), .Z(n2761) );
  IV U3539 ( .A(n2763), .Z(n2894) );
  XNOR U3540 ( .A(n2768), .B(n2899), .Z(n2769) );
  AND U3541 ( .A(n1852), .B(n1114), .Z(n2899) );
  XOR U3542 ( .A(n2903), .B(n2770), .Z(n2898) );
  NAND U3543 ( .A(n1176), .B(n1751), .Z(n2770) );
  IV U3544 ( .A(n2772), .Z(n2903) );
  XNOR U3545 ( .A(n2777), .B(n2778), .Z(n2774) );
  NAND U3546 ( .A(n1312), .B(n1566), .Z(n2778) );
  XNOR U3547 ( .A(n2776), .B(n2907), .Z(n2777) );
  AND U3548 ( .A(n1660), .B(n1242), .Z(n2907) );
  XNOR U3549 ( .A(n2801), .B(n2779), .Z(n2880) );
  XOR U3550 ( .A(n2914), .B(n2805), .Z(n2801) );
  XNOR U3551 ( .A(n2793), .B(n2916), .Z(n2794) );
  AND U3552 ( .A(n2792), .B(n740), .Z(n2916) );
  XOR U3553 ( .A(n2920), .B(n2795), .Z(n2915) );
  NAND U3554 ( .A(n774), .B(n2660), .Z(n2795) );
  IV U3555 ( .A(n2785), .Z(n2920) );
  XNOR U3556 ( .A(n2798), .B(n2799), .Z(n2789) );
  NAND U3557 ( .A(n854), .B(n2413), .Z(n2799) );
  XNOR U3558 ( .A(n2797), .B(n2924), .Z(n2798) );
  AND U3559 ( .A(n2538), .B(n814), .Z(n2924) );
  XNOR U3560 ( .A(n2804), .B(n2800), .Z(n2914) );
  AND U3561 ( .A(n2932), .B(n2933), .Z(n2931) );
  OR U3562 ( .A(n2934), .B(n2935), .Z(n2933) );
  AND U3563 ( .A(n2936), .B(n2937), .Z(n2932) );
  NANDN U3564 ( .B(n710), .A(n2938), .Z(n2937) );
  NANDN U3565 ( .B(n2939), .A(n2940), .Z(n2936) );
  XNOR U3566 ( .A(n2944), .B(n2830), .Z(n2821) );
  XNOR U3567 ( .A(n2809), .B(n2946), .Z(n2810) );
  AND U3568 ( .A(n1731), .B(n1194), .Z(n2946) );
  XOR U3569 ( .A(n2950), .B(n2811), .Z(n2945) );
  NAND U3570 ( .A(n1136), .B(n1825), .Z(n2811) );
  IV U3571 ( .A(n2813), .Z(n2950) );
  XNOR U3572 ( .A(n2818), .B(n2819), .Z(n2815) );
  NANDN U3573 ( .B(n1020), .A(n2030), .Z(n2819) );
  XNOR U3574 ( .A(n2817), .B(n2954), .Z(n2818) );
  AND U3575 ( .A(n1925), .B(n1079), .Z(n2954) );
  XNOR U3576 ( .A(n2829), .B(n2820), .Z(n2944) );
  XOR U3577 ( .A(n2961), .B(n2839), .Z(n2829) );
  XNOR U3578 ( .A(n2826), .B(n2827), .Z(n2839) );
  NAND U3579 ( .A(n1280), .B(n1638), .Z(n2827) );
  XNOR U3580 ( .A(n2825), .B(n2962), .Z(n2826) );
  AND U3581 ( .A(n1546), .B(n1348), .Z(n2962) );
  XNOR U3582 ( .A(n2838), .B(n2828), .Z(n2961) );
  XNOR U3583 ( .A(n2833), .B(n2970), .Z(n2834) );
  AND U3584 ( .A(n1383), .B(n1516), .Z(n2970) );
  XOR U3585 ( .A(n2974), .B(n2835), .Z(n2969) );
  NAND U3586 ( .A(n1428), .B(n1460), .Z(n2835) );
  IV U3587 ( .A(n2837), .Z(n2974) );
  XNOR U3588 ( .A(n2978), .B(n2856), .Z(n2846) );
  XNOR U3589 ( .A(n2843), .B(n2844), .Z(n2856) );
  NANDN U3590 ( .B(n835), .A(n2483), .Z(n2844) );
  XNOR U3591 ( .A(n2842), .B(n2979), .Z(n2843) );
  AND U3592 ( .A(n2362), .B(n874), .Z(n2979) );
  XNOR U3593 ( .A(n2855), .B(n2845), .Z(n2978) );
  XNOR U3594 ( .A(n2850), .B(n2987), .Z(n2851) );
  AND U3595 ( .A(n2135), .B(n982), .Z(n2987) );
  XOR U3596 ( .A(n2991), .B(n2852), .Z(n2986) );
  NAND U3597 ( .A(n928), .B(n2246), .Z(n2852) );
  IV U3598 ( .A(n2854), .Z(n2991) );
  XNOR U3599 ( .A(n2859), .B(n2996), .Z(n2860) );
  AND U3600 ( .A(n2607), .B(n806), .Z(n2996) );
  XOR U3601 ( .A(n3000), .B(n2861), .Z(n2995) );
  NAND U3602 ( .A(n770), .B(n2734), .Z(n2861) );
  IV U3603 ( .A(n2863), .Z(n3000) );
  XNOR U3604 ( .A(n2870), .B(n2871), .Z(n2865) );
  OR U3605 ( .A(n3004), .B(n709), .Z(n2871) );
  XNOR U3606 ( .A(n2869), .B(n3005), .Z(n2870) );
  ANDN U3607 ( .A(n742), .B(n2866), .Z(n3005) );
  ANDN U3608 ( .A(n3006), .B(n3007), .Z(n2869) );
  NANDN U3609 ( .B(n3008), .A(n3009), .Z(n3006) );
  XOR U3610 ( .A(n3011), .B(\_MxM/Y0[1] ), .Z(\_MxM/Y1[0] ) );
  XOR U3611 ( .A(n3012), .B(n3013), .Z(n3011) );
  XNOR U3612 ( .A(n3014), .B(n3010), .Z(n3012) );
  NANDN U3613 ( .B(n2879), .A(\_MxM/Y0[0] ), .Z(n3010) );
  NAND U3614 ( .A(n3015), .B(n667), .Z(n3014) );
  XOR U3615 ( .A(e_input[31]), .B(g_input[31]), .Z(n667) );
  XNOR U3616 ( .A(n2878), .B(n3013), .Z(n3015) );
  XOR U3617 ( .A(n2879), .B(n3013), .Z(n2878) );
  XOR U3618 ( .A(n2913), .B(n2912), .Z(n3013) );
  XNOR U3619 ( .A(n3016), .B(n2930), .Z(n2912) );
  XNOR U3620 ( .A(n3017), .B(n2897), .Z(n2887) );
  XNOR U3621 ( .A(n2884), .B(n2885), .Z(n2897) );
  NAND U3622 ( .A(n1114), .B(n1946), .Z(n2885) );
  XNOR U3623 ( .A(n2883), .B(n3018), .Z(n2884) );
  AND U3624 ( .A(n2047), .B(n1055), .Z(n3018) );
  XNOR U3625 ( .A(n2896), .B(n2886), .Z(n3017) );
  XNOR U3626 ( .A(n2891), .B(n3026), .Z(n2892) );
  AND U3627 ( .A(n2274), .B(n941), .Z(n3026) );
  XOR U3628 ( .A(n3030), .B(n2893), .Z(n3025) );
  NAND U3629 ( .A(n999), .B(n2160), .Z(n2893) );
  IV U3630 ( .A(n2895), .Z(n3030) );
  XNOR U3631 ( .A(n2900), .B(n3035), .Z(n2901) );
  AND U3632 ( .A(n1852), .B(n1176), .Z(n3035) );
  XOR U3633 ( .A(n3039), .B(n2902), .Z(n3034) );
  NAND U3634 ( .A(n1242), .B(n1751), .Z(n2902) );
  IV U3635 ( .A(n2904), .Z(n3039) );
  XNOR U3636 ( .A(n2909), .B(n2910), .Z(n2906) );
  NAND U3637 ( .A(n1383), .B(n1566), .Z(n2910) );
  XNOR U3638 ( .A(n2908), .B(n3043), .Z(n2909) );
  AND U3639 ( .A(n1660), .B(n1312), .Z(n3043) );
  XNOR U3640 ( .A(n2929), .B(n2911), .Z(n3016) );
  XOR U3641 ( .A(n3050), .B(n2943), .Z(n2929) );
  XNOR U3642 ( .A(n2917), .B(n3052), .Z(n2918) );
  AND U3643 ( .A(n2792), .B(n774), .Z(n3052) );
  XOR U3644 ( .A(n3056), .B(n2919), .Z(n3051) );
  NAND U3645 ( .A(n814), .B(n2660), .Z(n2919) );
  IV U3646 ( .A(n2921), .Z(n3056) );
  XNOR U3647 ( .A(n2926), .B(n2927), .Z(n2923) );
  NAND U3648 ( .A(n898), .B(n2413), .Z(n2927) );
  XNOR U3649 ( .A(n2925), .B(n3060), .Z(n2926) );
  AND U3650 ( .A(n2538), .B(n854), .Z(n3060) );
  XNOR U3651 ( .A(n2942), .B(n2928), .Z(n3050) );
  XNOR U3652 ( .A(n3067), .B(n2939), .Z(n2942) );
  XOR U3653 ( .A(n3068), .B(n2934), .Z(n2939) );
  NAND U3654 ( .A(n740), .B(n2938), .Z(n2934) );
  NANDN U3655 ( .B(n710), .A(n3070), .Z(n3069) );
  XNOR U3656 ( .A(n2940), .B(n2941), .Z(n3067) );
  XNOR U3657 ( .A(n3079), .B(n2968), .Z(n2959) );
  XNOR U3658 ( .A(n2947), .B(n3081), .Z(n2948) );
  AND U3659 ( .A(n1825), .B(n1194), .Z(n3081) );
  XOR U3660 ( .A(n3085), .B(n2949), .Z(n3080) );
  NAND U3661 ( .A(n1136), .B(n1925), .Z(n2949) );
  IV U3662 ( .A(n2951), .Z(n3085) );
  XNOR U3663 ( .A(n2956), .B(n2957), .Z(n2953) );
  NANDN U3664 ( .B(n1020), .A(n2135), .Z(n2957) );
  XNOR U3665 ( .A(n2955), .B(n3089), .Z(n2956) );
  AND U3666 ( .A(n2030), .B(n1079), .Z(n3089) );
  XNOR U3667 ( .A(n2967), .B(n2958), .Z(n3079) );
  XOR U3668 ( .A(n3096), .B(n2977), .Z(n2967) );
  XNOR U3669 ( .A(n2964), .B(n2965), .Z(n2977) );
  NAND U3670 ( .A(n1280), .B(n1731), .Z(n2965) );
  XNOR U3671 ( .A(n2963), .B(n3097), .Z(n2964) );
  AND U3672 ( .A(n1638), .B(n1348), .Z(n3097) );
  XNOR U3673 ( .A(n2976), .B(n2966), .Z(n3096) );
  XNOR U3674 ( .A(n2971), .B(n3105), .Z(n2972) );
  AND U3675 ( .A(n1460), .B(n1516), .Z(n3105) );
  XOR U3676 ( .A(n3109), .B(n2973), .Z(n3104) );
  NAND U3677 ( .A(n1428), .B(n1546), .Z(n2973) );
  IV U3678 ( .A(n2975), .Z(n3109) );
  XNOR U3679 ( .A(n3113), .B(n2994), .Z(n2984) );
  XNOR U3680 ( .A(n2981), .B(n2982), .Z(n2994) );
  NANDN U3681 ( .B(n835), .A(n2607), .Z(n2982) );
  XNOR U3682 ( .A(n2980), .B(n3114), .Z(n2981) );
  AND U3683 ( .A(n2483), .B(n874), .Z(n3114) );
  XNOR U3684 ( .A(n2993), .B(n2983), .Z(n3113) );
  XNOR U3685 ( .A(n2988), .B(n3122), .Z(n2989) );
  AND U3686 ( .A(n2246), .B(n982), .Z(n3122) );
  XOR U3687 ( .A(n3126), .B(n2990), .Z(n3121) );
  NAND U3688 ( .A(n928), .B(n2362), .Z(n2990) );
  IV U3689 ( .A(n2992), .Z(n3126) );
  XNOR U3690 ( .A(n2997), .B(n3131), .Z(n2998) );
  AND U3691 ( .A(n2734), .B(n806), .Z(n3131) );
  XOR U3692 ( .A(n3135), .B(n2999), .Z(n3130) );
  NANDN U3693 ( .B(n2866), .A(n770), .Z(n2999) );
  IV U3694 ( .A(n3001), .Z(n3135) );
  XNOR U3695 ( .A(n3008), .B(n3009), .Z(n3003) );
  NANDN U3696 ( .B(n709), .A(n3139), .Z(n3009) );
  ANDN U3697 ( .A(n742), .B(n3004), .Z(n3140) );
  NAND U3698 ( .A(n3141), .B(n3142), .Z(n3007) );
  NANDN U3699 ( .B(n3143), .A(n3144), .Z(n3141) );
  XOR U3700 ( .A(n3049), .B(n3048), .Z(n2879) );
  XNOR U3701 ( .A(n3145), .B(n3066), .Z(n3048) );
  XNOR U3702 ( .A(n3146), .B(n3033), .Z(n3023) );
  XNOR U3703 ( .A(n3020), .B(n3021), .Z(n3033) );
  NAND U3704 ( .A(n1176), .B(n1946), .Z(n3021) );
  XNOR U3705 ( .A(n3019), .B(n3147), .Z(n3020) );
  AND U3706 ( .A(n2047), .B(n1114), .Z(n3147) );
  XNOR U3707 ( .A(n3032), .B(n3022), .Z(n3146) );
  XNOR U3708 ( .A(n3027), .B(n3155), .Z(n3028) );
  AND U3709 ( .A(n2274), .B(n999), .Z(n3155) );
  XOR U3710 ( .A(n3159), .B(n3029), .Z(n3154) );
  NAND U3711 ( .A(n1055), .B(n2160), .Z(n3029) );
  IV U3712 ( .A(n3031), .Z(n3159) );
  XNOR U3713 ( .A(n3036), .B(n3164), .Z(n3037) );
  AND U3714 ( .A(n1852), .B(n1242), .Z(n3164) );
  XOR U3715 ( .A(n3168), .B(n3038), .Z(n3163) );
  NAND U3716 ( .A(n1312), .B(n1751), .Z(n3038) );
  IV U3717 ( .A(n3040), .Z(n3168) );
  XNOR U3718 ( .A(n3045), .B(n3046), .Z(n3042) );
  NAND U3719 ( .A(n1460), .B(n1566), .Z(n3046) );
  XNOR U3720 ( .A(n3044), .B(n3172), .Z(n3045) );
  AND U3721 ( .A(n1660), .B(n1383), .Z(n3172) );
  XNOR U3722 ( .A(n3065), .B(n3047), .Z(n3145) );
  XOR U3723 ( .A(n3176), .B(n3177), .Z(n3047) );
  XOR U3724 ( .A(n3178), .B(n3076), .Z(n3065) );
  XNOR U3725 ( .A(n3053), .B(n3180), .Z(n3054) );
  AND U3726 ( .A(n2792), .B(n814), .Z(n3180) );
  XOR U3727 ( .A(n3184), .B(n3055), .Z(n3179) );
  NAND U3728 ( .A(n854), .B(n2660), .Z(n3055) );
  IV U3729 ( .A(n3057), .Z(n3184) );
  XNOR U3730 ( .A(n3062), .B(n3063), .Z(n3059) );
  NAND U3731 ( .A(n941), .B(n2413), .Z(n3063) );
  XNOR U3732 ( .A(n3061), .B(n3188), .Z(n3062) );
  AND U3733 ( .A(n2538), .B(n898), .Z(n3188) );
  XNOR U3734 ( .A(n3075), .B(n3064), .Z(n3178) );
  XOR U3735 ( .A(n3192), .B(n3193), .Z(n3064) );
  AND U3736 ( .A(n3194), .B(n3195), .Z(n3193) );
  XNOR U3737 ( .A(n3196), .B(n3197), .Z(n3195) );
  XOR U3738 ( .A(n3198), .B(n3192), .Z(n3196) );
  XOR U3739 ( .A(n3152), .B(n3199), .Z(n3194) );
  XNOR U3740 ( .A(n3192), .B(n3153), .Z(n3199) );
  XNOR U3741 ( .A(n3165), .B(n3201), .Z(n3166) );
  AND U3742 ( .A(n1852), .B(n1312), .Z(n3201) );
  XOR U3743 ( .A(n3205), .B(n3167), .Z(n3200) );
  NAND U3744 ( .A(n1383), .B(n1751), .Z(n3167) );
  IV U3745 ( .A(n3169), .Z(n3205) );
  XNOR U3746 ( .A(n3174), .B(n3175), .Z(n3171) );
  NAND U3747 ( .A(n1566), .B(n1546), .Z(n3175) );
  XNOR U3748 ( .A(n3173), .B(n3209), .Z(n3174) );
  AND U3749 ( .A(n1660), .B(n1460), .Z(n3209) );
  XOR U3750 ( .A(n3213), .B(n3162), .Z(n3152) );
  XNOR U3751 ( .A(n3149), .B(n3150), .Z(n3162) );
  NAND U3752 ( .A(n1242), .B(n1946), .Z(n3150) );
  XNOR U3753 ( .A(n3148), .B(n3214), .Z(n3149) );
  AND U3754 ( .A(n2047), .B(n1176), .Z(n3214) );
  XNOR U3755 ( .A(n3161), .B(n3151), .Z(n3213) );
  XNOR U3756 ( .A(n3156), .B(n3222), .Z(n3157) );
  AND U3757 ( .A(n2274), .B(n1055), .Z(n3222) );
  XOR U3758 ( .A(n3226), .B(n3158), .Z(n3221) );
  NAND U3759 ( .A(n1114), .B(n2160), .Z(n3158) );
  IV U3760 ( .A(n3160), .Z(n3226) );
  XOR U3761 ( .A(n3230), .B(n3231), .Z(n3192) );
  AND U3762 ( .A(n3232), .B(n3233), .Z(n3231) );
  XNOR U3763 ( .A(n3234), .B(n3235), .Z(n3233) );
  XNOR U3764 ( .A(n3230), .B(n3236), .Z(n3235) );
  XOR U3765 ( .A(n3219), .B(n3237), .Z(n3232) );
  XNOR U3766 ( .A(n3230), .B(n3220), .Z(n3237) );
  XNOR U3767 ( .A(n3202), .B(n3239), .Z(n3203) );
  AND U3768 ( .A(n1852), .B(n1383), .Z(n3239) );
  XOR U3769 ( .A(n3243), .B(n3204), .Z(n3238) );
  NAND U3770 ( .A(n1460), .B(n1751), .Z(n3204) );
  IV U3771 ( .A(n3206), .Z(n3243) );
  XNOR U3772 ( .A(n3211), .B(n3212), .Z(n3208) );
  NAND U3773 ( .A(n1566), .B(n1638), .Z(n3212) );
  XNOR U3774 ( .A(n3210), .B(n3247), .Z(n3211) );
  AND U3775 ( .A(n1546), .B(n1660), .Z(n3247) );
  XOR U3776 ( .A(n3251), .B(n3229), .Z(n3219) );
  XNOR U3777 ( .A(n3216), .B(n3217), .Z(n3229) );
  NAND U3778 ( .A(n1312), .B(n1946), .Z(n3217) );
  XNOR U3779 ( .A(n3215), .B(n3252), .Z(n3216) );
  AND U3780 ( .A(n2047), .B(n1242), .Z(n3252) );
  XNOR U3781 ( .A(n3228), .B(n3218), .Z(n3251) );
  XNOR U3782 ( .A(n3223), .B(n3260), .Z(n3224) );
  AND U3783 ( .A(n2274), .B(n1114), .Z(n3260) );
  XOR U3784 ( .A(n3264), .B(n3225), .Z(n3259) );
  NAND U3785 ( .A(n1176), .B(n2160), .Z(n3225) );
  IV U3786 ( .A(n3227), .Z(n3264) );
  XOR U3787 ( .A(n3268), .B(n3269), .Z(n3230) );
  AND U3788 ( .A(n3270), .B(n3271), .Z(n3269) );
  XNOR U3789 ( .A(n3272), .B(n3273), .Z(n3271) );
  XNOR U3790 ( .A(n3268), .B(n3274), .Z(n3273) );
  XOR U3791 ( .A(n3257), .B(n3275), .Z(n3270) );
  XNOR U3792 ( .A(n3268), .B(n3258), .Z(n3275) );
  XNOR U3793 ( .A(n3240), .B(n3277), .Z(n3241) );
  AND U3794 ( .A(n1852), .B(n1460), .Z(n3277) );
  XOR U3795 ( .A(n3281), .B(n3242), .Z(n3276) );
  NAND U3796 ( .A(n1751), .B(n1546), .Z(n3242) );
  IV U3797 ( .A(n3244), .Z(n3281) );
  XNOR U3798 ( .A(n3249), .B(n3250), .Z(n3246) );
  NAND U3799 ( .A(n1566), .B(n1731), .Z(n3250) );
  XNOR U3800 ( .A(n3248), .B(n3285), .Z(n3249) );
  AND U3801 ( .A(n1638), .B(n1660), .Z(n3285) );
  XOR U3802 ( .A(n3289), .B(n3267), .Z(n3257) );
  XNOR U3803 ( .A(n3254), .B(n3255), .Z(n3267) );
  NAND U3804 ( .A(n1383), .B(n1946), .Z(n3255) );
  XNOR U3805 ( .A(n3253), .B(n3290), .Z(n3254) );
  AND U3806 ( .A(n2047), .B(n1312), .Z(n3290) );
  XNOR U3807 ( .A(n3266), .B(n3256), .Z(n3289) );
  XNOR U3808 ( .A(n3261), .B(n3298), .Z(n3262) );
  AND U3809 ( .A(n2274), .B(n1176), .Z(n3298) );
  XOR U3810 ( .A(n3302), .B(n3263), .Z(n3297) );
  NAND U3811 ( .A(n1242), .B(n2160), .Z(n3263) );
  IV U3812 ( .A(n3265), .Z(n3302) );
  XOR U3813 ( .A(n3306), .B(n3307), .Z(n3268) );
  AND U3814 ( .A(n3308), .B(n3309), .Z(n3307) );
  XNOR U3815 ( .A(n3310), .B(n3311), .Z(n3309) );
  XNOR U3816 ( .A(n3306), .B(n3312), .Z(n3311) );
  XOR U3817 ( .A(n3295), .B(n3313), .Z(n3308) );
  XNOR U3818 ( .A(n3306), .B(n3296), .Z(n3313) );
  XNOR U3819 ( .A(n3278), .B(n3315), .Z(n3279) );
  AND U3820 ( .A(n1546), .B(n1852), .Z(n3315) );
  XOR U3821 ( .A(n3319), .B(n3280), .Z(n3314) );
  NAND U3822 ( .A(n1751), .B(n1638), .Z(n3280) );
  IV U3823 ( .A(n3282), .Z(n3319) );
  XNOR U3824 ( .A(n3287), .B(n3288), .Z(n3284) );
  NAND U3825 ( .A(n1566), .B(n1825), .Z(n3288) );
  XNOR U3826 ( .A(n3286), .B(n3323), .Z(n3287) );
  AND U3827 ( .A(n1731), .B(n1660), .Z(n3323) );
  XOR U3828 ( .A(n3327), .B(n3305), .Z(n3295) );
  XNOR U3829 ( .A(n3292), .B(n3293), .Z(n3305) );
  NAND U3830 ( .A(n1460), .B(n1946), .Z(n3293) );
  XNOR U3831 ( .A(n3291), .B(n3328), .Z(n3292) );
  AND U3832 ( .A(n2047), .B(n1383), .Z(n3328) );
  XNOR U3833 ( .A(n3304), .B(n3294), .Z(n3327) );
  XNOR U3834 ( .A(n3299), .B(n3336), .Z(n3300) );
  AND U3835 ( .A(n2274), .B(n1242), .Z(n3336) );
  XOR U3836 ( .A(n3340), .B(n3301), .Z(n3335) );
  NAND U3837 ( .A(n1312), .B(n2160), .Z(n3301) );
  IV U3838 ( .A(n3303), .Z(n3340) );
  XOR U3839 ( .A(n3344), .B(n3345), .Z(n3306) );
  AND U3840 ( .A(n3346), .B(n3347), .Z(n3345) );
  XNOR U3841 ( .A(n3348), .B(n3349), .Z(n3347) );
  XNOR U3842 ( .A(n3344), .B(n3350), .Z(n3349) );
  XOR U3843 ( .A(n3333), .B(n3351), .Z(n3346) );
  XNOR U3844 ( .A(n3344), .B(n3334), .Z(n3351) );
  XNOR U3845 ( .A(n3316), .B(n3353), .Z(n3317) );
  AND U3846 ( .A(n1638), .B(n1852), .Z(n3353) );
  XOR U3847 ( .A(n3357), .B(n3318), .Z(n3352) );
  NAND U3848 ( .A(n1751), .B(n1731), .Z(n3318) );
  IV U3849 ( .A(n3320), .Z(n3357) );
  XNOR U3850 ( .A(n3325), .B(n3326), .Z(n3322) );
  NAND U3851 ( .A(n1566), .B(n1925), .Z(n3326) );
  XNOR U3852 ( .A(n3324), .B(n3361), .Z(n3325) );
  AND U3853 ( .A(n1825), .B(n1660), .Z(n3361) );
  XOR U3854 ( .A(n3365), .B(n3343), .Z(n3333) );
  XNOR U3855 ( .A(n3330), .B(n3331), .Z(n3343) );
  NAND U3856 ( .A(n1946), .B(n1546), .Z(n3331) );
  XNOR U3857 ( .A(n3329), .B(n3366), .Z(n3330) );
  AND U3858 ( .A(n2047), .B(n1460), .Z(n3366) );
  XNOR U3859 ( .A(n3342), .B(n3332), .Z(n3365) );
  XNOR U3860 ( .A(n3337), .B(n3374), .Z(n3338) );
  AND U3861 ( .A(n2274), .B(n1312), .Z(n3374) );
  XOR U3862 ( .A(n3378), .B(n3339), .Z(n3373) );
  NAND U3863 ( .A(n1383), .B(n2160), .Z(n3339) );
  IV U3864 ( .A(n3341), .Z(n3378) );
  XOR U3865 ( .A(n3382), .B(n3383), .Z(n3344) );
  AND U3866 ( .A(n3384), .B(n3385), .Z(n3383) );
  XNOR U3867 ( .A(n3386), .B(n3387), .Z(n3385) );
  XNOR U3868 ( .A(n3382), .B(n3388), .Z(n3387) );
  XOR U3869 ( .A(n3371), .B(n3389), .Z(n3384) );
  XNOR U3870 ( .A(n3382), .B(n3372), .Z(n3389) );
  XNOR U3871 ( .A(n3354), .B(n3391), .Z(n3355) );
  AND U3872 ( .A(n1731), .B(n1852), .Z(n3391) );
  XOR U3873 ( .A(n3395), .B(n3356), .Z(n3390) );
  NAND U3874 ( .A(n1751), .B(n1825), .Z(n3356) );
  IV U3875 ( .A(n3358), .Z(n3395) );
  XNOR U3876 ( .A(n3363), .B(n3364), .Z(n3360) );
  NAND U3877 ( .A(n1566), .B(n2030), .Z(n3364) );
  XNOR U3878 ( .A(n3362), .B(n3399), .Z(n3363) );
  AND U3879 ( .A(n1925), .B(n1660), .Z(n3399) );
  XOR U3880 ( .A(n3403), .B(n3381), .Z(n3371) );
  XNOR U3881 ( .A(n3368), .B(n3369), .Z(n3381) );
  NAND U3882 ( .A(n1946), .B(n1638), .Z(n3369) );
  XNOR U3883 ( .A(n3367), .B(n3404), .Z(n3368) );
  AND U3884 ( .A(n1546), .B(n2047), .Z(n3404) );
  XNOR U3885 ( .A(n3380), .B(n3370), .Z(n3403) );
  XNOR U3886 ( .A(n3375), .B(n3412), .Z(n3376) );
  AND U3887 ( .A(n2274), .B(n1383), .Z(n3412) );
  XOR U3888 ( .A(n3416), .B(n3377), .Z(n3411) );
  NAND U3889 ( .A(n1460), .B(n2160), .Z(n3377) );
  IV U3890 ( .A(n3379), .Z(n3416) );
  XOR U3891 ( .A(n3420), .B(n3421), .Z(n3382) );
  AND U3892 ( .A(n3422), .B(n3423), .Z(n3421) );
  XNOR U3893 ( .A(n3424), .B(n3425), .Z(n3423) );
  XNOR U3894 ( .A(n3420), .B(n3426), .Z(n3425) );
  XOR U3895 ( .A(n3409), .B(n3427), .Z(n3422) );
  XNOR U3896 ( .A(n3420), .B(n3410), .Z(n3427) );
  XNOR U3897 ( .A(n3392), .B(n3429), .Z(n3393) );
  AND U3898 ( .A(n1825), .B(n1852), .Z(n3429) );
  XOR U3899 ( .A(n3433), .B(n3394), .Z(n3428) );
  NAND U3900 ( .A(n1751), .B(n1925), .Z(n3394) );
  IV U3901 ( .A(n3396), .Z(n3433) );
  XNOR U3902 ( .A(n3401), .B(n3402), .Z(n3398) );
  NAND U3903 ( .A(n1566), .B(n2135), .Z(n3402) );
  XNOR U3904 ( .A(n3400), .B(n3437), .Z(n3401) );
  AND U3905 ( .A(n2030), .B(n1660), .Z(n3437) );
  XOR U3906 ( .A(n3441), .B(n3419), .Z(n3409) );
  XNOR U3907 ( .A(n3406), .B(n3407), .Z(n3419) );
  NAND U3908 ( .A(n1946), .B(n1731), .Z(n3407) );
  XNOR U3909 ( .A(n3405), .B(n3442), .Z(n3406) );
  AND U3910 ( .A(n1638), .B(n2047), .Z(n3442) );
  XNOR U3911 ( .A(n3418), .B(n3408), .Z(n3441) );
  XNOR U3912 ( .A(n3413), .B(n3450), .Z(n3414) );
  AND U3913 ( .A(n2274), .B(n1460), .Z(n3450) );
  XOR U3914 ( .A(n3454), .B(n3415), .Z(n3449) );
  NAND U3915 ( .A(n2160), .B(n1546), .Z(n3415) );
  IV U3916 ( .A(n3417), .Z(n3454) );
  XOR U3917 ( .A(n3458), .B(n3459), .Z(n3420) );
  AND U3918 ( .A(n3460), .B(n3461), .Z(n3459) );
  XNOR U3919 ( .A(n3462), .B(n3463), .Z(n3461) );
  XNOR U3920 ( .A(n3458), .B(n3464), .Z(n3463) );
  XOR U3921 ( .A(n3447), .B(n3465), .Z(n3460) );
  XNOR U3922 ( .A(n3458), .B(n3448), .Z(n3465) );
  XNOR U3923 ( .A(n3430), .B(n3467), .Z(n3431) );
  AND U3924 ( .A(n1925), .B(n1852), .Z(n3467) );
  XOR U3925 ( .A(n3471), .B(n3432), .Z(n3466) );
  NAND U3926 ( .A(n1751), .B(n2030), .Z(n3432) );
  IV U3927 ( .A(n3434), .Z(n3471) );
  XNOR U3928 ( .A(n3439), .B(n3440), .Z(n3436) );
  NAND U3929 ( .A(n1566), .B(n2246), .Z(n3440) );
  XNOR U3930 ( .A(n3438), .B(n3475), .Z(n3439) );
  AND U3931 ( .A(n2135), .B(n1660), .Z(n3475) );
  XOR U3932 ( .A(n3479), .B(n3457), .Z(n3447) );
  XNOR U3933 ( .A(n3444), .B(n3445), .Z(n3457) );
  NAND U3934 ( .A(n1946), .B(n1825), .Z(n3445) );
  XNOR U3935 ( .A(n3443), .B(n3480), .Z(n3444) );
  AND U3936 ( .A(n1731), .B(n2047), .Z(n3480) );
  XNOR U3937 ( .A(n3456), .B(n3446), .Z(n3479) );
  XNOR U3938 ( .A(n3451), .B(n3488), .Z(n3452) );
  AND U3939 ( .A(n1546), .B(n2274), .Z(n3488) );
  XOR U3940 ( .A(n3492), .B(n3453), .Z(n3487) );
  NAND U3941 ( .A(n2160), .B(n1638), .Z(n3453) );
  IV U3942 ( .A(n3455), .Z(n3492) );
  XOR U3943 ( .A(n3496), .B(n3497), .Z(n3458) );
  AND U3944 ( .A(n3498), .B(n3499), .Z(n3497) );
  XNOR U3945 ( .A(n3500), .B(n3501), .Z(n3499) );
  XNOR U3946 ( .A(n3496), .B(n3502), .Z(n3501) );
  XOR U3947 ( .A(n3485), .B(n3503), .Z(n3498) );
  XNOR U3948 ( .A(n3496), .B(n3486), .Z(n3503) );
  XNOR U3949 ( .A(n3468), .B(n3505), .Z(n3469) );
  AND U3950 ( .A(n2030), .B(n1852), .Z(n3505) );
  XOR U3951 ( .A(n3509), .B(n3470), .Z(n3504) );
  NAND U3952 ( .A(n1751), .B(n2135), .Z(n3470) );
  IV U3953 ( .A(n3472), .Z(n3509) );
  XNOR U3954 ( .A(n3477), .B(n3478), .Z(n3474) );
  NAND U3955 ( .A(n1566), .B(n2362), .Z(n3478) );
  XNOR U3956 ( .A(n3476), .B(n3513), .Z(n3477) );
  AND U3957 ( .A(n2246), .B(n1660), .Z(n3513) );
  XOR U3958 ( .A(n3517), .B(n3495), .Z(n3485) );
  XNOR U3959 ( .A(n3482), .B(n3483), .Z(n3495) );
  NAND U3960 ( .A(n1946), .B(n1925), .Z(n3483) );
  XNOR U3961 ( .A(n3481), .B(n3518), .Z(n3482) );
  AND U3962 ( .A(n1825), .B(n2047), .Z(n3518) );
  XNOR U3963 ( .A(n3494), .B(n3484), .Z(n3517) );
  XNOR U3964 ( .A(n3489), .B(n3526), .Z(n3490) );
  AND U3965 ( .A(n1638), .B(n2274), .Z(n3526) );
  XOR U3966 ( .A(n3530), .B(n3491), .Z(n3525) );
  NAND U3967 ( .A(n2160), .B(n1731), .Z(n3491) );
  IV U3968 ( .A(n3493), .Z(n3530) );
  XOR U3969 ( .A(n3534), .B(n3535), .Z(n3496) );
  AND U3970 ( .A(n3536), .B(n3537), .Z(n3535) );
  XNOR U3971 ( .A(n3538), .B(n3539), .Z(n3537) );
  XNOR U3972 ( .A(n3534), .B(n3540), .Z(n3539) );
  XOR U3973 ( .A(n3523), .B(n3541), .Z(n3536) );
  XNOR U3974 ( .A(n3534), .B(n3524), .Z(n3541) );
  XNOR U3975 ( .A(n3506), .B(n3543), .Z(n3507) );
  AND U3976 ( .A(n2135), .B(n1852), .Z(n3543) );
  XOR U3977 ( .A(n3547), .B(n3508), .Z(n3542) );
  NAND U3978 ( .A(n1751), .B(n2246), .Z(n3508) );
  IV U3979 ( .A(n3510), .Z(n3547) );
  XNOR U3980 ( .A(n3515), .B(n3516), .Z(n3512) );
  NAND U3981 ( .A(n1566), .B(n2483), .Z(n3516) );
  XNOR U3982 ( .A(n3514), .B(n3551), .Z(n3515) );
  AND U3983 ( .A(n2362), .B(n1660), .Z(n3551) );
  XOR U3984 ( .A(n3555), .B(n3533), .Z(n3523) );
  XNOR U3985 ( .A(n3520), .B(n3521), .Z(n3533) );
  NAND U3986 ( .A(n1946), .B(n2030), .Z(n3521) );
  XNOR U3987 ( .A(n3519), .B(n3556), .Z(n3520) );
  AND U3988 ( .A(n1925), .B(n2047), .Z(n3556) );
  XNOR U3989 ( .A(n3532), .B(n3522), .Z(n3555) );
  XNOR U3990 ( .A(n3527), .B(n3564), .Z(n3528) );
  AND U3991 ( .A(n1731), .B(n2274), .Z(n3564) );
  XOR U3992 ( .A(n3568), .B(n3529), .Z(n3563) );
  NAND U3993 ( .A(n2160), .B(n1825), .Z(n3529) );
  IV U3994 ( .A(n3531), .Z(n3568) );
  XOR U3995 ( .A(n3572), .B(n3573), .Z(n3534) );
  AND U3996 ( .A(n3574), .B(n3575), .Z(n3573) );
  XNOR U3997 ( .A(n3576), .B(n3577), .Z(n3575) );
  XNOR U3998 ( .A(n3572), .B(n3578), .Z(n3577) );
  XOR U3999 ( .A(n3561), .B(n3579), .Z(n3574) );
  XNOR U4000 ( .A(n3572), .B(n3562), .Z(n3579) );
  XNOR U4001 ( .A(n3544), .B(n3581), .Z(n3545) );
  AND U4002 ( .A(n2246), .B(n1852), .Z(n3581) );
  XOR U4003 ( .A(n3585), .B(n3546), .Z(n3580) );
  NAND U4004 ( .A(n1751), .B(n2362), .Z(n3546) );
  IV U4005 ( .A(n3548), .Z(n3585) );
  XNOR U4006 ( .A(n3553), .B(n3554), .Z(n3550) );
  NAND U4007 ( .A(n1566), .B(n2607), .Z(n3554) );
  XNOR U4008 ( .A(n3552), .B(n3589), .Z(n3553) );
  AND U4009 ( .A(n2483), .B(n1660), .Z(n3589) );
  XOR U4010 ( .A(n3593), .B(n3571), .Z(n3561) );
  XNOR U4011 ( .A(n3558), .B(n3559), .Z(n3571) );
  NAND U4012 ( .A(n1946), .B(n2135), .Z(n3559) );
  XNOR U4013 ( .A(n3557), .B(n3594), .Z(n3558) );
  AND U4014 ( .A(n2030), .B(n2047), .Z(n3594) );
  XNOR U4015 ( .A(n3570), .B(n3560), .Z(n3593) );
  XNOR U4016 ( .A(n3565), .B(n3602), .Z(n3566) );
  AND U4017 ( .A(n1825), .B(n2274), .Z(n3602) );
  XOR U4018 ( .A(n3606), .B(n3567), .Z(n3601) );
  NAND U4019 ( .A(n2160), .B(n1925), .Z(n3567) );
  IV U4020 ( .A(n3569), .Z(n3606) );
  XOR U4021 ( .A(n3610), .B(n3611), .Z(n3572) );
  AND U4022 ( .A(n3612), .B(n3613), .Z(n3611) );
  XNOR U4023 ( .A(n3614), .B(n3615), .Z(n3613) );
  XNOR U4024 ( .A(n3610), .B(n3616), .Z(n3615) );
  XOR U4025 ( .A(n3599), .B(n3617), .Z(n3612) );
  XNOR U4026 ( .A(n3610), .B(n3600), .Z(n3617) );
  XNOR U4027 ( .A(n3582), .B(n3619), .Z(n3583) );
  AND U4028 ( .A(n2362), .B(n1852), .Z(n3619) );
  XOR U4029 ( .A(n3623), .B(n3584), .Z(n3618) );
  NAND U4030 ( .A(n1751), .B(n2483), .Z(n3584) );
  IV U4031 ( .A(n3586), .Z(n3623) );
  XNOR U4032 ( .A(n3591), .B(n3592), .Z(n3588) );
  NAND U4033 ( .A(n1566), .B(n2734), .Z(n3592) );
  XNOR U4034 ( .A(n3590), .B(n3627), .Z(n3591) );
  AND U4035 ( .A(n2607), .B(n1660), .Z(n3627) );
  XOR U4036 ( .A(n3631), .B(n3609), .Z(n3599) );
  XNOR U4037 ( .A(n3596), .B(n3597), .Z(n3609) );
  NAND U4038 ( .A(n1946), .B(n2246), .Z(n3597) );
  XNOR U4039 ( .A(n3595), .B(n3632), .Z(n3596) );
  AND U4040 ( .A(n2135), .B(n2047), .Z(n3632) );
  XNOR U4041 ( .A(n3608), .B(n3598), .Z(n3631) );
  XNOR U4042 ( .A(n3603), .B(n3640), .Z(n3604) );
  AND U4043 ( .A(n1925), .B(n2274), .Z(n3640) );
  XOR U4044 ( .A(n3644), .B(n3605), .Z(n3639) );
  NAND U4045 ( .A(n2160), .B(n2030), .Z(n3605) );
  IV U4046 ( .A(n3607), .Z(n3644) );
  XOR U4047 ( .A(n3648), .B(n3649), .Z(n3610) );
  AND U4048 ( .A(n3650), .B(n3651), .Z(n3649) );
  XNOR U4049 ( .A(n3652), .B(n3653), .Z(n3651) );
  XNOR U4050 ( .A(n3648), .B(n3654), .Z(n3653) );
  XOR U4051 ( .A(n3637), .B(n3655), .Z(n3650) );
  XNOR U4052 ( .A(n3648), .B(n3638), .Z(n3655) );
  XNOR U4053 ( .A(n3620), .B(n3657), .Z(n3621) );
  AND U4054 ( .A(n2483), .B(n1852), .Z(n3657) );
  XOR U4055 ( .A(n3661), .B(n3622), .Z(n3656) );
  NAND U4056 ( .A(n1751), .B(n2607), .Z(n3622) );
  IV U4057 ( .A(n3624), .Z(n3661) );
  XNOR U4058 ( .A(n3629), .B(n3630), .Z(n3626) );
  NANDN U4059 ( .B(n2866), .A(n1566), .Z(n3630) );
  XNOR U4060 ( .A(n3628), .B(n3665), .Z(n3629) );
  AND U4061 ( .A(n2734), .B(n1660), .Z(n3665) );
  XOR U4062 ( .A(n3669), .B(n3647), .Z(n3637) );
  XNOR U4063 ( .A(n3634), .B(n3635), .Z(n3647) );
  NAND U4064 ( .A(n1946), .B(n2362), .Z(n3635) );
  XNOR U4065 ( .A(n3633), .B(n3670), .Z(n3634) );
  AND U4066 ( .A(n2246), .B(n2047), .Z(n3670) );
  XNOR U4067 ( .A(n3646), .B(n3636), .Z(n3669) );
  XNOR U4068 ( .A(n3641), .B(n3678), .Z(n3642) );
  AND U4069 ( .A(n2030), .B(n2274), .Z(n3678) );
  XOR U4070 ( .A(n3682), .B(n3643), .Z(n3677) );
  NAND U4071 ( .A(n2160), .B(n2135), .Z(n3643) );
  IV U4072 ( .A(n3645), .Z(n3682) );
  XOR U4073 ( .A(n3686), .B(n3687), .Z(n3648) );
  AND U4074 ( .A(n3688), .B(n3689), .Z(n3687) );
  XNOR U4075 ( .A(n3690), .B(n3691), .Z(n3689) );
  XNOR U4076 ( .A(n3686), .B(n3692), .Z(n3691) );
  XOR U4077 ( .A(n3675), .B(n3693), .Z(n3688) );
  XNOR U4078 ( .A(n3686), .B(n3676), .Z(n3693) );
  XNOR U4079 ( .A(n3658), .B(n3695), .Z(n3659) );
  AND U4080 ( .A(n2607), .B(n1852), .Z(n3695) );
  XOR U4081 ( .A(n3699), .B(n3660), .Z(n3694) );
  NAND U4082 ( .A(n1751), .B(n2734), .Z(n3660) );
  IV U4083 ( .A(n3662), .Z(n3699) );
  XNOR U4084 ( .A(n3667), .B(n3668), .Z(n3664) );
  NANDN U4085 ( .B(n3004), .A(n1566), .Z(n3668) );
  XNOR U4086 ( .A(n3666), .B(n3703), .Z(n3667) );
  ANDN U4087 ( .A(n1660), .B(n2866), .Z(n3703) );
  XOR U4088 ( .A(n3707), .B(n3685), .Z(n3675) );
  XNOR U4089 ( .A(n3672), .B(n3673), .Z(n3685) );
  NAND U4090 ( .A(n1946), .B(n2483), .Z(n3673) );
  XNOR U4091 ( .A(n3671), .B(n3708), .Z(n3672) );
  AND U4092 ( .A(n2362), .B(n2047), .Z(n3708) );
  XNOR U4093 ( .A(n3684), .B(n3674), .Z(n3707) );
  XNOR U4094 ( .A(n3679), .B(n3716), .Z(n3680) );
  AND U4095 ( .A(n2135), .B(n2274), .Z(n3716) );
  XOR U4096 ( .A(n3720), .B(n3681), .Z(n3715) );
  NAND U4097 ( .A(n2160), .B(n2246), .Z(n3681) );
  IV U4098 ( .A(n3683), .Z(n3720) );
  XOR U4099 ( .A(n3724), .B(n3725), .Z(n3686) );
  AND U4100 ( .A(n3726), .B(n3727), .Z(n3725) );
  XNOR U4101 ( .A(n3728), .B(n3729), .Z(n3727) );
  XNOR U4102 ( .A(n3724), .B(n3730), .Z(n3729) );
  XOR U4103 ( .A(n3713), .B(n3731), .Z(n3726) );
  XNOR U4104 ( .A(n3724), .B(n3714), .Z(n3731) );
  XNOR U4105 ( .A(n3696), .B(n3733), .Z(n3697) );
  AND U4106 ( .A(n2734), .B(n1852), .Z(n3733) );
  XOR U4107 ( .A(n3737), .B(n3698), .Z(n3732) );
  NANDN U4108 ( .B(n2866), .A(n1751), .Z(n3698) );
  IV U4109 ( .A(n3700), .Z(n3737) );
  XNOR U4110 ( .A(n3705), .B(n3706), .Z(n3702) );
  NAND U4111 ( .A(n1566), .B(n3139), .Z(n3706) );
  XNOR U4112 ( .A(n3704), .B(n3741), .Z(n3705) );
  ANDN U4113 ( .A(n1660), .B(n3004), .Z(n3741) );
  XOR U4114 ( .A(n3745), .B(n3723), .Z(n3713) );
  XNOR U4115 ( .A(n3710), .B(n3711), .Z(n3723) );
  NAND U4116 ( .A(n1946), .B(n2607), .Z(n3711) );
  XNOR U4117 ( .A(n3709), .B(n3746), .Z(n3710) );
  AND U4118 ( .A(n2483), .B(n2047), .Z(n3746) );
  XNOR U4119 ( .A(n3722), .B(n3712), .Z(n3745) );
  XNOR U4120 ( .A(n3717), .B(n3754), .Z(n3718) );
  AND U4121 ( .A(n2246), .B(n2274), .Z(n3754) );
  XOR U4122 ( .A(n3758), .B(n3719), .Z(n3753) );
  NAND U4123 ( .A(n2160), .B(n2362), .Z(n3719) );
  IV U4124 ( .A(n3721), .Z(n3758) );
  XNOR U4125 ( .A(n3763), .B(n3764), .Z(n3177) );
  XOR U4126 ( .A(n3765), .B(n3762), .Z(n3763) );
  XNOR U4127 ( .A(n3766), .B(n3761), .Z(n3751) );
  XNOR U4128 ( .A(n3748), .B(n3749), .Z(n3761) );
  NAND U4129 ( .A(n1946), .B(n2734), .Z(n3749) );
  XNOR U4130 ( .A(n3747), .B(n3767), .Z(n3748) );
  AND U4131 ( .A(n2607), .B(n2047), .Z(n3767) );
  XNOR U4132 ( .A(n3771), .B(n3768), .Z(n3770) );
  XNOR U4133 ( .A(n3760), .B(n3750), .Z(n3766) );
  XOR U4134 ( .A(n3772), .B(n3773), .Z(n3750) );
  XNOR U4135 ( .A(n3755), .B(n3775), .Z(n3756) );
  AND U4136 ( .A(n2362), .B(n2274), .Z(n3775) );
  XNOR U4137 ( .A(n3779), .B(n3776), .Z(n3778) );
  XOR U4138 ( .A(n3780), .B(n3757), .Z(n3774) );
  NAND U4139 ( .A(n2160), .B(n2483), .Z(n3757) );
  IV U4140 ( .A(n3759), .Z(n3780) );
  XNOR U4141 ( .A(n3781), .B(n3782), .Z(n3759) );
  AND U4142 ( .A(n3783), .B(n3784), .Z(n3782) );
  XOR U4143 ( .A(n3777), .B(n3785), .Z(n3784) );
  XNOR U4144 ( .A(n3779), .B(n3781), .Z(n3785) );
  NAND U4145 ( .A(n2160), .B(n2607), .Z(n3779) );
  XOR U4146 ( .A(n3776), .B(n3786), .Z(n3777) );
  AND U4147 ( .A(n2483), .B(n2274), .Z(n3786) );
  XNOR U4148 ( .A(n3790), .B(n3787), .Z(n3789) );
  XOR U4149 ( .A(n3769), .B(n3791), .Z(n3783) );
  XNOR U4150 ( .A(n3771), .B(n3781), .Z(n3791) );
  NANDN U4151 ( .B(n2866), .A(n1946), .Z(n3771) );
  XOR U4152 ( .A(n3768), .B(n3792), .Z(n3769) );
  AND U4153 ( .A(n2734), .B(n2047), .Z(n3792) );
  XNOR U4154 ( .A(n3796), .B(n3793), .Z(n3795) );
  XOR U4155 ( .A(n3797), .B(n3798), .Z(n3781) );
  AND U4156 ( .A(n3799), .B(n3800), .Z(n3798) );
  XOR U4157 ( .A(n3788), .B(n3801), .Z(n3800) );
  XNOR U4158 ( .A(n3790), .B(n3797), .Z(n3801) );
  NAND U4159 ( .A(n2160), .B(n2734), .Z(n3790) );
  XOR U4160 ( .A(n3787), .B(n3802), .Z(n3788) );
  AND U4161 ( .A(n2607), .B(n2274), .Z(n3802) );
  XNOR U4162 ( .A(n3806), .B(n3803), .Z(n3805) );
  XOR U4163 ( .A(n3794), .B(n3807), .Z(n3799) );
  XNOR U4164 ( .A(n3796), .B(n3797), .Z(n3807) );
  NANDN U4165 ( .B(n3004), .A(n1946), .Z(n3796) );
  XOR U4166 ( .A(n3793), .B(n3808), .Z(n3794) );
  ANDN U4167 ( .A(n2047), .B(n2866), .Z(n3808) );
  XNOR U4168 ( .A(n3812), .B(n3809), .Z(n3811) );
  XOR U4169 ( .A(n3813), .B(n3814), .Z(n3797) );
  AND U4170 ( .A(n3815), .B(n3816), .Z(n3814) );
  XOR U4171 ( .A(n3804), .B(n3817), .Z(n3816) );
  XNOR U4172 ( .A(n3806), .B(n3813), .Z(n3817) );
  NANDN U4173 ( .B(n2866), .A(n2160), .Z(n3806) );
  XOR U4174 ( .A(n3803), .B(n3818), .Z(n3804) );
  AND U4175 ( .A(n2734), .B(n2274), .Z(n3818) );
  XOR U4176 ( .A(n3810), .B(n3822), .Z(n3815) );
  XNOR U4177 ( .A(n3812), .B(n3813), .Z(n3822) );
  NAND U4178 ( .A(n1946), .B(n3139), .Z(n3812) );
  XOR U4179 ( .A(n3809), .B(n3823), .Z(n3810) );
  ANDN U4180 ( .A(n2047), .B(n3004), .Z(n3823) );
  NAND U4181 ( .A(n1946), .B(n3828), .Z(n3826) );
  XNOR U4182 ( .A(n3824), .B(n3829), .Z(n3825) );
  AND U4183 ( .A(n3139), .B(n2047), .Z(n3829) );
  AND U4184 ( .A(n3830), .B(g_input[0]), .Z(n3824) );
  NANDN U4185 ( .B(n1946), .A(n3831), .Z(n3830) );
  NAND U4186 ( .A(n3828), .B(n2047), .Z(n3831) );
  XNOR U4187 ( .A(n3819), .B(n3835), .Z(n3820) );
  ANDN U4188 ( .A(n2274), .B(n2866), .Z(n3835) );
  XOR U4189 ( .A(n3838), .B(n3836), .Z(n3837) );
  ANDN U4190 ( .A(n2274), .B(n3004), .Z(n3838) );
  AND U4191 ( .A(n3139), .B(n2160), .Z(n3839) );
  XOR U4192 ( .A(n3843), .B(n3821), .Z(n3834) );
  NANDN U4193 ( .B(n3004), .A(n2160), .Z(n3821) );
  IV U4194 ( .A(n3827), .Z(n3843) );
  NAND U4195 ( .A(n2160), .B(n3828), .Z(n3842) );
  XNOR U4196 ( .A(n3840), .B(n3844), .Z(n3841) );
  AND U4197 ( .A(n3139), .B(n2274), .Z(n3844) );
  AND U4198 ( .A(n3845), .B(g_input[0]), .Z(n3840) );
  NANDN U4199 ( .B(n2160), .A(n3846), .Z(n3845) );
  NAND U4200 ( .A(n3828), .B(n2274), .Z(n3846) );
  XNOR U4201 ( .A(n3734), .B(n3850), .Z(n3735) );
  ANDN U4202 ( .A(n1852), .B(n2866), .Z(n3850) );
  XOR U4203 ( .A(n3853), .B(n3851), .Z(n3852) );
  ANDN U4204 ( .A(n1852), .B(n3004), .Z(n3853) );
  AND U4205 ( .A(n3139), .B(n1751), .Z(n3854) );
  XOR U4206 ( .A(n3858), .B(n3736), .Z(n3849) );
  NANDN U4207 ( .B(n3004), .A(n1751), .Z(n3736) );
  IV U4208 ( .A(n3738), .Z(n3858) );
  NAND U4209 ( .A(n1751), .B(n3828), .Z(n3857) );
  XNOR U4210 ( .A(n3855), .B(n3859), .Z(n3856) );
  AND U4211 ( .A(n3139), .B(n1852), .Z(n3859) );
  AND U4212 ( .A(n3860), .B(g_input[0]), .Z(n3855) );
  NANDN U4213 ( .B(n1751), .A(n3861), .Z(n3860) );
  NAND U4214 ( .A(n3828), .B(n1852), .Z(n3861) );
  XNOR U4215 ( .A(n3743), .B(n3744), .Z(n3740) );
  NAND U4216 ( .A(n1566), .B(n3828), .Z(n3744) );
  XNOR U4217 ( .A(n3742), .B(n3864), .Z(n3743) );
  AND U4218 ( .A(n3139), .B(n1660), .Z(n3864) );
  AND U4219 ( .A(n3865), .B(g_input[0]), .Z(n3742) );
  NANDN U4220 ( .B(n1566), .A(n3866), .Z(n3865) );
  NAND U4221 ( .A(n3828), .B(n1660), .Z(n3866) );
  XOR U4222 ( .A(n3869), .B(n3870), .Z(n3762) );
  XNOR U4223 ( .A(n3871), .B(n3078), .Z(n3075) );
  NAND U4224 ( .A(n774), .B(n2938), .Z(n3073) );
  XNOR U4225 ( .A(n3071), .B(n3872), .Z(n3072) );
  AND U4226 ( .A(n3070), .B(n740), .Z(n3872) );
  XNOR U4227 ( .A(n3077), .B(n3074), .Z(n3871) );
  XNOR U4228 ( .A(n3181), .B(n3878), .Z(n3182) );
  AND U4229 ( .A(n2792), .B(n854), .Z(n3878) );
  XOR U4230 ( .A(n3882), .B(n3183), .Z(n3877) );
  NAND U4231 ( .A(n898), .B(n2660), .Z(n3183) );
  IV U4232 ( .A(n3185), .Z(n3882) );
  XNOR U4233 ( .A(n3190), .B(n3191), .Z(n3187) );
  NAND U4234 ( .A(n999), .B(n2413), .Z(n3191) );
  XNOR U4235 ( .A(n3189), .B(n3886), .Z(n3190) );
  AND U4236 ( .A(n2538), .B(n941), .Z(n3886) );
  XOR U4237 ( .A(n3890), .B(n3891), .Z(n3198) );
  XNOR U4238 ( .A(n3892), .B(n3876), .Z(n3890) );
  XOR U4239 ( .A(n3894), .B(n3895), .Z(n3236) );
  XNOR U4240 ( .A(n3896), .B(n3893), .Z(n3894) );
  XNOR U4241 ( .A(n3879), .B(n3898), .Z(n3880) );
  AND U4242 ( .A(n2792), .B(n898), .Z(n3898) );
  XOR U4243 ( .A(n3902), .B(n3881), .Z(n3897) );
  NAND U4244 ( .A(n941), .B(n2660), .Z(n3881) );
  IV U4245 ( .A(n3883), .Z(n3902) );
  XNOR U4246 ( .A(n3888), .B(n3889), .Z(n3885) );
  NAND U4247 ( .A(n1055), .B(n2413), .Z(n3889) );
  XNOR U4248 ( .A(n3887), .B(n3906), .Z(n3888) );
  AND U4249 ( .A(n2538), .B(n999), .Z(n3906) );
  XOR U4250 ( .A(n3911), .B(n3912), .Z(n3274) );
  XNOR U4251 ( .A(n3913), .B(n3910), .Z(n3911) );
  XNOR U4252 ( .A(n3899), .B(n3915), .Z(n3900) );
  AND U4253 ( .A(n2792), .B(n941), .Z(n3915) );
  XOR U4254 ( .A(n3919), .B(n3901), .Z(n3914) );
  NAND U4255 ( .A(n999), .B(n2660), .Z(n3901) );
  IV U4256 ( .A(n3903), .Z(n3919) );
  XNOR U4257 ( .A(n3908), .B(n3909), .Z(n3905) );
  NAND U4258 ( .A(n1114), .B(n2413), .Z(n3909) );
  XNOR U4259 ( .A(n3907), .B(n3923), .Z(n3908) );
  AND U4260 ( .A(n2538), .B(n1055), .Z(n3923) );
  XOR U4261 ( .A(n3928), .B(n3929), .Z(n3312) );
  XNOR U4262 ( .A(n3930), .B(n3927), .Z(n3928) );
  XNOR U4263 ( .A(n3916), .B(n3932), .Z(n3917) );
  AND U4264 ( .A(n2792), .B(n999), .Z(n3932) );
  XOR U4265 ( .A(n3936), .B(n3918), .Z(n3931) );
  NAND U4266 ( .A(n1055), .B(n2660), .Z(n3918) );
  IV U4267 ( .A(n3920), .Z(n3936) );
  XNOR U4268 ( .A(n3925), .B(n3926), .Z(n3922) );
  NAND U4269 ( .A(n1176), .B(n2413), .Z(n3926) );
  XNOR U4270 ( .A(n3924), .B(n3940), .Z(n3925) );
  AND U4271 ( .A(n2538), .B(n1114), .Z(n3940) );
  XOR U4272 ( .A(n3945), .B(n3946), .Z(n3350) );
  XNOR U4273 ( .A(n3947), .B(n3944), .Z(n3945) );
  XNOR U4274 ( .A(n3933), .B(n3949), .Z(n3934) );
  AND U4275 ( .A(n2792), .B(n1055), .Z(n3949) );
  XOR U4276 ( .A(n3953), .B(n3935), .Z(n3948) );
  NAND U4277 ( .A(n1114), .B(n2660), .Z(n3935) );
  IV U4278 ( .A(n3937), .Z(n3953) );
  XNOR U4279 ( .A(n3942), .B(n3943), .Z(n3939) );
  NAND U4280 ( .A(n1242), .B(n2413), .Z(n3943) );
  XNOR U4281 ( .A(n3941), .B(n3957), .Z(n3942) );
  AND U4282 ( .A(n2538), .B(n1176), .Z(n3957) );
  XOR U4283 ( .A(n3962), .B(n3963), .Z(n3388) );
  XNOR U4284 ( .A(n3964), .B(n3961), .Z(n3962) );
  XNOR U4285 ( .A(n3950), .B(n3966), .Z(n3951) );
  AND U4286 ( .A(n2792), .B(n1114), .Z(n3966) );
  XOR U4287 ( .A(n3970), .B(n3952), .Z(n3965) );
  NAND U4288 ( .A(n1176), .B(n2660), .Z(n3952) );
  IV U4289 ( .A(n3954), .Z(n3970) );
  XNOR U4290 ( .A(n3959), .B(n3960), .Z(n3956) );
  NAND U4291 ( .A(n1312), .B(n2413), .Z(n3960) );
  XNOR U4292 ( .A(n3958), .B(n3974), .Z(n3959) );
  AND U4293 ( .A(n2538), .B(n1242), .Z(n3974) );
  XOR U4294 ( .A(n3979), .B(n3980), .Z(n3426) );
  XNOR U4295 ( .A(n3981), .B(n3978), .Z(n3979) );
  XNOR U4296 ( .A(n3967), .B(n3983), .Z(n3968) );
  AND U4297 ( .A(n2792), .B(n1176), .Z(n3983) );
  XOR U4298 ( .A(n3987), .B(n3969), .Z(n3982) );
  NAND U4299 ( .A(n1242), .B(n2660), .Z(n3969) );
  IV U4300 ( .A(n3971), .Z(n3987) );
  XNOR U4301 ( .A(n3976), .B(n3977), .Z(n3973) );
  NAND U4302 ( .A(n1383), .B(n2413), .Z(n3977) );
  XNOR U4303 ( .A(n3975), .B(n3991), .Z(n3976) );
  AND U4304 ( .A(n2538), .B(n1312), .Z(n3991) );
  XOR U4305 ( .A(n3996), .B(n3997), .Z(n3464) );
  XNOR U4306 ( .A(n3998), .B(n3995), .Z(n3996) );
  XNOR U4307 ( .A(n3984), .B(n4000), .Z(n3985) );
  AND U4308 ( .A(n2792), .B(n1242), .Z(n4000) );
  XOR U4309 ( .A(n4004), .B(n3986), .Z(n3999) );
  NAND U4310 ( .A(n1312), .B(n2660), .Z(n3986) );
  IV U4311 ( .A(n3988), .Z(n4004) );
  XNOR U4312 ( .A(n3993), .B(n3994), .Z(n3990) );
  NAND U4313 ( .A(n1460), .B(n2413), .Z(n3994) );
  XNOR U4314 ( .A(n3992), .B(n4008), .Z(n3993) );
  AND U4315 ( .A(n2538), .B(n1383), .Z(n4008) );
  XOR U4316 ( .A(n4013), .B(n4014), .Z(n3502) );
  XNOR U4317 ( .A(n4015), .B(n4012), .Z(n4013) );
  XNOR U4318 ( .A(n4001), .B(n4017), .Z(n4002) );
  AND U4319 ( .A(n2792), .B(n1312), .Z(n4017) );
  XOR U4320 ( .A(n4021), .B(n4003), .Z(n4016) );
  NAND U4321 ( .A(n1383), .B(n2660), .Z(n4003) );
  IV U4322 ( .A(n4005), .Z(n4021) );
  XNOR U4323 ( .A(n4010), .B(n4011), .Z(n4007) );
  NAND U4324 ( .A(n1546), .B(n2413), .Z(n4011) );
  XNOR U4325 ( .A(n4009), .B(n4025), .Z(n4010) );
  AND U4326 ( .A(n2538), .B(n1460), .Z(n4025) );
  XOR U4327 ( .A(n4030), .B(n4031), .Z(n3540) );
  XNOR U4328 ( .A(n4032), .B(n4029), .Z(n4030) );
  XNOR U4329 ( .A(n4018), .B(n4034), .Z(n4019) );
  AND U4330 ( .A(n2792), .B(n1383), .Z(n4034) );
  XOR U4331 ( .A(n4038), .B(n4020), .Z(n4033) );
  NAND U4332 ( .A(n1460), .B(n2660), .Z(n4020) );
  IV U4333 ( .A(n4022), .Z(n4038) );
  XNOR U4334 ( .A(n4027), .B(n4028), .Z(n4024) );
  NAND U4335 ( .A(n1638), .B(n2413), .Z(n4028) );
  XNOR U4336 ( .A(n4026), .B(n4042), .Z(n4027) );
  AND U4337 ( .A(n2538), .B(n1546), .Z(n4042) );
  XOR U4338 ( .A(n4047), .B(n4048), .Z(n3578) );
  XNOR U4339 ( .A(n4049), .B(n4046), .Z(n4047) );
  XNOR U4340 ( .A(n4035), .B(n4051), .Z(n4036) );
  AND U4341 ( .A(n2792), .B(n1460), .Z(n4051) );
  XOR U4342 ( .A(n4055), .B(n4037), .Z(n4050) );
  NAND U4343 ( .A(n1546), .B(n2660), .Z(n4037) );
  IV U4344 ( .A(n4039), .Z(n4055) );
  XNOR U4345 ( .A(n4044), .B(n4045), .Z(n4041) );
  NAND U4346 ( .A(n1731), .B(n2413), .Z(n4045) );
  XNOR U4347 ( .A(n4043), .B(n4059), .Z(n4044) );
  AND U4348 ( .A(n2538), .B(n1638), .Z(n4059) );
  XOR U4349 ( .A(n4064), .B(n4065), .Z(n3616) );
  XNOR U4350 ( .A(n4066), .B(n4063), .Z(n4064) );
  XNOR U4351 ( .A(n4052), .B(n4068), .Z(n4053) );
  AND U4352 ( .A(n2792), .B(n1546), .Z(n4068) );
  XOR U4353 ( .A(n4072), .B(n4054), .Z(n4067) );
  NAND U4354 ( .A(n1638), .B(n2660), .Z(n4054) );
  IV U4355 ( .A(n4056), .Z(n4072) );
  XNOR U4356 ( .A(n4061), .B(n4062), .Z(n4058) );
  NAND U4357 ( .A(n1825), .B(n2413), .Z(n4062) );
  XNOR U4358 ( .A(n4060), .B(n4076), .Z(n4061) );
  AND U4359 ( .A(n2538), .B(n1731), .Z(n4076) );
  XOR U4360 ( .A(n4081), .B(n4082), .Z(n3654) );
  XNOR U4361 ( .A(n4083), .B(n4080), .Z(n4081) );
  XNOR U4362 ( .A(n4069), .B(n4085), .Z(n4070) );
  AND U4363 ( .A(n2792), .B(n1638), .Z(n4085) );
  XOR U4364 ( .A(n4089), .B(n4071), .Z(n4084) );
  NAND U4365 ( .A(n1731), .B(n2660), .Z(n4071) );
  IV U4366 ( .A(n4073), .Z(n4089) );
  XNOR U4367 ( .A(n4078), .B(n4079), .Z(n4075) );
  NAND U4368 ( .A(n1925), .B(n2413), .Z(n4079) );
  XNOR U4369 ( .A(n4077), .B(n4093), .Z(n4078) );
  AND U4370 ( .A(n2538), .B(n1825), .Z(n4093) );
  XOR U4371 ( .A(n4098), .B(n4099), .Z(n3692) );
  XNOR U4372 ( .A(n4100), .B(n4097), .Z(n4098) );
  XNOR U4373 ( .A(n4086), .B(n4102), .Z(n4087) );
  AND U4374 ( .A(n2792), .B(n1731), .Z(n4102) );
  XOR U4375 ( .A(n4106), .B(n4088), .Z(n4101) );
  NAND U4376 ( .A(n1825), .B(n2660), .Z(n4088) );
  IV U4377 ( .A(n4090), .Z(n4106) );
  XNOR U4378 ( .A(n4095), .B(n4096), .Z(n4092) );
  NAND U4379 ( .A(n2030), .B(n2413), .Z(n4096) );
  XNOR U4380 ( .A(n4094), .B(n4110), .Z(n4095) );
  AND U4381 ( .A(n2538), .B(n1925), .Z(n4110) );
  XOR U4382 ( .A(n4115), .B(n4116), .Z(n3730) );
  XNOR U4383 ( .A(n4117), .B(n4114), .Z(n4115) );
  XNOR U4384 ( .A(n4103), .B(n4119), .Z(n4104) );
  AND U4385 ( .A(n2792), .B(n1825), .Z(n4119) );
  XOR U4386 ( .A(n4123), .B(n4105), .Z(n4118) );
  NAND U4387 ( .A(n1925), .B(n2660), .Z(n4105) );
  IV U4388 ( .A(n4107), .Z(n4123) );
  XNOR U4389 ( .A(n4112), .B(n4113), .Z(n4109) );
  NAND U4390 ( .A(n2135), .B(n2413), .Z(n4113) );
  XNOR U4391 ( .A(n4111), .B(n4127), .Z(n4112) );
  AND U4392 ( .A(n2538), .B(n2030), .Z(n4127) );
  XOR U4393 ( .A(n4132), .B(n4133), .Z(n3765) );
  XNOR U4394 ( .A(n4134), .B(n4131), .Z(n4132) );
  XNOR U4395 ( .A(n4120), .B(n4136), .Z(n4121) );
  AND U4396 ( .A(n2792), .B(n1925), .Z(n4136) );
  XOR U4397 ( .A(n4140), .B(n4122), .Z(n4135) );
  NAND U4398 ( .A(n2030), .B(n2660), .Z(n4122) );
  IV U4399 ( .A(n4124), .Z(n4140) );
  XNOR U4400 ( .A(n4129), .B(n4130), .Z(n4126) );
  NAND U4401 ( .A(n2246), .B(n2413), .Z(n4130) );
  XNOR U4402 ( .A(n4128), .B(n4144), .Z(n4129) );
  AND U4403 ( .A(n2538), .B(n2135), .Z(n4144) );
  XOR U4404 ( .A(n4148), .B(n4149), .Z(n4131) );
  AND U4405 ( .A(n4150), .B(n4151), .Z(n4149) );
  XOR U4406 ( .A(n4152), .B(n4153), .Z(n4151) );
  XOR U4407 ( .A(n4148), .B(n4154), .Z(n4153) );
  XOR U4408 ( .A(n4142), .B(n4155), .Z(n4150) );
  XOR U4409 ( .A(n4148), .B(n4143), .Z(n4155) );
  NAND U4410 ( .A(n2413), .B(n2362), .Z(n4147) );
  XNOR U4411 ( .A(n4145), .B(n4156), .Z(n4146) );
  AND U4412 ( .A(n2538), .B(n2246), .Z(n4156) );
  XNOR U4413 ( .A(n4137), .B(n4161), .Z(n4138) );
  AND U4414 ( .A(n2792), .B(n2030), .Z(n4161) );
  XOR U4415 ( .A(n4165), .B(n4139), .Z(n4160) );
  NAND U4416 ( .A(n2135), .B(n2660), .Z(n4139) );
  IV U4417 ( .A(n4141), .Z(n4165) );
  XOR U4418 ( .A(n4169), .B(n4170), .Z(n4148) );
  AND U4419 ( .A(n4171), .B(n4172), .Z(n4170) );
  XOR U4420 ( .A(n4173), .B(n4174), .Z(n4172) );
  XOR U4421 ( .A(n4169), .B(n4175), .Z(n4174) );
  XOR U4422 ( .A(n4167), .B(n4176), .Z(n4171) );
  XOR U4423 ( .A(n4169), .B(n4168), .Z(n4176) );
  NAND U4424 ( .A(n2413), .B(n2483), .Z(n4159) );
  XNOR U4425 ( .A(n4157), .B(n4177), .Z(n4158) );
  AND U4426 ( .A(n2362), .B(n2538), .Z(n4177) );
  XNOR U4427 ( .A(n4162), .B(n4182), .Z(n4163) );
  AND U4428 ( .A(n2792), .B(n2135), .Z(n4182) );
  XOR U4429 ( .A(n4186), .B(n4164), .Z(n4181) );
  NAND U4430 ( .A(n2246), .B(n2660), .Z(n4164) );
  IV U4431 ( .A(n4166), .Z(n4186) );
  XOR U4432 ( .A(n4190), .B(n4191), .Z(n4169) );
  AND U4433 ( .A(n4192), .B(n4193), .Z(n4191) );
  XOR U4434 ( .A(n4194), .B(n4195), .Z(n4193) );
  XOR U4435 ( .A(n4190), .B(n4196), .Z(n4195) );
  XOR U4436 ( .A(n4188), .B(n4197), .Z(n4192) );
  XOR U4437 ( .A(n4190), .B(n4189), .Z(n4197) );
  NAND U4438 ( .A(n2413), .B(n2607), .Z(n4180) );
  XNOR U4439 ( .A(n4178), .B(n4198), .Z(n4179) );
  AND U4440 ( .A(n2483), .B(n2538), .Z(n4198) );
  XNOR U4441 ( .A(n4183), .B(n4203), .Z(n4184) );
  AND U4442 ( .A(n2792), .B(n2246), .Z(n4203) );
  XOR U4443 ( .A(n4207), .B(n4185), .Z(n4202) );
  NAND U4444 ( .A(n2660), .B(n2362), .Z(n4185) );
  IV U4445 ( .A(n4187), .Z(n4207) );
  XOR U4446 ( .A(n4211), .B(n4212), .Z(n4190) );
  AND U4447 ( .A(n4213), .B(n4214), .Z(n4212) );
  XOR U4448 ( .A(n4215), .B(n4216), .Z(n4214) );
  XOR U4449 ( .A(n4211), .B(n4217), .Z(n4216) );
  XOR U4450 ( .A(n4209), .B(n4218), .Z(n4213) );
  XOR U4451 ( .A(n4211), .B(n4210), .Z(n4218) );
  NAND U4452 ( .A(n2413), .B(n2734), .Z(n4201) );
  XNOR U4453 ( .A(n4199), .B(n4219), .Z(n4200) );
  AND U4454 ( .A(n2607), .B(n2538), .Z(n4219) );
  XNOR U4455 ( .A(n4204), .B(n4224), .Z(n4205) );
  AND U4456 ( .A(n2362), .B(n2792), .Z(n4224) );
  XOR U4457 ( .A(n4228), .B(n4206), .Z(n4223) );
  NAND U4458 ( .A(n2660), .B(n2483), .Z(n4206) );
  IV U4459 ( .A(n4208), .Z(n4228) );
  XOR U4460 ( .A(n4232), .B(n4233), .Z(n4211) );
  AND U4461 ( .A(n4234), .B(n4235), .Z(n4233) );
  XOR U4462 ( .A(n4236), .B(n4237), .Z(n4235) );
  XOR U4463 ( .A(n4232), .B(n4238), .Z(n4237) );
  XOR U4464 ( .A(n4230), .B(n4239), .Z(n4234) );
  XOR U4465 ( .A(n4232), .B(n4231), .Z(n4239) );
  NANDN U4466 ( .B(n2866), .A(n2413), .Z(n4222) );
  XNOR U4467 ( .A(n4220), .B(n4240), .Z(n4221) );
  AND U4468 ( .A(n2734), .B(n2538), .Z(n4240) );
  XNOR U4469 ( .A(n4225), .B(n4245), .Z(n4226) );
  AND U4470 ( .A(n2483), .B(n2792), .Z(n4245) );
  XOR U4471 ( .A(n4249), .B(n4227), .Z(n4244) );
  NAND U4472 ( .A(n2660), .B(n2607), .Z(n4227) );
  IV U4473 ( .A(n4229), .Z(n4249) );
  XOR U4474 ( .A(n4253), .B(n4254), .Z(n4232) );
  AND U4475 ( .A(n4255), .B(n4256), .Z(n4254) );
  XOR U4476 ( .A(n4257), .B(n4258), .Z(n4256) );
  XOR U4477 ( .A(n4253), .B(n4259), .Z(n4258) );
  XOR U4478 ( .A(n4251), .B(n4260), .Z(n4255) );
  XOR U4479 ( .A(n4253), .B(n4252), .Z(n4260) );
  NANDN U4480 ( .B(n3004), .A(n2413), .Z(n4243) );
  XNOR U4481 ( .A(n4241), .B(n4261), .Z(n4242) );
  ANDN U4482 ( .A(n2538), .B(n2866), .Z(n4261) );
  XNOR U4483 ( .A(n4246), .B(n4266), .Z(n4247) );
  AND U4484 ( .A(n2607), .B(n2792), .Z(n4266) );
  XOR U4485 ( .A(n4270), .B(n4248), .Z(n4265) );
  NAND U4486 ( .A(n2660), .B(n2734), .Z(n4248) );
  IV U4487 ( .A(n4250), .Z(n4270) );
  XOR U4488 ( .A(n4274), .B(n4275), .Z(n4253) );
  AND U4489 ( .A(n4276), .B(n4277), .Z(n4275) );
  XOR U4490 ( .A(n4278), .B(n4279), .Z(n4277) );
  XOR U4491 ( .A(n4274), .B(n4280), .Z(n4279) );
  XOR U4492 ( .A(n4272), .B(n4281), .Z(n4276) );
  XOR U4493 ( .A(n4274), .B(n4273), .Z(n4281) );
  NAND U4494 ( .A(n2413), .B(n3139), .Z(n4264) );
  XNOR U4495 ( .A(n4262), .B(n4282), .Z(n4263) );
  ANDN U4496 ( .A(n2538), .B(n3004), .Z(n4282) );
  XNOR U4497 ( .A(n4267), .B(n4287), .Z(n4268) );
  AND U4498 ( .A(n2734), .B(n2792), .Z(n4287) );
  XOR U4499 ( .A(n4291), .B(n4269), .Z(n4286) );
  NANDN U4500 ( .B(n2866), .A(n2660), .Z(n4269) );
  IV U4501 ( .A(n4271), .Z(n4291) );
  XOR U4502 ( .A(n4296), .B(n4297), .Z(n3870) );
  XNOR U4503 ( .A(n4298), .B(n4295), .Z(n4296) );
  XNOR U4504 ( .A(n4288), .B(n4300), .Z(n4289) );
  ANDN U4505 ( .A(n2792), .B(n2866), .Z(n4300) );
  XOR U4506 ( .A(n4303), .B(n4301), .Z(n4302) );
  ANDN U4507 ( .A(n2792), .B(n3004), .Z(n4303) );
  AND U4508 ( .A(n3139), .B(n2660), .Z(n4304) );
  XOR U4509 ( .A(n4308), .B(n4290), .Z(n4299) );
  NANDN U4510 ( .B(n3004), .A(n2660), .Z(n4290) );
  IV U4511 ( .A(n4292), .Z(n4308) );
  NAND U4512 ( .A(n2660), .B(n3828), .Z(n4307) );
  XNOR U4513 ( .A(n4305), .B(n4309), .Z(n4306) );
  AND U4514 ( .A(n3139), .B(n2792), .Z(n4309) );
  AND U4515 ( .A(n4310), .B(g_input[0]), .Z(n4305) );
  NANDN U4516 ( .B(n2660), .A(n4311), .Z(n4310) );
  NAND U4517 ( .A(n3828), .B(n2792), .Z(n4311) );
  XNOR U4518 ( .A(n4284), .B(n4285), .Z(n4294) );
  NAND U4519 ( .A(n2413), .B(n3828), .Z(n4285) );
  XNOR U4520 ( .A(n4283), .B(n4314), .Z(n4284) );
  AND U4521 ( .A(n3139), .B(n2538), .Z(n4314) );
  AND U4522 ( .A(n4315), .B(g_input[0]), .Z(n4283) );
  NANDN U4523 ( .B(n2413), .A(n4316), .Z(n4315) );
  NAND U4524 ( .A(n3828), .B(n2538), .Z(n4316) );
  XOR U4525 ( .A(n4319), .B(n4320), .Z(n4295) );
  AND U4526 ( .A(n4322), .B(n4323), .Z(n4321) );
  NANDN U4527 ( .B(n710), .A(n4324), .Z(n4323) );
  OR U4528 ( .A(n4325), .B(n4326), .Z(n4322) );
  XNOR U4529 ( .A(n4328), .B(n4327), .Z(n3892) );
  XNOR U4530 ( .A(n4329), .B(n4325), .Z(n4328) );
  NAND U4531 ( .A(n740), .B(n4324), .Z(n4325) );
  NANDN U4532 ( .B(n710), .A(e_input[0]), .Z(n4330) );
  NANDN U4533 ( .B(n4331), .A(n4332), .Z(n710) );
  AND U4534 ( .A(n4333), .B(g_input[31]), .Z(n4332) );
  NAND U4535 ( .A(n814), .B(n2938), .Z(n3875) );
  XNOR U4536 ( .A(n3873), .B(n4337), .Z(n3874) );
  AND U4537 ( .A(n3070), .B(n774), .Z(n4337) );
  NAND U4538 ( .A(n854), .B(n2938), .Z(n4340) );
  XNOR U4539 ( .A(n4338), .B(n4342), .Z(n4339) );
  AND U4540 ( .A(n3070), .B(n814), .Z(n4342) );
  XNOR U4541 ( .A(n4334), .B(n4347), .Z(n4335) );
  AND U4542 ( .A(n740), .B(e_input[0]), .Z(n4347) );
  XNOR U4543 ( .A(n4333), .B(g_input[30]), .Z(n4331) );
  NOR U4544 ( .A(n4348), .B(n4349), .Z(n4333) );
  XOR U4545 ( .A(n4353), .B(n4336), .Z(n4346) );
  NAND U4546 ( .A(n774), .B(n4324), .Z(n4336) );
  IV U4547 ( .A(n4341), .Z(n4353) );
  NAND U4548 ( .A(n898), .B(n2938), .Z(n4345) );
  XNOR U4549 ( .A(n4343), .B(n4355), .Z(n4344) );
  AND U4550 ( .A(n3070), .B(n854), .Z(n4355) );
  XNOR U4551 ( .A(n4350), .B(n4360), .Z(n4351) );
  AND U4552 ( .A(n774), .B(e_input[0]), .Z(n4360) );
  XOR U4553 ( .A(n4348), .B(g_input[29]), .Z(n4349) );
  NANDN U4554 ( .B(n4361), .A(n4362), .Z(n4348) );
  XOR U4555 ( .A(n4366), .B(n4352), .Z(n4359) );
  NAND U4556 ( .A(n814), .B(n4324), .Z(n4352) );
  IV U4557 ( .A(n4354), .Z(n4366) );
  NAND U4558 ( .A(n941), .B(n2938), .Z(n4358) );
  XNOR U4559 ( .A(n4356), .B(n4368), .Z(n4357) );
  AND U4560 ( .A(n3070), .B(n898), .Z(n4368) );
  XNOR U4561 ( .A(n4363), .B(n4373), .Z(n4364) );
  AND U4562 ( .A(n814), .B(e_input[0]), .Z(n4373) );
  XNOR U4563 ( .A(n4362), .B(g_input[28]), .Z(n4361) );
  NOR U4564 ( .A(n4374), .B(n4375), .Z(n4362) );
  XOR U4565 ( .A(n4379), .B(n4365), .Z(n4372) );
  NAND U4566 ( .A(n854), .B(n4324), .Z(n4365) );
  IV U4567 ( .A(n4367), .Z(n4379) );
  NAND U4568 ( .A(n999), .B(n2938), .Z(n4371) );
  XNOR U4569 ( .A(n4369), .B(n4381), .Z(n4370) );
  AND U4570 ( .A(n3070), .B(n941), .Z(n4381) );
  XNOR U4571 ( .A(n4376), .B(n4386), .Z(n4377) );
  AND U4572 ( .A(n854), .B(e_input[0]), .Z(n4386) );
  XOR U4573 ( .A(n4374), .B(g_input[27]), .Z(n4375) );
  NANDN U4574 ( .B(n4387), .A(n4388), .Z(n4374) );
  XOR U4575 ( .A(n4392), .B(n4378), .Z(n4385) );
  NAND U4576 ( .A(n898), .B(n4324), .Z(n4378) );
  IV U4577 ( .A(n4380), .Z(n4392) );
  NAND U4578 ( .A(n1055), .B(n2938), .Z(n4384) );
  XNOR U4579 ( .A(n4382), .B(n4394), .Z(n4383) );
  AND U4580 ( .A(n3070), .B(n999), .Z(n4394) );
  XNOR U4581 ( .A(n4389), .B(n4399), .Z(n4390) );
  AND U4582 ( .A(n898), .B(e_input[0]), .Z(n4399) );
  XNOR U4583 ( .A(n4388), .B(g_input[26]), .Z(n4387) );
  NOR U4584 ( .A(n4400), .B(n4401), .Z(n4388) );
  XOR U4585 ( .A(n4405), .B(n4391), .Z(n4398) );
  NAND U4586 ( .A(n941), .B(n4324), .Z(n4391) );
  IV U4587 ( .A(n4393), .Z(n4405) );
  NAND U4588 ( .A(n1114), .B(n2938), .Z(n4397) );
  XNOR U4589 ( .A(n4395), .B(n4407), .Z(n4396) );
  AND U4590 ( .A(n3070), .B(n1055), .Z(n4407) );
  XNOR U4591 ( .A(n4402), .B(n4412), .Z(n4403) );
  AND U4592 ( .A(n941), .B(e_input[0]), .Z(n4412) );
  XOR U4593 ( .A(n4400), .B(g_input[25]), .Z(n4401) );
  NANDN U4594 ( .B(n4413), .A(n4414), .Z(n4400) );
  XOR U4595 ( .A(n4418), .B(n4404), .Z(n4411) );
  NAND U4596 ( .A(n999), .B(n4324), .Z(n4404) );
  IV U4597 ( .A(n4406), .Z(n4418) );
  NAND U4598 ( .A(n1176), .B(n2938), .Z(n4410) );
  XNOR U4599 ( .A(n4408), .B(n4420), .Z(n4409) );
  AND U4600 ( .A(n3070), .B(n1114), .Z(n4420) );
  XNOR U4601 ( .A(n4415), .B(n4425), .Z(n4416) );
  AND U4602 ( .A(n999), .B(e_input[0]), .Z(n4425) );
  XNOR U4603 ( .A(n4414), .B(g_input[24]), .Z(n4413) );
  NOR U4604 ( .A(n4426), .B(n4427), .Z(n4414) );
  XOR U4605 ( .A(n4431), .B(n4417), .Z(n4424) );
  NAND U4606 ( .A(n1055), .B(n4324), .Z(n4417) );
  IV U4607 ( .A(n4419), .Z(n4431) );
  NAND U4608 ( .A(n1242), .B(n2938), .Z(n4423) );
  XNOR U4609 ( .A(n4421), .B(n4433), .Z(n4422) );
  AND U4610 ( .A(n3070), .B(n1176), .Z(n4433) );
  XNOR U4611 ( .A(n4428), .B(n4438), .Z(n4429) );
  AND U4612 ( .A(n1055), .B(e_input[0]), .Z(n4438) );
  XOR U4613 ( .A(n4426), .B(g_input[23]), .Z(n4427) );
  NANDN U4614 ( .B(n4439), .A(n4440), .Z(n4426) );
  XOR U4615 ( .A(n4444), .B(n4430), .Z(n4437) );
  NAND U4616 ( .A(n1114), .B(n4324), .Z(n4430) );
  IV U4617 ( .A(n4432), .Z(n4444) );
  NAND U4618 ( .A(n1312), .B(n2938), .Z(n4436) );
  XNOR U4619 ( .A(n4434), .B(n4446), .Z(n4435) );
  AND U4620 ( .A(n3070), .B(n1242), .Z(n4446) );
  XNOR U4621 ( .A(n4441), .B(n4451), .Z(n4442) );
  AND U4622 ( .A(n1114), .B(e_input[0]), .Z(n4451) );
  XNOR U4623 ( .A(n4440), .B(g_input[22]), .Z(n4439) );
  NOR U4624 ( .A(n4452), .B(n4453), .Z(n4440) );
  XOR U4625 ( .A(n4457), .B(n4443), .Z(n4450) );
  NAND U4626 ( .A(n1176), .B(n4324), .Z(n4443) );
  IV U4627 ( .A(n4445), .Z(n4457) );
  NAND U4628 ( .A(n1383), .B(n2938), .Z(n4449) );
  XNOR U4629 ( .A(n4447), .B(n4459), .Z(n4448) );
  AND U4630 ( .A(n3070), .B(n1312), .Z(n4459) );
  XNOR U4631 ( .A(n4454), .B(n4464), .Z(n4455) );
  AND U4632 ( .A(n1176), .B(e_input[0]), .Z(n4464) );
  XOR U4633 ( .A(n4452), .B(g_input[21]), .Z(n4453) );
  NANDN U4634 ( .B(n4465), .A(n4466), .Z(n4452) );
  XOR U4635 ( .A(n4470), .B(n4456), .Z(n4463) );
  NAND U4636 ( .A(n1242), .B(n4324), .Z(n4456) );
  IV U4637 ( .A(n4458), .Z(n4470) );
  NAND U4638 ( .A(n1460), .B(n2938), .Z(n4462) );
  XNOR U4639 ( .A(n4460), .B(n4472), .Z(n4461) );
  AND U4640 ( .A(n3070), .B(n1383), .Z(n4472) );
  XNOR U4641 ( .A(n4467), .B(n4477), .Z(n4468) );
  AND U4642 ( .A(n1242), .B(e_input[0]), .Z(n4477) );
  XNOR U4643 ( .A(n4466), .B(g_input[20]), .Z(n4465) );
  NOR U4644 ( .A(n4478), .B(n4479), .Z(n4466) );
  XOR U4645 ( .A(n4483), .B(n4469), .Z(n4476) );
  NAND U4646 ( .A(n1312), .B(n4324), .Z(n4469) );
  IV U4647 ( .A(n4471), .Z(n4483) );
  NAND U4648 ( .A(n1546), .B(n2938), .Z(n4475) );
  XNOR U4649 ( .A(n4473), .B(n4485), .Z(n4474) );
  AND U4650 ( .A(n3070), .B(n1460), .Z(n4485) );
  XNOR U4651 ( .A(n4480), .B(n4490), .Z(n4481) );
  AND U4652 ( .A(n1312), .B(e_input[0]), .Z(n4490) );
  XOR U4653 ( .A(n4478), .B(g_input[19]), .Z(n4479) );
  NANDN U4654 ( .B(n4491), .A(n4492), .Z(n4478) );
  XOR U4655 ( .A(n4496), .B(n4482), .Z(n4489) );
  NAND U4656 ( .A(n1383), .B(n4324), .Z(n4482) );
  IV U4657 ( .A(n4484), .Z(n4496) );
  NAND U4658 ( .A(n1638), .B(n2938), .Z(n4488) );
  XNOR U4659 ( .A(n4486), .B(n4498), .Z(n4487) );
  AND U4660 ( .A(n3070), .B(n1546), .Z(n4498) );
  XNOR U4661 ( .A(n4493), .B(n4503), .Z(n4494) );
  AND U4662 ( .A(n1383), .B(e_input[0]), .Z(n4503) );
  XNOR U4663 ( .A(n4492), .B(g_input[18]), .Z(n4491) );
  NOR U4664 ( .A(n4504), .B(n4505), .Z(n4492) );
  XOR U4665 ( .A(n4509), .B(n4495), .Z(n4502) );
  NAND U4666 ( .A(n1460), .B(n4324), .Z(n4495) );
  IV U4667 ( .A(n4497), .Z(n4509) );
  XOR U4668 ( .A(n4510), .B(n4511), .Z(n4497) );
  AND U4669 ( .A(n4117), .B(n4512), .Z(n4511) );
  XNOR U4670 ( .A(n4510), .B(n4116), .Z(n4512) );
  NAND U4671 ( .A(n1731), .B(n2938), .Z(n4501) );
  XNOR U4672 ( .A(n4499), .B(n4513), .Z(n4500) );
  AND U4673 ( .A(n3070), .B(n1638), .Z(n4513) );
  XNOR U4674 ( .A(n4506), .B(n4518), .Z(n4507) );
  AND U4675 ( .A(n1460), .B(e_input[0]), .Z(n4518) );
  XOR U4676 ( .A(n4504), .B(g_input[17]), .Z(n4505) );
  NANDN U4677 ( .B(n4519), .A(n4520), .Z(n4504) );
  XOR U4678 ( .A(n4524), .B(n4508), .Z(n4517) );
  NAND U4679 ( .A(n1546), .B(n4324), .Z(n4508) );
  IV U4680 ( .A(n4510), .Z(n4524) );
  XOR U4681 ( .A(n4525), .B(n4526), .Z(n4510) );
  AND U4682 ( .A(n4134), .B(n4527), .Z(n4526) );
  XNOR U4683 ( .A(n4525), .B(n4133), .Z(n4527) );
  NAND U4684 ( .A(n1825), .B(n2938), .Z(n4516) );
  XNOR U4685 ( .A(n4514), .B(n4528), .Z(n4515) );
  AND U4686 ( .A(n3070), .B(n1731), .Z(n4528) );
  XNOR U4687 ( .A(n4521), .B(n4533), .Z(n4522) );
  AND U4688 ( .A(n1546), .B(e_input[0]), .Z(n4533) );
  XOR U4689 ( .A(n4537), .B(n4523), .Z(n4532) );
  NAND U4690 ( .A(n1638), .B(n4324), .Z(n4523) );
  IV U4691 ( .A(n4525), .Z(n4537) );
  NAND U4692 ( .A(n1925), .B(n2938), .Z(n4531) );
  XNOR U4693 ( .A(n4529), .B(n4539), .Z(n4530) );
  AND U4694 ( .A(n3070), .B(n1825), .Z(n4539) );
  XNOR U4695 ( .A(n4534), .B(n4544), .Z(n4535) );
  AND U4696 ( .A(n1638), .B(e_input[0]), .Z(n4544) );
  XOR U4697 ( .A(n4548), .B(n4536), .Z(n4543) );
  NAND U4698 ( .A(n1731), .B(n4324), .Z(n4536) );
  IV U4699 ( .A(n4538), .Z(n4548) );
  NAND U4700 ( .A(n2030), .B(n2938), .Z(n4542) );
  XNOR U4701 ( .A(n4540), .B(n4550), .Z(n4541) );
  AND U4702 ( .A(n3070), .B(n1925), .Z(n4550) );
  XNOR U4703 ( .A(n4545), .B(n4555), .Z(n4546) );
  AND U4704 ( .A(n1731), .B(e_input[0]), .Z(n4555) );
  XOR U4705 ( .A(n4559), .B(n4547), .Z(n4554) );
  NAND U4706 ( .A(n1825), .B(n4324), .Z(n4547) );
  IV U4707 ( .A(n4549), .Z(n4559) );
  NAND U4708 ( .A(n2135), .B(n2938), .Z(n4553) );
  XNOR U4709 ( .A(n4551), .B(n4561), .Z(n4552) );
  AND U4710 ( .A(n3070), .B(n2030), .Z(n4561) );
  XNOR U4711 ( .A(n4556), .B(n4566), .Z(n4557) );
  AND U4712 ( .A(n1825), .B(e_input[0]), .Z(n4566) );
  XOR U4713 ( .A(n4570), .B(n4558), .Z(n4565) );
  NAND U4714 ( .A(n1925), .B(n4324), .Z(n4558) );
  IV U4715 ( .A(n4560), .Z(n4570) );
  NAND U4716 ( .A(n2246), .B(n2938), .Z(n4564) );
  XNOR U4717 ( .A(n4562), .B(n4572), .Z(n4563) );
  AND U4718 ( .A(n3070), .B(n2135), .Z(n4572) );
  XNOR U4719 ( .A(n4567), .B(n4577), .Z(n4568) );
  AND U4720 ( .A(n1925), .B(e_input[0]), .Z(n4577) );
  XOR U4721 ( .A(n4581), .B(n4569), .Z(n4576) );
  NAND U4722 ( .A(n2030), .B(n4324), .Z(n4569) );
  IV U4723 ( .A(n4571), .Z(n4581) );
  NAND U4724 ( .A(n2362), .B(n2938), .Z(n4575) );
  XNOR U4725 ( .A(n4573), .B(n4583), .Z(n4574) );
  AND U4726 ( .A(n3070), .B(n2246), .Z(n4583) );
  XNOR U4727 ( .A(n4578), .B(n4588), .Z(n4579) );
  AND U4728 ( .A(n2030), .B(e_input[0]), .Z(n4588) );
  XOR U4729 ( .A(n4592), .B(n4580), .Z(n4587) );
  NAND U4730 ( .A(n2135), .B(n4324), .Z(n4580) );
  IV U4731 ( .A(n4582), .Z(n4592) );
  NAND U4732 ( .A(n2483), .B(n2938), .Z(n4586) );
  XNOR U4733 ( .A(n4584), .B(n4594), .Z(n4585) );
  AND U4734 ( .A(n3070), .B(n2362), .Z(n4594) );
  XNOR U4735 ( .A(n4589), .B(n4599), .Z(n4590) );
  AND U4736 ( .A(n2135), .B(e_input[0]), .Z(n4599) );
  XOR U4737 ( .A(n4603), .B(n4591), .Z(n4598) );
  NAND U4738 ( .A(n2246), .B(n4324), .Z(n4591) );
  IV U4739 ( .A(n4593), .Z(n4603) );
  NAND U4740 ( .A(n2607), .B(n2938), .Z(n4597) );
  XNOR U4741 ( .A(n4595), .B(n4605), .Z(n4596) );
  AND U4742 ( .A(n3070), .B(n2483), .Z(n4605) );
  XNOR U4743 ( .A(n4600), .B(n4610), .Z(n4601) );
  AND U4744 ( .A(n2246), .B(e_input[0]), .Z(n4610) );
  XOR U4745 ( .A(n4614), .B(n4602), .Z(n4609) );
  NAND U4746 ( .A(n2362), .B(n4324), .Z(n4602) );
  IV U4747 ( .A(n4604), .Z(n4614) );
  NAND U4748 ( .A(n2734), .B(n2938), .Z(n4608) );
  XNOR U4749 ( .A(n4606), .B(n4616), .Z(n4607) );
  AND U4750 ( .A(n3070), .B(n2607), .Z(n4616) );
  XNOR U4751 ( .A(n4620), .B(n4617), .Z(n4619) );
  XNOR U4752 ( .A(n4611), .B(n4622), .Z(n4612) );
  AND U4753 ( .A(n2362), .B(e_input[0]), .Z(n4622) );
  XNOR U4754 ( .A(n4626), .B(n4623), .Z(n4625) );
  XOR U4755 ( .A(n4627), .B(n4613), .Z(n4621) );
  NAND U4756 ( .A(n2483), .B(n4324), .Z(n4613) );
  IV U4757 ( .A(n4615), .Z(n4627) );
  XNOR U4758 ( .A(n4628), .B(n4629), .Z(n4615) );
  AND U4759 ( .A(n4630), .B(n4631), .Z(n4629) );
  XOR U4760 ( .A(n4624), .B(n4632), .Z(n4631) );
  XNOR U4761 ( .A(n4626), .B(n4628), .Z(n4632) );
  NAND U4762 ( .A(n2607), .B(n4324), .Z(n4626) );
  XOR U4763 ( .A(n4623), .B(n4633), .Z(n4624) );
  AND U4764 ( .A(n2483), .B(e_input[0]), .Z(n4633) );
  XNOR U4765 ( .A(n4637), .B(n4634), .Z(n4636) );
  XOR U4766 ( .A(n4618), .B(n4638), .Z(n4630) );
  XNOR U4767 ( .A(n4620), .B(n4628), .Z(n4638) );
  NANDN U4768 ( .B(n2866), .A(n2938), .Z(n4620) );
  XOR U4769 ( .A(n4617), .B(n4639), .Z(n4618) );
  AND U4770 ( .A(n3070), .B(n2734), .Z(n4639) );
  XNOR U4771 ( .A(n4643), .B(n4640), .Z(n4642) );
  XOR U4772 ( .A(n4644), .B(n4645), .Z(n4628) );
  AND U4773 ( .A(n4646), .B(n4647), .Z(n4645) );
  XOR U4774 ( .A(n4635), .B(n4648), .Z(n4647) );
  XNOR U4775 ( .A(n4637), .B(n4644), .Z(n4648) );
  NAND U4776 ( .A(n2734), .B(n4324), .Z(n4637) );
  XOR U4777 ( .A(n4634), .B(n4649), .Z(n4635) );
  AND U4778 ( .A(n2607), .B(e_input[0]), .Z(n4649) );
  XNOR U4779 ( .A(n4653), .B(n4650), .Z(n4652) );
  XOR U4780 ( .A(n4641), .B(n4654), .Z(n4646) );
  XNOR U4781 ( .A(n4643), .B(n4644), .Z(n4654) );
  NANDN U4782 ( .B(n3004), .A(n2938), .Z(n4643) );
  XOR U4783 ( .A(n4640), .B(n4655), .Z(n4641) );
  ANDN U4784 ( .A(n3070), .B(n2866), .Z(n4655) );
  XNOR U4785 ( .A(n4659), .B(n4656), .Z(n4658) );
  XOR U4786 ( .A(n4660), .B(n4661), .Z(n4644) );
  AND U4787 ( .A(n4662), .B(n4663), .Z(n4661) );
  XOR U4788 ( .A(n4651), .B(n4664), .Z(n4663) );
  XNOR U4789 ( .A(n4653), .B(n4660), .Z(n4664) );
  NANDN U4790 ( .B(n2866), .A(n4324), .Z(n4653) );
  XOR U4791 ( .A(n4650), .B(n4665), .Z(n4651) );
  AND U4792 ( .A(n2734), .B(e_input[0]), .Z(n4665) );
  XOR U4793 ( .A(n4657), .B(n4669), .Z(n4662) );
  XNOR U4794 ( .A(n4659), .B(n4660), .Z(n4669) );
  NAND U4795 ( .A(n2938), .B(n3139), .Z(n4659) );
  XOR U4796 ( .A(n4656), .B(n4670), .Z(n4657) );
  ANDN U4797 ( .A(n3070), .B(n3004), .Z(n4670) );
  NAND U4798 ( .A(n2938), .B(n3828), .Z(n4673) );
  XNOR U4799 ( .A(n4671), .B(n4675), .Z(n4672) );
  AND U4800 ( .A(n3139), .B(n3070), .Z(n4675) );
  AND U4801 ( .A(n4676), .B(g_input[0]), .Z(n4671) );
  NANDN U4802 ( .B(n2938), .A(n4677), .Z(n4676) );
  NAND U4803 ( .A(n3828), .B(n3070), .Z(n4677) );
  XNOR U4804 ( .A(n4666), .B(n4681), .Z(n4667) );
  ANDN U4805 ( .A(e_input[0]), .B(n2866), .Z(n4681) );
  XOR U4806 ( .A(n4684), .B(n4682), .Z(n4683) );
  ANDN U4807 ( .A(e_input[0]), .B(n3004), .Z(n4684) );
  AND U4808 ( .A(n4324), .B(n3139), .Z(n4685) );
  XOR U4809 ( .A(n4689), .B(n4668), .Z(n4680) );
  NANDN U4810 ( .B(n3004), .A(n4324), .Z(n4668) );
  IV U4811 ( .A(n4674), .Z(n4689) );
  NAND U4812 ( .A(n4324), .B(n3828), .Z(n4688) );
  XNOR U4813 ( .A(n4686), .B(n4690), .Z(n4687) );
  AND U4814 ( .A(n3139), .B(e_input[0]), .Z(n4690) );
  AND U4815 ( .A(n4691), .B(g_input[0]), .Z(n4686) );
  NANDN U4816 ( .B(n4324), .A(n4692), .Z(n4691) );
  NAND U4817 ( .A(n3828), .B(e_input[0]), .Z(n4692) );
  XNOR U4818 ( .A(n4694), .B(n3103), .Z(n3094) );
  XNOR U4819 ( .A(n3082), .B(n4696), .Z(n3083) );
  AND U4820 ( .A(n1925), .B(n1194), .Z(n4696) );
  XOR U4821 ( .A(n4700), .B(n3084), .Z(n4695) );
  NAND U4822 ( .A(n1136), .B(n2030), .Z(n3084) );
  IV U4823 ( .A(n3086), .Z(n4700) );
  XNOR U4824 ( .A(n3091), .B(n3092), .Z(n3088) );
  NANDN U4825 ( .B(n1020), .A(n2246), .Z(n3092) );
  XNOR U4826 ( .A(n3090), .B(n4704), .Z(n3091) );
  AND U4827 ( .A(n2135), .B(n1079), .Z(n4704) );
  XNOR U4828 ( .A(n3102), .B(n3093), .Z(n4694) );
  XOR U4829 ( .A(n4708), .B(n4709), .Z(n3093) );
  XOR U4830 ( .A(n4710), .B(n3112), .Z(n3102) );
  XNOR U4831 ( .A(n3099), .B(n3100), .Z(n3112) );
  NAND U4832 ( .A(n1280), .B(n1825), .Z(n3100) );
  XNOR U4833 ( .A(n3098), .B(n4711), .Z(n3099) );
  AND U4834 ( .A(n1731), .B(n1348), .Z(n4711) );
  XNOR U4835 ( .A(n3111), .B(n3101), .Z(n4710) );
  XOR U4836 ( .A(n4715), .B(n4716), .Z(n3101) );
  AND U4837 ( .A(n4717), .B(n4718), .Z(n4716) );
  XOR U4838 ( .A(n4719), .B(n4720), .Z(n4718) );
  XOR U4839 ( .A(n4715), .B(n4721), .Z(n4720) );
  XOR U4840 ( .A(n4702), .B(n4722), .Z(n4717) );
  XOR U4841 ( .A(n4715), .B(n4703), .Z(n4722) );
  NANDN U4842 ( .B(n1020), .A(n2362), .Z(n4707) );
  XNOR U4843 ( .A(n4705), .B(n4723), .Z(n4706) );
  AND U4844 ( .A(n2246), .B(n1079), .Z(n4723) );
  XNOR U4845 ( .A(n4697), .B(n4728), .Z(n4698) );
  AND U4846 ( .A(n2030), .B(n1194), .Z(n4728) );
  XOR U4847 ( .A(n4732), .B(n4699), .Z(n4727) );
  NAND U4848 ( .A(n1136), .B(n2135), .Z(n4699) );
  IV U4849 ( .A(n4701), .Z(n4732) );
  XOR U4850 ( .A(n4736), .B(n4737), .Z(n4715) );
  AND U4851 ( .A(n4738), .B(n4739), .Z(n4737) );
  XOR U4852 ( .A(n4740), .B(n4741), .Z(n4739) );
  XOR U4853 ( .A(n4736), .B(n4742), .Z(n4741) );
  XOR U4854 ( .A(n4734), .B(n4743), .Z(n4738) );
  XOR U4855 ( .A(n4736), .B(n4735), .Z(n4743) );
  NANDN U4856 ( .B(n1020), .A(n2483), .Z(n4726) );
  XNOR U4857 ( .A(n4724), .B(n4744), .Z(n4725) );
  AND U4858 ( .A(n2362), .B(n1079), .Z(n4744) );
  XNOR U4859 ( .A(n4729), .B(n4749), .Z(n4730) );
  AND U4860 ( .A(n2135), .B(n1194), .Z(n4749) );
  XOR U4861 ( .A(n4753), .B(n4731), .Z(n4748) );
  NAND U4862 ( .A(n1136), .B(n2246), .Z(n4731) );
  IV U4863 ( .A(n4733), .Z(n4753) );
  XOR U4864 ( .A(n4757), .B(n4758), .Z(n4736) );
  AND U4865 ( .A(n4759), .B(n4760), .Z(n4758) );
  XOR U4866 ( .A(n4761), .B(n4762), .Z(n4760) );
  XOR U4867 ( .A(n4757), .B(n4763), .Z(n4762) );
  XOR U4868 ( .A(n4755), .B(n4764), .Z(n4759) );
  XOR U4869 ( .A(n4757), .B(n4756), .Z(n4764) );
  NANDN U4870 ( .B(n1020), .A(n2607), .Z(n4747) );
  XNOR U4871 ( .A(n4745), .B(n4765), .Z(n4746) );
  AND U4872 ( .A(n2483), .B(n1079), .Z(n4765) );
  XNOR U4873 ( .A(n4750), .B(n4770), .Z(n4751) );
  AND U4874 ( .A(n2246), .B(n1194), .Z(n4770) );
  XOR U4875 ( .A(n4774), .B(n4752), .Z(n4769) );
  NAND U4876 ( .A(n1136), .B(n2362), .Z(n4752) );
  IV U4877 ( .A(n4754), .Z(n4774) );
  XOR U4878 ( .A(n4778), .B(n4779), .Z(n4757) );
  AND U4879 ( .A(n4780), .B(n4781), .Z(n4779) );
  XOR U4880 ( .A(n4782), .B(n4783), .Z(n4781) );
  XOR U4881 ( .A(n4778), .B(n4784), .Z(n4783) );
  XOR U4882 ( .A(n4776), .B(n4785), .Z(n4780) );
  XOR U4883 ( .A(n4778), .B(n4777), .Z(n4785) );
  NANDN U4884 ( .B(n1020), .A(n2734), .Z(n4768) );
  XNOR U4885 ( .A(n4766), .B(n4786), .Z(n4767) );
  AND U4886 ( .A(n2607), .B(n1079), .Z(n4786) );
  XNOR U4887 ( .A(n4771), .B(n4791), .Z(n4772) );
  AND U4888 ( .A(n2362), .B(n1194), .Z(n4791) );
  XOR U4889 ( .A(n4795), .B(n4773), .Z(n4790) );
  NAND U4890 ( .A(n1136), .B(n2483), .Z(n4773) );
  IV U4891 ( .A(n4775), .Z(n4795) );
  XOR U4892 ( .A(n4799), .B(n4800), .Z(n4778) );
  AND U4893 ( .A(n4801), .B(n4802), .Z(n4800) );
  XOR U4894 ( .A(n4803), .B(n4804), .Z(n4802) );
  XOR U4895 ( .A(n4799), .B(n4805), .Z(n4804) );
  XOR U4896 ( .A(n4797), .B(n4806), .Z(n4801) );
  XOR U4897 ( .A(n4799), .B(n4798), .Z(n4806) );
  OR U4898 ( .A(n1020), .B(n2866), .Z(n4789) );
  XNOR U4899 ( .A(n4787), .B(n4807), .Z(n4788) );
  AND U4900 ( .A(n2734), .B(n1079), .Z(n4807) );
  XNOR U4901 ( .A(n4792), .B(n4812), .Z(n4793) );
  AND U4902 ( .A(n2483), .B(n1194), .Z(n4812) );
  XOR U4903 ( .A(n4816), .B(n4794), .Z(n4811) );
  NAND U4904 ( .A(n1136), .B(n2607), .Z(n4794) );
  IV U4905 ( .A(n4796), .Z(n4816) );
  XOR U4906 ( .A(n4820), .B(n4821), .Z(n4799) );
  AND U4907 ( .A(n4822), .B(n4823), .Z(n4821) );
  XOR U4908 ( .A(n4824), .B(n4825), .Z(n4823) );
  XOR U4909 ( .A(n4820), .B(n4826), .Z(n4825) );
  XOR U4910 ( .A(n4818), .B(n4827), .Z(n4822) );
  XOR U4911 ( .A(n4820), .B(n4819), .Z(n4827) );
  OR U4912 ( .A(n1020), .B(n3004), .Z(n4810) );
  XNOR U4913 ( .A(n4808), .B(n4828), .Z(n4809) );
  ANDN U4914 ( .A(n1079), .B(n2866), .Z(n4828) );
  XNOR U4915 ( .A(n4813), .B(n4833), .Z(n4814) );
  AND U4916 ( .A(n2607), .B(n1194), .Z(n4833) );
  XOR U4917 ( .A(n4837), .B(n4815), .Z(n4832) );
  NAND U4918 ( .A(n1136), .B(n2734), .Z(n4815) );
  IV U4919 ( .A(n4817), .Z(n4837) );
  XOR U4920 ( .A(n4841), .B(n4842), .Z(n4820) );
  AND U4921 ( .A(n4843), .B(n4844), .Z(n4842) );
  XOR U4922 ( .A(n4845), .B(n4846), .Z(n4844) );
  XOR U4923 ( .A(n4841), .B(n4847), .Z(n4846) );
  XOR U4924 ( .A(n4839), .B(n4848), .Z(n4843) );
  XOR U4925 ( .A(n4841), .B(n4840), .Z(n4848) );
  NANDN U4926 ( .B(n1020), .A(n3139), .Z(n4831) );
  XNOR U4927 ( .A(n4829), .B(n4849), .Z(n4830) );
  ANDN U4928 ( .A(n1079), .B(n3004), .Z(n4849) );
  XNOR U4929 ( .A(n4834), .B(n4854), .Z(n4835) );
  AND U4930 ( .A(n2734), .B(n1194), .Z(n4854) );
  XOR U4931 ( .A(n4858), .B(n4836), .Z(n4853) );
  NANDN U4932 ( .B(n2866), .A(n1136), .Z(n4836) );
  IV U4933 ( .A(n4838), .Z(n4858) );
  XOR U4934 ( .A(n4863), .B(n4864), .Z(n4709) );
  XNOR U4935 ( .A(n4865), .B(n4862), .Z(n4863) );
  XNOR U4936 ( .A(n4855), .B(n4867), .Z(n4856) );
  ANDN U4937 ( .A(n1194), .B(n2866), .Z(n4867) );
  XOR U4938 ( .A(n4870), .B(n4868), .Z(n4869) );
  ANDN U4939 ( .A(n1194), .B(n3004), .Z(n4870) );
  AND U4940 ( .A(n3139), .B(n1136), .Z(n4871) );
  XOR U4941 ( .A(n4875), .B(n4857), .Z(n4866) );
  NANDN U4942 ( .B(n3004), .A(n1136), .Z(n4857) );
  IV U4943 ( .A(n4859), .Z(n4875) );
  NAND U4944 ( .A(n1136), .B(n3828), .Z(n4874) );
  XNOR U4945 ( .A(n4872), .B(n4876), .Z(n4873) );
  AND U4946 ( .A(n3139), .B(n1194), .Z(n4876) );
  AND U4947 ( .A(n4877), .B(g_input[0]), .Z(n4872) );
  NANDN U4948 ( .B(n1136), .A(n4878), .Z(n4877) );
  NAND U4949 ( .A(n3828), .B(n1194), .Z(n4878) );
  XNOR U4950 ( .A(n4851), .B(n4852), .Z(n4861) );
  NANDN U4951 ( .B(n1020), .A(n3828), .Z(n4852) );
  XNOR U4952 ( .A(n4850), .B(n4881), .Z(n4851) );
  AND U4953 ( .A(n3139), .B(n1079), .Z(n4881) );
  AND U4954 ( .A(n4882), .B(g_input[0]), .Z(n4850) );
  NAND U4955 ( .A(n4883), .B(n1020), .Z(n4882) );
  NAND U4956 ( .A(n3828), .B(n1079), .Z(n4883) );
  XOR U4957 ( .A(n4886), .B(n4887), .Z(n4862) );
  XNOR U4958 ( .A(n3106), .B(n4889), .Z(n3107) );
  AND U4959 ( .A(n1546), .B(n1516), .Z(n4889) );
  XNOR U4960 ( .A(n4520), .B(g_input[16]), .Z(n4519) );
  NOR U4961 ( .A(n4890), .B(n4891), .Z(n4520) );
  XOR U4962 ( .A(n4895), .B(n3108), .Z(n4888) );
  NAND U4963 ( .A(n1428), .B(n1638), .Z(n3108) );
  IV U4964 ( .A(n3110), .Z(n4895) );
  NAND U4965 ( .A(n1280), .B(n1925), .Z(n4714) );
  XNOR U4966 ( .A(n4712), .B(n4897), .Z(n4713) );
  AND U4967 ( .A(n1825), .B(n1348), .Z(n4897) );
  XNOR U4968 ( .A(n4892), .B(n4902), .Z(n4893) );
  AND U4969 ( .A(n1638), .B(n1516), .Z(n4902) );
  XOR U4970 ( .A(n4890), .B(g_input[15]), .Z(n4891) );
  NANDN U4971 ( .B(n4903), .A(n4904), .Z(n4890) );
  XOR U4972 ( .A(n4908), .B(n4894), .Z(n4901) );
  NAND U4973 ( .A(n1428), .B(n1731), .Z(n4894) );
  IV U4974 ( .A(n4896), .Z(n4908) );
  NAND U4975 ( .A(n1280), .B(n2030), .Z(n4900) );
  XNOR U4976 ( .A(n4898), .B(n4910), .Z(n4899) );
  AND U4977 ( .A(n1925), .B(n1348), .Z(n4910) );
  XNOR U4978 ( .A(n4905), .B(n4915), .Z(n4906) );
  AND U4979 ( .A(n1731), .B(n1516), .Z(n4915) );
  XNOR U4980 ( .A(n4904), .B(g_input[14]), .Z(n4903) );
  NOR U4981 ( .A(n4916), .B(n4917), .Z(n4904) );
  XOR U4982 ( .A(n4921), .B(n4907), .Z(n4914) );
  NAND U4983 ( .A(n1428), .B(n1825), .Z(n4907) );
  IV U4984 ( .A(n4909), .Z(n4921) );
  NAND U4985 ( .A(n1280), .B(n2135), .Z(n4913) );
  XNOR U4986 ( .A(n4911), .B(n4923), .Z(n4912) );
  AND U4987 ( .A(n2030), .B(n1348), .Z(n4923) );
  XNOR U4988 ( .A(n4918), .B(n4928), .Z(n4919) );
  AND U4989 ( .A(n1825), .B(n1516), .Z(n4928) );
  XOR U4990 ( .A(n4916), .B(g_input[13]), .Z(n4917) );
  NANDN U4991 ( .B(n4929), .A(n4930), .Z(n4916) );
  XOR U4992 ( .A(n4934), .B(n4920), .Z(n4927) );
  NAND U4993 ( .A(n1428), .B(n1925), .Z(n4920) );
  IV U4994 ( .A(n4922), .Z(n4934) );
  NAND U4995 ( .A(n1280), .B(n2246), .Z(n4926) );
  XNOR U4996 ( .A(n4924), .B(n4936), .Z(n4925) );
  AND U4997 ( .A(n2135), .B(n1348), .Z(n4936) );
  XNOR U4998 ( .A(n4931), .B(n4941), .Z(n4932) );
  AND U4999 ( .A(n1925), .B(n1516), .Z(n4941) );
  XNOR U5000 ( .A(n4930), .B(g_input[12]), .Z(n4929) );
  NOR U5001 ( .A(n4942), .B(n4943), .Z(n4930) );
  XOR U5002 ( .A(n4947), .B(n4933), .Z(n4940) );
  NAND U5003 ( .A(n1428), .B(n2030), .Z(n4933) );
  IV U5004 ( .A(n4935), .Z(n4947) );
  NAND U5005 ( .A(n1280), .B(n2362), .Z(n4939) );
  XNOR U5006 ( .A(n4937), .B(n4949), .Z(n4938) );
  AND U5007 ( .A(n2246), .B(n1348), .Z(n4949) );
  XNOR U5008 ( .A(n4944), .B(n4954), .Z(n4945) );
  AND U5009 ( .A(n2030), .B(n1516), .Z(n4954) );
  XOR U5010 ( .A(n4942), .B(g_input[11]), .Z(n4943) );
  NANDN U5011 ( .B(n4955), .A(n4956), .Z(n4942) );
  XOR U5012 ( .A(n4960), .B(n4946), .Z(n4953) );
  NAND U5013 ( .A(n1428), .B(n2135), .Z(n4946) );
  IV U5014 ( .A(n4948), .Z(n4960) );
  NAND U5015 ( .A(n1280), .B(n2483), .Z(n4952) );
  XNOR U5016 ( .A(n4950), .B(n4962), .Z(n4951) );
  AND U5017 ( .A(n2362), .B(n1348), .Z(n4962) );
  XNOR U5018 ( .A(n4957), .B(n4967), .Z(n4958) );
  AND U5019 ( .A(n2135), .B(n1516), .Z(n4967) );
  XNOR U5020 ( .A(n4956), .B(g_input[10]), .Z(n4955) );
  NOR U5021 ( .A(n4968), .B(n4969), .Z(n4956) );
  XOR U5022 ( .A(n4973), .B(n4959), .Z(n4966) );
  NAND U5023 ( .A(n1428), .B(n2246), .Z(n4959) );
  IV U5024 ( .A(n4961), .Z(n4973) );
  NAND U5025 ( .A(n1280), .B(n2607), .Z(n4965) );
  XNOR U5026 ( .A(n4963), .B(n4975), .Z(n4964) );
  AND U5027 ( .A(n2483), .B(n1348), .Z(n4975) );
  XNOR U5028 ( .A(n4970), .B(n4980), .Z(n4971) );
  AND U5029 ( .A(n2246), .B(n1516), .Z(n4980) );
  XOR U5030 ( .A(n4968), .B(g_input[9]), .Z(n4969) );
  NANDN U5031 ( .B(n4981), .A(n4982), .Z(n4968) );
  XOR U5032 ( .A(n4986), .B(n4972), .Z(n4979) );
  NAND U5033 ( .A(n1428), .B(n2362), .Z(n4972) );
  IV U5034 ( .A(n4974), .Z(n4986) );
  NAND U5035 ( .A(n1280), .B(n2734), .Z(n4978) );
  XNOR U5036 ( .A(n4976), .B(n4988), .Z(n4977) );
  AND U5037 ( .A(n2607), .B(n1348), .Z(n4988) );
  XNOR U5038 ( .A(n4992), .B(n4989), .Z(n4991) );
  XNOR U5039 ( .A(n4983), .B(n4994), .Z(n4984) );
  AND U5040 ( .A(n2362), .B(n1516), .Z(n4994) );
  XNOR U5041 ( .A(n4998), .B(n4995), .Z(n4997) );
  XOR U5042 ( .A(n4999), .B(n4985), .Z(n4993) );
  NAND U5043 ( .A(n1428), .B(n2483), .Z(n4985) );
  IV U5044 ( .A(n4987), .Z(n4999) );
  XNOR U5045 ( .A(n5000), .B(n5001), .Z(n4987) );
  AND U5046 ( .A(n5002), .B(n5003), .Z(n5001) );
  XOR U5047 ( .A(n4996), .B(n5004), .Z(n5003) );
  XNOR U5048 ( .A(n4998), .B(n5000), .Z(n5004) );
  NAND U5049 ( .A(n1428), .B(n2607), .Z(n4998) );
  XOR U5050 ( .A(n4995), .B(n5005), .Z(n4996) );
  AND U5051 ( .A(n2483), .B(n1516), .Z(n5005) );
  XNOR U5052 ( .A(n5009), .B(n5006), .Z(n5008) );
  XOR U5053 ( .A(n4990), .B(n5010), .Z(n5002) );
  XNOR U5054 ( .A(n4992), .B(n5000), .Z(n5010) );
  NANDN U5055 ( .B(n2866), .A(n1280), .Z(n4992) );
  XOR U5056 ( .A(n4989), .B(n5011), .Z(n4990) );
  AND U5057 ( .A(n2734), .B(n1348), .Z(n5011) );
  XNOR U5058 ( .A(n5015), .B(n5012), .Z(n5014) );
  XOR U5059 ( .A(n5016), .B(n5017), .Z(n5000) );
  AND U5060 ( .A(n5018), .B(n5019), .Z(n5017) );
  XOR U5061 ( .A(n5007), .B(n5020), .Z(n5019) );
  XNOR U5062 ( .A(n5009), .B(n5016), .Z(n5020) );
  NAND U5063 ( .A(n1428), .B(n2734), .Z(n5009) );
  XOR U5064 ( .A(n5006), .B(n5021), .Z(n5007) );
  AND U5065 ( .A(n2607), .B(n1516), .Z(n5021) );
  XNOR U5066 ( .A(n5025), .B(n5022), .Z(n5024) );
  XOR U5067 ( .A(n5013), .B(n5026), .Z(n5018) );
  XNOR U5068 ( .A(n5015), .B(n5016), .Z(n5026) );
  NANDN U5069 ( .B(n3004), .A(n1280), .Z(n5015) );
  XOR U5070 ( .A(n5012), .B(n5027), .Z(n5013) );
  ANDN U5071 ( .A(n1348), .B(n2866), .Z(n5027) );
  XNOR U5072 ( .A(n5031), .B(n5028), .Z(n5030) );
  XOR U5073 ( .A(n5032), .B(n5033), .Z(n5016) );
  AND U5074 ( .A(n5034), .B(n5035), .Z(n5033) );
  XOR U5075 ( .A(n5023), .B(n5036), .Z(n5035) );
  XNOR U5076 ( .A(n5025), .B(n5032), .Z(n5036) );
  NANDN U5077 ( .B(n2866), .A(n1428), .Z(n5025) );
  XOR U5078 ( .A(n5022), .B(n5037), .Z(n5023) );
  AND U5079 ( .A(n2734), .B(n1516), .Z(n5037) );
  XOR U5080 ( .A(n5029), .B(n5041), .Z(n5034) );
  XNOR U5081 ( .A(n5031), .B(n5032), .Z(n5041) );
  NAND U5082 ( .A(n1280), .B(n3139), .Z(n5031) );
  XOR U5083 ( .A(n5028), .B(n5042), .Z(n5029) );
  ANDN U5084 ( .A(n1348), .B(n3004), .Z(n5042) );
  NAND U5085 ( .A(n1280), .B(n3828), .Z(n5045) );
  XNOR U5086 ( .A(n5043), .B(n5047), .Z(n5044) );
  AND U5087 ( .A(n3139), .B(n1348), .Z(n5047) );
  AND U5088 ( .A(n5048), .B(g_input[0]), .Z(n5043) );
  NANDN U5089 ( .B(n1280), .A(n5049), .Z(n5048) );
  NAND U5090 ( .A(n3828), .B(n1348), .Z(n5049) );
  XNOR U5091 ( .A(n5038), .B(n5053), .Z(n5039) );
  ANDN U5092 ( .A(n1516), .B(n2866), .Z(n5053) );
  XOR U5093 ( .A(n5056), .B(n5054), .Z(n5055) );
  ANDN U5094 ( .A(n1516), .B(n3004), .Z(n5056) );
  AND U5095 ( .A(n3139), .B(n1428), .Z(n5057) );
  XOR U5096 ( .A(n5061), .B(n5040), .Z(n5052) );
  NANDN U5097 ( .B(n3004), .A(n1428), .Z(n5040) );
  IV U5098 ( .A(n5046), .Z(n5061) );
  NAND U5099 ( .A(n1428), .B(n3828), .Z(n5060) );
  XNOR U5100 ( .A(n5058), .B(n5062), .Z(n5059) );
  AND U5101 ( .A(n3139), .B(n1516), .Z(n5062) );
  AND U5102 ( .A(n5063), .B(g_input[0]), .Z(n5058) );
  NANDN U5103 ( .B(n1428), .A(n5064), .Z(n5063) );
  NAND U5104 ( .A(n3828), .B(n1516), .Z(n5064) );
  XNOR U5105 ( .A(n5067), .B(n3129), .Z(n3119) );
  XNOR U5106 ( .A(n3116), .B(n3117), .Z(n3129) );
  NANDN U5107 ( .B(n835), .A(n2734), .Z(n3117) );
  XNOR U5108 ( .A(n3115), .B(n5068), .Z(n3116) );
  AND U5109 ( .A(n2607), .B(n874), .Z(n5068) );
  XNOR U5110 ( .A(n5072), .B(n5069), .Z(n5071) );
  XNOR U5111 ( .A(n3128), .B(n3118), .Z(n5067) );
  XOR U5112 ( .A(n5073), .B(n5074), .Z(n3118) );
  XNOR U5113 ( .A(n3123), .B(n5076), .Z(n3124) );
  AND U5114 ( .A(n2362), .B(n982), .Z(n5076) );
  XNOR U5115 ( .A(n4982), .B(g_input[8]), .Z(n4981) );
  NOR U5116 ( .A(n5077), .B(n5078), .Z(n4982) );
  XNOR U5117 ( .A(n5082), .B(n5079), .Z(n5081) );
  XOR U5118 ( .A(n5083), .B(n3125), .Z(n5075) );
  NAND U5119 ( .A(n928), .B(n2483), .Z(n3125) );
  IV U5120 ( .A(n3127), .Z(n5083) );
  XNOR U5121 ( .A(n5084), .B(n5085), .Z(n3127) );
  AND U5122 ( .A(n5086), .B(n5087), .Z(n5085) );
  XOR U5123 ( .A(n5080), .B(n5088), .Z(n5087) );
  XNOR U5124 ( .A(n5082), .B(n5084), .Z(n5088) );
  NAND U5125 ( .A(n928), .B(n2607), .Z(n5082) );
  XOR U5126 ( .A(n5079), .B(n5089), .Z(n5080) );
  AND U5127 ( .A(n2483), .B(n982), .Z(n5089) );
  XOR U5128 ( .A(n5077), .B(g_input[7]), .Z(n5078) );
  NANDN U5129 ( .B(n5090), .A(n5091), .Z(n5077) );
  XNOR U5130 ( .A(n5095), .B(n5092), .Z(n5094) );
  XOR U5131 ( .A(n5070), .B(n5096), .Z(n5086) );
  XNOR U5132 ( .A(n5072), .B(n5084), .Z(n5096) );
  OR U5133 ( .A(n835), .B(n2866), .Z(n5072) );
  XOR U5134 ( .A(n5069), .B(n5097), .Z(n5070) );
  AND U5135 ( .A(n2734), .B(n874), .Z(n5097) );
  XNOR U5136 ( .A(n5101), .B(n5098), .Z(n5100) );
  XOR U5137 ( .A(n5102), .B(n5103), .Z(n5084) );
  AND U5138 ( .A(n5104), .B(n5105), .Z(n5103) );
  XOR U5139 ( .A(n5093), .B(n5106), .Z(n5105) );
  XNOR U5140 ( .A(n5095), .B(n5102), .Z(n5106) );
  NAND U5141 ( .A(n928), .B(n2734), .Z(n5095) );
  XOR U5142 ( .A(n5092), .B(n5107), .Z(n5093) );
  AND U5143 ( .A(n2607), .B(n982), .Z(n5107) );
  XNOR U5144 ( .A(n5091), .B(g_input[6]), .Z(n5090) );
  NOR U5145 ( .A(n5108), .B(n5109), .Z(n5091) );
  XNOR U5146 ( .A(n5113), .B(n5110), .Z(n5112) );
  XOR U5147 ( .A(n5099), .B(n5114), .Z(n5104) );
  XNOR U5148 ( .A(n5101), .B(n5102), .Z(n5114) );
  OR U5149 ( .A(n835), .B(n3004), .Z(n5101) );
  XOR U5150 ( .A(n5098), .B(n5115), .Z(n5099) );
  ANDN U5151 ( .A(n874), .B(n2866), .Z(n5115) );
  XNOR U5152 ( .A(n5119), .B(n5116), .Z(n5118) );
  XOR U5153 ( .A(n5120), .B(n5121), .Z(n5102) );
  AND U5154 ( .A(n5122), .B(n5123), .Z(n5121) );
  XOR U5155 ( .A(n5111), .B(n5124), .Z(n5123) );
  XNOR U5156 ( .A(n5113), .B(n5120), .Z(n5124) );
  NANDN U5157 ( .B(n2866), .A(n928), .Z(n5113) );
  XOR U5158 ( .A(n5110), .B(n5125), .Z(n5111) );
  AND U5159 ( .A(n2734), .B(n982), .Z(n5125) );
  XOR U5160 ( .A(n5108), .B(g_input[5]), .Z(n5109) );
  NANDN U5161 ( .B(n5126), .A(n5127), .Z(n5108) );
  XOR U5162 ( .A(n5117), .B(n5131), .Z(n5122) );
  XNOR U5163 ( .A(n5119), .B(n5120), .Z(n5131) );
  NANDN U5164 ( .B(n835), .A(n3139), .Z(n5119) );
  XOR U5165 ( .A(n5116), .B(n5132), .Z(n5117) );
  ANDN U5166 ( .A(n874), .B(n3004), .Z(n5132) );
  NANDN U5167 ( .B(n835), .A(n3828), .Z(n5135) );
  XNOR U5168 ( .A(n5133), .B(n5137), .Z(n5134) );
  AND U5169 ( .A(n3139), .B(n874), .Z(n5137) );
  AND U5170 ( .A(n5138), .B(g_input[0]), .Z(n5133) );
  NAND U5171 ( .A(n5139), .B(n835), .Z(n5138) );
  NAND U5172 ( .A(n3828), .B(n874), .Z(n5139) );
  XNOR U5173 ( .A(n5128), .B(n5143), .Z(n5129) );
  ANDN U5174 ( .A(n982), .B(n2866), .Z(n5143) );
  XOR U5175 ( .A(n5146), .B(n5144), .Z(n5145) );
  ANDN U5176 ( .A(n982), .B(n3004), .Z(n5146) );
  AND U5177 ( .A(n3139), .B(n928), .Z(n5147) );
  XOR U5178 ( .A(n5151), .B(n5130), .Z(n5142) );
  NANDN U5179 ( .B(n3004), .A(n928), .Z(n5130) );
  IV U5180 ( .A(n5136), .Z(n5151) );
  NAND U5181 ( .A(n928), .B(n3828), .Z(n5150) );
  XNOR U5182 ( .A(n5148), .B(n5152), .Z(n5149) );
  AND U5183 ( .A(n3139), .B(n982), .Z(n5152) );
  AND U5184 ( .A(n5153), .B(g_input[0]), .Z(n5148) );
  NANDN U5185 ( .B(n928), .A(n5154), .Z(n5153) );
  NAND U5186 ( .A(n3828), .B(n982), .Z(n5154) );
  XNOR U5187 ( .A(n3132), .B(n5158), .Z(n3133) );
  ANDN U5188 ( .A(n806), .B(n2866), .Z(n5158) );
  XNOR U5189 ( .A(n5127), .B(g_input[4]), .Z(n5126) );
  NOR U5190 ( .A(n5159), .B(n5160), .Z(n5127) );
  XOR U5191 ( .A(n5163), .B(n5161), .Z(n5162) );
  ANDN U5192 ( .A(n806), .B(n3004), .Z(n5163) );
  AND U5193 ( .A(n3139), .B(n770), .Z(n5164) );
  XOR U5194 ( .A(n5168), .B(n3134), .Z(n5157) );
  NANDN U5195 ( .B(n3004), .A(n770), .Z(n3134) );
  NANDN U5196 ( .B(n5169), .A(n5170), .Z(n5159) );
  IV U5197 ( .A(n3136), .Z(n5168) );
  NAND U5198 ( .A(n770), .B(n3828), .Z(n5167) );
  XNOR U5199 ( .A(n5165), .B(n5171), .Z(n5166) );
  AND U5200 ( .A(n3139), .B(n806), .Z(n5171) );
  AND U5201 ( .A(n5172), .B(g_input[0]), .Z(n5165) );
  NANDN U5202 ( .B(n770), .A(n5173), .Z(n5172) );
  NAND U5203 ( .A(n3828), .B(n806), .Z(n5173) );
  XNOR U5204 ( .A(n3143), .B(n3144), .Z(n3138) );
  NANDN U5205 ( .B(n709), .A(n3828), .Z(n3144) );
  XNOR U5206 ( .A(n3142), .B(n5176), .Z(n3143) );
  AND U5207 ( .A(n3139), .B(n742), .Z(n5176) );
  XNOR U5208 ( .A(n5170), .B(g_input[2]), .Z(n5169) );
  AND U5209 ( .A(n5178), .B(g_input[0]), .Z(n3142) );
  NAND U5210 ( .A(n5179), .B(n709), .Z(n5178) );
  NANDN U5211 ( .B(n5180), .A(n5181), .Z(n709) );
  ANDN U5212 ( .A(e_input[31]), .B(n5182), .Z(n5181) );
  NAND U5213 ( .A(n3828), .B(n742), .Z(n5179) );
  XOR U5214 ( .A(n5182), .B(e_input[30]), .Z(n5180) );
  OR U5215 ( .A(n5175), .B(n5183), .Z(n5182) );
  XOR U5216 ( .A(n5183), .B(e_input[29]), .Z(n5175) );
  OR U5217 ( .A(n5174), .B(n5184), .Z(n5183) );
  XOR U5218 ( .A(n5184), .B(e_input[28]), .Z(n5174) );
  OR U5219 ( .A(n5140), .B(n5185), .Z(n5184) );
  XOR U5220 ( .A(n5185), .B(e_input[27]), .Z(n5140) );
  OR U5221 ( .A(n5141), .B(n5186), .Z(n5185) );
  XOR U5222 ( .A(n5186), .B(e_input[26]), .Z(n5141) );
  OR U5223 ( .A(n5156), .B(n5187), .Z(n5186) );
  XOR U5224 ( .A(n5187), .B(e_input[25]), .Z(n5156) );
  OR U5225 ( .A(n5155), .B(n5188), .Z(n5187) );
  XOR U5226 ( .A(n5188), .B(e_input[24]), .Z(n5155) );
  OR U5227 ( .A(n4884), .B(n5189), .Z(n5188) );
  XOR U5228 ( .A(n5189), .B(e_input[23]), .Z(n4884) );
  OR U5229 ( .A(n4885), .B(n5190), .Z(n5189) );
  XOR U5230 ( .A(n5190), .B(e_input[22]), .Z(n4885) );
  OR U5231 ( .A(n4880), .B(n5191), .Z(n5190) );
  XOR U5232 ( .A(n5191), .B(e_input[21]), .Z(n4880) );
  OR U5233 ( .A(n4879), .B(n5192), .Z(n5191) );
  XOR U5234 ( .A(n5192), .B(e_input[20]), .Z(n4879) );
  OR U5235 ( .A(n5051), .B(n5193), .Z(n5192) );
  XOR U5236 ( .A(n5193), .B(e_input[19]), .Z(n5051) );
  OR U5237 ( .A(n5050), .B(n5194), .Z(n5193) );
  XOR U5238 ( .A(n5194), .B(e_input[18]), .Z(n5050) );
  OR U5239 ( .A(n5066), .B(n5195), .Z(n5194) );
  XOR U5240 ( .A(n5195), .B(e_input[17]), .Z(n5066) );
  OR U5241 ( .A(n5065), .B(n5196), .Z(n5195) );
  XOR U5242 ( .A(n5196), .B(e_input[16]), .Z(n5065) );
  OR U5243 ( .A(n3868), .B(n5197), .Z(n5196) );
  XOR U5244 ( .A(n5197), .B(e_input[15]), .Z(n3868) );
  OR U5245 ( .A(n3867), .B(n5198), .Z(n5197) );
  XOR U5246 ( .A(n5198), .B(e_input[14]), .Z(n3867) );
  OR U5247 ( .A(n3863), .B(n5199), .Z(n5198) );
  XOR U5248 ( .A(n5199), .B(e_input[13]), .Z(n3863) );
  OR U5249 ( .A(n3862), .B(n5200), .Z(n5199) );
  XOR U5250 ( .A(n5200), .B(e_input[12]), .Z(n3862) );
  OR U5251 ( .A(n3833), .B(n5201), .Z(n5200) );
  XOR U5252 ( .A(n5201), .B(e_input[11]), .Z(n3833) );
  OR U5253 ( .A(n3832), .B(n5202), .Z(n5201) );
  XOR U5254 ( .A(n5202), .B(e_input[10]), .Z(n3832) );
  OR U5255 ( .A(n3848), .B(n5203), .Z(n5202) );
  XOR U5256 ( .A(n5203), .B(e_input[9]), .Z(n3848) );
  OR U5257 ( .A(n3847), .B(n5204), .Z(n5203) );
  XOR U5258 ( .A(n5204), .B(e_input[8]), .Z(n3847) );
  OR U5259 ( .A(n4318), .B(n5205), .Z(n5204) );
  XOR U5260 ( .A(n5205), .B(e_input[7]), .Z(n4318) );
  OR U5261 ( .A(n4317), .B(n5206), .Z(n5205) );
  XOR U5262 ( .A(n5206), .B(e_input[6]), .Z(n4317) );
  OR U5263 ( .A(n4313), .B(n5207), .Z(n5206) );
  XOR U5264 ( .A(n5207), .B(e_input[5]), .Z(n4313) );
  OR U5265 ( .A(n4312), .B(n5208), .Z(n5207) );
  XOR U5266 ( .A(n5208), .B(e_input[4]), .Z(n4312) );
  OR U5267 ( .A(n4679), .B(n5209), .Z(n5208) );
  XOR U5268 ( .A(n5209), .B(e_input[3]), .Z(n4679) );
  OR U5269 ( .A(n4678), .B(n5210), .Z(n5209) );
  XOR U5270 ( .A(n5210), .B(e_input[2]), .Z(n4678) );
  NANDN U5271 ( .B(e_input[0]), .A(n4693), .Z(n5210) );
  XNOR U5272 ( .A(e_input[0]), .B(e_input[1]), .Z(n4693) );
  XOR U5273 ( .A(g_input[0]), .B(g_input[1]), .Z(n5177) );
  AND U5274 ( .A(n5211), .B(n5212), .Z(\_MxM/N17 ) );
  XOR U5275 ( .A(\_MxM/n[6] ), .B(\_MxM/add_43/carry[6] ), .Z(n5212) );
  AND U5276 ( .A(\_MxM/N9 ), .B(n5211), .Z(\_MxM/N16 ) );
  AND U5277 ( .A(\_MxM/N8 ), .B(n5211), .Z(\_MxM/N15 ) );
  AND U5278 ( .A(\_MxM/N7 ), .B(n5211), .Z(\_MxM/N14 ) );
  AND U5279 ( .A(\_MxM/N6 ), .B(n5211), .Z(\_MxM/N13 ) );
  AND U5280 ( .A(\_MxM/N5 ), .B(n5211), .Z(\_MxM/N12 ) );
  NAND U5281 ( .A(n5213), .B(n5214), .Z(n5211) );
  ANDN U5282 ( .A(n5215), .B(n650), .Z(n5214) );
  OR U5283 ( .A(\_MxM/n[4] ), .B(\_MxM/n[3] ), .Z(n650) );
  NOR U5284 ( .A(\_MxM/N11 ), .B(\_MxM/n[2] ), .Z(n5215) );
  AND U5285 ( .A(\_MxM/n[6] ), .B(n5216), .Z(n5213) );
  AND U5286 ( .A(\_MxM/n[5] ), .B(\_MxM/n[1] ), .Z(n5216) );
  IV U5287 ( .A(\_MxM/n[0] ), .Z(\_MxM/N11 ) );
endmodule

