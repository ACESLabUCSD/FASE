
module MxM_W32_N1000 ( clk, rst, A, X, Y );
  input [31:0] A;
  input [31:0] X;
  output [31:0] Y;
  input clk, rst;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, \add_25/carry[9] , \add_25/carry[8] ,
         \add_25/carry[7] , \add_25/carry[6] , \add_25/carry[5] ,
         \add_25/carry[4] , \add_25/carry[3] , \add_25/carry[2] , n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649;
  wire   [31:0] Y0;
  wire   [9:0] n;

  DFF \n_reg[0]  ( .D(n372), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[0]) );
  DFF \n_reg[1]  ( .D(n371), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[1]) );
  DFF \n_reg[2]  ( .D(n370), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[2]) );
  DFF \n_reg[3]  ( .D(n369), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[3]) );
  DFF \n_reg[4]  ( .D(n368), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[4]) );
  DFF \n_reg[5]  ( .D(n367), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[5]) );
  DFF \n_reg[6]  ( .D(n366), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[6]) );
  DFF \n_reg[7]  ( .D(n365), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[7]) );
  DFF \n_reg[8]  ( .D(n364), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[8]) );
  DFF \n_reg[9]  ( .D(n363), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(n[9]) );
  DFF \Y0_reg[0]  ( .D(n362), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[0]) );
  DFF \Y0_reg[1]  ( .D(n361), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[1]) );
  DFF \Y0_reg[2]  ( .D(n360), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[2]) );
  DFF \Y0_reg[3]  ( .D(n359), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[3]) );
  DFF \Y0_reg[4]  ( .D(n358), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[4]) );
  DFF \Y0_reg[5]  ( .D(n357), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[5]) );
  DFF \Y0_reg[6]  ( .D(n356), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[6]) );
  DFF \Y0_reg[7]  ( .D(n355), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[7]) );
  DFF \Y0_reg[8]  ( .D(n354), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[8]) );
  DFF \Y0_reg[9]  ( .D(n353), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[9]) );
  DFF \Y0_reg[10]  ( .D(n352), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[10]) );
  DFF \Y0_reg[11]  ( .D(n351), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[11]) );
  DFF \Y0_reg[12]  ( .D(n350), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[12]) );
  DFF \Y0_reg[13]  ( .D(n349), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[13]) );
  DFF \Y0_reg[14]  ( .D(n348), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[14]) );
  DFF \Y0_reg[15]  ( .D(n347), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[15]) );
  DFF \Y0_reg[16]  ( .D(n346), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[16]) );
  DFF \Y0_reg[17]  ( .D(n345), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[17]) );
  DFF \Y0_reg[18]  ( .D(n344), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[18]) );
  DFF \Y0_reg[19]  ( .D(n343), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[19]) );
  DFF \Y0_reg[20]  ( .D(n342), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[20]) );
  DFF \Y0_reg[21]  ( .D(n341), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[21]) );
  DFF \Y0_reg[22]  ( .D(n340), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[22]) );
  DFF \Y0_reg[23]  ( .D(n339), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[23]) );
  DFF \Y0_reg[24]  ( .D(n338), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[24]) );
  DFF \Y0_reg[25]  ( .D(n337), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[25]) );
  DFF \Y0_reg[26]  ( .D(n336), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[26]) );
  DFF \Y0_reg[27]  ( .D(n335), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[27]) );
  DFF \Y0_reg[28]  ( .D(n334), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[28]) );
  DFF \Y0_reg[29]  ( .D(n333), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[29]) );
  DFF \Y0_reg[30]  ( .D(n332), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[30]) );
  DFF \Y0_reg[31]  ( .D(n331), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y0[31]) );
  DFF \Y_reg[31]  ( .D(n330), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[31]) );
  DFF \Y_reg[30]  ( .D(n329), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[30]) );
  DFF \Y_reg[29]  ( .D(n328), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[29]) );
  DFF \Y_reg[28]  ( .D(n327), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[28]) );
  DFF \Y_reg[27]  ( .D(n326), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[27]) );
  DFF \Y_reg[26]  ( .D(n325), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[26]) );
  DFF \Y_reg[25]  ( .D(n324), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[25]) );
  DFF \Y_reg[24]  ( .D(n323), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[24]) );
  DFF \Y_reg[23]  ( .D(n322), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[23]) );
  DFF \Y_reg[22]  ( .D(n321), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[22]) );
  DFF \Y_reg[21]  ( .D(n320), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[21]) );
  DFF \Y_reg[20]  ( .D(n319), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[20]) );
  DFF \Y_reg[19]  ( .D(n318), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[19]) );
  DFF \Y_reg[18]  ( .D(n317), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[18]) );
  DFF \Y_reg[17]  ( .D(n316), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[17]) );
  DFF \Y_reg[16]  ( .D(n315), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[16]) );
  DFF \Y_reg[15]  ( .D(n314), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[15]) );
  DFF \Y_reg[14]  ( .D(n313), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[14]) );
  DFF \Y_reg[13]  ( .D(n312), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[13]) );
  DFF \Y_reg[12]  ( .D(n311), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[12]) );
  DFF \Y_reg[11]  ( .D(n310), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[11]) );
  DFF \Y_reg[10]  ( .D(n309), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[10]) );
  DFF \Y_reg[9]  ( .D(n308), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[9]) );
  DFF \Y_reg[8]  ( .D(n307), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[8]) );
  DFF \Y_reg[7]  ( .D(n306), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[7]) );
  DFF \Y_reg[6]  ( .D(n305), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[6]) );
  DFF \Y_reg[5]  ( .D(n304), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[5]) );
  DFF \Y_reg[4]  ( .D(n303), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[4]) );
  DFF \Y_reg[3]  ( .D(n302), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[3]) );
  DFF \Y_reg[2]  ( .D(n301), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[2]) );
  DFF \Y_reg[1]  ( .D(n300), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[1]) );
  DFF \Y_reg[0]  ( .D(n299), .CLK(clk), .RST(1'b0), .I(1'b0), .Q(Y[0]) );
  HADDER \add_25/U1_1_1  ( .IN0(n[1]), .IN1(n[0]), .COUT(\add_25/carry[2] ), 
        .SUM(N8) );
  HADDER \add_25/U1_1_2  ( .IN0(n[2]), .IN1(\add_25/carry[2] ), .COUT(
        \add_25/carry[3] ), .SUM(N9) );
  HADDER \add_25/U1_1_3  ( .IN0(n[3]), .IN1(\add_25/carry[3] ), .COUT(
        \add_25/carry[4] ), .SUM(N10) );
  HADDER \add_25/U1_1_4  ( .IN0(n[4]), .IN1(\add_25/carry[4] ), .COUT(
        \add_25/carry[5] ), .SUM(N11) );
  HADDER \add_25/U1_1_5  ( .IN0(n[5]), .IN1(\add_25/carry[5] ), .COUT(
        \add_25/carry[6] ), .SUM(N12) );
  HADDER \add_25/U1_1_6  ( .IN0(n[6]), .IN1(\add_25/carry[6] ), .COUT(
        \add_25/carry[7] ), .SUM(N13) );
  HADDER \add_25/U1_1_7  ( .IN0(n[7]), .IN1(\add_25/carry[7] ), .COUT(
        \add_25/carry[8] ), .SUM(N14) );
  HADDER \add_25/U1_1_8  ( .IN0(n[8]), .IN1(\add_25/carry[8] ), .COUT(
        \add_25/carry[9] ), .SUM(N15) );
  MUX U375 ( .IN0(n4080), .IN1(n373), .SEL(n4081), .F(n4034) );
  IV U376 ( .A(n4082), .Z(n373) );
  MUX U377 ( .IN0(n3908), .IN1(n3910), .SEL(n3909), .F(n3862) );
  MUX U378 ( .IN0(n4681), .IN1(n4683), .SEL(n4682), .F(n4657) );
  MUX U379 ( .IN0(n3733), .IN1(n3735), .SEL(n3734), .F(n3687) );
  XNOR U380 ( .A(n4669), .B(n4668), .Z(n4684) );
  XNOR U381 ( .A(n5052), .B(n5050), .Z(n5057) );
  MUX U382 ( .IN0(n3637), .IN1(n3639), .SEL(n3638), .F(n3594) );
  MUX U383 ( .IN0(n5385), .IN1(n5387), .SEL(n5386), .F(n5373) );
  MUX U384 ( .IN0(n5243), .IN1(n374), .SEL(n5244), .F(n5223) );
  IV U385 ( .A(n5245), .Z(n374) );
  MUX U386 ( .IN0(n5392), .IN1(n375), .SEL(n5393), .F(n5380) );
  IV U387 ( .A(n5394), .Z(n375) );
  MUX U388 ( .IN0(n4602), .IN1(n376), .SEL(n4603), .F(n4582) );
  IV U389 ( .A(n4604), .Z(n376) );
  XNOR U390 ( .A(n3590), .B(n3589), .Z(n3626) );
  MUX U391 ( .IN0(n5007), .IN1(n377), .SEL(n5008), .F(n4997) );
  IV U392 ( .A(n5009), .Z(n377) );
  XNOR U393 ( .A(n3615), .B(n3613), .Z(n3650) );
  XNOR U394 ( .A(n4778), .B(n4776), .Z(n4785) );
  NANDN U395 ( .B(n1666), .A(n3391), .Z(n390) );
  MUX U396 ( .IN0(n3467), .IN1(n3469), .SEL(n3468), .F(n3428) );
  MUX U397 ( .IN0(n3460), .IN1(n378), .SEL(n3461), .F(n3421) );
  IV U398 ( .A(n3462), .Z(n378) );
  MUX U399 ( .IN0(n3472), .IN1(n3474), .SEL(n3473), .F(n3401) );
  MUX U400 ( .IN0(n1377), .IN1(n379), .SEL(n1378), .F(n1308) );
  IV U401 ( .A(n1379), .Z(n379) );
  MUX U402 ( .IN0(n1674), .IN1(n1676), .SEL(n1675), .F(n1590) );
  MUX U403 ( .IN0(n1729), .IN1(n380), .SEL(n1730), .F(n1638) );
  IV U404 ( .A(n1731), .Z(n380) );
  MUX U405 ( .IN0(n1777), .IN1(n381), .SEL(n1778), .F(n1682) );
  IV U406 ( .A(n1779), .Z(n381) );
  MUX U407 ( .IN0(n1882), .IN1(n382), .SEL(n1883), .F(n1785) );
  IV U408 ( .A(n1884), .Z(n382) );
  MUX U409 ( .IN0(n2141), .IN1(n2143), .SEL(n2142), .F(n2040) );
  MUX U410 ( .IN0(n2257), .IN1(n383), .SEL(n2258), .F(n2149) );
  IV U411 ( .A(n2259), .Z(n383) );
  MUX U412 ( .IN0(n2430), .IN1(n384), .SEL(n2431), .F(n2321) );
  IV U413 ( .A(n2432), .Z(n384) );
  MUX U414 ( .IN0(A[29]), .IN1(n4754), .SEL(A[31]), .F(n385) );
  IV U415 ( .A(n385), .Z(n1001) );
  MUX U416 ( .IN0(n386), .IN1(n4742), .SEL(A[31]), .F(n957) );
  IV U417 ( .A(A[30]), .Z(n386) );
  MUX U418 ( .IN0(n5304), .IN1(n5306), .SEL(n5305), .F(n5280) );
  MUX U419 ( .IN0(n5054), .IN1(n5056), .SEL(n5055), .F(n5039) );
  XNOR U420 ( .A(n5426), .B(n5424), .Z(n5431) );
  MUX U421 ( .IN0(n4637), .IN1(n4639), .SEL(n4638), .F(n4617) );
  MUX U422 ( .IN0(n4642), .IN1(n387), .SEL(n4643), .F(n4622) );
  IV U423 ( .A(n4644), .Z(n387) );
  XNOR U424 ( .A(n5292), .B(n5291), .Z(n5307) );
  MUX U425 ( .IN0(n5373), .IN1(n5375), .SEL(n5374), .F(n5361) );
  MUX U426 ( .IN0(n5223), .IN1(n388), .SEL(n5224), .F(n5203) );
  IV U427 ( .A(n5225), .Z(n388) );
  MUX U428 ( .IN0(n5380), .IN1(n389), .SEL(n5381), .F(n5368) );
  IV U429 ( .A(n5382), .Z(n389) );
  MUX U430 ( .IN0(n3552), .IN1(n3554), .SEL(n3553), .F(n3507) );
  XNOR U431 ( .A(n5010), .B(n5009), .Z(n5015) );
  MUX U432 ( .IN0(n5002), .IN1(n5004), .SEL(n5003), .F(n4992) );
  MUX U433 ( .IN0(n5497), .IN1(n390), .SEL(n5498), .F(n5486) );
  XNOR U434 ( .A(n3503), .B(n3502), .Z(n3541) );
  MUX U435 ( .IN0(n4987), .IN1(n391), .SEL(n4988), .F(n4974) );
  IV U436 ( .A(n4989), .Z(n391) );
  MUX U437 ( .IN0(n3421), .IN1(n392), .SEL(n3422), .F(n3291) );
  IV U438 ( .A(n3423), .Z(n392) );
  MUX U439 ( .IN0(n1529), .IN1(n393), .SEL(n1530), .F(n1449) );
  IV U440 ( .A(n1531), .Z(n393) );
  MUX U441 ( .IN0(n1590), .IN1(n1592), .SEL(n1591), .F(n1509) );
  MUX U442 ( .IN0(n1647), .IN1(n1649), .SEL(n1648), .F(n1565) );
  MUX U443 ( .IN0(n1962), .IN1(n1964), .SEL(n1963), .F(n1866) );
  MUX U444 ( .IN0(n1970), .IN1(n394), .SEL(n1971), .F(n1874) );
  IV U445 ( .A(n1972), .Z(n394) );
  MUX U446 ( .IN0(n1978), .IN1(n395), .SEL(n1979), .F(n1882) );
  IV U447 ( .A(n1980), .Z(n395) );
  MUX U448 ( .IN0(n2025), .IN1(n396), .SEL(n2026), .F(n1925) );
  IV U449 ( .A(n2027), .Z(n396) );
  MUX U450 ( .IN0(n2222), .IN1(n2224), .SEL(n2223), .F(n2114) );
  MUX U451 ( .IN0(n2364), .IN1(n397), .SEL(n2365), .F(n2257) );
  IV U452 ( .A(n2366), .Z(n397) );
  MUX U453 ( .IN0(n2544), .IN1(n398), .SEL(n2545), .F(n2430) );
  IV U454 ( .A(n2546), .Z(n398) );
  MUX U455 ( .IN0(n3170), .IN1(n399), .SEL(n3171), .F(n3045) );
  IV U456 ( .A(n3172), .Z(n399) );
  MUX U457 ( .IN0(n1077), .IN1(n400), .SEL(n1078), .F(n1031) );
  IV U458 ( .A(n1079), .Z(n400) );
  MUX U459 ( .IN0(n3324), .IN1(n3326), .SEL(n3325), .F(n3186) );
  MUX U460 ( .IN0(n401), .IN1(n1112), .SEL(n1111), .F(n1074) );
  IV U461 ( .A(n1110), .Z(n401) );
  MUX U462 ( .IN0(n4088), .IN1(n4090), .SEL(n4089), .F(n4044) );
  MUX U463 ( .IN0(n5066), .IN1(n5068), .SEL(n5067), .F(n5054) );
  XNOR U464 ( .A(n5064), .B(n5063), .Z(n5069) );
  MUX U465 ( .IN0(n5258), .IN1(n5260), .SEL(n5259), .F(n5238) );
  MUX U466 ( .IN0(n5406), .IN1(n402), .SEL(n5407), .F(n5392) );
  IV U467 ( .A(n5408), .Z(n402) );
  MUX U468 ( .IN0(n4617), .IN1(n4619), .SEL(n4618), .F(n4597) );
  MUX U469 ( .IN0(n4622), .IN1(n403), .SEL(n4623), .F(n4602) );
  IV U470 ( .A(n4624), .Z(n403) );
  MUX U471 ( .IN0(n3601), .IN1(n3603), .SEL(n3602), .F(n3557) );
  XNOR U472 ( .A(n5226), .B(n5225), .Z(n5241) );
  MUX U473 ( .IN0(n5361), .IN1(n5363), .SEL(n5362), .F(n5349) );
  XNOR U474 ( .A(n5371), .B(n5370), .Z(n5376) );
  NANDN U475 ( .B(n2422), .A(n3391), .Z(n416) );
  MUX U476 ( .IN0(n4997), .IN1(n404), .SEL(n4998), .F(n4987) );
  IV U477 ( .A(n4999), .Z(n404) );
  MUX U478 ( .IN0(n4992), .IN1(n4994), .SEL(n4993), .F(n4982) );
  XNOR U479 ( .A(n3463), .B(n3462), .Z(n3496) );
  MUX U480 ( .IN0(n1769), .IN1(n1771), .SEL(n1770), .F(n1674) );
  MUX U481 ( .IN0(n2066), .IN1(n405), .SEL(n2067), .F(n1970) );
  IV U482 ( .A(n2068), .Z(n405) );
  MUX U483 ( .IN0(n2074), .IN1(n406), .SEL(n2075), .F(n1978) );
  IV U484 ( .A(n2076), .Z(n406) );
  MUX U485 ( .IN0(n2032), .IN1(n2034), .SEL(n2033), .F(n1934) );
  MUX U486 ( .IN0(n2040), .IN1(n2042), .SEL(n2041), .F(n1942) );
  MUX U487 ( .IN0(n2126), .IN1(n407), .SEL(n2127), .F(n2025) );
  IV U488 ( .A(n2128), .Z(n407) );
  MUX U489 ( .IN0(n2159), .IN1(n2161), .SEL(n2160), .F(n2058) );
  MUX U490 ( .IN0(n2330), .IN1(n2332), .SEL(n2331), .F(n2222) );
  MUX U491 ( .IN0(n2472), .IN1(n408), .SEL(n2473), .F(n2364) );
  IV U492 ( .A(n2474), .Z(n408) );
  MUX U493 ( .IN0(n2640), .IN1(n2642), .SEL(n2641), .F(n2521) );
  MUX U494 ( .IN0(n2778), .IN1(n409), .SEL(n2779), .F(n2658) );
  IV U495 ( .A(n2780), .Z(n409) );
  MUX U496 ( .IN0(n3307), .IN1(n410), .SEL(n3308), .F(n3170) );
  IV U497 ( .A(n3309), .Z(n410) );
  MUX U498 ( .IN0(n1103), .IN1(n1105), .SEL(n1104), .F(n1061) );
  MUX U499 ( .IN0(n993), .IN1(n411), .SEL(n994), .F(n947) );
  IV U500 ( .A(n995), .Z(n411) );
  MUX U501 ( .IN0(n412), .IN1(n1339), .SEL(n1338), .F(n1274) );
  IV U502 ( .A(n1337), .Z(n412) );
  MUX U503 ( .IN0(n5428), .IN1(n5430), .SEL(n5429), .F(n5411) );
  MUX U504 ( .IN0(n5309), .IN1(n413), .SEL(n5310), .F(n5287) );
  IV U505 ( .A(n5311), .Z(n413) );
  MUX U506 ( .IN0(n5127), .IN1(n5129), .SEL(n5128), .F(n5111) );
  MUX U507 ( .IN0(n5238), .IN1(n5240), .SEL(n5239), .F(n5218) );
  MUX U508 ( .IN0(n5012), .IN1(n5014), .SEL(n5013), .F(n5002) );
  XNOR U509 ( .A(n4794), .B(n4793), .Z(n4801) );
  MUX U510 ( .IN0(n4577), .IN1(n4579), .SEL(n4578), .F(n4557) );
  XNOR U511 ( .A(n4605), .B(n4604), .Z(n4620) );
  MUX U512 ( .IN0(n5203), .IN1(n414), .SEL(n5204), .F(n5183) );
  IV U513 ( .A(n5205), .Z(n414) );
  MUX U514 ( .IN0(n5368), .IN1(n415), .SEL(n5369), .F(n5356) );
  IV U515 ( .A(n5370), .Z(n415) );
  MUX U516 ( .IN0(n4173), .IN1(n416), .SEL(n4174), .F(n4162) );
  MUX U517 ( .IN0(n5349), .IN1(n5351), .SEL(n5350), .F(n5166) );
  MUX U518 ( .IN0(n4538), .IN1(n417), .SEL(n4539), .F(n4517) );
  IV U519 ( .A(n4540), .Z(n417) );
  XNOR U520 ( .A(n4990), .B(n4989), .Z(n4995) );
  MUX U521 ( .IN0(n3428), .IN1(n3430), .SEL(n3429), .F(n3298) );
  MUX U522 ( .IN0(n1838), .IN1(n1840), .SEL(n1839), .F(n1736) );
  MUX U523 ( .IN0(n1874), .IN1(n418), .SEL(n1875), .F(n1777) );
  IV U524 ( .A(n1876), .Z(n418) );
  MUX U525 ( .IN0(n1866), .IN1(n1868), .SEL(n1867), .F(n1769) );
  MUX U526 ( .IN0(n2175), .IN1(n419), .SEL(n2176), .F(n2074) );
  IV U527 ( .A(n2177), .Z(n419) );
  MUX U528 ( .IN0(n2348), .IN1(n2350), .SEL(n2349), .F(n2241) );
  MUX U529 ( .IN0(n2341), .IN1(n420), .SEL(n2342), .F(n2234) );
  IV U530 ( .A(n2343), .Z(n420) );
  MUX U531 ( .IN0(n2380), .IN1(n421), .SEL(n2381), .F(n2273) );
  IV U532 ( .A(n2382), .Z(n421) );
  MUX U533 ( .IN0(n2437), .IN1(n2439), .SEL(n2438), .F(n2330) );
  MUX U534 ( .IN0(n2591), .IN1(n422), .SEL(n2592), .F(n2472) );
  IV U535 ( .A(n2593), .Z(n422) );
  MUX U536 ( .IN0(n3008), .IN1(n3010), .SEL(n3009), .F(n2884) );
  MUX U537 ( .IN0(n3016), .IN1(n423), .SEL(n3017), .F(n2892) );
  IV U538 ( .A(n3018), .Z(n423) );
  MUX U539 ( .IN0(A[28]), .IN1(n4771), .SEL(A[31]), .F(n424) );
  IV U540 ( .A(n424), .Z(n1041) );
  MUX U541 ( .IN0(n1061), .IN1(n1063), .SEL(n1062), .F(n1020) );
  XNOR U542 ( .A(n1342), .B(n1339), .Z(n1402) );
  MUX U543 ( .IN0(n5491), .IN1(n5493), .SEL(n5492), .F(n5475) );
  MUX U544 ( .IN0(n425), .IN1(n5106), .SEL(n5107), .F(n5092) );
  IV U545 ( .A(n5108), .Z(n425) );
  XNOR U546 ( .A(n4625), .B(n4624), .Z(n4640) );
  MUX U547 ( .IN0(n5569), .IN1(n426), .SEL(n5570), .F(n5551) );
  IV U548 ( .A(n5571), .Z(n426) );
  MUX U549 ( .IN0(n5218), .IN1(n5220), .SEL(n5219), .F(n5198) );
  MUX U550 ( .IN0(n4557), .IN1(n4559), .SEL(n4558), .F(n4545) );
  NANDN U551 ( .B(n2917), .A(n3391), .Z(n439) );
  MUX U552 ( .IN0(n4562), .IN1(n427), .SEL(n4563), .F(n4538) );
  IV U553 ( .A(n4564), .Z(n427) );
  XNOR U554 ( .A(n4272), .B(n4270), .Z(n4285) );
  XNOR U555 ( .A(n5206), .B(n5205), .Z(n5221) );
  MUX U556 ( .IN0(n5356), .IN1(n428), .SEL(n5357), .F(n5344) );
  IV U557 ( .A(n5358), .Z(n428) );
  MUX U558 ( .IN0(n4982), .IN1(n4984), .SEL(n4983), .F(n4965) );
  MUX U559 ( .IN0(n5152), .IN1(n429), .SEL(n5153), .F(n3338) );
  IV U560 ( .A(n5154), .Z(n429) );
  MUX U561 ( .IN0(n1785), .IN1(n430), .SEL(n1786), .F(n1692) );
  IV U562 ( .A(n1787), .Z(n430) );
  MUX U563 ( .IN0(n1934), .IN1(n1936), .SEL(n1935), .F(n1838) );
  MUX U564 ( .IN0(n2058), .IN1(n2060), .SEL(n2059), .F(n1962) );
  MUX U565 ( .IN0(n2234), .IN1(n431), .SEL(n2235), .F(n2126) );
  IV U566 ( .A(n2236), .Z(n431) );
  MUX U567 ( .IN0(n2388), .IN1(n432), .SEL(n2389), .F(n2281) );
  IV U568 ( .A(n2390), .Z(n432) );
  MUX U569 ( .IN0(n2488), .IN1(n433), .SEL(n2489), .F(n2380) );
  IV U570 ( .A(n2490), .Z(n433) );
  MUX U571 ( .IN0(n2583), .IN1(n2585), .SEL(n2584), .F(n2464) );
  MUX U572 ( .IN0(n2575), .IN1(n2577), .SEL(n2576), .F(n2456) );
  MUX U573 ( .IN0(n2665), .IN1(n2667), .SEL(n2666), .F(n2551) );
  MUX U574 ( .IN0(n2958), .IN1(n434), .SEL(n2959), .F(n2833) );
  IV U575 ( .A(n2960), .Z(n434) );
  MUX U576 ( .IN0(n1042), .IN1(n1044), .SEL(n1043), .F(n1002) );
  MUX U577 ( .IN0(n1414), .IN1(n1416), .SEL(n1415), .F(n1346) );
  MUX U578 ( .IN0(A[25]), .IN1(n4820), .SEL(A[31]), .F(n435) );
  IV U579 ( .A(n435), .Z(n1186) );
  MUX U580 ( .IN0(n2413), .IN1(n2415), .SEL(n2414), .F(n2308) );
  XNOR U581 ( .A(n1173), .B(n1172), .Z(n1228) );
  XNOR U582 ( .A(n662), .B(n1663), .Z(n1586) );
  AND U583 ( .A(n942), .B(n944), .Z(n913) );
  MUX U584 ( .IN0(n5122), .IN1(n436), .SEL(n5123), .F(n5106) );
  IV U585 ( .A(n5124), .Z(n436) );
  XNOR U586 ( .A(n5268), .B(n5267), .Z(n5285) );
  MUX U587 ( .IN0(n4167), .IN1(n4169), .SEL(n4168), .F(n4153) );
  MUX U588 ( .IN0(n4582), .IN1(n437), .SEL(n4583), .F(n4562) );
  IV U589 ( .A(n4584), .Z(n437) );
  XNOR U590 ( .A(n3548), .B(n3547), .Z(n3583) );
  MUX U591 ( .IN0(n438), .IN1(n5551), .SEL(n5552), .F(n5535) );
  IV U592 ( .A(n5553), .Z(n438) );
  MUX U593 ( .IN0(n5198), .IN1(n5200), .SEL(n5199), .F(n5178) );
  MUX U594 ( .IN0(n4700), .IN1(n439), .SEL(n4701), .F(n4686) );
  XNOR U595 ( .A(n5000), .B(n4999), .Z(n5005) );
  MUX U596 ( .IN0(n5183), .IN1(n440), .SEL(n5184), .F(n5152) );
  IV U597 ( .A(n5185), .Z(n440) );
  XNOR U598 ( .A(n3530), .B(n3528), .Z(n3565) );
  MUX U599 ( .IN0(n5344), .IN1(n441), .SEL(n5345), .F(n3361) );
  IV U600 ( .A(n5346), .Z(n441) );
  MUX U601 ( .IN0(n2281), .IN1(n442), .SEL(n2282), .F(n2175) );
  IV U602 ( .A(n2283), .Z(n442) );
  MUX U603 ( .IN0(n2719), .IN1(n2721), .SEL(n2720), .F(n2599) );
  MUX U604 ( .IN0(n2849), .IN1(n443), .SEL(n2850), .F(n2727) );
  IV U605 ( .A(n2851), .Z(n443) );
  MUX U606 ( .IN0(n2857), .IN1(n444), .SEL(n2858), .F(n2735) );
  IV U607 ( .A(n2859), .Z(n444) );
  MUX U608 ( .IN0(A[22]), .IN1(n4871), .SEL(A[31]), .F(n445) );
  IV U609 ( .A(n445), .Z(n1385) );
  MUX U610 ( .IN0(A[24]), .IN1(n4837), .SEL(A[31]), .F(n446) );
  IV U611 ( .A(n446), .Z(n1250) );
  MUX U612 ( .IN0(A[17]), .IN1(n4956), .SEL(A[31]), .F(n447) );
  IV U613 ( .A(n447), .Z(n1793) );
  MUX U614 ( .IN0(A[19]), .IN1(n4922), .SEL(A[31]), .F(n448) );
  IV U615 ( .A(n448), .Z(n1618) );
  MUX U616 ( .IN0(A[26]), .IN1(n4804), .SEL(A[31]), .F(n449) );
  IV U617 ( .A(n449), .Z(n1127) );
  MUX U618 ( .IN0(A[27]), .IN1(n4788), .SEL(A[31]), .F(n450) );
  IV U619 ( .A(n450), .Z(n1085) );
  MUX U620 ( .IN0(n1247), .IN1(n1245), .SEL(n1246), .F(n1181) );
  MUX U621 ( .IN0(n2924), .IN1(n2926), .SEL(n2925), .F(n2798) );
  XNOR U622 ( .A(n1410), .B(n1409), .Z(n1476) );
  XOR U623 ( .A(n1754), .B(n1669), .Z(n1670) );
  ANDN U624 ( .A(n964), .B(n944), .Z(n933) );
  XNOR U625 ( .A(n5395), .B(n5394), .Z(n5402) );
  MUX U626 ( .IN0(n4162), .IN1(n451), .SEL(n4163), .F(n4148) );
  IV U627 ( .A(n4164), .Z(n451) );
  MUX U628 ( .IN0(n5137), .IN1(n5139), .SEL(n5138), .F(n5133) );
  MUX U629 ( .IN0(n452), .IN1(n5470), .SEL(n5471), .F(n5456) );
  IV U630 ( .A(n5472), .Z(n452) );
  MUX U631 ( .IN0(n453), .IN1(n5092), .SEL(n5093), .F(n5083) );
  IV U632 ( .A(n5094), .Z(n453) );
  XNOR U633 ( .A(n4585), .B(n4584), .Z(n4600) );
  NANDN U634 ( .B(n5583), .A(n3391), .Z(n469) );
  MUX U635 ( .IN0(n5178), .IN1(n5180), .SEL(n5179), .F(n5159) );
  XNOR U636 ( .A(n5359), .B(n5358), .Z(n5364) );
  XNOR U637 ( .A(n5186), .B(n5185), .Z(n5201) );
  XNOR U638 ( .A(n3424), .B(n3423), .Z(n3458) );
  MUX U639 ( .IN0(n2273), .IN1(n454), .SEL(n2274), .F(n2167) );
  IV U640 ( .A(n2275), .Z(n454) );
  MUX U641 ( .IN0(n2568), .IN1(n455), .SEL(n2569), .F(n2449) );
  IV U642 ( .A(n2570), .Z(n455) );
  MUX U643 ( .IN0(n2760), .IN1(n2762), .SEL(n2761), .F(n2640) );
  MUX U644 ( .IN0(n2982), .IN1(n456), .SEL(n2983), .F(n2857) );
  IV U645 ( .A(n2984), .Z(n456) );
  MUX U646 ( .IN0(A[12]), .IN1(n5379), .SEL(A[31]), .F(n457) );
  IV U647 ( .A(n457), .Z(n2289) );
  MUX U648 ( .IN0(n3177), .IN1(n3179), .SEL(n3178), .F(n3052) );
  MUX U649 ( .IN0(A[20]), .IN1(n4905), .SEL(A[31]), .F(n458) );
  IV U650 ( .A(n458), .Z(n1537) );
  MUX U651 ( .IN0(n3146), .IN1(n459), .SEL(n3147), .F(n3016) );
  IV U652 ( .A(n3148), .Z(n459) );
  MUX U653 ( .IN0(A[15]), .IN1(n5343), .SEL(A[31]), .F(n460) );
  IV U654 ( .A(n460), .Z(n1986) );
  MUX U655 ( .IN0(A[23]), .IN1(n4854), .SEL(A[31]), .F(n461) );
  IV U656 ( .A(n461), .Z(n1318) );
  MUX U657 ( .IN0(A[21]), .IN1(n4888), .SEL(A[31]), .F(n462) );
  IV U658 ( .A(n462), .Z(n1459) );
  MUX U659 ( .IN0(n1159), .IN1(n1161), .SEL(n1160), .F(n1103) );
  MUX U660 ( .IN0(n1315), .IN1(n1313), .SEL(n1314), .F(n1245) );
  MUX U661 ( .IN0(n1374), .IN1(n1372), .SEL(n1373), .F(n1303) );
  MUX U662 ( .IN0(n1563), .IN1(n1561), .SEL(n1562), .F(n1483) );
  MUX U663 ( .IN0(n463), .IN1(n1697), .SEL(n1698), .F(n1613) );
  IV U664 ( .A(n1699), .Z(n463) );
  MUX U665 ( .IN0(n2328), .IN1(n2326), .SEL(n2327), .F(n2218) );
  MUX U666 ( .IN0(n464), .IN1(n2618), .SEL(n2619), .F(n2499) );
  IV U667 ( .A(n2620), .Z(n464) );
  MUX U668 ( .IN0(n1038), .IN1(n1036), .SEL(n1037), .F(n996) );
  MUX U669 ( .IN0(n1346), .IN1(n1348), .SEL(n1347), .F(n1277) );
  MUX U670 ( .IN0(n465), .IN1(n1514), .SEL(n1515), .F(n1434) );
  IV U671 ( .A(n1516), .Z(n465) );
  XOR U672 ( .A(n720), .B(n2003), .Z(n1907) );
  MUX U673 ( .IN0(n2308), .IN1(n2310), .SEL(n2309), .F(n2201) );
  ANDN U674 ( .A(n933), .B(n915), .Z(n904) );
  AND U675 ( .A(n973), .B(n975), .Z(n942) );
  MUX U676 ( .IN0(n1725), .IN1(n1723), .SEL(n1724), .F(n1632) );
  MUX U677 ( .IN0(n5486), .IN1(n466), .SEL(n5487), .F(n5470) );
  IV U678 ( .A(n5488), .Z(n466) );
  MUX U679 ( .IN0(n4597), .IN1(n4599), .SEL(n4598), .F(n4577) );
  MUX U680 ( .IN0(n5574), .IN1(n5576), .SEL(n5575), .F(n5556) );
  XNOR U681 ( .A(n5383), .B(n5382), .Z(n5388) );
  MUX U682 ( .IN0(n467), .IN1(n4148), .SEL(n4149), .F(n4134) );
  IV U683 ( .A(n4150), .Z(n467) );
  MUX U684 ( .IN0(n468), .IN1(n5083), .SEL(n5084), .F(n5071) );
  IV U685 ( .A(n5085), .Z(n468) );
  MUX U686 ( .IN0(n5580), .IN1(n469), .SEL(n5581), .F(n5569) );
  MUX U687 ( .IN0(n5159), .IN1(n5161), .SEL(n5160), .F(n3345) );
  MUX U688 ( .IN0(n2496), .IN1(n470), .SEL(n2497), .F(n2388) );
  IV U689 ( .A(n2498), .Z(n470) );
  MUX U690 ( .IN0(n2464), .IN1(n2466), .SEL(n2465), .F(n2356) );
  MUX U691 ( .IN0(n2658), .IN1(n471), .SEL(n2659), .F(n2544) );
  IV U692 ( .A(n2660), .Z(n471) );
  MUX U693 ( .IN0(n2833), .IN1(n472), .SEL(n2834), .F(n2711) );
  IV U694 ( .A(n2835), .Z(n472) );
  MUX U695 ( .IN0(n2785), .IN1(n2787), .SEL(n2786), .F(n2665) );
  MUX U696 ( .IN0(n3098), .IN1(n3100), .SEL(n3099), .F(n2966) );
  MUX U697 ( .IN0(n3106), .IN1(n473), .SEL(n3107), .F(n2974) );
  IV U698 ( .A(n3108), .Z(n473) );
  MUX U699 ( .IN0(A[16]), .IN1(n4973), .SEL(A[31]), .F(n474) );
  IV U700 ( .A(n474), .Z(n1890) );
  MUX U701 ( .IN0(A[18]), .IN1(n4939), .SEL(A[31]), .F(n475) );
  IV U702 ( .A(n475), .Z(n1702) );
  MUX U703 ( .IN0(A[14]), .IN1(n5355), .SEL(A[31]), .F(n476) );
  IV U704 ( .A(n476), .Z(n2082) );
  MUX U705 ( .IN0(n3138), .IN1(n3140), .SEL(n3139), .F(n3008) );
  MUX U706 ( .IN0(A[13]), .IN1(n5367), .SEL(A[31]), .F(n477) );
  IV U707 ( .A(n477), .Z(n2183) );
  MUX U708 ( .IN0(n3283), .IN1(n478), .SEL(n3284), .F(n3146) );
  IV U709 ( .A(n3285), .Z(n478) );
  XNOR U710 ( .A(n3441), .B(n3440), .Z(n4220) );
  MUX U711 ( .IN0(n1178), .IN1(n479), .SEL(n1179), .F(n1119) );
  IV U712 ( .A(n1180), .Z(n479) );
  MUX U713 ( .IN0(n1412), .IN1(n1410), .SEL(n1411), .F(n1342) );
  MUX U714 ( .IN0(n480), .IN1(n1454), .SEL(n1455), .F(n1380) );
  IV U715 ( .A(n1456), .Z(n480) );
  MUX U716 ( .IN0(n2114), .IN1(n2116), .SEL(n2115), .F(n2013) );
  MUX U717 ( .IN0(n1734), .IN1(n1732), .SEL(n1733), .F(n1643) );
  MUX U718 ( .IN0(n1782), .IN1(n1780), .SEL(n1781), .F(n1687) );
  MUX U719 ( .IN0(n2278), .IN1(n2276), .SEL(n2277), .F(n2170) );
  MUX U720 ( .IN0(n2239), .IN1(n2237), .SEL(n2238), .F(n2129) );
  MUX U721 ( .IN0(n2262), .IN1(n2260), .SEL(n2261), .F(n2154) );
  MUX U722 ( .IN0(n2693), .IN1(n2691), .SEL(n2692), .F(n2571) );
  MUX U723 ( .IN0(n2854), .IN1(n2852), .SEL(n2853), .F(n2730) );
  MUX U724 ( .IN0(n481), .IN1(n2860), .SEL(n2861), .F(n2738) );
  IV U725 ( .A(n2862), .Z(n481) );
  MUX U726 ( .IN0(n1071), .IN1(n1069), .SEL(n1070), .F(n1026) );
  MUX U727 ( .IN0(n1082), .IN1(n1080), .SEL(n1081), .F(n1036) );
  XNOR U728 ( .A(n1235), .B(n1234), .Z(n1296) );
  MUX U729 ( .IN0(n482), .IN1(n1677), .SEL(n1678), .F(n1593) );
  IV U730 ( .A(n1679), .Z(n482) );
  XNOR U731 ( .A(n1755), .B(n1765), .Z(n1854) );
  MUX U732 ( .IN0(n2208), .IN1(n483), .SEL(n2209), .F(n2097) );
  IV U733 ( .A(n2210), .Z(n483) );
  XOR U734 ( .A(n946), .B(n923), .Z(n920) );
  MUX U735 ( .IN0(n1020), .IN1(n1022), .SEL(n1021), .F(n484) );
  IV U736 ( .A(n484), .Z(n986) );
  AND U737 ( .A(n1054), .B(n1056), .Z(n1014) );
  NOR U738 ( .A(n1721), .B(n1722), .Z(n1720) );
  NANDN U739 ( .B(n892), .A(n904), .Z(n872) );
  MUX U740 ( .IN0(n907), .IN1(Y0[29]), .SEL(n908), .F(n884) );
  MUX U741 ( .IN0(n4504), .IN1(n4502), .SEL(n4503), .F(n4481) );
  MUX U742 ( .IN0(n5440), .IN1(n5317), .SEL(n5318), .F(n5426) );
  MUX U743 ( .IN0(n5500), .IN1(n5502), .SEL(n5501), .F(n5497) );
  MUX U744 ( .IN0(n485), .IN1(n5097), .SEL(n5098), .F(n5078) );
  IV U745 ( .A(n5099), .Z(n485) );
  MUX U746 ( .IN0(n486), .IN1(n5456), .SEL(n5457), .F(n5447) );
  IV U747 ( .A(n5458), .Z(n486) );
  NANDN U748 ( .B(n5324), .A(n3391), .Z(n507) );
  MUX U749 ( .IN0(n4545), .IN1(n4547), .SEL(n4546), .F(n4527) );
  XNOR U750 ( .A(n4565), .B(n4564), .Z(n4580) );
  MUX U751 ( .IN0(n487), .IN1(n5524), .SEL(n5525), .F(n3377) );
  IV U752 ( .A(n5526), .Z(n487) );
  XNOR U753 ( .A(n5347), .B(n5346), .Z(n5352) );
  XNOR U754 ( .A(n5076), .B(n5075), .Z(n5081) );
  MUX U755 ( .IN0(n2241), .IN1(n2243), .SEL(n2242), .F(n2133) );
  MUX U756 ( .IN0(n2356), .IN1(n2358), .SEL(n2357), .F(n2249) );
  MUX U757 ( .IN0(n2599), .IN1(n2601), .SEL(n2600), .F(n2480) );
  MUX U758 ( .IN0(n2607), .IN1(n488), .SEL(n2608), .F(n2488) );
  IV U759 ( .A(n2609), .Z(n488) );
  MUX U760 ( .IN0(n2551), .IN1(n2553), .SEL(n2552), .F(n2437) );
  MUX U761 ( .IN0(n2688), .IN1(n489), .SEL(n2689), .F(n2568) );
  IV U762 ( .A(n2690), .Z(n489) );
  MUX U763 ( .IN0(n2884), .IN1(n2886), .SEL(n2885), .F(n2760) );
  MUX U764 ( .IN0(n2892), .IN1(n490), .SEL(n2893), .F(n2768) );
  IV U765 ( .A(n2894), .Z(n490) );
  MUX U766 ( .IN0(n3031), .IN1(n3033), .SEL(n3032), .F(n2907) );
  MUX U767 ( .IN0(n3082), .IN1(n3084), .SEL(n3083), .F(n2950) );
  MUX U768 ( .IN0(n3090), .IN1(n491), .SEL(n3091), .F(n2958) );
  IV U769 ( .A(n3092), .Z(n491) );
  MUX U770 ( .IN0(n3206), .IN1(n3208), .SEL(n3207), .F(n3074) );
  MUX U771 ( .IN0(n3199), .IN1(n492), .SEL(n3200), .F(n3067) );
  IV U772 ( .A(n3201), .Z(n492) );
  MUX U773 ( .IN0(n3246), .IN1(n493), .SEL(n3247), .F(n3114) );
  IV U774 ( .A(n3248), .Z(n493) );
  MUX U775 ( .IN0(n3154), .IN1(n494), .SEL(n3155), .F(n3024) );
  IV U776 ( .A(n3156), .Z(n494) );
  MUX U777 ( .IN0(n5157), .IN1(n5155), .SEL(n5156), .F(n3341) );
  MUX U778 ( .IN0(n3426), .IN1(n3424), .SEL(n3425), .F(n3294) );
  XNOR U779 ( .A(n3416), .B(n3415), .Z(n3478) );
  MUX U780 ( .IN0(n1086), .IN1(n1088), .SEL(n1087), .F(n1042) );
  MUX U781 ( .IN0(n1689), .IN1(n1687), .SEL(n1688), .F(n1603) );
  MUX U782 ( .IN0(n495), .IN1(n2077), .SEL(n2078), .F(n1981) );
  IV U783 ( .A(n2079), .Z(n495) );
  MUX U784 ( .IN0(n2055), .IN1(n2053), .SEL(n2054), .F(n1957) );
  MUX U785 ( .IN0(n2346), .IN1(n2344), .SEL(n2345), .F(n2237) );
  MUX U786 ( .IN0(n2385), .IN1(n2383), .SEL(n2384), .F(n2276) );
  MUX U787 ( .IN0(n2425), .IN1(n2427), .SEL(n2426), .F(n496) );
  IV U788 ( .A(n496), .Z(n2315) );
  MUX U789 ( .IN0(n2596), .IN1(n2594), .SEL(n2595), .F(n2475) );
  MUX U790 ( .IN0(n2783), .IN1(n2781), .SEL(n2782), .F(n2661) );
  MUX U791 ( .IN0(n497), .IN1(n2985), .SEL(n2986), .F(n2860) );
  IV U792 ( .A(n2987), .Z(n497) );
  MUX U793 ( .IN0(n2979), .IN1(n2977), .SEL(n2978), .F(n2852) );
  MUX U794 ( .IN0(n2940), .IN1(n2938), .SEL(n2939), .F(n2813) );
  MUX U795 ( .IN0(n2922), .IN1(n2920), .SEL(n2921), .F(n498) );
  IV U796 ( .A(n498), .Z(n2792) );
  MUX U797 ( .IN0(n3021), .IN1(n3019), .SEL(n3020), .F(n2895) );
  XNOR U798 ( .A(n3310), .B(n3309), .Z(n3434) );
  MUX U799 ( .IN0(n998), .IN1(n996), .SEL(n997), .F(n952) );
  MUX U800 ( .IN0(n1183), .IN1(n1181), .SEL(n1182), .F(n1122) );
  MUX U801 ( .IN0(n1354), .IN1(n1352), .SEL(n1353), .F(n1283) );
  MUX U802 ( .IN0(n499), .IN1(n1362), .SEL(n1363), .F(n1293) );
  IV U803 ( .A(n1364), .Z(n499) );
  XNOR U804 ( .A(n1483), .B(n1482), .Z(n1554) );
  MUX U805 ( .IN0(n500), .IN1(n1772), .SEL(n1773), .F(n1677) );
  IV U806 ( .A(n1774), .Z(n500) );
  XNOR U807 ( .A(n2100), .B(n2009), .Z(n2010) );
  MUX U808 ( .IN0(n2312), .IN1(n501), .SEL(n2313), .F(n2208) );
  IV U809 ( .A(n2314), .Z(n501) );
  MUX U810 ( .IN0(n2798), .IN1(n2800), .SEL(n2799), .F(n2680) );
  ANDN U811 ( .A(n979), .B(n983), .Z(n982) );
  MUX U812 ( .IN0(n502), .IN1(n1213), .SEL(n1214), .F(n1154) );
  IV U813 ( .A(n1215), .Z(n502) );
  ANDN U814 ( .A(n1919), .B(n1921), .Z(n1810) );
  MUX U815 ( .IN0(n550), .IN1(n2560), .SEL(n2559), .F(n2443) );
  NANDN U816 ( .B(n965), .A(n966), .Z(n934) );
  AND U817 ( .A(n1014), .B(n1016), .Z(n973) );
  NANDN U818 ( .B(n1134), .A(n1135), .Z(n1090) );
  AND U819 ( .A(n1332), .B(n1334), .Z(n1264) );
  MUX U820 ( .IN0(n1825), .IN1(n503), .SEL(n1824), .F(n1723) );
  IV U821 ( .A(n1823), .Z(n503) );
  AND U822 ( .A(n880), .B(n881), .Z(n875) );
  MUX U823 ( .IN0(n936), .IN1(Y0[28]), .SEL(n937), .F(n907) );
  MUX U824 ( .IN0(n4111), .IN1(n4109), .SEL(n4110), .F(n4067) );
  MUX U825 ( .IN0(n4176), .IN1(n4178), .SEL(n4177), .F(n4173) );
  MUX U826 ( .IN0(n504), .IN1(n5461), .SEL(n5462), .F(n5442) );
  IV U827 ( .A(n5463), .Z(n504) );
  MUX U828 ( .IN0(n505), .IN1(n4134), .SEL(n4135), .F(n4125) );
  IV U829 ( .A(n4136), .Z(n505) );
  MUX U830 ( .IN0(n506), .IN1(n5078), .SEL(n5079), .F(n5066) );
  IV U831 ( .A(n5080), .Z(n506) );
  MUX U832 ( .IN0(n5321), .IN1(n507), .SEL(n5322), .F(n5309) );
  MUX U833 ( .IN0(n508), .IN1(n5447), .SEL(n5448), .F(n5435) );
  IV U834 ( .A(n5449), .Z(n508) );
  XNOR U835 ( .A(n4541), .B(n4540), .Z(n4560) );
  MUX U836 ( .IN0(n2133), .IN1(n2135), .SEL(n2134), .F(n2032) );
  MUX U837 ( .IN0(n2167), .IN1(n509), .SEL(n2168), .F(n2066) );
  IV U838 ( .A(n2169), .Z(n509) );
  MUX U839 ( .IN0(n2615), .IN1(n510), .SEL(n2616), .F(n2496) );
  IV U840 ( .A(n2617), .Z(n510) );
  MUX U841 ( .IN0(n2727), .IN1(n511), .SEL(n2728), .F(n2607) );
  IV U842 ( .A(n2729), .Z(n511) );
  MUX U843 ( .IN0(n2703), .IN1(n2705), .SEL(n2704), .F(n2583) );
  MUX U844 ( .IN0(n2817), .IN1(n2819), .SEL(n2818), .F(n2695) );
  MUX U845 ( .IN0(n2810), .IN1(n512), .SEL(n2811), .F(n2688) );
  IV U846 ( .A(n2812), .Z(n512) );
  MUX U847 ( .IN0(n2966), .IN1(n2968), .SEL(n2967), .F(n2841) );
  MUX U848 ( .IN0(n2900), .IN1(n513), .SEL(n2901), .F(n2778) );
  IV U849 ( .A(n2902), .Z(n513) );
  MUX U850 ( .IN0(n3214), .IN1(n3216), .SEL(n3215), .F(n3082) );
  MUX U851 ( .IN0(n3222), .IN1(n514), .SEL(n3223), .F(n3090) );
  IV U852 ( .A(n3224), .Z(n514) );
  MUX U853 ( .IN0(n3377), .IN1(n515), .SEL(n3378), .F(n3238) );
  IV U854 ( .A(n3379), .Z(n515) );
  MUX U855 ( .IN0(n3338), .IN1(n516), .SEL(n3339), .F(n3199) );
  IV U856 ( .A(n3340), .Z(n516) );
  MUX U857 ( .IN0(n3275), .IN1(n3277), .SEL(n3276), .F(n3138) );
  MUX U858 ( .IN0(n5347), .IN1(n5173), .SEL(n5175), .F(n3364) );
  MUX U859 ( .IN0(n1128), .IN1(n1130), .SEL(n1129), .F(n1086) );
  MUX U860 ( .IN0(n1932), .IN1(n1930), .SEL(n1931), .F(n1834) );
  MUX U861 ( .IN0(n1975), .IN1(n1973), .SEL(n1974), .F(n1877) );
  MUX U862 ( .IN0(n517), .IN1(n1981), .SEL(n1982), .F(n1885) );
  IV U863 ( .A(n1983), .Z(n517) );
  MUX U864 ( .IN0(n2369), .IN1(n2367), .SEL(n2368), .F(n2260) );
  MUX U865 ( .IN0(n518), .IN1(n2391), .SEL(n2392), .F(n2284) );
  IV U866 ( .A(n2393), .Z(n518) );
  MUX U867 ( .IN0(n2493), .IN1(n2491), .SEL(n2492), .F(n2383) );
  MUX U868 ( .IN0(n2454), .IN1(n2452), .SEL(n2453), .F(n2344) );
  MUX U869 ( .IN0(n2549), .IN1(n2547), .SEL(n2548), .F(n2433) );
  MUX U870 ( .IN0(n2963), .IN1(n2961), .SEL(n2962), .F(n2836) );
  MUX U871 ( .IN0(n2897), .IN1(n2895), .SEL(n2896), .F(n2773) );
  MUX U872 ( .IN0(n3111), .IN1(n3109), .SEL(n3110), .F(n2977) );
  MUX U873 ( .IN0(n519), .IN1(n3117), .SEL(n3118), .F(n2985) );
  IV U874 ( .A(n3119), .Z(n519) );
  MUX U875 ( .IN0(n3072), .IN1(n3070), .SEL(n3071), .F(n2938) );
  MUX U876 ( .IN0(n3159), .IN1(n3157), .SEL(n3158), .F(n3027) );
  XNOR U877 ( .A(n3286), .B(n3285), .Z(n3409) );
  MUX U878 ( .IN0(n1116), .IN1(n1114), .SEL(n1115), .F(n1069) );
  XNOR U879 ( .A(n1181), .B(n1180), .Z(n1238) );
  MUX U880 ( .IN0(n1422), .IN1(n1424), .SEL(n1423), .F(n1352) );
  XNOR U881 ( .A(n1372), .B(n1371), .Z(n1437) );
  XNOR U882 ( .A(n1532), .B(n1531), .Z(n1606) );
  XNOR U883 ( .A(n1561), .B(n1560), .Z(n1636) );
  MUX U884 ( .IN0(n2013), .IN1(n2015), .SEL(n2014), .F(n1912) );
  MUX U885 ( .IN0(n520), .IN1(n1751), .SEL(n1752), .F(n1660) );
  IV U886 ( .A(n1753), .Z(n520) );
  XNOR U887 ( .A(n2101), .B(n2111), .Z(n2211) );
  XOR U888 ( .A(n2529), .B(n2425), .Z(n2426) );
  MUX U889 ( .IN0(n521), .IN1(n2722), .SEL(n2723), .F(n2602) );
  IV U890 ( .A(n2724), .Z(n521) );
  MUX U891 ( .IN0(n2794), .IN1(n522), .SEL(n2793), .F(n2678) );
  IV U892 ( .A(n2792), .Z(n522) );
  MUX U893 ( .IN0(n989), .IN1(n523), .SEL(n988), .F(n961) );
  IV U894 ( .A(n987), .Z(n523) );
  XNOR U895 ( .A(n1152), .B(n1151), .Z(n1205) );
  AND U896 ( .A(n1542), .B(n1544), .Z(n1464) );
  MUX U897 ( .IN0(n524), .IN1(n1650), .SEL(n1651), .F(n1570) );
  IV U898 ( .A(n1652), .Z(n524) );
  MUX U899 ( .IN0(n2804), .IN1(n2806), .SEL(n2805), .F(n2682) );
  NANDN U900 ( .B(n1006), .A(n1007), .Z(n965) );
  ANDN U901 ( .A(n1045), .B(n1016), .Z(n1005) );
  NANDN U902 ( .B(n1193), .A(n1194), .Z(n1134) );
  NAND U903 ( .A(n1810), .B(n1809), .Z(n1721) );
  MUX U904 ( .IN0(n525), .IN1(n2333), .SEL(n2334), .F(n2225) );
  IV U905 ( .A(n2335), .Z(n525) );
  ANDN U906 ( .A(n1473), .B(n1474), .Z(n1399) );
  MUX U907 ( .IN0(Y0[3]), .IN1(n2995), .SEL(n2996), .F(n2872) );
  MUX U908 ( .IN0(n872), .IN1(n874), .SEL(n873), .F(n526) );
  IV U909 ( .A(n526), .Z(n871) );
  MUX U910 ( .IN0(n967), .IN1(Y0[27]), .SEL(n968), .F(n936) );
  MUX U911 ( .IN0(n1136), .IN1(Y0[23]), .SEL(n1137), .F(n1092) );
  MUX U912 ( .IN0(n1393), .IN1(Y0[19]), .SEL(n1394), .F(n1326) );
  MUX U913 ( .IN0(n1710), .IN1(Y0[15]), .SEL(n1711), .F(n1626) );
  MUX U914 ( .IN0(n2090), .IN1(Y0[11]), .SEL(n2091), .F(n1994) );
  MUX U915 ( .IN0(n2512), .IN1(Y0[7]), .SEL(n2513), .F(n2404) );
  MUX U916 ( .IN0(n4980), .IN1(n4534), .SEL(n4535), .F(n4963) );
  MUX U917 ( .IN0(n527), .IN1(n4511), .SEL(n4076), .F(n4490) );
  IV U918 ( .A(n4074), .Z(n527) );
  MUX U919 ( .IN0(n3950), .IN1(n3948), .SEL(n3949), .F(n3904) );
  MUX U920 ( .IN0(n4671), .IN1(n4669), .SEL(n4670), .F(n4645) );
  XNOR U921 ( .A(n5246), .B(n5245), .Z(n5261) );
  MUX U922 ( .IN0(n4703), .IN1(n4705), .SEL(n4704), .F(n4700) );
  MUX U923 ( .IN0(n528), .IN1(n4139), .SEL(n4140), .F(n4118) );
  IV U924 ( .A(n4141), .Z(n528) );
  NANDN U925 ( .B(n2006), .A(n3391), .Z(n560) );
  MUX U926 ( .IN0(n529), .IN1(n5515), .SEL(n5516), .F(n3369) );
  IV U927 ( .A(n5517), .Z(n529) );
  MUX U928 ( .IN0(n5166), .IN1(n5168), .SEL(n5167), .F(n3353) );
  MUX U929 ( .IN0(n4229), .IN1(n4227), .SEL(n4228), .F(n3441) );
  MUX U930 ( .IN0(n2249), .IN1(n2251), .SEL(n2250), .F(n2141) );
  MUX U931 ( .IN0(n2372), .IN1(n2374), .SEL(n2373), .F(n2265) );
  MUX U932 ( .IN0(n2456), .IN1(n2458), .SEL(n2457), .F(n2348) );
  MUX U933 ( .IN0(n2449), .IN1(n530), .SEL(n2450), .F(n2341) );
  IV U934 ( .A(n2451), .Z(n530) );
  MUX U935 ( .IN0(n2711), .IN1(n531), .SEL(n2712), .F(n2591) );
  IV U936 ( .A(n2713), .Z(n531) );
  MUX U937 ( .IN0(n2825), .IN1(n2827), .SEL(n2826), .F(n2703) );
  MUX U938 ( .IN0(n2841), .IN1(n2843), .SEL(n2842), .F(n2719) );
  MUX U939 ( .IN0(n2974), .IN1(n532), .SEL(n2975), .F(n2849) );
  IV U940 ( .A(n2976), .Z(n532) );
  MUX U941 ( .IN0(n2935), .IN1(n533), .SEL(n2936), .F(n2810) );
  IV U942 ( .A(n2937), .Z(n533) );
  MUX U943 ( .IN0(n3024), .IN1(n534), .SEL(n3025), .F(n2900) );
  IV U944 ( .A(n3026), .Z(n534) );
  MUX U945 ( .IN0(n3114), .IN1(n535), .SEL(n3115), .F(n2982) );
  IV U946 ( .A(n3116), .Z(n535) );
  MUX U947 ( .IN0(n3074), .IN1(n3076), .SEL(n3075), .F(n2942) );
  MUX U948 ( .IN0(A[8]), .IN1(n5434), .SEL(A[31]), .F(n536) );
  IV U949 ( .A(n536), .Z(n2743) );
  MUX U950 ( .IN0(n3361), .IN1(n537), .SEL(n3362), .F(n3222) );
  IV U951 ( .A(n3363), .Z(n537) );
  MUX U952 ( .IN0(n3314), .IN1(n3316), .SEL(n3315), .F(n3177) );
  MUX U953 ( .IN0(n1237), .IN1(n1235), .SEL(n1236), .F(n1173) );
  MUX U954 ( .IN0(n2131), .IN1(n2129), .SEL(n2130), .F(n2028) );
  MUX U955 ( .IN0(n2172), .IN1(n2170), .SEL(n2171), .F(n2069) );
  MUX U956 ( .IN0(n2103), .IN1(n2101), .SEL(n2102), .F(n2009) );
  MUX U957 ( .IN0(n538), .IN1(n2284), .SEL(n2285), .F(n2178) );
  IV U958 ( .A(n2286), .Z(n538) );
  MUX U959 ( .IN0(n2477), .IN1(n2475), .SEL(n2476), .F(n2367) );
  MUX U960 ( .IN0(n2573), .IN1(n2571), .SEL(n2572), .F(n2452) );
  MUX U961 ( .IN0(n2612), .IN1(n2610), .SEL(n2611), .F(n2491) );
  MUX U962 ( .IN0(n2532), .IN1(n2530), .SEL(n2531), .F(n2425) );
  MUX U963 ( .IN0(n2663), .IN1(n2661), .SEL(n2662), .F(n2547) );
  MUX U964 ( .IN0(n539), .IN1(n2738), .SEL(n2739), .F(n2618) );
  IV U965 ( .A(n2740), .Z(n539) );
  MUX U966 ( .IN0(n3041), .IN1(n3039), .SEL(n3040), .F(n2920) );
  MUX U967 ( .IN0(n3095), .IN1(n3093), .SEL(n3094), .F(n2961) );
  MUX U968 ( .IN0(n3204), .IN1(n3202), .SEL(n3203), .F(n3070) );
  MUX U969 ( .IN0(n3243), .IN1(n3241), .SEL(n3242), .F(n3109) );
  MUX U970 ( .IN0(n540), .IN1(n3249), .SEL(n3250), .F(n3117) );
  IV U971 ( .A(n3251), .Z(n540) );
  MUX U972 ( .IN0(n3151), .IN1(n3149), .SEL(n3150), .F(n3019) );
  MUX U973 ( .IN0(n3296), .IN1(n3294), .SEL(n3295), .F(n3157) );
  MUX U974 ( .IN0(n1002), .IN1(n1004), .SEL(n1003), .F(n958) );
  MUX U975 ( .IN0(n1124), .IN1(n1122), .SEL(n1123), .F(n1080) );
  XNOR U976 ( .A(n1313), .B(n1312), .Z(n1375) );
  XNOR U977 ( .A(n1524), .B(n1523), .Z(n1596) );
  XNOR U978 ( .A(n1613), .B(n1612), .Z(n1690) );
  XNOR U979 ( .A(n1643), .B(n1642), .Z(n1727) );
  MUX U980 ( .IN0(n541), .IN1(n1869), .SEL(n1870), .F(n1772) );
  IV U981 ( .A(n1871), .Z(n541) );
  XNOR U982 ( .A(n1861), .B(n1860), .Z(n1950) );
  MUX U983 ( .IN0(n2416), .IN1(n542), .SEL(n2417), .F(n2312) );
  IV U984 ( .A(n2418), .Z(n542) );
  MUX U985 ( .IN0(n543), .IN1(n2483), .SEL(n2484), .F(n2375) );
  IV U986 ( .A(n2485), .Z(n543) );
  MUX U987 ( .IN0(n544), .IN1(n2706), .SEL(n2707), .F(n2586) );
  IV U988 ( .A(n2708), .Z(n544) );
  MUX U989 ( .IN0(n545), .IN1(n2969), .SEL(n2970), .F(n2844) );
  IV U990 ( .A(n2971), .Z(n545) );
  MUX U991 ( .IN0(n546), .IN1(n2887), .SEL(n2888), .F(n2763) );
  IV U992 ( .A(n2889), .Z(n546) );
  MUX U993 ( .IN0(n547), .IN1(n949), .SEL(n948), .F(n923) );
  IV U994 ( .A(n947), .Z(n547) );
  AND U995 ( .A(n985), .B(n986), .Z(n981) );
  MUX U996 ( .IN0(n1272), .IN1(n1270), .SEL(n1271), .F(n1210) );
  MUX U997 ( .IN0(n548), .IN1(n1417), .SEL(n1418), .F(n1349) );
  IV U998 ( .A(n1419), .Z(n548) );
  AND U999 ( .A(n1623), .B(n1625), .Z(n1542) );
  MUX U1000 ( .IN0(n1912), .IN1(n1914), .SEL(n1913), .F(n1821) );
  MUX U1001 ( .IN0(n549), .IN1(n2136), .SEL(n2137), .F(n2035) );
  IV U1002 ( .A(n2138), .Z(n549) );
  ANDN U1003 ( .A(n2120), .B(n2122), .Z(n2019) );
  AND U1004 ( .A(n2401), .B(n2403), .Z(n2294) );
  MUX U1005 ( .IN0(n2684), .IN1(n2682), .SEL(n2683), .F(n550) );
  IV U1006 ( .A(n550), .Z(n2558) );
  NANDN U1007 ( .B(n1046), .A(n1047), .Z(n1006) );
  MUX U1008 ( .IN0(n1133), .IN1(n551), .SEL(n1132), .F(n1089) );
  IV U1009 ( .A(n1131), .Z(n551) );
  AND U1010 ( .A(n1201), .B(n1203), .Z(n1190) );
  NANDN U1011 ( .B(n1256), .A(n1257), .Z(n1193) );
  MUX U1012 ( .IN0(n552), .IN1(n1916), .SEL(n1917), .F(n1823) );
  IV U1013 ( .A(n1918), .Z(n552) );
  MUX U1014 ( .IN0(n553), .IN1(n2440), .SEL(n2441), .F(n2333) );
  IV U1015 ( .A(n2442), .Z(n553) );
  MUX U1016 ( .IN0(n2912), .IN1(n580), .SEL(n2911), .F(n554) );
  IV U1017 ( .A(n554), .Z(n2788) );
  AND U1018 ( .A(n913), .B(n915), .Z(n890) );
  ANDN U1019 ( .A(n1551), .B(n1552), .Z(n1473) );
  NAND U1020 ( .A(n861), .B(n863), .Z(n860) );
  MUX U1021 ( .IN0(n1008), .IN1(Y0[26]), .SEL(n1009), .F(n967) );
  MUX U1022 ( .IN0(n1195), .IN1(Y0[22]), .SEL(n1196), .F(n1136) );
  MUX U1023 ( .IN0(n1467), .IN1(Y0[18]), .SEL(n1468), .F(n1393) );
  MUX U1024 ( .IN0(n1801), .IN1(Y0[14]), .SEL(n1802), .F(n1710) );
  MUX U1025 ( .IN0(n2191), .IN1(Y0[10]), .SEL(n2192), .F(n2090) );
  MUX U1026 ( .IN0(n2631), .IN1(Y0[6]), .SEL(n2632), .F(n2512) );
  MUX U1027 ( .IN0(n4525), .IN1(n4523), .SEL(n4524), .F(n4502) );
  MUX U1028 ( .IN0(n4100), .IN1(n4098), .SEL(n4099), .F(n555) );
  IV U1029 ( .A(n555), .Z(n4056) );
  MUX U1030 ( .IN0(n4023), .IN1(n4021), .SEL(n4022), .F(n3975) );
  MUX U1031 ( .IN0(n4946), .IN1(n4492), .SEL(n4493), .F(n4929) );
  MUX U1032 ( .IN0(n556), .IN1(n4427), .SEL(n3894), .F(n4406) );
  IV U1033 ( .A(n3892), .Z(n556) );
  MUX U1034 ( .IN0(n5076), .IN1(n4696), .SEL(n4697), .F(n5064) );
  MUX U1035 ( .IN0(n5314), .IN1(n5312), .SEL(n5313), .F(n5292) );
  XNOR U1036 ( .A(n4645), .B(n4644), .Z(n4662) );
  MUX U1037 ( .IN0(n557), .IN1(n4343), .SEL(n3712), .F(n4322) );
  IV U1038 ( .A(n3710), .Z(n557) );
  MUX U1039 ( .IN0(n5022), .IN1(n4612), .SEL(n4614), .F(n5010) );
  MUX U1040 ( .IN0(n5584), .IN1(n5586), .SEL(n5585), .F(n5580) );
  MUX U1041 ( .IN0(n5228), .IN1(n5226), .SEL(n5227), .F(n5206) );
  MUX U1042 ( .IN0(n558), .IN1(n5540), .SEL(n5541), .F(n5515) );
  IV U1043 ( .A(n5542), .Z(n558) );
  MUX U1044 ( .IN0(n559), .IN1(n5442), .SEL(n5443), .F(n5428) );
  IV U1045 ( .A(n5444), .Z(n559) );
  MUX U1046 ( .IN0(n4194), .IN1(n560), .SEL(n4195), .F(n4080) );
  MUX U1047 ( .IN0(n561), .IN1(n4260), .SEL(n3539), .F(n4239) );
  IV U1048 ( .A(n3537), .Z(n561) );
  MUX U1049 ( .IN0(n2265), .IN1(n2267), .SEL(n2266), .F(n2159) );
  MUX U1050 ( .IN0(n3238), .IN1(n562), .SEL(n3239), .F(n3106) );
  IV U1051 ( .A(n3240), .Z(n562) );
  MUX U1052 ( .IN0(A[7]), .IN1(n5523), .SEL(A[31]), .F(n563) );
  IV U1053 ( .A(n563), .Z(n2865) );
  MUX U1054 ( .IN0(A[11]), .IN1(n5391), .SEL(A[31]), .F(n564) );
  IV U1055 ( .A(n564), .Z(n2396) );
  MUX U1056 ( .IN0(n3298), .IN1(n3300), .SEL(n3299), .F(n3161) );
  MUX U1057 ( .IN0(n3291), .IN1(n565), .SEL(n3292), .F(n3154) );
  IV U1058 ( .A(n3293), .Z(n565) );
  MUX U1059 ( .IN0(n3418), .IN1(n3416), .SEL(n3417), .F(n3286) );
  MUX U1060 ( .IN0(n1187), .IN1(n1189), .SEL(n1188), .F(n1128) );
  MUX U1061 ( .IN0(n1605), .IN1(n1603), .SEL(n1604), .F(n1524) );
  MUX U1062 ( .IN0(n1757), .IN1(n1755), .SEL(n1756), .F(n1669) );
  MUX U1063 ( .IN0(n2156), .IN1(n2154), .SEL(n2155), .F(n2053) );
  MUX U1064 ( .IN0(n2716), .IN1(n2714), .SEL(n2715), .F(n2594) );
  MUX U1065 ( .IN0(n2815), .IN1(n2813), .SEL(n2814), .F(n2691) );
  MUX U1066 ( .IN0(n3029), .IN1(n3027), .SEL(n3028), .F(n2903) );
  MUX U1067 ( .IN0(n3227), .IN1(n3225), .SEL(n3226), .F(n3093) );
  MUX U1068 ( .IN0(n566), .IN1(n3388), .SEL(n3389), .F(n3249) );
  IV U1069 ( .A(n3390), .Z(n566) );
  MUX U1070 ( .IN0(n3382), .IN1(n3380), .SEL(n3381), .F(n3241) );
  MUX U1071 ( .IN0(n3343), .IN1(n3341), .SEL(n3342), .F(n3202) );
  XNOR U1072 ( .A(n1245), .B(n1244), .Z(n1306) );
  XNOR U1073 ( .A(n1303), .B(n1302), .Z(n1365) );
  XNOR U1074 ( .A(n1454), .B(n1453), .Z(n1527) );
  MUX U1075 ( .IN0(n1583), .IN1(n567), .SEL(n1584), .F(n1504) );
  IV U1076 ( .A(n1585), .Z(n567) );
  XNOR U1077 ( .A(n1697), .B(n1696), .Z(n1783) );
  XNOR U1078 ( .A(n1732), .B(n1731), .Z(n1827) );
  XNOR U1079 ( .A(n1877), .B(n1876), .Z(n1968) );
  MUX U1080 ( .IN0(n568), .IN1(n2061), .SEL(n2062), .F(n1965) );
  IV U1081 ( .A(n2063), .Z(n568) );
  XNOR U1082 ( .A(n1981), .B(n1980), .Z(n2072) );
  XNOR U1083 ( .A(n2028), .B(n2027), .Z(n2124) );
  MUX U1084 ( .IN0(n569), .IN1(n2252), .SEL(n2253), .F(n2144) );
  IV U1085 ( .A(n2254), .Z(n569) );
  XNOR U1086 ( .A(n2276), .B(n2275), .Z(n2378) );
  XNOR U1087 ( .A(n2284), .B(n2283), .Z(n2386) );
  XNOR U1088 ( .A(n2433), .B(n2432), .Z(n2542) );
  XNOR U1089 ( .A(n2610), .B(n2609), .Z(n2725) );
  XNOR U1090 ( .A(n2618), .B(n2617), .Z(n2733) );
  XNOR U1091 ( .A(n2653), .B(n2652), .Z(n2766) );
  MUX U1092 ( .IN0(n570), .IN1(n2953), .SEL(n2954), .F(n2828) );
  IV U1093 ( .A(n2955), .Z(n570) );
  XNOR U1094 ( .A(n3039), .B(n3049), .Z(n3168) );
  MUX U1095 ( .IN0(n571), .IN1(n3141), .SEL(n3142), .F(n3011) );
  IV U1096 ( .A(n3143), .Z(n571) );
  XNOR U1097 ( .A(n952), .B(n949), .Z(n990) );
  MUX U1098 ( .IN0(n1028), .IN1(n1026), .SEL(n1027), .F(n979) );
  MUX U1099 ( .IN0(n572), .IN1(n1064), .SEL(n1065), .F(n1023) );
  IV U1100 ( .A(n1066), .Z(n572) );
  AND U1101 ( .A(n1283), .B(n1285), .Z(n1216) );
  MUX U1102 ( .IN0(n573), .IN1(n1492), .SEL(n1493), .F(n1417) );
  IV U1103 ( .A(n1494), .Z(n573) );
  MUX U1104 ( .IN0(n1908), .IN1(n720), .SEL(n1907), .F(n1820) );
  AND U1105 ( .A(n1991), .B(n1993), .Z(n1895) );
  ANDN U1106 ( .A(n2228), .B(n2230), .Z(n2120) );
  MUX U1107 ( .IN0(n574), .IN1(n2351), .SEL(n2352), .F(n2244) );
  IV U1108 ( .A(n2353), .Z(n574) );
  AND U1109 ( .A(n2628), .B(n2630), .Z(n2509) );
  MUX U1110 ( .IN0(n575), .IN1(n2820), .SEL(n2821), .F(n2698) );
  IV U1111 ( .A(n2822), .Z(n575) );
  MUX U1112 ( .IN0(n576), .IN1(n2931), .SEL(n2930), .F(n2804) );
  IV U1113 ( .A(n2929), .Z(n576) );
  NANDN U1114 ( .B(n934), .A(n935), .Z(n905) );
  ANDN U1115 ( .A(n1089), .B(n1056), .Z(n1045) );
  NANDN U1116 ( .B(n1090), .A(n1091), .Z(n1046) );
  MUX U1117 ( .IN0(n1212), .IN1(n1210), .SEL(n1211), .F(n577) );
  IV U1118 ( .A(n577), .Z(n1150) );
  OR U1119 ( .A(n1391), .B(n1392), .Z(n1324) );
  MUX U1120 ( .IN0(n578), .IN1(n2016), .SEL(n2017), .F(n1916) );
  IV U1121 ( .A(n2018), .Z(n578) );
  MUX U1122 ( .IN0(n579), .IN1(n2554), .SEL(n2555), .F(n2440) );
  IV U1123 ( .A(n2556), .Z(n579) );
  MUX U1124 ( .IN0(n3036), .IN1(n613), .SEL(n3035), .F(n580) );
  IV U1125 ( .A(n580), .Z(n2910) );
  AND U1126 ( .A(n1190), .B(n1192), .Z(n1098) );
  MUX U1127 ( .IN0(n581), .IN1(n1632), .SEL(n1633), .F(n1551) );
  IV U1128 ( .A(n1634), .Z(n581) );
  ANDN U1129 ( .A(n865), .B(n866), .Z(n857) );
  MUX U1130 ( .IN0(n1048), .IN1(Y0[25]), .SEL(n1049), .F(n1008) );
  MUX U1131 ( .IN0(n1258), .IN1(Y0[21]), .SEL(n1259), .F(n1195) );
  MUX U1132 ( .IN0(n1545), .IN1(Y0[17]), .SEL(n1546), .F(n1467) );
  MUX U1133 ( .IN0(n1898), .IN1(Y0[13]), .SEL(n1899), .F(n1801) );
  MUX U1134 ( .IN0(n2297), .IN1(Y0[9]), .SEL(n2298), .F(n2191) );
  MUX U1135 ( .IN0(n2751), .IN1(Y0[5]), .SEL(n2752), .F(n2631) );
  MUX U1136 ( .IN0(n884), .IN1(Y0[30]), .SEL(n885), .F(n850) );
  MUX U1137 ( .IN0(n3431), .IN1(n4112), .SEL(n3432), .F(n582) );
  IV U1138 ( .A(n582), .Z(n4070) );
  MUX U1139 ( .IN0(n583), .IN1(n4056), .SEL(n4057), .F(n4010) );
  IV U1140 ( .A(n4058), .Z(n583) );
  MUX U1141 ( .IN0(n4462), .IN1(n4460), .SEL(n4461), .F(n4439) );
  MUX U1142 ( .IN0(n3977), .IN1(n3975), .SEL(n3976), .F(n3929) );
  MUX U1143 ( .IN0(n584), .IN1(n3874), .SEL(n3875), .F(n3828) );
  IV U1144 ( .A(n3876), .Z(n584) );
  MUX U1145 ( .IN0(n4878), .IN1(n4408), .SEL(n4409), .F(n4861) );
  MUX U1146 ( .IN0(n3768), .IN1(n3766), .SEL(n3767), .F(n3722) );
  MUX U1147 ( .IN0(n4378), .IN1(n4376), .SEL(n4377), .F(n4355) );
  MUX U1148 ( .IN0(n3795), .IN1(n3793), .SEL(n3794), .F(n3747) );
  MUX U1149 ( .IN0(n5162), .IN1(n5315), .SEL(n5163), .F(n585) );
  IV U1150 ( .A(n585), .Z(n5295) );
  MUX U1151 ( .IN0(n586), .IN1(n3692), .SEL(n3693), .F(n3647) );
  IV U1152 ( .A(n3694), .Z(n586) );
  MUX U1153 ( .IN0(n4810), .IN1(n4324), .SEL(n4325), .F(n4794) );
  MUX U1154 ( .IN0(n5395), .IN1(n5253), .SEL(n5255), .F(n5383) );
  MUX U1155 ( .IN0(n3592), .IN1(n3590), .SEL(n3591), .F(n3548) );
  MUX U1156 ( .IN0(n5133), .IN1(n587), .SEL(n5134), .F(n5122) );
  IV U1157 ( .A(n5136), .Z(n587) );
  MUX U1158 ( .IN0(n4294), .IN1(n4292), .SEL(n4293), .F(n4272) );
  MUX U1159 ( .IN0(n3617), .IN1(n3615), .SEL(n3616), .F(n3572) );
  MUX U1160 ( .IN0(n5325), .IN1(n5327), .SEL(n5326), .F(n5321) );
  MUX U1161 ( .IN0(n4587), .IN1(n4585), .SEL(n4586), .F(n4565) );
  NANDN U1162 ( .B(n5604), .A(n3391), .Z(n622) );
  MUX U1163 ( .IN0(n588), .IN1(n3519), .SEL(n3520), .F(n3475) );
  IV U1164 ( .A(n3521), .Z(n588) );
  MUX U1165 ( .IN0(n2695), .IN1(n2697), .SEL(n2696), .F(n2575) );
  MUX U1166 ( .IN0(n3067), .IN1(n589), .SEL(n3068), .F(n2935) );
  IV U1167 ( .A(n3069), .Z(n589) );
  MUX U1168 ( .IN0(A[10]), .IN1(n5405), .SEL(A[31]), .F(n590) );
  IV U1169 ( .A(n590), .Z(n2504) );
  MUX U1170 ( .IN0(A[6]), .IN1(n5534), .SEL(A[31]), .F(n591) );
  IV U1171 ( .A(n591), .Z(n2990) );
  MUX U1172 ( .IN0(A[5]), .IN1(n5550), .SEL(A[31]), .F(n592) );
  IV U1173 ( .A(n592), .Z(n3122) );
  MUX U1174 ( .IN0(n4744), .IN1(n4241), .SEL(n4242), .F(n4724) );
  XNOR U1175 ( .A(n4980), .B(n4978), .Z(n4985) );
  MUX U1176 ( .IN0(n3443), .IN1(n3441), .SEL(n3442), .F(n3310) );
  MUX U1177 ( .IN0(n1119), .IN1(n593), .SEL(n1120), .F(n1077) );
  IV U1178 ( .A(n1121), .Z(n593) );
  MUX U1179 ( .IN0(n662), .IN1(n1587), .SEL(n1586), .F(n1498) );
  MUX U1180 ( .IN0(n1959), .IN1(n1957), .SEL(n1958), .F(n1861) );
  MUX U1181 ( .IN0(n594), .IN1(n2178), .SEL(n2179), .F(n2077) );
  IV U1182 ( .A(n2180), .Z(n594) );
  MUX U1183 ( .IN0(n2838), .IN1(n2836), .SEL(n2837), .F(n2714) );
  MUX U1184 ( .IN0(n2775), .IN1(n2773), .SEL(n2774), .F(n2653) );
  MUX U1185 ( .IN0(n2905), .IN1(n2903), .SEL(n2904), .F(n2781) );
  MUX U1186 ( .IN0(n3366), .IN1(n3364), .SEL(n3365), .F(n3225) );
  MUX U1187 ( .IN0(n3288), .IN1(n3286), .SEL(n3287), .F(n3149) );
  XNOR U1188 ( .A(n3380), .B(n3379), .Z(n5520) );
  XNOR U1189 ( .A(n3341), .B(n3340), .Z(n5150) );
  XNOR U1190 ( .A(n3294), .B(n3293), .Z(n3419) );
  MUX U1191 ( .IN0(n1344), .IN1(n1342), .SEL(n1343), .F(n1270) );
  MUX U1192 ( .IN0(n1175), .IN1(n1173), .SEL(n1174), .F(n1114) );
  XNOR U1193 ( .A(n1380), .B(n1379), .Z(n1447) );
  MUX U1194 ( .IN0(n1506), .IN1(n595), .SEL(n1505), .F(n1422) );
  IV U1195 ( .A(n1504), .Z(n595) );
  XNOR U1196 ( .A(n1444), .B(n1443), .Z(n1517) );
  XNOR U1197 ( .A(n1780), .B(n1779), .Z(n1872) );
  XNOR U1198 ( .A(n1788), .B(n1787), .Z(n1880) );
  XNOR U1199 ( .A(n1834), .B(n1833), .Z(n1923) );
  MUX U1200 ( .IN0(n596), .IN1(n2043), .SEL(n2044), .F(n1947) );
  IV U1201 ( .A(n2045), .Z(n596) );
  XNOR U1202 ( .A(n2069), .B(n2068), .Z(n2165) );
  MUX U1203 ( .IN0(n597), .IN1(n2268), .SEL(n2269), .F(n2162) );
  IV U1204 ( .A(n2270), .Z(n597) );
  XNOR U1205 ( .A(n2237), .B(n2236), .Z(n2339) );
  XNOR U1206 ( .A(n2326), .B(n2325), .Z(n2428) );
  XNOR U1207 ( .A(n2367), .B(n2366), .Z(n2470) );
  MUX U1208 ( .IN0(n598), .IN1(n2586), .SEL(n2587), .F(n2467) );
  IV U1209 ( .A(n2588), .Z(n598) );
  MUX U1210 ( .IN0(n599), .IN1(n2643), .SEL(n2644), .F(n2526) );
  IV U1211 ( .A(n2645), .Z(n599) );
  XNOR U1212 ( .A(n2691), .B(n2690), .Z(n2808) );
  XNOR U1213 ( .A(n2730), .B(n2729), .Z(n2847) );
  XNOR U1214 ( .A(n2738), .B(n2737), .Z(n2855) );
  XNOR U1215 ( .A(n3038), .B(n2920), .Z(n2921) );
  MUX U1216 ( .IN0(n600), .IN1(n3217), .SEL(n3218), .F(n3085) );
  IV U1217 ( .A(n3219), .Z(n600) );
  MUX U1218 ( .IN0(n3235), .IN1(n670), .SEL(n3234), .F(n601) );
  IV U1219 ( .A(n601), .Z(n3101) );
  MUX U1220 ( .IN0(n602), .IN1(n3193), .SEL(n3194), .F(n3060) );
  IV U1221 ( .A(n3195), .Z(n602) );
  MUX U1222 ( .IN0(n958), .IN1(n960), .SEL(n959), .F(n928) );
  XNOR U1223 ( .A(n996), .B(n995), .Z(n1029) );
  MUX U1224 ( .IN0(n603), .IN1(n1106), .SEL(n1107), .F(n1064) );
  IV U1225 ( .A(n1108), .Z(n603) );
  MUX U1226 ( .IN0(n604), .IN1(n1280), .SEL(n1281), .F(n1213) );
  IV U1227 ( .A(n1282), .Z(n604) );
  MUX U1228 ( .IN0(n605), .IN1(n1570), .SEL(n1571), .F(n1492) );
  IV U1229 ( .A(n1572), .Z(n605) );
  AND U1230 ( .A(n1798), .B(n1800), .Z(n1707) );
  MUX U1231 ( .IN0(n606), .IN1(n1937), .SEL(n1938), .F(n1841) );
  IV U1232 ( .A(n1939), .Z(n606) );
  XNOR U1233 ( .A(n1819), .B(n1820), .Z(n1816) );
  AND U1234 ( .A(n2019), .B(n2021), .Z(n1919) );
  AND U1235 ( .A(n2188), .B(n2190), .Z(n2087) );
  MUX U1236 ( .IN0(n607), .IN1(n2459), .SEL(n2460), .F(n2351) );
  IV U1237 ( .A(n2461), .Z(n607) );
  AND U1238 ( .A(n2748), .B(n2750), .Z(n2628) );
  MUX U1239 ( .IN0(n608), .IN1(n2945), .SEL(n2946), .F(n2820) );
  IV U1240 ( .A(n2947), .Z(n608) );
  MUX U1241 ( .IN0(n609), .IN1(n3057), .SEL(n3058), .F(n2929) );
  IV U1242 ( .A(n3059), .Z(n609) );
  NAND U1243 ( .A(n923), .B(n922), .Z(n917) );
  XNOR U1244 ( .A(n961), .B(n986), .Z(n977) );
  ANDN U1245 ( .A(n1098), .B(n1099), .Z(n1054) );
  AND U1246 ( .A(n1146), .B(n1147), .Z(n1145) );
  ANDN U1247 ( .A(n1399), .B(n1400), .Z(n1332) );
  NAND U1248 ( .A(n1464), .B(n1466), .Z(n1391) );
  MUX U1249 ( .IN0(n610), .IN1(n2225), .SEL(n2226), .F(n2117) );
  IV U1250 ( .A(n2227), .Z(n610) );
  MUX U1251 ( .IN0(n611), .IN1(n2443), .SEL(n2444), .F(n2336) );
  IV U1252 ( .A(n2445), .Z(n611) );
  MUX U1253 ( .IN0(n612), .IN1(n2668), .SEL(n2669), .F(n2554) );
  IV U1254 ( .A(n2670), .Z(n612) );
  MUX U1255 ( .IN0(n3166), .IN1(n644), .SEL(n3165), .F(n613) );
  IV U1256 ( .A(n613), .Z(n3034) );
  XNOR U1257 ( .A(n934), .B(n939), .Z(n935) );
  XNOR U1258 ( .A(n1046), .B(n1051), .Z(n1047) );
  XNOR U1259 ( .A(n1193), .B(n1198), .Z(n1194) );
  XOR U1260 ( .A(n1632), .B(n1721), .Z(n1716) );
  XNOR U1261 ( .A(n3303), .B(n3302), .Z(n3134) );
  MUX U1262 ( .IN0(n1092), .IN1(Y0[24]), .SEL(n1093), .F(n1048) );
  MUX U1263 ( .IN0(n1326), .IN1(Y0[20]), .SEL(n1327), .F(n1258) );
  MUX U1264 ( .IN0(n1626), .IN1(Y0[16]), .SEL(n1627), .F(n1545) );
  MUX U1265 ( .IN0(n1994), .IN1(Y0[12]), .SEL(n1995), .F(n1898) );
  MUX U1266 ( .IN0(n2404), .IN1(Y0[8]), .SEL(n2405), .F(n2297) );
  MUX U1267 ( .IN0(Y0[4]), .IN1(n2872), .SEL(n2873), .F(n2751) );
  XNOR U1268 ( .A(n884), .B(n888), .Z(n886) );
  MUX U1269 ( .IN0(n4042), .IN1(n4040), .SEL(n4041), .F(n3994) );
  MUX U1270 ( .IN0(n4963), .IN1(n4513), .SEL(n4514), .F(n4946) );
  MUX U1271 ( .IN0(n614), .IN1(n4490), .SEL(n4030), .F(n4469) );
  IV U1272 ( .A(n4028), .Z(n614) );
  MUX U1273 ( .IN0(n4441), .IN1(n4439), .SEL(n4440), .F(n4418) );
  MUX U1274 ( .IN0(n3931), .IN1(n3929), .SEL(n3930), .F(n3885) );
  MUX U1275 ( .IN0(n615), .IN1(n3964), .SEL(n3965), .F(n3918) );
  IV U1276 ( .A(n3966), .Z(n615) );
  MUX U1277 ( .IN0(n3860), .IN1(n3858), .SEL(n3859), .F(n3812) );
  MUX U1278 ( .IN0(n4895), .IN1(n4429), .SEL(n4430), .F(n4878) );
  MUX U1279 ( .IN0(n4693), .IN1(n4691), .SEL(n4692), .F(n4669) );
  MUX U1280 ( .IN0(n616), .IN1(n4406), .SEL(n3848), .F(n4385) );
  IV U1281 ( .A(n3846), .Z(n616) );
  MUX U1282 ( .IN0(n5064), .IN1(n4676), .SEL(n4678), .F(n5052) );
  MUX U1283 ( .IN0(n4357), .IN1(n4355), .SEL(n4356), .F(n4334) );
  MUX U1284 ( .IN0(n3749), .IN1(n3747), .SEL(n3748), .F(n3703) );
  MUX U1285 ( .IN0(n617), .IN1(n3782), .SEL(n3783), .F(n3736) );
  IV U1286 ( .A(n3784), .Z(n617) );
  MUX U1287 ( .IN0(n3678), .IN1(n3676), .SEL(n3677), .F(n3633) );
  MUX U1288 ( .IN0(n4827), .IN1(n4345), .SEL(n4346), .F(n4810) );
  MUX U1289 ( .IN0(n5130), .IN1(n4716), .SEL(n4717), .F(n618) );
  IV U1290 ( .A(n618), .Z(n5116) );
  MUX U1291 ( .IN0(n5248), .IN1(n5246), .SEL(n5247), .F(n5226) );
  MUX U1292 ( .IN0(n4607), .IN1(n4605), .SEL(n4606), .F(n4585) );
  MUX U1293 ( .IN0(n619), .IN1(n4322), .SEL(n3666), .F(n4301) );
  IV U1294 ( .A(n3664), .Z(n619) );
  MUX U1295 ( .IN0(n5383), .IN1(n5233), .SEL(n5235), .F(n5371) );
  MUX U1296 ( .IN0(n4197), .IN1(n4199), .SEL(n4198), .F(n4194) );
  MUX U1297 ( .IN0(n5010), .IN1(n4592), .SEL(n4594), .F(n5000) );
  MUX U1298 ( .IN0(n4274), .IN1(n4272), .SEL(n4273), .F(n4251) );
  MUX U1299 ( .IN0(n3574), .IN1(n3572), .SEL(n3573), .F(n3530) );
  MUX U1300 ( .IN0(n620), .IN1(n3604), .SEL(n3605), .F(n3562) );
  IV U1301 ( .A(n3606), .Z(n620) );
  MUX U1302 ( .IN0(n3505), .IN1(n3503), .SEL(n3504), .F(n3463) );
  MUX U1303 ( .IN0(n621), .IN1(n4118), .SEL(n4119), .F(n4093) );
  IV U1304 ( .A(n4120), .Z(n621) );
  XNOR U1305 ( .A(n5599), .B(A[3]), .Z(n5600) );
  MUX U1306 ( .IN0(n4761), .IN1(n4262), .SEL(n4263), .F(n4744) );
  MUX U1307 ( .IN0(n5601), .IN1(n622), .SEL(n5602), .F(n3385) );
  MUX U1308 ( .IN0(n2480), .IN1(n2482), .SEL(n2481), .F(n2372) );
  MUX U1309 ( .IN0(n2735), .IN1(n623), .SEL(n2736), .F(n2615) );
  IV U1310 ( .A(n2737), .Z(n623) );
  MUX U1311 ( .IN0(n2950), .IN1(n2952), .SEL(n2951), .F(n2825) );
  MUX U1312 ( .IN0(n2907), .IN1(n2909), .SEL(n2908), .F(n2785) );
  MUX U1313 ( .IN0(n3230), .IN1(n3232), .SEL(n3231), .F(n3098) );
  XNOR U1314 ( .A(n5440), .B(n5439), .Z(n5445) );
  XNOR U1315 ( .A(n5155), .B(n5154), .Z(n5181) );
  XNOR U1316 ( .A(n4523), .B(n4521), .Z(n4536) );
  MUX U1317 ( .IN0(n624), .IN1(n4239), .SEL(n3494), .F(n4219) );
  IV U1318 ( .A(n3492), .Z(n624) );
  MUX U1319 ( .IN0(n1305), .IN1(n1303), .SEL(n1304), .F(n1235) );
  MUX U1320 ( .IN0(n1382), .IN1(n1380), .SEL(n1381), .F(n1313) );
  MUX U1321 ( .IN0(n625), .IN1(n5507), .SEL(X[31]), .F(n1501) );
  IV U1322 ( .A(X[19]), .Z(n625) );
  MUX U1323 ( .IN0(n626), .IN1(n1788), .SEL(n1789), .F(n1697) );
  IV U1324 ( .A(n1790), .Z(n626) );
  MUX U1325 ( .IN0(n627), .IN1(n4204), .SEL(X[31]), .F(n2006) );
  IV U1326 ( .A(X[13]), .Z(n627) );
  MUX U1327 ( .IN0(n2030), .IN1(n2028), .SEL(n2029), .F(n1930) );
  MUX U1328 ( .IN0(n2220), .IN1(n2218), .SEL(n2219), .F(n2101) );
  MUX U1329 ( .IN0(n628), .IN1(n2499), .SEL(n2500), .F(n2391) );
  IV U1330 ( .A(n2501), .Z(n628) );
  MUX U1331 ( .IN0(n2732), .IN1(n2730), .SEL(n2731), .F(n2610) );
  MUX U1332 ( .IN0(n3312), .IN1(n3310), .SEL(n3311), .F(n3173) );
  XNOR U1333 ( .A(n3364), .B(n3363), .Z(n5340) );
  MUX U1334 ( .IN0(n629), .IN1(n3406), .SEL(n3407), .F(n3278) );
  IV U1335 ( .A(n3408), .Z(n629) );
  XOR U1336 ( .A(n1336), .B(n1274), .Z(n1271) );
  MUX U1337 ( .IN0(n630), .IN1(n1434), .SEL(n1435), .F(n1362) );
  IV U1338 ( .A(n1436), .Z(n630) );
  ANDN U1339 ( .A(n1498), .B(n1497), .Z(n1425) );
  XNOR U1340 ( .A(n1603), .B(n1602), .Z(n1680) );
  MUX U1341 ( .IN0(n1660), .IN1(n631), .SEL(n1661), .F(n1583) );
  IV U1342 ( .A(n1662), .Z(n631) );
  XNOR U1343 ( .A(n1973), .B(n1972), .Z(n2064) );
  XNOR U1344 ( .A(n1957), .B(n1956), .Z(n2046) );
  MUX U1345 ( .IN0(n632), .IN1(n2144), .SEL(n2145), .F(n2043) );
  IV U1346 ( .A(n2146), .Z(n632) );
  MUX U1347 ( .IN0(n633), .IN1(n2162), .SEL(n2163), .F(n2061) );
  IV U1348 ( .A(n2164), .Z(n633) );
  XNOR U1349 ( .A(n2077), .B(n2076), .Z(n2173) );
  XNOR U1350 ( .A(n2260), .B(n2259), .Z(n2362) );
  MUX U1351 ( .IN0(n634), .IN1(n2602), .SEL(n2603), .F(n2483) );
  IV U1352 ( .A(n2604), .Z(n634) );
  XNOR U1353 ( .A(n2530), .B(n2540), .Z(n2646) );
  XNOR U1354 ( .A(n2547), .B(n2546), .Z(n2656) );
  XNOR U1355 ( .A(n2571), .B(n2570), .Z(n2686) );
  XNOR U1356 ( .A(n2594), .B(n2593), .Z(n2709) );
  MUX U1357 ( .IN0(n635), .IN1(n2828), .SEL(n2829), .F(n2706) );
  IV U1358 ( .A(n2830), .Z(n635) );
  XNOR U1359 ( .A(n2903), .B(n2902), .Z(n3022) );
  XNOR U1360 ( .A(n2895), .B(n2894), .Z(n3014) );
  XNOR U1361 ( .A(n2961), .B(n2960), .Z(n3088) );
  XNOR U1362 ( .A(n3070), .B(n3069), .Z(n3197) );
  XNOR U1363 ( .A(n3109), .B(n3108), .Z(n3236) );
  XNOR U1364 ( .A(n3117), .B(n3116), .Z(n3244) );
  MUX U1365 ( .IN0(n963), .IN1(n961), .SEL(n962), .F(n931) );
  NAND U1366 ( .A(n1074), .B(n1073), .Z(n1067) );
  XNOR U1367 ( .A(n1036), .B(n1035), .Z(n1075) );
  MUX U1368 ( .IN0(n636), .IN1(n1162), .SEL(n1163), .F(n1106) );
  IV U1369 ( .A(n1164), .Z(n636) );
  AND U1370 ( .A(n1707), .B(n1709), .Z(n1623) );
  MUX U1371 ( .IN0(n637), .IN1(n1741), .SEL(n1742), .F(n1650) );
  IV U1372 ( .A(n1743), .Z(n637) );
  MUX U1373 ( .IN0(n638), .IN1(n2244), .SEL(n2245), .F(n2136) );
  IV U1374 ( .A(n2246), .Z(n638) );
  AND U1375 ( .A(n2294), .B(n2296), .Z(n2188) );
  MUX U1376 ( .IN0(n639), .IN1(n2698), .SEL(n2699), .F(n2578) );
  IV U1377 ( .A(n2700), .Z(n639) );
  XNOR U1378 ( .A(n2679), .B(n2678), .Z(n2676) );
  ANDN U1379 ( .A(n2870), .B(n2871), .Z(n2748) );
  MUX U1380 ( .IN0(n3060), .IN1(n3183), .SEL(n3062), .F(n2927) );
  MUX U1381 ( .IN0(n3211), .IN1(n733), .SEL(n3210), .F(n640) );
  IV U1382 ( .A(n640), .Z(n3077) );
  MUX U1383 ( .IN0(n641), .IN1(n3180), .SEL(n3181), .F(n3057) );
  IV U1384 ( .A(n3182), .Z(n641) );
  ANDN U1385 ( .A(n1005), .B(n975), .Z(n964) );
  MUX U1386 ( .IN0(n1207), .IN1(n1209), .SEL(n1208), .F(n642) );
  IV U1387 ( .A(n642), .Z(n1152) );
  AND U1388 ( .A(n1264), .B(n1266), .Z(n1201) );
  XOR U1389 ( .A(n1216), .B(n1213), .Z(n1267) );
  NANDN U1390 ( .B(n1324), .A(n1325), .Z(n1256) );
  XNOR U1391 ( .A(n2001), .B(n2002), .Z(n2021) );
  MUX U1392 ( .IN0(n643), .IN1(n2788), .SEL(n2789), .F(n2668) );
  IV U1393 ( .A(n2790), .Z(n643) );
  MUX U1394 ( .IN0(n3303), .IN1(n3301), .SEL(n3302), .F(n644) );
  IV U1395 ( .A(n644), .Z(n3164) );
  MUX U1396 ( .IN0(n901), .IN1(n899), .SEL(n900), .F(n645) );
  IV U1397 ( .A(n645), .Z(n878) );
  NANDN U1398 ( .B(n905), .A(n906), .Z(n862) );
  XOR U1399 ( .A(n1494), .B(n1493), .Z(n1474) );
  XOR U1400 ( .A(n1723), .B(n1722), .Z(n1807) );
  XOR U1401 ( .A(n2336), .B(n2333), .Z(n2410) );
  AND U1402 ( .A(n890), .B(n892), .Z(n865) );
  MUX U1403 ( .IN0(n3259), .IN1(Y0[1]), .SEL(n3260), .F(n3127) );
  XNOR U1404 ( .A(n936), .B(n940), .Z(n938) );
  XNOR U1405 ( .A(n1048), .B(n1052), .Z(n1050) );
  XNOR U1406 ( .A(n1195), .B(n1199), .Z(n1197) );
  XNOR U1407 ( .A(n1393), .B(n1397), .Z(n1395) );
  XNOR U1408 ( .A(n1626), .B(n1630), .Z(n1628) );
  XNOR U1409 ( .A(n1898), .B(n1902), .Z(n1900) );
  XNOR U1410 ( .A(n2191), .B(n2195), .Z(n2193) );
  XNOR U1411 ( .A(n2512), .B(n2516), .Z(n2514) );
  MUX U1412 ( .IN0(n646), .IN1(n4532), .SEL(n4115), .F(n4511) );
  IV U1413 ( .A(n4114), .Z(n646) );
  MUX U1414 ( .IN0(n3996), .IN1(n3994), .SEL(n3995), .F(n3948) );
  MUX U1415 ( .IN0(n4483), .IN1(n4481), .SEL(n4482), .F(n4460) );
  MUX U1416 ( .IN0(n4929), .IN1(n4471), .SEL(n4472), .F(n4912) );
  MUX U1417 ( .IN0(n647), .IN1(n3918), .SEL(n3919), .F(n3874) );
  IV U1418 ( .A(n3920), .Z(n647) );
  MUX U1419 ( .IN0(n648), .IN1(n4448), .SEL(n3938), .F(n4427) );
  IV U1420 ( .A(n3936), .Z(n648) );
  MUX U1421 ( .IN0(n3814), .IN1(n3812), .SEL(n3813), .F(n3766) );
  MUX U1422 ( .IN0(n4399), .IN1(n4397), .SEL(n4398), .F(n4376) );
  MUX U1423 ( .IN0(n3841), .IN1(n3839), .SEL(n3840), .F(n3793) );
  MUX U1424 ( .IN0(n4861), .IN1(n4387), .SEL(n4388), .F(n4844) );
  MUX U1425 ( .IN0(n4210), .IN1(n4694), .SEL(n4211), .F(n649) );
  IV U1426 ( .A(n649), .Z(n4672) );
  MUX U1427 ( .IN0(n5052), .IN1(n4652), .SEL(n4654), .F(n5037) );
  MUX U1428 ( .IN0(n4647), .IN1(n4645), .SEL(n4646), .F(n4625) );
  MUX U1429 ( .IN0(n650), .IN1(n3736), .SEL(n3737), .F(n3692) );
  IV U1430 ( .A(n3738), .Z(n650) );
  MUX U1431 ( .IN0(n651), .IN1(n4364), .SEL(n3756), .F(n4343) );
  IV U1432 ( .A(n3754), .Z(n651) );
  MUX U1433 ( .IN0(n5270), .IN1(n5268), .SEL(n5269), .F(n5246) );
  MUX U1434 ( .IN0(n5409), .IN1(n5275), .SEL(n5277), .F(n5395) );
  MUX U1435 ( .IN0(n3635), .IN1(n3633), .SEL(n3634), .F(n3590) );
  MUX U1436 ( .IN0(n4315), .IN1(n4313), .SEL(n4314), .F(n4292) );
  MUX U1437 ( .IN0(n3659), .IN1(n3657), .SEL(n3658), .F(n3615) );
  MUX U1438 ( .IN0(n4794), .IN1(n4303), .SEL(n4304), .F(n4778) );
  MUX U1439 ( .IN0(A[1]), .IN1(n5616), .SEL(A[31]), .F(n652) );
  IV U1440 ( .A(n652), .Z(n4184) );
  MUX U1441 ( .IN0(n653), .IN1(n5535), .SEL(n5536), .F(n5524) );
  IV U1442 ( .A(n5537), .Z(n653) );
  MUX U1443 ( .IN0(n5000), .IN1(n4572), .SEL(n4574), .F(n4990) );
  MUX U1444 ( .IN0(n4567), .IN1(n4565), .SEL(n4566), .F(n4541) );
  MUX U1445 ( .IN0(n654), .IN1(n3562), .SEL(n3563), .F(n3519) );
  IV U1446 ( .A(n3564), .Z(n654) );
  MUX U1447 ( .IN0(n655), .IN1(n4281), .SEL(n3581), .F(n4260) );
  IV U1448 ( .A(n3579), .Z(n655) );
  XNOR U1449 ( .A(n5522), .B(A[7]), .Z(n5523) );
  XNOR U1450 ( .A(n5390), .B(A[11]), .Z(n5391) );
  XNOR U1451 ( .A(n5342), .B(A[15]), .Z(n5343) );
  XNOR U1452 ( .A(n4853), .B(A[23]), .Z(n4854) );
  XNOR U1453 ( .A(n4921), .B(A[19]), .Z(n4922) );
  MUX U1454 ( .IN0(A[2]), .IN1(n5609), .SEL(A[31]), .F(n656) );
  IV U1455 ( .A(n656), .Z(n4181) );
  MUX U1456 ( .IN0(n5188), .IN1(n5186), .SEL(n5187), .F(n5155) );
  MUX U1457 ( .IN0(n5359), .IN1(n5193), .SEL(n5195), .F(n5347) );
  MUX U1458 ( .IN0(n3465), .IN1(n3463), .SEL(n3464), .F(n3424) );
  MUX U1459 ( .IN0(n3487), .IN1(n3485), .SEL(n3486), .F(n3416) );
  XNOR U1460 ( .A(n4787), .B(A[27]), .Z(n4788) );
  MUX U1461 ( .IN0(n657), .IN1(n4191), .SEL(X[31]), .F(n2422) );
  IV U1462 ( .A(X[9]), .Z(n657) );
  MUX U1463 ( .IN0(n2942), .IN1(n2944), .SEL(n2943), .F(n2817) );
  MUX U1464 ( .IN0(n3161), .IN1(n3163), .SEL(n3162), .F(n3031) );
  MUX U1465 ( .IN0(A[4]), .IN1(n5568), .SEL(A[31]), .F(n3120) );
  MUX U1466 ( .IN0(n3385), .IN1(n658), .SEL(n3386), .F(n3246) );
  IV U1467 ( .A(n3387), .Z(n658) );
  MUX U1468 ( .IN0(A[9]), .IN1(n5419), .SEL(A[31]), .F(n659) );
  IV U1469 ( .A(n659), .Z(n2623) );
  MUX U1470 ( .IN0(n3353), .IN1(n3355), .SEL(n3354), .F(n3214) );
  MUX U1471 ( .IN0(X[1]), .IN1(n5148), .SEL(X[31]), .F(n660) );
  IV U1472 ( .A(n660), .Z(n4721) );
  XNOR U1473 ( .A(n4109), .B(n4107), .Z(n4123) );
  MUX U1474 ( .IN0(n1446), .IN1(n1444), .SEL(n1445), .F(n1372) );
  MUX U1475 ( .IN0(n661), .IN1(n1613), .SEL(n1614), .F(n1532) );
  IV U1476 ( .A(n1615), .Z(n661) );
  MUX U1477 ( .IN0(n1645), .IN1(n1643), .SEL(n1644), .F(n1561) );
  MUX U1478 ( .IN0(n1669), .IN1(n1671), .SEL(n1670), .F(n662) );
  MUX U1479 ( .IN0(n2071), .IN1(n2069), .SEL(n2070), .F(n1973) );
  MUX U1480 ( .IN0(n2655), .IN1(n2653), .SEL(n2654), .F(n2530) );
  MUX U1481 ( .IN0(n3175), .IN1(n3173), .SEL(n3174), .F(n3039) );
  MUX U1482 ( .IN0(n4724), .IN1(n4237), .SEL(n4238), .F(n663) );
  IV U1483 ( .A(n663), .Z(n3331) );
  XNOR U1484 ( .A(n5318), .B(n5315), .Z(n5316) );
  XNOR U1485 ( .A(n5621), .B(X[30]), .Z(n5619) );
  MUX U1486 ( .IN0(n664), .IN1(n1225), .SEL(n1226), .F(n1162) );
  IV U1487 ( .A(n1227), .Z(n664) );
  XNOR U1488 ( .A(n1687), .B(n1686), .Z(n1775) );
  MUX U1489 ( .IN0(n665), .IN1(n1851), .SEL(n1852), .F(n1751) );
  IV U1490 ( .A(n1853), .Z(n665) );
  MUX U1491 ( .IN0(n666), .IN1(n1965), .SEL(n1966), .F(n1869) );
  IV U1492 ( .A(n1967), .Z(n666) );
  XNOR U1493 ( .A(n1885), .B(n1884), .Z(n1976) );
  XNOR U1494 ( .A(n1930), .B(n1929), .Z(n2023) );
  XNOR U1495 ( .A(n2053), .B(n2052), .Z(n2147) );
  XNOR U1496 ( .A(n2218), .B(n2217), .Z(n2319) );
  XNOR U1497 ( .A(n2383), .B(n2382), .Z(n2486) );
  XNOR U1498 ( .A(n2391), .B(n2390), .Z(n2494) );
  XNOR U1499 ( .A(n2344), .B(n2343), .Z(n2447) );
  MUX U1500 ( .IN0(n667), .IN1(n2467), .SEL(n2468), .F(n2359) );
  IV U1501 ( .A(n2469), .Z(n667) );
  XNOR U1502 ( .A(n2714), .B(n2713), .Z(n2831) );
  MUX U1503 ( .IN0(n668), .IN1(n2844), .SEL(n2845), .F(n2722) );
  IV U1504 ( .A(n2846), .Z(n668) );
  XNOR U1505 ( .A(n2661), .B(n2660), .Z(n2776) );
  MUX U1506 ( .IN0(n669), .IN1(n2763), .SEL(n2764), .F(n2643) );
  IV U1507 ( .A(n2765), .Z(n669) );
  XNOR U1508 ( .A(n2977), .B(n2976), .Z(n3104) );
  XNOR U1509 ( .A(n2985), .B(n2984), .Z(n3112) );
  XNOR U1510 ( .A(n2938), .B(n2937), .Z(n3065) );
  XNOR U1511 ( .A(n3093), .B(n3092), .Z(n3220) );
  XNOR U1512 ( .A(n3027), .B(n3026), .Z(n3152) );
  XNOR U1513 ( .A(n3019), .B(n3018), .Z(n3144) );
  MUX U1514 ( .IN0(n3374), .IN1(n3372), .SEL(n3373), .F(n670) );
  IV U1515 ( .A(n670), .Z(n3233) );
  MUX U1516 ( .IN0(n671), .IN1(n3356), .SEL(n3357), .F(n3217) );
  IV U1517 ( .A(n3358), .Z(n671) );
  MUX U1518 ( .IN0(n672), .IN1(n3278), .SEL(n3279), .F(n3141) );
  IV U1519 ( .A(n3280), .Z(n672) );
  MUX U1520 ( .IN0(n3328), .IN1(n673), .SEL(n3329), .F(n3193) );
  IV U1521 ( .A(n3330), .Z(n673) );
  MUX U1522 ( .IN0(n954), .IN1(n952), .SEL(n953), .F(n919) );
  MUX U1523 ( .IN0(n674), .IN1(n1023), .SEL(n1024), .F(n987) );
  IV U1524 ( .A(n1025), .Z(n674) );
  XNOR U1525 ( .A(n1080), .B(n1079), .Z(n1117) );
  XNOR U1526 ( .A(n1114), .B(n1112), .Z(n1165) );
  AND U1527 ( .A(n1216), .B(n1217), .Z(n1146) );
  MUX U1528 ( .IN0(n675), .IN1(n1349), .SEL(n1350), .F(n1280) );
  IV U1529 ( .A(n1351), .Z(n675) );
  XOR U1530 ( .A(n1422), .B(n1426), .Z(n1495) );
  XNOR U1531 ( .A(n1908), .B(n1907), .Z(n1906) );
  MUX U1532 ( .IN0(n676), .IN1(n2035), .SEL(n2036), .F(n1937) );
  IV U1533 ( .A(n2037), .Z(n676) );
  AND U1534 ( .A(n2087), .B(n2089), .Z(n1991) );
  MUX U1535 ( .IN0(n677), .IN1(n2099), .SEL(n2098), .F(n2002) );
  IV U1536 ( .A(n2097), .Z(n677) );
  AND U1537 ( .A(n2509), .B(n2511), .Z(n2401) );
  MUX U1538 ( .IN0(n678), .IN1(n2578), .SEL(n2579), .F(n2459) );
  IV U1539 ( .A(n2580), .Z(n678) );
  MUX U1540 ( .IN0(n679), .IN1(n3077), .SEL(n3078), .F(n2945) );
  IV U1541 ( .A(n3079), .Z(n679) );
  MUX U1542 ( .IN0(n928), .IN1(n930), .SEL(n929), .F(n896) );
  AND U1543 ( .A(n1151), .B(n1152), .Z(n1148) );
  MUX U1544 ( .IN0(n680), .IN1(n2117), .SEL(n2118), .F(n2016) );
  IV U1545 ( .A(n2119), .Z(n680) );
  XOR U1546 ( .A(n2557), .B(n2443), .Z(n2444) );
  XNOR U1547 ( .A(n2804), .B(n2802), .Z(n2913) );
  NANDN U1548 ( .B(n903), .A(n902), .Z(n874) );
  XNOR U1549 ( .A(n905), .B(n910), .Z(n906) );
  XNOR U1550 ( .A(n1006), .B(n1011), .Z(n1007) );
  XNOR U1551 ( .A(n1134), .B(n1099), .Z(n1135) );
  XNOR U1552 ( .A(n1324), .B(n1329), .Z(n1325) );
  XOR U1553 ( .A(n1572), .B(n1571), .Z(n1552) );
  MUX U1554 ( .IN0(Y0[2]), .IN1(n3127), .SEL(n3128), .F(n2995) );
  XOR U1555 ( .A(n1725), .B(n1724), .Z(n1804) );
  XOR U1556 ( .A(n2335), .B(n2334), .Z(n2407) );
  XOR U1557 ( .A(n2670), .B(n2669), .Z(n2754) );
  XNOR U1558 ( .A(n3000), .B(n2879), .Z(n2880) );
  XOR U1559 ( .A(n3166), .B(n3165), .Z(n3269) );
  XNOR U1560 ( .A(n967), .B(n971), .Z(n969) );
  XNOR U1561 ( .A(n1092), .B(n1096), .Z(n1094) );
  XNOR U1562 ( .A(n1258), .B(n1262), .Z(n1260) );
  XNOR U1563 ( .A(n1467), .B(n1471), .Z(n1469) );
  XNOR U1564 ( .A(n1710), .B(n1714), .Z(n1712) );
  XNOR U1565 ( .A(n1994), .B(n1998), .Z(n1996) );
  XNOR U1566 ( .A(n2297), .B(n2301), .Z(n2299) );
  XNOR U1567 ( .A(n2631), .B(n2635), .Z(n2633) );
  XOR U1568 ( .A(n850), .B(n851), .Z(n737) );
  MUX U1569 ( .IN0(n4086), .IN1(n4084), .SEL(n4085), .F(n4040) );
  MUX U1570 ( .IN0(n4069), .IN1(n4067), .SEL(n4068), .F(n4021) );
  MUX U1571 ( .IN0(n681), .IN1(n4010), .SEL(n4011), .F(n3964) );
  IV U1572 ( .A(n4012), .Z(n681) );
  MUX U1573 ( .IN0(n3906), .IN1(n3904), .SEL(n3905), .F(n3858) );
  MUX U1574 ( .IN0(n682), .IN1(n4469), .SEL(n3984), .F(n4448) );
  IV U1575 ( .A(n3982), .Z(n682) );
  MUX U1576 ( .IN0(n4912), .IN1(n4450), .SEL(n4451), .F(n4895) );
  MUX U1577 ( .IN0(n4420), .IN1(n4418), .SEL(n4419), .F(n4397) );
  MUX U1578 ( .IN0(n3887), .IN1(n3885), .SEL(n3886), .F(n3839) );
  MUX U1579 ( .IN0(n683), .IN1(n3828), .SEL(n3829), .F(n3782) );
  IV U1580 ( .A(n3830), .Z(n683) );
  MUX U1581 ( .IN0(n3724), .IN1(n3722), .SEL(n3723), .F(n3676) );
  MUX U1582 ( .IN0(n684), .IN1(n4385), .SEL(n3802), .F(n4364) );
  IV U1583 ( .A(n3800), .Z(n684) );
  MUX U1584 ( .IN0(n4844), .IN1(n4366), .SEL(n4367), .F(n4827) );
  MUX U1585 ( .IN0(n5294), .IN1(n5292), .SEL(n5293), .F(n5268) );
  MUX U1586 ( .IN0(n5426), .IN1(n5299), .SEL(n5301), .F(n5409) );
  MUX U1587 ( .IN0(n4336), .IN1(n4334), .SEL(n4335), .F(n4313) );
  MUX U1588 ( .IN0(n3705), .IN1(n3703), .SEL(n3704), .F(n3657) );
  MUX U1589 ( .IN0(n5037), .IN1(n4632), .SEL(n4634), .F(n5022) );
  MUX U1590 ( .IN0(n4627), .IN1(n4625), .SEL(n4626), .F(n4605) );
  MUX U1591 ( .IN0(n5494), .IN1(n5338), .SEL(n5339), .F(n685) );
  IV U1592 ( .A(n685), .Z(n5480) );
  MUX U1593 ( .IN0(n4170), .IN1(n4121), .SEL(n4122), .F(n686) );
  IV U1594 ( .A(n686), .Z(n4156) );
  MUX U1595 ( .IN0(n687), .IN1(n4153), .SEL(n4154), .F(n4139) );
  IV U1596 ( .A(n4155), .Z(n687) );
  MUX U1597 ( .IN0(n688), .IN1(n3647), .SEL(n3648), .F(n3604) );
  IV U1598 ( .A(n3649), .Z(n688) );
  MUX U1599 ( .IN0(n5577), .IN1(n5518), .SEL(n5519), .F(n689) );
  IV U1600 ( .A(n689), .Z(n5561) );
  MUX U1601 ( .IN0(n3550), .IN1(n3548), .SEL(n3549), .F(n3503) );
  MUX U1602 ( .IN0(n690), .IN1(n4301), .SEL(n3624), .F(n4281) );
  IV U1603 ( .A(n3622), .Z(n690) );
  MUX U1604 ( .IN0(n4778), .IN1(n4283), .SEL(n4284), .F(n4761) );
  MUX U1605 ( .IN0(n5605), .IN1(n5607), .SEL(n5606), .F(n5601) );
  MUX U1606 ( .IN0(n5208), .IN1(n5206), .SEL(n5207), .F(n5186) );
  MUX U1607 ( .IN0(n5371), .IN1(n5213), .SEL(n5215), .F(n5359) );
  MUX U1608 ( .IN0(n691), .IN1(n4125), .SEL(n4126), .F(n4103) );
  IV U1609 ( .A(n4127), .Z(n691) );
  MUX U1610 ( .IN0(n4253), .IN1(n4251), .SEL(n4252), .F(n4227) );
  MUX U1611 ( .IN0(n3532), .IN1(n3530), .SEL(n3531), .F(n3485) );
  XNOR U1612 ( .A(n5549), .B(A[5]), .Z(n5550) );
  XNOR U1613 ( .A(n5418), .B(A[9]), .Z(n5419) );
  MUX U1614 ( .IN0(n692), .IN1(n5332), .SEL(X[31]), .F(n5324) );
  IV U1615 ( .A(X[21]), .Z(n692) );
  XNOR U1616 ( .A(n5366), .B(A[13]), .Z(n5367) );
  XNOR U1617 ( .A(n4955), .B(A[17]), .Z(n4956) );
  XNOR U1618 ( .A(n4887), .B(A[21]), .Z(n4888) );
  AND U1619 ( .A(n5617), .B(A[0]), .Z(n3395) );
  MUX U1620 ( .IN0(n4543), .IN1(n4541), .SEL(n4542), .F(n4523) );
  MUX U1621 ( .IN0(n4990), .IN1(n4552), .SEL(n4554), .F(n4980) );
  MUX U1622 ( .IN0(n693), .IN1(n5596), .SEL(X[31]), .F(n5583) );
  IV U1623 ( .A(X[25]), .Z(n693) );
  XNOR U1624 ( .A(n4819), .B(A[25]), .Z(n4820) );
  MUX U1625 ( .IN0(n694), .IN1(n5614), .SEL(X[31]), .F(n5604) );
  IV U1626 ( .A(X[29]), .Z(n694) );
  MUX U1627 ( .IN0(A[3]), .IN1(n5600), .SEL(A[31]), .F(n3252) );
  MUX U1628 ( .IN0(n3369), .IN1(n3371), .SEL(n3370), .F(n3230) );
  MUX U1629 ( .IN0(n3345), .IN1(n3347), .SEL(n3346), .F(n3206) );
  MUX U1630 ( .IN0(X[20]), .IN1(n695), .SEL(X[31]), .F(n1404) );
  IV U1631 ( .A(n5331), .Z(n695) );
  MUX U1632 ( .IN0(X[16]), .IN1(n696), .SEL(X[31]), .F(n1766) );
  IV U1633 ( .A(n5511), .Z(n696) );
  MUX U1634 ( .IN0(X[8]), .IN1(n697), .SEL(X[31]), .F(n2541) );
  IV U1635 ( .A(n4190), .Z(n697) );
  MUX U1636 ( .IN0(X[12]), .IN1(n698), .SEL(X[31]), .F(n2112) );
  IV U1637 ( .A(n4203), .Z(n698) );
  MUX U1638 ( .IN0(X[4]), .IN1(n699), .SEL(X[31]), .F(n3050) );
  IV U1639 ( .A(n4709), .Z(n699) );
  XNOR U1640 ( .A(n4697), .B(n4694), .Z(n4695) );
  MUX U1641 ( .IN0(n700), .IN1(n3475), .SEL(n3476), .F(n3406) );
  IV U1642 ( .A(n3477), .Z(n700) );
  MUX U1643 ( .IN0(n701), .IN1(n5590), .SEL(X[31]), .F(n1019) );
  IV U1644 ( .A(X[27]), .Z(n701) );
  MUX U1645 ( .IN0(X[26]), .IN1(n702), .SEL(X[31]), .F(n1060) );
  IV U1646 ( .A(n5591), .Z(n702) );
  MUX U1647 ( .IN0(X[24]), .IN1(n703), .SEL(X[31]), .F(n1167) );
  IV U1648 ( .A(n5595), .Z(n703) );
  MUX U1649 ( .IN0(X[28]), .IN1(n704), .SEL(X[31]), .F(n992) );
  IV U1650 ( .A(n5613), .Z(n704) );
  MUX U1651 ( .IN0(n1485), .IN1(n1483), .SEL(n1484), .F(n1410) );
  MUX U1652 ( .IN0(n705), .IN1(n1532), .SEL(n1533), .F(n1454) );
  IV U1653 ( .A(n1534), .Z(n705) );
  MUX U1654 ( .IN0(n1526), .IN1(n1524), .SEL(n1525), .F(n1444) );
  MUX U1655 ( .IN0(X[18]), .IN1(n706), .SEL(X[31]), .F(n1582) );
  IV U1656 ( .A(n5506), .Z(n706) );
  MUX U1657 ( .IN0(n707), .IN1(n5512), .SEL(X[31]), .F(n1666) );
  IV U1658 ( .A(X[17]), .Z(n707) );
  MUX U1659 ( .IN0(n1863), .IN1(n1861), .SEL(n1862), .F(n1755) );
  MUX U1660 ( .IN0(n1836), .IN1(n1834), .SEL(n1835), .F(n1732) );
  MUX U1661 ( .IN0(n1879), .IN1(n1877), .SEL(n1878), .F(n1780) );
  MUX U1662 ( .IN0(n708), .IN1(n1885), .SEL(n1886), .F(n1788) );
  IV U1663 ( .A(n1887), .Z(n708) );
  XNOR U1664 ( .A(n4753), .B(A[29]), .Z(n4754) );
  MUX U1665 ( .IN0(n709), .IN1(n4186), .SEL(X[31]), .F(n2205) );
  IV U1666 ( .A(X[11]), .Z(n709) );
  MUX U1667 ( .IN0(X[10]), .IN1(n710), .SEL(X[31]), .F(n2311) );
  IV U1668 ( .A(n4185), .Z(n710) );
  MUX U1669 ( .IN0(n2435), .IN1(n2433), .SEL(n2434), .F(n2326) );
  MUX U1670 ( .IN0(X[6]), .IN1(n711), .SEL(X[31]), .F(n2801) );
  IV U1671 ( .A(n4714), .Z(n711) );
  MUX U1672 ( .IN0(n712), .IN1(n4710), .SEL(X[31]), .F(n2917) );
  IV U1673 ( .A(X[5]), .Z(n712) );
  MUX U1674 ( .IN0(n713), .IN1(n5144), .SEL(X[31]), .F(n3190) );
  IV U1675 ( .A(X[3]), .Z(n713) );
  MUX U1676 ( .IN0(X[2]), .IN1(n714), .SEL(X[31]), .F(n3327) );
  IV U1677 ( .A(n5143), .Z(n714) );
  MUX U1678 ( .IN0(n4219), .IN1(n715), .SEL(n3456), .F(n3328) );
  IV U1679 ( .A(n3455), .Z(n715) );
  MUX U1680 ( .IN0(X[22]), .IN1(n716), .SEL(X[31]), .F(n1276) );
  IV U1681 ( .A(n5337), .Z(n716) );
  MUX U1682 ( .IN0(n717), .IN1(n5336), .SEL(X[31]), .F(n1206) );
  IV U1683 ( .A(X[23]), .Z(n717) );
  MUX U1684 ( .IN0(n718), .IN1(n1293), .SEL(n1294), .F(n1225) );
  IV U1685 ( .A(n1295), .Z(n718) );
  MUX U1686 ( .IN0(n719), .IN1(n1593), .SEL(n1594), .F(n1514) );
  IV U1687 ( .A(n1595), .Z(n719) );
  MUX U1688 ( .IN0(n2011), .IN1(n2009), .SEL(n2010), .F(n720) );
  MUX U1689 ( .IN0(X[14]), .IN1(n721), .SEL(X[31]), .F(n1915) );
  IV U1690 ( .A(n4208), .Z(n721) );
  MUX U1691 ( .IN0(n722), .IN1(n1947), .SEL(n1948), .F(n1851) );
  IV U1692 ( .A(n1949), .Z(n722) );
  XNOR U1693 ( .A(n2170), .B(n2169), .Z(n2271) );
  XNOR U1694 ( .A(n2178), .B(n2177), .Z(n2279) );
  XNOR U1695 ( .A(n2129), .B(n2128), .Z(n2232) );
  XNOR U1696 ( .A(n2154), .B(n2153), .Z(n2255) );
  MUX U1697 ( .IN0(n723), .IN1(n2359), .SEL(n2360), .F(n2252) );
  IV U1698 ( .A(n2361), .Z(n723) );
  MUX U1699 ( .IN0(n724), .IN1(n2375), .SEL(n2376), .F(n2268) );
  IV U1700 ( .A(n2377), .Z(n724) );
  MUX U1701 ( .IN0(n2315), .IN1(n2419), .SEL(n2317), .F(n2207) );
  XNOR U1702 ( .A(n2475), .B(n2474), .Z(n2589) );
  XNOR U1703 ( .A(n2452), .B(n2451), .Z(n2566) );
  XNOR U1704 ( .A(n2491), .B(n2490), .Z(n2605) );
  XNOR U1705 ( .A(n2499), .B(n2498), .Z(n2613) );
  MUX U1706 ( .IN0(n725), .IN1(n2526), .SEL(n2527), .F(n2416) );
  IV U1707 ( .A(n2528), .Z(n725) );
  MUX U1708 ( .IN0(n726), .IN1(n4715), .SEL(X[31]), .F(n2675) );
  IV U1709 ( .A(X[7]), .Z(n726) );
  XNOR U1710 ( .A(n2860), .B(n2859), .Z(n2980) );
  XNOR U1711 ( .A(n2852), .B(n2851), .Z(n2972) );
  XNOR U1712 ( .A(n2813), .B(n2812), .Z(n2933) );
  XNOR U1713 ( .A(n2836), .B(n2835), .Z(n2956) );
  XNOR U1714 ( .A(n2773), .B(n2772), .Z(n2890) );
  XNOR U1715 ( .A(n2781), .B(n2780), .Z(n2898) );
  MUX U1716 ( .IN0(n727), .IN1(n3011), .SEL(n3012), .F(n2887) );
  IV U1717 ( .A(n3013), .Z(n727) );
  MUX U1718 ( .IN0(n728), .IN1(n3101), .SEL(n3102), .F(n2969) );
  IV U1719 ( .A(n3103), .Z(n728) );
  MUX U1720 ( .IN0(n729), .IN1(n3085), .SEL(n3086), .F(n2953) );
  IV U1721 ( .A(n3087), .Z(n729) );
  XNOR U1722 ( .A(n3249), .B(n3248), .Z(n3383) );
  XNOR U1723 ( .A(n3241), .B(n3240), .Z(n3375) );
  XNOR U1724 ( .A(n3202), .B(n3201), .Z(n3336) );
  XNOR U1725 ( .A(n3225), .B(n3224), .Z(n3359) );
  XNOR U1726 ( .A(n3149), .B(n3148), .Z(n3281) );
  XNOR U1727 ( .A(n3157), .B(n3156), .Z(n3289) );
  MUX U1728 ( .IN0(n3331), .IN1(n4718), .SEL(n3333), .F(n3192) );
  XNOR U1729 ( .A(n3173), .B(n3172), .Z(n3305) );
  MUX U1730 ( .IN0(X[30]), .IN1(n730), .SEL(X[31]), .F(n926) );
  IV U1731 ( .A(n5619), .Z(n730) );
  XNOR U1732 ( .A(n1069), .B(n1073), .Z(n1109) );
  NAND U1733 ( .A(n1274), .B(n1273), .Z(n1268) );
  MUX U1734 ( .IN0(n1277), .IN1(n1279), .SEL(n1278), .F(n1207) );
  XNOR U1735 ( .A(n1122), .B(n1121), .Z(n1176) );
  NAND U1736 ( .A(n1425), .B(n1426), .Z(n1420) );
  MUX U1737 ( .IN0(n731), .IN1(n1841), .SEL(n1842), .F(n1741) );
  IV U1738 ( .A(n1843), .Z(n731) );
  MUX U1739 ( .IN0(n732), .IN1(n4209), .SEL(X[31]), .F(n1814) );
  IV U1740 ( .A(X[15]), .Z(n732) );
  AND U1741 ( .A(n1895), .B(n1897), .Z(n1798) );
  ANDN U1742 ( .A(n2336), .B(n2337), .Z(n2228) );
  MUX U1743 ( .IN0(n3350), .IN1(n3348), .SEL(n3349), .F(n733) );
  IV U1744 ( .A(n733), .Z(n3209) );
  MUX U1745 ( .IN0(n734), .IN1(n3317), .SEL(n3318), .F(n3180) );
  IV U1746 ( .A(n3319), .Z(n734) );
  MUX U1747 ( .IN0(n921), .IN1(n919), .SEL(n920), .F(n899) );
  ANDN U1748 ( .A(n931), .B(n932), .Z(n902) );
  MUX U1749 ( .IN0(n735), .IN1(n1154), .SEL(n1155), .F(n1131) );
  IV U1750 ( .A(n1156), .Z(n735) );
  XNOR U1751 ( .A(n1816), .B(n1815), .Z(n1809) );
  XNOR U1752 ( .A(n2682), .B(n2677), .Z(n2791) );
  MUX U1753 ( .IN0(n896), .IN1(n898), .SEL(n897), .F(n736) );
  IV U1754 ( .A(n736), .Z(n881) );
  XNOR U1755 ( .A(n965), .B(n970), .Z(n966) );
  XNOR U1756 ( .A(n1090), .B(n1095), .Z(n1091) );
  XNOR U1757 ( .A(n1256), .B(n1261), .Z(n1257) );
  XOR U1758 ( .A(n1419), .B(n1418), .Z(n1400) );
  XOR U1759 ( .A(n1652), .B(n1651), .Z(n1634) );
  XOR U1760 ( .A(n1918), .B(n1917), .Z(n1997) );
  XOR U1761 ( .A(n2119), .B(n2118), .Z(n2194) );
  XOR U1762 ( .A(n2227), .B(n2226), .Z(n2300) );
  XOR U1763 ( .A(n2442), .B(n2441), .Z(n2515) );
  XOR U1764 ( .A(n2556), .B(n2555), .Z(n2634) );
  XOR U1765 ( .A(n2790), .B(n2789), .Z(n2876) );
  XOR U1766 ( .A(n2912), .B(n2911), .Z(n3000) );
  XOR U1767 ( .A(n3036), .B(n3035), .Z(n3130) );
  AND U1768 ( .A(Y0[0]), .B(n3134), .Z(n3259) );
  XNOR U1769 ( .A(n907), .B(n911), .Z(n909) );
  XNOR U1770 ( .A(n1008), .B(n1012), .Z(n1010) );
  XNOR U1771 ( .A(n1136), .B(n1139), .Z(n1138) );
  XNOR U1772 ( .A(n1326), .B(n1330), .Z(n1328) );
  XNOR U1773 ( .A(n1545), .B(n1549), .Z(n1547) );
  XNOR U1774 ( .A(n1801), .B(n1805), .Z(n1803) );
  XNOR U1775 ( .A(n2090), .B(n2094), .Z(n2092) );
  XNOR U1776 ( .A(n2404), .B(n2408), .Z(n2406) );
  XNOR U1777 ( .A(n2751), .B(n2755), .Z(n2753) );
  MUX U1778 ( .IN0(n737), .IN1(n842), .SEL(n848), .F(n845) );
  ANDN U1779 ( .A(n738), .B(n[0]), .Z(n372) );
  AND U1780 ( .A(N8), .B(n738), .Z(n371) );
  AND U1781 ( .A(N9), .B(n738), .Z(n370) );
  AND U1782 ( .A(N10), .B(n738), .Z(n369) );
  AND U1783 ( .A(N11), .B(n738), .Z(n368) );
  AND U1784 ( .A(N12), .B(n738), .Z(n367) );
  AND U1785 ( .A(N13), .B(n738), .Z(n366) );
  AND U1786 ( .A(N14), .B(n738), .Z(n365) );
  AND U1787 ( .A(N15), .B(n738), .Z(n364) );
  AND U1788 ( .A(n738), .B(n739), .Z(n363) );
  XOR U1789 ( .A(n[9]), .B(\add_25/carry[9] ), .Z(n739) );
  ANDN U1790 ( .A(n740), .B(rst), .Z(n738) );
  NAND U1791 ( .A(n741), .B(n742), .Z(n740) );
  AND U1792 ( .A(n743), .B(n744), .Z(n742) );
  AND U1793 ( .A(n[1]), .B(n745), .Z(n744) );
  AND U1794 ( .A(n746), .B(n[0]), .Z(n745) );
  AND U1795 ( .A(n[5]), .B(n[2]), .Z(n743) );
  AND U1796 ( .A(n747), .B(n748), .Z(n741) );
  AND U1797 ( .A(n[6]), .B(n[7]), .Z(n748) );
  AND U1798 ( .A(n[8]), .B(n[9]), .Z(n747) );
  NAND U1799 ( .A(n749), .B(n750), .Z(n362) );
  NAND U1800 ( .A(n751), .B(n752), .Z(n750) );
  NAND U1801 ( .A(Y0[0]), .B(rst), .Z(n749) );
  NAND U1802 ( .A(n753), .B(n754), .Z(n361) );
  NAND U1803 ( .A(n755), .B(n752), .Z(n754) );
  NAND U1804 ( .A(Y0[1]), .B(rst), .Z(n753) );
  NAND U1805 ( .A(n756), .B(n757), .Z(n360) );
  NAND U1806 ( .A(n758), .B(n752), .Z(n757) );
  NAND U1807 ( .A(Y0[2]), .B(rst), .Z(n756) );
  NAND U1808 ( .A(n759), .B(n760), .Z(n359) );
  NAND U1809 ( .A(n761), .B(n752), .Z(n760) );
  NAND U1810 ( .A(Y0[3]), .B(rst), .Z(n759) );
  NAND U1811 ( .A(n762), .B(n763), .Z(n358) );
  NAND U1812 ( .A(n764), .B(n752), .Z(n763) );
  NAND U1813 ( .A(Y0[4]), .B(rst), .Z(n762) );
  NAND U1814 ( .A(n765), .B(n766), .Z(n357) );
  NAND U1815 ( .A(n767), .B(n752), .Z(n766) );
  NAND U1816 ( .A(rst), .B(Y0[5]), .Z(n765) );
  NAND U1817 ( .A(n768), .B(n769), .Z(n356) );
  NAND U1818 ( .A(n770), .B(n752), .Z(n769) );
  NAND U1819 ( .A(rst), .B(Y0[6]), .Z(n768) );
  NAND U1820 ( .A(n771), .B(n772), .Z(n355) );
  NAND U1821 ( .A(n773), .B(n752), .Z(n772) );
  NAND U1822 ( .A(rst), .B(Y0[7]), .Z(n771) );
  NAND U1823 ( .A(n774), .B(n775), .Z(n354) );
  NAND U1824 ( .A(n776), .B(n752), .Z(n775) );
  NAND U1825 ( .A(rst), .B(Y0[8]), .Z(n774) );
  NAND U1826 ( .A(n777), .B(n778), .Z(n353) );
  NAND U1827 ( .A(n779), .B(n752), .Z(n778) );
  NAND U1828 ( .A(rst), .B(Y0[9]), .Z(n777) );
  NAND U1829 ( .A(n780), .B(n781), .Z(n352) );
  NAND U1830 ( .A(n782), .B(n752), .Z(n781) );
  NAND U1831 ( .A(rst), .B(Y0[10]), .Z(n780) );
  NAND U1832 ( .A(n783), .B(n784), .Z(n351) );
  NAND U1833 ( .A(n785), .B(n752), .Z(n784) );
  NAND U1834 ( .A(rst), .B(Y0[11]), .Z(n783) );
  NAND U1835 ( .A(n786), .B(n787), .Z(n350) );
  NAND U1836 ( .A(n788), .B(n752), .Z(n787) );
  NAND U1837 ( .A(rst), .B(Y0[12]), .Z(n786) );
  NAND U1838 ( .A(n789), .B(n790), .Z(n349) );
  NAND U1839 ( .A(n791), .B(n752), .Z(n790) );
  NAND U1840 ( .A(rst), .B(Y0[13]), .Z(n789) );
  NAND U1841 ( .A(n792), .B(n793), .Z(n348) );
  NAND U1842 ( .A(n794), .B(n752), .Z(n793) );
  NAND U1843 ( .A(rst), .B(Y0[14]), .Z(n792) );
  NAND U1844 ( .A(n795), .B(n796), .Z(n347) );
  NAND U1845 ( .A(n797), .B(n752), .Z(n796) );
  NAND U1846 ( .A(rst), .B(Y0[15]), .Z(n795) );
  NAND U1847 ( .A(n798), .B(n799), .Z(n346) );
  NAND U1848 ( .A(n800), .B(n752), .Z(n799) );
  NAND U1849 ( .A(rst), .B(Y0[16]), .Z(n798) );
  NAND U1850 ( .A(n801), .B(n802), .Z(n345) );
  NAND U1851 ( .A(n803), .B(n752), .Z(n802) );
  NAND U1852 ( .A(rst), .B(Y0[17]), .Z(n801) );
  NAND U1853 ( .A(n804), .B(n805), .Z(n344) );
  NAND U1854 ( .A(n806), .B(n752), .Z(n805) );
  NAND U1855 ( .A(rst), .B(Y0[18]), .Z(n804) );
  NAND U1856 ( .A(n807), .B(n808), .Z(n343) );
  NAND U1857 ( .A(n809), .B(n752), .Z(n808) );
  NAND U1858 ( .A(rst), .B(Y0[19]), .Z(n807) );
  NAND U1859 ( .A(n810), .B(n811), .Z(n342) );
  NAND U1860 ( .A(n812), .B(n752), .Z(n811) );
  NAND U1861 ( .A(rst), .B(Y0[20]), .Z(n810) );
  NAND U1862 ( .A(n813), .B(n814), .Z(n341) );
  NAND U1863 ( .A(n815), .B(n752), .Z(n814) );
  NAND U1864 ( .A(rst), .B(Y0[21]), .Z(n813) );
  NAND U1865 ( .A(n816), .B(n817), .Z(n340) );
  NAND U1866 ( .A(n818), .B(n752), .Z(n817) );
  NAND U1867 ( .A(rst), .B(Y0[22]), .Z(n816) );
  NAND U1868 ( .A(n819), .B(n820), .Z(n339) );
  NAND U1869 ( .A(n821), .B(n752), .Z(n820) );
  NAND U1870 ( .A(rst), .B(Y0[23]), .Z(n819) );
  NAND U1871 ( .A(n822), .B(n823), .Z(n338) );
  NAND U1872 ( .A(n824), .B(n752), .Z(n823) );
  NAND U1873 ( .A(rst), .B(Y0[24]), .Z(n822) );
  NAND U1874 ( .A(n825), .B(n826), .Z(n337) );
  NAND U1875 ( .A(n827), .B(n752), .Z(n826) );
  NAND U1876 ( .A(rst), .B(Y0[25]), .Z(n825) );
  NAND U1877 ( .A(n828), .B(n829), .Z(n336) );
  NAND U1878 ( .A(n830), .B(n752), .Z(n829) );
  NAND U1879 ( .A(rst), .B(Y0[26]), .Z(n828) );
  NAND U1880 ( .A(n831), .B(n832), .Z(n335) );
  NAND U1881 ( .A(n833), .B(n752), .Z(n832) );
  NAND U1882 ( .A(rst), .B(Y0[27]), .Z(n831) );
  NAND U1883 ( .A(n834), .B(n835), .Z(n334) );
  NAND U1884 ( .A(n836), .B(n752), .Z(n835) );
  NAND U1885 ( .A(rst), .B(Y0[28]), .Z(n834) );
  NAND U1886 ( .A(n837), .B(n838), .Z(n333) );
  NAND U1887 ( .A(n839), .B(n752), .Z(n838) );
  NAND U1888 ( .A(rst), .B(Y0[29]), .Z(n837) );
  NAND U1889 ( .A(n840), .B(n841), .Z(n332) );
  NAND U1890 ( .A(n842), .B(n752), .Z(n841) );
  NAND U1891 ( .A(rst), .B(Y0[30]), .Z(n840) );
  NAND U1892 ( .A(n843), .B(n844), .Z(n331) );
  NAND U1893 ( .A(n845), .B(n752), .Z(n844) );
  NOR U1894 ( .A(rst), .B(n846), .Z(n752) );
  NAND U1895 ( .A(Y0[31]), .B(rst), .Z(n843) );
  MUX U1896 ( .IN0(Y[31]), .IN1(n845), .SEL(n847), .F(n330) );
  XNOR U1897 ( .A(Y0[31]), .B(n849), .Z(n848) );
  AND U1898 ( .A(n852), .B(n853), .Z(n851) );
  XNOR U1899 ( .A(Y0[31]), .B(n854), .Z(n853) );
  MUX U1900 ( .IN0(Y[30]), .IN1(n842), .SEL(n847), .F(n329) );
  XOR U1901 ( .A(n852), .B(Y0[31]), .Z(n842) );
  XOR U1902 ( .A(n854), .B(n849), .Z(n852) );
  XOR U1903 ( .A(n855), .B(n856), .Z(n849) );
  XOR U1904 ( .A(n857), .B(n858), .Z(n856) );
  AND U1905 ( .A(n859), .B(n860), .Z(n858) );
  XOR U1906 ( .A(n867), .B(n865), .Z(n855) );
  XOR U1907 ( .A(n868), .B(n869), .Z(n867) );
  XOR U1908 ( .A(n870), .B(n871), .Z(n869) );
  XOR U1909 ( .A(n875), .B(n876), .Z(n870) );
  ANDN U1910 ( .A(n877), .B(n878), .Z(n876) );
  XOR U1911 ( .A(n882), .B(n883), .Z(n868) );
  XOR U1912 ( .A(n872), .B(n874), .Z(n883) );
  XOR U1913 ( .A(n881), .B(n878), .Z(n882) );
  IV U1914 ( .A(n850), .Z(n854) );
  MUX U1915 ( .IN0(Y[29]), .IN1(n839), .SEL(n847), .F(n328) );
  XOR U1916 ( .A(n885), .B(Y0[30]), .Z(n839) );
  XNOR U1917 ( .A(n886), .B(n887), .Z(n885) );
  AND U1918 ( .A(n859), .B(n889), .Z(n888) );
  XNOR U1919 ( .A(n863), .B(n887), .Z(n889) );
  XOR U1920 ( .A(n861), .B(n887), .Z(n863) );
  XNOR U1921 ( .A(n866), .B(n864), .Z(n887) );
  IV U1922 ( .A(n865), .Z(n864) );
  XNOR U1923 ( .A(n872), .B(n873), .Z(n866) );
  XNOR U1924 ( .A(n874), .B(n877), .Z(n873) );
  XNOR U1925 ( .A(n878), .B(n893), .Z(n877) );
  XOR U1926 ( .A(n879), .B(n880), .Z(n893) );
  NAND U1927 ( .A(n894), .B(n895), .Z(n880) );
  IV U1928 ( .A(n881), .Z(n879) );
  IV U1929 ( .A(n862), .Z(n861) );
  MUX U1930 ( .IN0(Y[28]), .IN1(n836), .SEL(n847), .F(n327) );
  XOR U1931 ( .A(n908), .B(Y0[29]), .Z(n836) );
  XNOR U1932 ( .A(n909), .B(n910), .Z(n908) );
  AND U1933 ( .A(n859), .B(n912), .Z(n911) );
  XNOR U1934 ( .A(n906), .B(n910), .Z(n912) );
  XNOR U1935 ( .A(n892), .B(n891), .Z(n910) );
  IV U1936 ( .A(n890), .Z(n891) );
  XOR U1937 ( .A(n904), .B(n903), .Z(n892) );
  XOR U1938 ( .A(n902), .B(n916), .Z(n903) );
  XNOR U1939 ( .A(n901), .B(n900), .Z(n916) );
  XNOR U1940 ( .A(n917), .B(n918), .Z(n900) );
  IV U1941 ( .A(n899), .Z(n918) );
  XNOR U1942 ( .A(n897), .B(n898), .Z(n901) );
  NAND U1943 ( .A(n924), .B(n895), .Z(n898) );
  XNOR U1944 ( .A(n896), .B(n925), .Z(n897) );
  ANDN U1945 ( .A(n926), .B(n927), .Z(n925) );
  MUX U1946 ( .IN0(Y[27]), .IN1(n833), .SEL(n847), .F(n326) );
  XOR U1947 ( .A(n937), .B(Y0[28]), .Z(n833) );
  XNOR U1948 ( .A(n938), .B(n939), .Z(n937) );
  AND U1949 ( .A(n859), .B(n941), .Z(n940) );
  XNOR U1950 ( .A(n935), .B(n939), .Z(n941) );
  XNOR U1951 ( .A(n915), .B(n914), .Z(n939) );
  IV U1952 ( .A(n913), .Z(n914) );
  XOR U1953 ( .A(n933), .B(n932), .Z(n915) );
  XOR U1954 ( .A(n931), .B(n945), .Z(n932) );
  XNOR U1955 ( .A(n921), .B(n920), .Z(n945) );
  XOR U1956 ( .A(n950), .B(n922), .Z(n946) );
  AND U1957 ( .A(n951), .B(n894), .Z(n922) );
  IV U1958 ( .A(n919), .Z(n950) );
  XNOR U1959 ( .A(n929), .B(n930), .Z(n921) );
  NAND U1960 ( .A(n955), .B(n895), .Z(n930) );
  XNOR U1961 ( .A(n928), .B(n956), .Z(n929) );
  ANDN U1962 ( .A(n926), .B(n957), .Z(n956) );
  MUX U1963 ( .IN0(Y[26]), .IN1(n830), .SEL(n847), .F(n325) );
  XOR U1964 ( .A(n968), .B(Y0[27]), .Z(n830) );
  XNOR U1965 ( .A(n969), .B(n970), .Z(n968) );
  AND U1966 ( .A(n859), .B(n972), .Z(n971) );
  XNOR U1967 ( .A(n966), .B(n970), .Z(n972) );
  XNOR U1968 ( .A(n944), .B(n943), .Z(n970) );
  IV U1969 ( .A(n942), .Z(n943) );
  XNOR U1970 ( .A(n964), .B(n976), .Z(n944) );
  XOR U1971 ( .A(n963), .B(n962), .Z(n976) );
  XOR U1972 ( .A(n977), .B(n978), .Z(n962) );
  XOR U1973 ( .A(n979), .B(n980), .Z(n978) );
  XOR U1974 ( .A(n981), .B(n982), .Z(n980) );
  XNOR U1975 ( .A(n954), .B(n953), .Z(n963) );
  XOR U1976 ( .A(n990), .B(n948), .Z(n953) );
  XNOR U1977 ( .A(n947), .B(n991), .Z(n948) );
  ANDN U1978 ( .A(n992), .B(n927), .Z(n991) );
  AND U1979 ( .A(n924), .B(n951), .Z(n949) );
  XNOR U1980 ( .A(n959), .B(n960), .Z(n954) );
  NAND U1981 ( .A(n999), .B(n895), .Z(n960) );
  XNOR U1982 ( .A(n958), .B(n1000), .Z(n959) );
  ANDN U1983 ( .A(n926), .B(n1001), .Z(n1000) );
  MUX U1984 ( .IN0(Y[25]), .IN1(n827), .SEL(n847), .F(n324) );
  XOR U1985 ( .A(n1009), .B(Y0[26]), .Z(n827) );
  XNOR U1986 ( .A(n1010), .B(n1011), .Z(n1009) );
  AND U1987 ( .A(n859), .B(n1013), .Z(n1012) );
  XNOR U1988 ( .A(n1007), .B(n1011), .Z(n1013) );
  XNOR U1989 ( .A(n975), .B(n974), .Z(n1011) );
  IV U1990 ( .A(n973), .Z(n974) );
  XOR U1991 ( .A(n1005), .B(n1017), .Z(n975) );
  XNOR U1992 ( .A(n989), .B(n988), .Z(n1017) );
  XOR U1993 ( .A(n1018), .B(n983), .Z(n988) );
  XOR U1994 ( .A(n984), .B(n985), .Z(n983) );
  NANDN U1995 ( .B(n1019), .A(n894), .Z(n985) );
  IV U1996 ( .A(n986), .Z(n984) );
  XOR U1997 ( .A(n979), .B(n987), .Z(n1018) );
  XNOR U1998 ( .A(n998), .B(n997), .Z(n989) );
  XOR U1999 ( .A(n1029), .B(n994), .Z(n997) );
  XNOR U2000 ( .A(n993), .B(n1030), .Z(n994) );
  ANDN U2001 ( .A(n992), .B(n957), .Z(n1030) );
  XOR U2002 ( .A(n1031), .B(n1032), .Z(n993) );
  AND U2003 ( .A(n1033), .B(n1034), .Z(n1032) );
  XNOR U2004 ( .A(n1035), .B(n1031), .Z(n1034) );
  AND U2005 ( .A(n955), .B(n951), .Z(n995) );
  XNOR U2006 ( .A(n1003), .B(n1004), .Z(n998) );
  NAND U2007 ( .A(n1039), .B(n895), .Z(n1004) );
  XNOR U2008 ( .A(n1002), .B(n1040), .Z(n1003) );
  ANDN U2009 ( .A(n926), .B(n1041), .Z(n1040) );
  MUX U2010 ( .IN0(Y[24]), .IN1(n824), .SEL(n847), .F(n323) );
  XOR U2011 ( .A(n1049), .B(Y0[25]), .Z(n824) );
  XNOR U2012 ( .A(n1050), .B(n1051), .Z(n1049) );
  AND U2013 ( .A(n859), .B(n1053), .Z(n1052) );
  XNOR U2014 ( .A(n1047), .B(n1051), .Z(n1053) );
  XNOR U2015 ( .A(n1016), .B(n1015), .Z(n1051) );
  IV U2016 ( .A(n1014), .Z(n1015) );
  XOR U2017 ( .A(n1045), .B(n1057), .Z(n1016) );
  XNOR U2018 ( .A(n1025), .B(n1024), .Z(n1057) );
  XOR U2019 ( .A(n1058), .B(n1028), .Z(n1024) );
  XNOR U2020 ( .A(n1021), .B(n1022), .Z(n1028) );
  NANDN U2021 ( .B(n1019), .A(n924), .Z(n1022) );
  XNOR U2022 ( .A(n1020), .B(n1059), .Z(n1021) );
  ANDN U2023 ( .A(n1060), .B(n927), .Z(n1059) );
  XNOR U2024 ( .A(n1027), .B(n1023), .Z(n1058) );
  XNOR U2025 ( .A(n1067), .B(n1068), .Z(n1027) );
  IV U2026 ( .A(n1026), .Z(n1068) );
  XNOR U2027 ( .A(n1038), .B(n1037), .Z(n1025) );
  XOR U2028 ( .A(n1075), .B(n1033), .Z(n1037) );
  XNOR U2029 ( .A(n1031), .B(n1076), .Z(n1033) );
  ANDN U2030 ( .A(n992), .B(n1001), .Z(n1076) );
  AND U2031 ( .A(n999), .B(n951), .Z(n1035) );
  XNOR U2032 ( .A(n1043), .B(n1044), .Z(n1038) );
  NAND U2033 ( .A(n1083), .B(n895), .Z(n1044) );
  XNOR U2034 ( .A(n1042), .B(n1084), .Z(n1043) );
  ANDN U2035 ( .A(n926), .B(n1085), .Z(n1084) );
  MUX U2036 ( .IN0(Y[23]), .IN1(n821), .SEL(n847), .F(n322) );
  XOR U2037 ( .A(n1093), .B(Y0[24]), .Z(n821) );
  XNOR U2038 ( .A(n1094), .B(n1095), .Z(n1093) );
  AND U2039 ( .A(n859), .B(n1097), .Z(n1096) );
  XNOR U2040 ( .A(n1091), .B(n1095), .Z(n1097) );
  XNOR U2041 ( .A(n1056), .B(n1055), .Z(n1095) );
  IV U2042 ( .A(n1054), .Z(n1055) );
  XOR U2043 ( .A(n1089), .B(n1100), .Z(n1056) );
  XNOR U2044 ( .A(n1066), .B(n1065), .Z(n1100) );
  XOR U2045 ( .A(n1101), .B(n1071), .Z(n1065) );
  XNOR U2046 ( .A(n1062), .B(n1063), .Z(n1071) );
  NANDN U2047 ( .B(n1019), .A(n955), .Z(n1063) );
  XNOR U2048 ( .A(n1061), .B(n1102), .Z(n1062) );
  ANDN U2049 ( .A(n1060), .B(n957), .Z(n1102) );
  XNOR U2050 ( .A(n1070), .B(n1064), .Z(n1101) );
  XNOR U2051 ( .A(n1109), .B(n1072), .Z(n1070) );
  IV U2052 ( .A(n1074), .Z(n1072) );
  AND U2053 ( .A(n1113), .B(n894), .Z(n1073) );
  XNOR U2054 ( .A(n1082), .B(n1081), .Z(n1066) );
  XOR U2055 ( .A(n1117), .B(n1078), .Z(n1081) );
  XNOR U2056 ( .A(n1077), .B(n1118), .Z(n1078) );
  ANDN U2057 ( .A(n992), .B(n1041), .Z(n1118) );
  AND U2058 ( .A(n1039), .B(n951), .Z(n1079) );
  XNOR U2059 ( .A(n1087), .B(n1088), .Z(n1082) );
  NAND U2060 ( .A(n1125), .B(n895), .Z(n1088) );
  XNOR U2061 ( .A(n1086), .B(n1126), .Z(n1087) );
  ANDN U2062 ( .A(n926), .B(n1127), .Z(n1126) );
  MUX U2063 ( .IN0(Y[22]), .IN1(n818), .SEL(n847), .F(n321) );
  XOR U2064 ( .A(n1137), .B(Y0[23]), .Z(n818) );
  XNOR U2065 ( .A(n1138), .B(n1099), .Z(n1137) );
  AND U2066 ( .A(n859), .B(n1140), .Z(n1139) );
  XNOR U2067 ( .A(n1135), .B(n1099), .Z(n1140) );
  XOR U2068 ( .A(n1098), .B(n1141), .Z(n1099) );
  XNOR U2069 ( .A(n1133), .B(n1132), .Z(n1141) );
  XOR U2070 ( .A(n1142), .B(n1143), .Z(n1132) );
  XOR U2071 ( .A(n1144), .B(n1145), .Z(n1143) );
  XOR U2072 ( .A(n1148), .B(n1149), .Z(n1144) );
  ANDN U2073 ( .A(n1147), .B(n1150), .Z(n1149) );
  XNOR U2074 ( .A(n1153), .B(n1131), .Z(n1142) );
  XOR U2075 ( .A(n1152), .B(n1150), .Z(n1153) );
  XNOR U2076 ( .A(n1108), .B(n1107), .Z(n1133) );
  XOR U2077 ( .A(n1157), .B(n1116), .Z(n1107) );
  XNOR U2078 ( .A(n1104), .B(n1105), .Z(n1116) );
  NANDN U2079 ( .B(n1019), .A(n999), .Z(n1105) );
  XNOR U2080 ( .A(n1103), .B(n1158), .Z(n1104) );
  ANDN U2081 ( .A(n1060), .B(n1001), .Z(n1158) );
  XNOR U2082 ( .A(n1115), .B(n1106), .Z(n1157) );
  XOR U2083 ( .A(n1165), .B(n1111), .Z(n1115) );
  XNOR U2084 ( .A(n1110), .B(n1166), .Z(n1111) );
  ANDN U2085 ( .A(n1167), .B(n927), .Z(n1166) );
  XOR U2086 ( .A(n1168), .B(n1169), .Z(n1110) );
  AND U2087 ( .A(n1170), .B(n1171), .Z(n1169) );
  XNOR U2088 ( .A(n1172), .B(n1168), .Z(n1171) );
  AND U2089 ( .A(n924), .B(n1113), .Z(n1112) );
  XNOR U2090 ( .A(n1124), .B(n1123), .Z(n1108) );
  XOR U2091 ( .A(n1176), .B(n1120), .Z(n1123) );
  XNOR U2092 ( .A(n1119), .B(n1177), .Z(n1120) );
  ANDN U2093 ( .A(n992), .B(n1085), .Z(n1177) );
  AND U2094 ( .A(n1083), .B(n951), .Z(n1121) );
  XNOR U2095 ( .A(n1129), .B(n1130), .Z(n1124) );
  NAND U2096 ( .A(n1184), .B(n895), .Z(n1130) );
  XNOR U2097 ( .A(n1128), .B(n1185), .Z(n1129) );
  ANDN U2098 ( .A(n926), .B(n1186), .Z(n1185) );
  MUX U2099 ( .IN0(Y[21]), .IN1(n815), .SEL(n847), .F(n320) );
  XOR U2100 ( .A(n1196), .B(Y0[22]), .Z(n815) );
  XNOR U2101 ( .A(n1197), .B(n1198), .Z(n1196) );
  AND U2102 ( .A(n859), .B(n1200), .Z(n1199) );
  XNOR U2103 ( .A(n1194), .B(n1198), .Z(n1200) );
  XNOR U2104 ( .A(n1192), .B(n1191), .Z(n1198) );
  IV U2105 ( .A(n1190), .Z(n1191) );
  XNOR U2106 ( .A(n1156), .B(n1155), .Z(n1192) );
  XOR U2107 ( .A(n1204), .B(n1147), .Z(n1155) );
  XNOR U2108 ( .A(n1150), .B(n1205), .Z(n1147) );
  NANDN U2109 ( .B(n1206), .A(n894), .Z(n1151) );
  XOR U2110 ( .A(n1146), .B(n1154), .Z(n1204) );
  XNOR U2111 ( .A(n1164), .B(n1163), .Z(n1156) );
  XOR U2112 ( .A(n1218), .B(n1175), .Z(n1163) );
  XNOR U2113 ( .A(n1160), .B(n1161), .Z(n1175) );
  NANDN U2114 ( .B(n1019), .A(n1039), .Z(n1161) );
  XNOR U2115 ( .A(n1159), .B(n1219), .Z(n1160) );
  ANDN U2116 ( .A(n1060), .B(n1041), .Z(n1219) );
  XOR U2117 ( .A(n1220), .B(n1221), .Z(n1159) );
  AND U2118 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U2119 ( .A(n1224), .B(n1220), .Z(n1223) );
  XNOR U2120 ( .A(n1174), .B(n1162), .Z(n1218) );
  XOR U2121 ( .A(n1228), .B(n1170), .Z(n1174) );
  XNOR U2122 ( .A(n1168), .B(n1229), .Z(n1170) );
  ANDN U2123 ( .A(n1167), .B(n957), .Z(n1229) );
  XOR U2124 ( .A(n1230), .B(n1231), .Z(n1168) );
  AND U2125 ( .A(n1232), .B(n1233), .Z(n1231) );
  XNOR U2126 ( .A(n1234), .B(n1230), .Z(n1233) );
  AND U2127 ( .A(n955), .B(n1113), .Z(n1172) );
  XNOR U2128 ( .A(n1183), .B(n1182), .Z(n1164) );
  XOR U2129 ( .A(n1238), .B(n1179), .Z(n1182) );
  XNOR U2130 ( .A(n1178), .B(n1239), .Z(n1179) );
  ANDN U2131 ( .A(n992), .B(n1127), .Z(n1239) );
  XOR U2132 ( .A(n1240), .B(n1241), .Z(n1178) );
  AND U2133 ( .A(n1242), .B(n1243), .Z(n1241) );
  XNOR U2134 ( .A(n1244), .B(n1240), .Z(n1243) );
  AND U2135 ( .A(n1125), .B(n951), .Z(n1180) );
  XNOR U2136 ( .A(n1188), .B(n1189), .Z(n1183) );
  NAND U2137 ( .A(n1248), .B(n895), .Z(n1189) );
  XNOR U2138 ( .A(n1187), .B(n1249), .Z(n1188) );
  ANDN U2139 ( .A(n926), .B(n1250), .Z(n1249) );
  XOR U2140 ( .A(n1251), .B(n1252), .Z(n1187) );
  AND U2141 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U2142 ( .A(n1255), .B(n1251), .Z(n1254) );
  MUX U2143 ( .IN0(Y[20]), .IN1(n812), .SEL(n847), .F(n319) );
  XOR U2144 ( .A(n1259), .B(Y0[21]), .Z(n812) );
  XNOR U2145 ( .A(n1260), .B(n1261), .Z(n1259) );
  AND U2146 ( .A(n859), .B(n1263), .Z(n1262) );
  XNOR U2147 ( .A(n1257), .B(n1261), .Z(n1263) );
  XNOR U2148 ( .A(n1203), .B(n1202), .Z(n1261) );
  IV U2149 ( .A(n1201), .Z(n1202) );
  XNOR U2150 ( .A(n1215), .B(n1214), .Z(n1203) );
  XOR U2151 ( .A(n1267), .B(n1217), .Z(n1214) );
  XNOR U2152 ( .A(n1212), .B(n1211), .Z(n1217) );
  XNOR U2153 ( .A(n1268), .B(n1269), .Z(n1211) );
  IV U2154 ( .A(n1210), .Z(n1269) );
  XNOR U2155 ( .A(n1208), .B(n1209), .Z(n1212) );
  NANDN U2156 ( .B(n1206), .A(n924), .Z(n1209) );
  XNOR U2157 ( .A(n1207), .B(n1275), .Z(n1208) );
  ANDN U2158 ( .A(n1276), .B(n927), .Z(n1275) );
  XNOR U2159 ( .A(n1227), .B(n1226), .Z(n1215) );
  XOR U2160 ( .A(n1286), .B(n1237), .Z(n1226) );
  XNOR U2161 ( .A(n1222), .B(n1224), .Z(n1237) );
  NANDN U2162 ( .B(n1019), .A(n1083), .Z(n1224) );
  XNOR U2163 ( .A(n1220), .B(n1287), .Z(n1222) );
  ANDN U2164 ( .A(n1060), .B(n1085), .Z(n1287) );
  XOR U2165 ( .A(n1288), .B(n1289), .Z(n1220) );
  AND U2166 ( .A(n1290), .B(n1291), .Z(n1289) );
  XOR U2167 ( .A(n1292), .B(n1288), .Z(n1291) );
  XNOR U2168 ( .A(n1236), .B(n1225), .Z(n1286) );
  XOR U2169 ( .A(n1296), .B(n1232), .Z(n1236) );
  XNOR U2170 ( .A(n1230), .B(n1297), .Z(n1232) );
  ANDN U2171 ( .A(n1167), .B(n1001), .Z(n1297) );
  XOR U2172 ( .A(n1298), .B(n1299), .Z(n1230) );
  AND U2173 ( .A(n1300), .B(n1301), .Z(n1299) );
  XNOR U2174 ( .A(n1302), .B(n1298), .Z(n1301) );
  AND U2175 ( .A(n999), .B(n1113), .Z(n1234) );
  XNOR U2176 ( .A(n1247), .B(n1246), .Z(n1227) );
  XOR U2177 ( .A(n1306), .B(n1242), .Z(n1246) );
  XNOR U2178 ( .A(n1240), .B(n1307), .Z(n1242) );
  ANDN U2179 ( .A(n992), .B(n1186), .Z(n1307) );
  XOR U2180 ( .A(n1308), .B(n1309), .Z(n1240) );
  AND U2181 ( .A(n1310), .B(n1311), .Z(n1309) );
  XNOR U2182 ( .A(n1312), .B(n1308), .Z(n1311) );
  AND U2183 ( .A(n1184), .B(n951), .Z(n1244) );
  XNOR U2184 ( .A(n1253), .B(n1255), .Z(n1247) );
  NAND U2185 ( .A(n1316), .B(n895), .Z(n1255) );
  XNOR U2186 ( .A(n1251), .B(n1317), .Z(n1253) );
  ANDN U2187 ( .A(n926), .B(n1318), .Z(n1317) );
  XOR U2188 ( .A(n1319), .B(n1320), .Z(n1251) );
  AND U2189 ( .A(n1321), .B(n1322), .Z(n1320) );
  XOR U2190 ( .A(n1323), .B(n1319), .Z(n1322) );
  MUX U2191 ( .IN0(Y[19]), .IN1(n809), .SEL(n847), .F(n318) );
  XOR U2192 ( .A(n1327), .B(Y0[20]), .Z(n809) );
  XNOR U2193 ( .A(n1328), .B(n1329), .Z(n1327) );
  AND U2194 ( .A(n859), .B(n1331), .Z(n1330) );
  XNOR U2195 ( .A(n1325), .B(n1329), .Z(n1331) );
  XNOR U2196 ( .A(n1266), .B(n1265), .Z(n1329) );
  IV U2197 ( .A(n1264), .Z(n1265) );
  XNOR U2198 ( .A(n1282), .B(n1281), .Z(n1266) );
  XOR U2199 ( .A(n1335), .B(n1285), .Z(n1281) );
  XNOR U2200 ( .A(n1272), .B(n1271), .Z(n1285) );
  XOR U2201 ( .A(n1340), .B(n1273), .Z(n1336) );
  AND U2202 ( .A(n1341), .B(n894), .Z(n1273) );
  IV U2203 ( .A(n1270), .Z(n1340) );
  XNOR U2204 ( .A(n1278), .B(n1279), .Z(n1272) );
  NANDN U2205 ( .B(n1206), .A(n955), .Z(n1279) );
  XNOR U2206 ( .A(n1277), .B(n1345), .Z(n1278) );
  ANDN U2207 ( .A(n1276), .B(n957), .Z(n1345) );
  XNOR U2208 ( .A(n1284), .B(n1280), .Z(n1335) );
  IV U2209 ( .A(n1283), .Z(n1284) );
  XNOR U2210 ( .A(n1295), .B(n1294), .Z(n1282) );
  XOR U2211 ( .A(n1355), .B(n1305), .Z(n1294) );
  XNOR U2212 ( .A(n1290), .B(n1292), .Z(n1305) );
  NANDN U2213 ( .B(n1019), .A(n1125), .Z(n1292) );
  XNOR U2214 ( .A(n1288), .B(n1356), .Z(n1290) );
  ANDN U2215 ( .A(n1060), .B(n1127), .Z(n1356) );
  XOR U2216 ( .A(n1357), .B(n1358), .Z(n1288) );
  AND U2217 ( .A(n1359), .B(n1360), .Z(n1358) );
  XOR U2218 ( .A(n1361), .B(n1357), .Z(n1360) );
  XNOR U2219 ( .A(n1304), .B(n1293), .Z(n1355) );
  XOR U2220 ( .A(n1365), .B(n1300), .Z(n1304) );
  XNOR U2221 ( .A(n1298), .B(n1366), .Z(n1300) );
  ANDN U2222 ( .A(n1167), .B(n1041), .Z(n1366) );
  XOR U2223 ( .A(n1367), .B(n1368), .Z(n1298) );
  AND U2224 ( .A(n1369), .B(n1370), .Z(n1368) );
  XNOR U2225 ( .A(n1371), .B(n1367), .Z(n1370) );
  AND U2226 ( .A(n1039), .B(n1113), .Z(n1302) );
  XNOR U2227 ( .A(n1315), .B(n1314), .Z(n1295) );
  XOR U2228 ( .A(n1375), .B(n1310), .Z(n1314) );
  XNOR U2229 ( .A(n1308), .B(n1376), .Z(n1310) );
  ANDN U2230 ( .A(n992), .B(n1250), .Z(n1376) );
  AND U2231 ( .A(n1248), .B(n951), .Z(n1312) );
  XNOR U2232 ( .A(n1321), .B(n1323), .Z(n1315) );
  NAND U2233 ( .A(n1383), .B(n895), .Z(n1323) );
  XNOR U2234 ( .A(n1319), .B(n1384), .Z(n1321) );
  ANDN U2235 ( .A(n926), .B(n1385), .Z(n1384) );
  XOR U2236 ( .A(n1386), .B(n1387), .Z(n1319) );
  AND U2237 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR U2238 ( .A(n1390), .B(n1386), .Z(n1389) );
  MUX U2239 ( .IN0(Y[18]), .IN1(n806), .SEL(n847), .F(n317) );
  XOR U2240 ( .A(n1394), .B(Y0[19]), .Z(n806) );
  XNOR U2241 ( .A(n1395), .B(n1396), .Z(n1394) );
  AND U2242 ( .A(n859), .B(n1398), .Z(n1397) );
  XOR U2243 ( .A(n1392), .B(n1396), .Z(n1398) );
  XOR U2244 ( .A(n1391), .B(n1396), .Z(n1392) );
  XNOR U2245 ( .A(n1334), .B(n1333), .Z(n1396) );
  IV U2246 ( .A(n1332), .Z(n1333) );
  XNOR U2247 ( .A(n1351), .B(n1350), .Z(n1334) );
  XOR U2248 ( .A(n1401), .B(n1354), .Z(n1350) );
  XNOR U2249 ( .A(n1344), .B(n1343), .Z(n1354) );
  XOR U2250 ( .A(n1402), .B(n1338), .Z(n1343) );
  XNOR U2251 ( .A(n1337), .B(n1403), .Z(n1338) );
  ANDN U2252 ( .A(n1404), .B(n927), .Z(n1403) );
  XOR U2253 ( .A(n1405), .B(n1406), .Z(n1337) );
  AND U2254 ( .A(n1407), .B(n1408), .Z(n1406) );
  XNOR U2255 ( .A(n1409), .B(n1405), .Z(n1408) );
  AND U2256 ( .A(n924), .B(n1341), .Z(n1339) );
  XNOR U2257 ( .A(n1347), .B(n1348), .Z(n1344) );
  NANDN U2258 ( .B(n1206), .A(n999), .Z(n1348) );
  XNOR U2259 ( .A(n1346), .B(n1413), .Z(n1347) );
  ANDN U2260 ( .A(n1276), .B(n1001), .Z(n1413) );
  XNOR U2261 ( .A(n1353), .B(n1349), .Z(n1401) );
  XNOR U2262 ( .A(n1420), .B(n1421), .Z(n1353) );
  IV U2263 ( .A(n1352), .Z(n1421) );
  XNOR U2264 ( .A(n1364), .B(n1363), .Z(n1351) );
  XOR U2265 ( .A(n1427), .B(n1374), .Z(n1363) );
  XNOR U2266 ( .A(n1359), .B(n1361), .Z(n1374) );
  NANDN U2267 ( .B(n1019), .A(n1184), .Z(n1361) );
  XNOR U2268 ( .A(n1357), .B(n1428), .Z(n1359) );
  ANDN U2269 ( .A(n1060), .B(n1186), .Z(n1428) );
  XOR U2270 ( .A(n1429), .B(n1430), .Z(n1357) );
  AND U2271 ( .A(n1431), .B(n1432), .Z(n1430) );
  XOR U2272 ( .A(n1433), .B(n1429), .Z(n1432) );
  XNOR U2273 ( .A(n1373), .B(n1362), .Z(n1427) );
  XOR U2274 ( .A(n1437), .B(n1369), .Z(n1373) );
  XNOR U2275 ( .A(n1367), .B(n1438), .Z(n1369) );
  ANDN U2276 ( .A(n1167), .B(n1085), .Z(n1438) );
  XOR U2277 ( .A(n1439), .B(n1440), .Z(n1367) );
  AND U2278 ( .A(n1441), .B(n1442), .Z(n1440) );
  XNOR U2279 ( .A(n1443), .B(n1439), .Z(n1442) );
  AND U2280 ( .A(n1083), .B(n1113), .Z(n1371) );
  XNOR U2281 ( .A(n1382), .B(n1381), .Z(n1364) );
  XOR U2282 ( .A(n1447), .B(n1378), .Z(n1381) );
  XNOR U2283 ( .A(n1377), .B(n1448), .Z(n1378) );
  ANDN U2284 ( .A(n992), .B(n1318), .Z(n1448) );
  XOR U2285 ( .A(n1449), .B(n1450), .Z(n1377) );
  AND U2286 ( .A(n1451), .B(n1452), .Z(n1450) );
  XNOR U2287 ( .A(n1453), .B(n1449), .Z(n1452) );
  AND U2288 ( .A(n1316), .B(n951), .Z(n1379) );
  XNOR U2289 ( .A(n1388), .B(n1390), .Z(n1382) );
  NAND U2290 ( .A(n1457), .B(n895), .Z(n1390) );
  XNOR U2291 ( .A(n1386), .B(n1458), .Z(n1388) );
  ANDN U2292 ( .A(n926), .B(n1459), .Z(n1458) );
  NANDN U2293 ( .B(n1460), .A(n1461), .Z(n1386) );
  NAND U2294 ( .A(n1462), .B(n1463), .Z(n1461) );
  MUX U2295 ( .IN0(Y[17]), .IN1(n803), .SEL(n847), .F(n316) );
  XOR U2296 ( .A(n1468), .B(Y0[18]), .Z(n803) );
  XOR U2297 ( .A(n1469), .B(n1470), .Z(n1468) );
  AND U2298 ( .A(n859), .B(n1472), .Z(n1471) );
  XOR U2299 ( .A(n1466), .B(n1470), .Z(n1472) );
  XOR U2300 ( .A(n1465), .B(n1470), .Z(n1466) );
  XOR U2301 ( .A(n1400), .B(n1399), .Z(n1470) );
  XNOR U2302 ( .A(n1475), .B(n1424), .Z(n1418) );
  XNOR U2303 ( .A(n1412), .B(n1411), .Z(n1424) );
  XOR U2304 ( .A(n1476), .B(n1407), .Z(n1411) );
  XNOR U2305 ( .A(n1405), .B(n1477), .Z(n1407) );
  ANDN U2306 ( .A(n1404), .B(n957), .Z(n1477) );
  XOR U2307 ( .A(n1478), .B(n1479), .Z(n1405) );
  AND U2308 ( .A(n1480), .B(n1481), .Z(n1479) );
  XNOR U2309 ( .A(n1482), .B(n1478), .Z(n1481) );
  AND U2310 ( .A(n955), .B(n1341), .Z(n1409) );
  XNOR U2311 ( .A(n1415), .B(n1416), .Z(n1412) );
  NANDN U2312 ( .B(n1206), .A(n1039), .Z(n1416) );
  XNOR U2313 ( .A(n1414), .B(n1486), .Z(n1415) );
  ANDN U2314 ( .A(n1276), .B(n1041), .Z(n1486) );
  XOR U2315 ( .A(n1487), .B(n1488), .Z(n1414) );
  AND U2316 ( .A(n1489), .B(n1490), .Z(n1488) );
  XOR U2317 ( .A(n1491), .B(n1487), .Z(n1490) );
  XNOR U2318 ( .A(n1423), .B(n1417), .Z(n1475) );
  XOR U2319 ( .A(n1495), .B(n1425), .Z(n1423) );
  NAND U2320 ( .A(n1499), .B(n1500), .Z(n1426) );
  NANDN U2321 ( .B(n1501), .A(n894), .Z(n1500) );
  NANDN U2322 ( .B(n1502), .A(n1503), .Z(n1499) );
  XNOR U2323 ( .A(n1436), .B(n1435), .Z(n1419) );
  XOR U2324 ( .A(n1507), .B(n1446), .Z(n1435) );
  XNOR U2325 ( .A(n1431), .B(n1433), .Z(n1446) );
  NANDN U2326 ( .B(n1019), .A(n1248), .Z(n1433) );
  XNOR U2327 ( .A(n1429), .B(n1508), .Z(n1431) );
  ANDN U2328 ( .A(n1060), .B(n1250), .Z(n1508) );
  XOR U2329 ( .A(n1509), .B(n1510), .Z(n1429) );
  AND U2330 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U2331 ( .A(n1513), .B(n1509), .Z(n1512) );
  XNOR U2332 ( .A(n1445), .B(n1434), .Z(n1507) );
  XOR U2333 ( .A(n1517), .B(n1441), .Z(n1445) );
  XNOR U2334 ( .A(n1439), .B(n1518), .Z(n1441) );
  ANDN U2335 ( .A(n1167), .B(n1127), .Z(n1518) );
  XOR U2336 ( .A(n1519), .B(n1520), .Z(n1439) );
  AND U2337 ( .A(n1521), .B(n1522), .Z(n1520) );
  XNOR U2338 ( .A(n1523), .B(n1519), .Z(n1522) );
  AND U2339 ( .A(n1125), .B(n1113), .Z(n1443) );
  XOR U2340 ( .A(n1456), .B(n1455), .Z(n1436) );
  XOR U2341 ( .A(n1527), .B(n1451), .Z(n1455) );
  XNOR U2342 ( .A(n1449), .B(n1528), .Z(n1451) );
  ANDN U2343 ( .A(n992), .B(n1385), .Z(n1528) );
  AND U2344 ( .A(n1383), .B(n951), .Z(n1453) );
  XOR U2345 ( .A(n1463), .B(n1462), .Z(n1456) );
  NAND U2346 ( .A(n1535), .B(n895), .Z(n1462) );
  XNOR U2347 ( .A(n1460), .B(n1536), .Z(n1463) );
  ANDN U2348 ( .A(n926), .B(n1537), .Z(n1536) );
  NANDN U2349 ( .B(n1538), .A(n1539), .Z(n1460) );
  NAND U2350 ( .A(n1540), .B(n1541), .Z(n1539) );
  IV U2351 ( .A(n1464), .Z(n1465) );
  MUX U2352 ( .IN0(Y[16]), .IN1(n800), .SEL(n847), .F(n315) );
  XOR U2353 ( .A(n1546), .B(Y0[17]), .Z(n800) );
  XOR U2354 ( .A(n1547), .B(n1548), .Z(n1546) );
  AND U2355 ( .A(n859), .B(n1550), .Z(n1549) );
  XOR U2356 ( .A(n1544), .B(n1548), .Z(n1550) );
  XOR U2357 ( .A(n1543), .B(n1548), .Z(n1544) );
  XOR U2358 ( .A(n1474), .B(n1473), .Z(n1548) );
  XNOR U2359 ( .A(n1553), .B(n1506), .Z(n1493) );
  XNOR U2360 ( .A(n1485), .B(n1484), .Z(n1506) );
  XOR U2361 ( .A(n1554), .B(n1480), .Z(n1484) );
  XNOR U2362 ( .A(n1478), .B(n1555), .Z(n1480) );
  ANDN U2363 ( .A(n1404), .B(n1001), .Z(n1555) );
  XOR U2364 ( .A(n1556), .B(n1557), .Z(n1478) );
  AND U2365 ( .A(n1558), .B(n1559), .Z(n1557) );
  XNOR U2366 ( .A(n1560), .B(n1556), .Z(n1559) );
  AND U2367 ( .A(n999), .B(n1341), .Z(n1482) );
  XNOR U2368 ( .A(n1489), .B(n1491), .Z(n1485) );
  NANDN U2369 ( .B(n1206), .A(n1083), .Z(n1491) );
  XNOR U2370 ( .A(n1487), .B(n1564), .Z(n1489) );
  ANDN U2371 ( .A(n1276), .B(n1085), .Z(n1564) );
  XOR U2372 ( .A(n1565), .B(n1566), .Z(n1487) );
  AND U2373 ( .A(n1567), .B(n1568), .Z(n1566) );
  XOR U2374 ( .A(n1569), .B(n1565), .Z(n1568) );
  XOR U2375 ( .A(n1505), .B(n1492), .Z(n1553) );
  XNOR U2376 ( .A(n1573), .B(n1497), .Z(n1505) );
  XNOR U2377 ( .A(n1574), .B(n1503), .Z(n1497) );
  AND U2378 ( .A(n924), .B(n1575), .Z(n1503) );
  NAND U2379 ( .A(n1576), .B(n1502), .Z(n1574) );
  XOR U2380 ( .A(n1577), .B(n1578), .Z(n1502) );
  AND U2381 ( .A(n1579), .B(n1580), .Z(n1578) );
  XOR U2382 ( .A(n1581), .B(n1577), .Z(n1580) );
  NANDN U2383 ( .B(n927), .A(n1582), .Z(n1576) );
  XNOR U2384 ( .A(n1496), .B(n1504), .Z(n1573) );
  IV U2385 ( .A(n1498), .Z(n1496) );
  XNOR U2386 ( .A(n1516), .B(n1515), .Z(n1494) );
  XOR U2387 ( .A(n1588), .B(n1526), .Z(n1515) );
  XNOR U2388 ( .A(n1511), .B(n1513), .Z(n1526) );
  NANDN U2389 ( .B(n1019), .A(n1316), .Z(n1513) );
  XNOR U2390 ( .A(n1509), .B(n1589), .Z(n1511) );
  ANDN U2391 ( .A(n1060), .B(n1318), .Z(n1589) );
  XNOR U2392 ( .A(n1525), .B(n1514), .Z(n1588) );
  XOR U2393 ( .A(n1596), .B(n1521), .Z(n1525) );
  XNOR U2394 ( .A(n1519), .B(n1597), .Z(n1521) );
  ANDN U2395 ( .A(n1167), .B(n1186), .Z(n1597) );
  XOR U2396 ( .A(n1598), .B(n1599), .Z(n1519) );
  AND U2397 ( .A(n1600), .B(n1601), .Z(n1599) );
  XNOR U2398 ( .A(n1602), .B(n1598), .Z(n1601) );
  AND U2399 ( .A(n1184), .B(n1113), .Z(n1523) );
  XOR U2400 ( .A(n1534), .B(n1533), .Z(n1516) );
  XOR U2401 ( .A(n1606), .B(n1530), .Z(n1533) );
  XNOR U2402 ( .A(n1529), .B(n1607), .Z(n1530) );
  ANDN U2403 ( .A(n992), .B(n1459), .Z(n1607) );
  XOR U2404 ( .A(n1608), .B(n1609), .Z(n1529) );
  AND U2405 ( .A(n1610), .B(n1611), .Z(n1609) );
  XNOR U2406 ( .A(n1612), .B(n1608), .Z(n1611) );
  AND U2407 ( .A(n1457), .B(n951), .Z(n1531) );
  XOR U2408 ( .A(n1541), .B(n1540), .Z(n1534) );
  NAND U2409 ( .A(n1616), .B(n895), .Z(n1540) );
  XNOR U2410 ( .A(n1538), .B(n1617), .Z(n1541) );
  ANDN U2411 ( .A(n926), .B(n1618), .Z(n1617) );
  NAND U2412 ( .A(n1619), .B(n1620), .Z(n1538) );
  NAND U2413 ( .A(n1621), .B(n1622), .Z(n1619) );
  IV U2414 ( .A(n1542), .Z(n1543) );
  MUX U2415 ( .IN0(Y[15]), .IN1(n797), .SEL(n847), .F(n314) );
  XOR U2416 ( .A(n1627), .B(Y0[16]), .Z(n797) );
  XOR U2417 ( .A(n1628), .B(n1629), .Z(n1627) );
  AND U2418 ( .A(n859), .B(n1631), .Z(n1630) );
  XOR U2419 ( .A(n1625), .B(n1629), .Z(n1631) );
  XOR U2420 ( .A(n1624), .B(n1629), .Z(n1625) );
  XOR U2421 ( .A(n1552), .B(n1551), .Z(n1629) );
  XNOR U2422 ( .A(n1635), .B(n1585), .Z(n1571) );
  XNOR U2423 ( .A(n1563), .B(n1562), .Z(n1585) );
  XOR U2424 ( .A(n1636), .B(n1558), .Z(n1562) );
  XNOR U2425 ( .A(n1556), .B(n1637), .Z(n1558) );
  ANDN U2426 ( .A(n1404), .B(n1041), .Z(n1637) );
  XOR U2427 ( .A(n1638), .B(n1639), .Z(n1556) );
  AND U2428 ( .A(n1640), .B(n1641), .Z(n1639) );
  XNOR U2429 ( .A(n1642), .B(n1638), .Z(n1641) );
  AND U2430 ( .A(n1039), .B(n1341), .Z(n1560) );
  XNOR U2431 ( .A(n1567), .B(n1569), .Z(n1563) );
  NANDN U2432 ( .B(n1206), .A(n1125), .Z(n1569) );
  XNOR U2433 ( .A(n1565), .B(n1646), .Z(n1567) );
  ANDN U2434 ( .A(n1276), .B(n1127), .Z(n1646) );
  XNOR U2435 ( .A(n1584), .B(n1570), .Z(n1635) );
  XOR U2436 ( .A(n1653), .B(n1587), .Z(n1584) );
  XNOR U2437 ( .A(n1579), .B(n1581), .Z(n1587) );
  NAND U2438 ( .A(n955), .B(n1575), .Z(n1581) );
  XNOR U2439 ( .A(n1577), .B(n1654), .Z(n1579) );
  ANDN U2440 ( .A(n1582), .B(n957), .Z(n1654) );
  XOR U2441 ( .A(n1655), .B(n1656), .Z(n1577) );
  AND U2442 ( .A(n1657), .B(n1658), .Z(n1656) );
  XOR U2443 ( .A(n1659), .B(n1655), .Z(n1658) );
  XNOR U2444 ( .A(n1586), .B(n1583), .Z(n1653) );
  AND U2445 ( .A(n1664), .B(n1665), .Z(n1663) );
  NANDN U2446 ( .B(n1666), .A(n894), .Z(n1665) );
  NANDN U2447 ( .B(n1667), .A(n1668), .Z(n1664) );
  XNOR U2448 ( .A(n1595), .B(n1594), .Z(n1572) );
  XOR U2449 ( .A(n1672), .B(n1605), .Z(n1594) );
  XNOR U2450 ( .A(n1591), .B(n1592), .Z(n1605) );
  NANDN U2451 ( .B(n1019), .A(n1383), .Z(n1592) );
  XNOR U2452 ( .A(n1590), .B(n1673), .Z(n1591) );
  ANDN U2453 ( .A(n1060), .B(n1385), .Z(n1673) );
  XNOR U2454 ( .A(n1604), .B(n1593), .Z(n1672) );
  XOR U2455 ( .A(n1680), .B(n1600), .Z(n1604) );
  XNOR U2456 ( .A(n1598), .B(n1681), .Z(n1600) );
  ANDN U2457 ( .A(n1167), .B(n1250), .Z(n1681) );
  XOR U2458 ( .A(n1682), .B(n1683), .Z(n1598) );
  AND U2459 ( .A(n1684), .B(n1685), .Z(n1683) );
  XNOR U2460 ( .A(n1686), .B(n1682), .Z(n1685) );
  AND U2461 ( .A(n1248), .B(n1113), .Z(n1602) );
  XOR U2462 ( .A(n1615), .B(n1614), .Z(n1595) );
  XOR U2463 ( .A(n1690), .B(n1610), .Z(n1614) );
  XNOR U2464 ( .A(n1608), .B(n1691), .Z(n1610) );
  ANDN U2465 ( .A(n992), .B(n1537), .Z(n1691) );
  XOR U2466 ( .A(n1692), .B(n1693), .Z(n1608) );
  AND U2467 ( .A(n1694), .B(n1695), .Z(n1693) );
  XNOR U2468 ( .A(n1696), .B(n1692), .Z(n1695) );
  AND U2469 ( .A(n1535), .B(n951), .Z(n1612) );
  XOR U2470 ( .A(n1622), .B(n1621), .Z(n1615) );
  NAND U2471 ( .A(n1700), .B(n895), .Z(n1621) );
  XOR U2472 ( .A(n1620), .B(n1701), .Z(n1622) );
  ANDN U2473 ( .A(n926), .B(n1702), .Z(n1701) );
  ANDN U2474 ( .A(n1703), .B(n1704), .Z(n1620) );
  NAND U2475 ( .A(n1705), .B(n1706), .Z(n1703) );
  IV U2476 ( .A(n1623), .Z(n1624) );
  MUX U2477 ( .IN0(Y[14]), .IN1(n794), .SEL(n847), .F(n313) );
  XOR U2478 ( .A(n1711), .B(Y0[15]), .Z(n794) );
  XOR U2479 ( .A(n1712), .B(n1713), .Z(n1711) );
  AND U2480 ( .A(n859), .B(n1715), .Z(n1714) );
  XOR U2481 ( .A(n1709), .B(n1713), .Z(n1715) );
  XOR U2482 ( .A(n1708), .B(n1713), .Z(n1709) );
  XNOR U2483 ( .A(n1634), .B(n1633), .Z(n1713) );
  XOR U2484 ( .A(n1716), .B(n1717), .Z(n1633) );
  XOR U2485 ( .A(n1718), .B(n1719), .Z(n1717) );
  XOR U2486 ( .A(n1720), .B(n1718), .Z(n1719) );
  XNOR U2487 ( .A(n1726), .B(n1662), .Z(n1651) );
  XNOR U2488 ( .A(n1645), .B(n1644), .Z(n1662) );
  XOR U2489 ( .A(n1727), .B(n1640), .Z(n1644) );
  XNOR U2490 ( .A(n1638), .B(n1728), .Z(n1640) );
  ANDN U2491 ( .A(n1404), .B(n1085), .Z(n1728) );
  AND U2492 ( .A(n1083), .B(n1341), .Z(n1642) );
  XNOR U2493 ( .A(n1648), .B(n1649), .Z(n1645) );
  NANDN U2494 ( .B(n1206), .A(n1184), .Z(n1649) );
  XNOR U2495 ( .A(n1647), .B(n1735), .Z(n1648) );
  ANDN U2496 ( .A(n1276), .B(n1186), .Z(n1735) );
  XOR U2497 ( .A(n1736), .B(n1737), .Z(n1647) );
  AND U2498 ( .A(n1738), .B(n1739), .Z(n1737) );
  XOR U2499 ( .A(n1740), .B(n1736), .Z(n1739) );
  XNOR U2500 ( .A(n1661), .B(n1650), .Z(n1726) );
  XOR U2501 ( .A(n1744), .B(n1671), .Z(n1661) );
  XNOR U2502 ( .A(n1657), .B(n1659), .Z(n1671) );
  NAND U2503 ( .A(n999), .B(n1575), .Z(n1659) );
  XNOR U2504 ( .A(n1655), .B(n1745), .Z(n1657) );
  ANDN U2505 ( .A(n1582), .B(n1001), .Z(n1745) );
  XOR U2506 ( .A(n1746), .B(n1747), .Z(n1655) );
  AND U2507 ( .A(n1748), .B(n1749), .Z(n1747) );
  XOR U2508 ( .A(n1750), .B(n1746), .Z(n1749) );
  XNOR U2509 ( .A(n1670), .B(n1660), .Z(n1744) );
  XOR U2510 ( .A(n1758), .B(n1668), .Z(n1754) );
  AND U2511 ( .A(n924), .B(n1759), .Z(n1668) );
  NAND U2512 ( .A(n1760), .B(n1667), .Z(n1758) );
  XOR U2513 ( .A(n1761), .B(n1762), .Z(n1667) );
  AND U2514 ( .A(n1763), .B(n1764), .Z(n1762) );
  XNOR U2515 ( .A(n1765), .B(n1761), .Z(n1764) );
  NANDN U2516 ( .B(n927), .A(n1766), .Z(n1760) );
  XNOR U2517 ( .A(n1679), .B(n1678), .Z(n1652) );
  XOR U2518 ( .A(n1767), .B(n1689), .Z(n1678) );
  XNOR U2519 ( .A(n1675), .B(n1676), .Z(n1689) );
  NANDN U2520 ( .B(n1019), .A(n1457), .Z(n1676) );
  XNOR U2521 ( .A(n1674), .B(n1768), .Z(n1675) );
  ANDN U2522 ( .A(n1060), .B(n1459), .Z(n1768) );
  XNOR U2523 ( .A(n1688), .B(n1677), .Z(n1767) );
  XOR U2524 ( .A(n1775), .B(n1684), .Z(n1688) );
  XNOR U2525 ( .A(n1682), .B(n1776), .Z(n1684) );
  ANDN U2526 ( .A(n1167), .B(n1318), .Z(n1776) );
  AND U2527 ( .A(n1316), .B(n1113), .Z(n1686) );
  XOR U2528 ( .A(n1699), .B(n1698), .Z(n1679) );
  XOR U2529 ( .A(n1783), .B(n1694), .Z(n1698) );
  XNOR U2530 ( .A(n1692), .B(n1784), .Z(n1694) );
  ANDN U2531 ( .A(n992), .B(n1618), .Z(n1784) );
  AND U2532 ( .A(n1616), .B(n951), .Z(n1696) );
  XOR U2533 ( .A(n1706), .B(n1705), .Z(n1699) );
  NAND U2534 ( .A(n1791), .B(n895), .Z(n1705) );
  XNOR U2535 ( .A(n1704), .B(n1792), .Z(n1706) );
  ANDN U2536 ( .A(n926), .B(n1793), .Z(n1792) );
  NAND U2537 ( .A(n1794), .B(n1795), .Z(n1704) );
  NAND U2538 ( .A(n1796), .B(n1797), .Z(n1794) );
  IV U2539 ( .A(n1707), .Z(n1708) );
  MUX U2540 ( .IN0(Y[13]), .IN1(n791), .SEL(n847), .F(n312) );
  XOR U2541 ( .A(n1802), .B(Y0[14]), .Z(n791) );
  XOR U2542 ( .A(n1803), .B(n1804), .Z(n1802) );
  AND U2543 ( .A(n859), .B(n1806), .Z(n1805) );
  XOR U2544 ( .A(n1800), .B(n1804), .Z(n1806) );
  XOR U2545 ( .A(n1799), .B(n1804), .Z(n1800) );
  XOR U2546 ( .A(n1807), .B(n1721), .Z(n1724) );
  NAND U2547 ( .A(n1718), .B(n1811), .Z(n1722) );
  AND U2548 ( .A(n1812), .B(n1813), .Z(n1811) );
  NANDN U2549 ( .B(n1814), .A(n894), .Z(n1813) );
  NANDN U2550 ( .B(n1815), .A(n1816), .Z(n1812) );
  AND U2551 ( .A(n1817), .B(n1818), .Z(n1718) );
  NANDN U2552 ( .B(n1819), .A(n1820), .Z(n1818) );
  OR U2553 ( .A(n1821), .B(n1822), .Z(n1817) );
  XNOR U2554 ( .A(n1743), .B(n1742), .Z(n1725) );
  XOR U2555 ( .A(n1826), .B(n1753), .Z(n1742) );
  XNOR U2556 ( .A(n1734), .B(n1733), .Z(n1753) );
  XOR U2557 ( .A(n1827), .B(n1730), .Z(n1733) );
  XNOR U2558 ( .A(n1729), .B(n1828), .Z(n1730) );
  ANDN U2559 ( .A(n1404), .B(n1127), .Z(n1828) );
  XOR U2560 ( .A(n1829), .B(n1830), .Z(n1729) );
  AND U2561 ( .A(n1831), .B(n1832), .Z(n1830) );
  XNOR U2562 ( .A(n1833), .B(n1829), .Z(n1832) );
  AND U2563 ( .A(n1125), .B(n1341), .Z(n1731) );
  XNOR U2564 ( .A(n1738), .B(n1740), .Z(n1734) );
  NANDN U2565 ( .B(n1206), .A(n1248), .Z(n1740) );
  XNOR U2566 ( .A(n1736), .B(n1837), .Z(n1738) );
  ANDN U2567 ( .A(n1276), .B(n1250), .Z(n1837) );
  XNOR U2568 ( .A(n1752), .B(n1741), .Z(n1826) );
  XOR U2569 ( .A(n1844), .B(n1757), .Z(n1752) );
  XNOR U2570 ( .A(n1748), .B(n1750), .Z(n1757) );
  NAND U2571 ( .A(n1039), .B(n1575), .Z(n1750) );
  XNOR U2572 ( .A(n1746), .B(n1845), .Z(n1748) );
  ANDN U2573 ( .A(n1582), .B(n1041), .Z(n1845) );
  XOR U2574 ( .A(n1846), .B(n1847), .Z(n1746) );
  AND U2575 ( .A(n1848), .B(n1849), .Z(n1847) );
  XOR U2576 ( .A(n1850), .B(n1846), .Z(n1849) );
  XNOR U2577 ( .A(n1756), .B(n1751), .Z(n1844) );
  XOR U2578 ( .A(n1854), .B(n1763), .Z(n1756) );
  XNOR U2579 ( .A(n1761), .B(n1855), .Z(n1763) );
  ANDN U2580 ( .A(n1766), .B(n957), .Z(n1855) );
  XOR U2581 ( .A(n1856), .B(n1857), .Z(n1761) );
  AND U2582 ( .A(n1858), .B(n1859), .Z(n1857) );
  XNOR U2583 ( .A(n1860), .B(n1856), .Z(n1859) );
  AND U2584 ( .A(n955), .B(n1759), .Z(n1765) );
  XNOR U2585 ( .A(n1774), .B(n1773), .Z(n1743) );
  XOR U2586 ( .A(n1864), .B(n1782), .Z(n1773) );
  XNOR U2587 ( .A(n1770), .B(n1771), .Z(n1782) );
  NANDN U2588 ( .B(n1019), .A(n1535), .Z(n1771) );
  XNOR U2589 ( .A(n1769), .B(n1865), .Z(n1770) );
  ANDN U2590 ( .A(n1060), .B(n1537), .Z(n1865) );
  XNOR U2591 ( .A(n1781), .B(n1772), .Z(n1864) );
  XOR U2592 ( .A(n1872), .B(n1778), .Z(n1781) );
  XNOR U2593 ( .A(n1777), .B(n1873), .Z(n1778) );
  ANDN U2594 ( .A(n1167), .B(n1385), .Z(n1873) );
  AND U2595 ( .A(n1383), .B(n1113), .Z(n1779) );
  XOR U2596 ( .A(n1790), .B(n1789), .Z(n1774) );
  XOR U2597 ( .A(n1880), .B(n1786), .Z(n1789) );
  XNOR U2598 ( .A(n1785), .B(n1881), .Z(n1786) );
  ANDN U2599 ( .A(n992), .B(n1702), .Z(n1881) );
  AND U2600 ( .A(n1700), .B(n951), .Z(n1787) );
  XOR U2601 ( .A(n1797), .B(n1796), .Z(n1790) );
  NAND U2602 ( .A(n1888), .B(n895), .Z(n1796) );
  XOR U2603 ( .A(n1795), .B(n1889), .Z(n1797) );
  ANDN U2604 ( .A(n926), .B(n1890), .Z(n1889) );
  ANDN U2605 ( .A(n1891), .B(n1892), .Z(n1795) );
  NAND U2606 ( .A(n1893), .B(n1894), .Z(n1891) );
  IV U2607 ( .A(n1798), .Z(n1799) );
  MUX U2608 ( .IN0(Y[12]), .IN1(n788), .SEL(n847), .F(n311) );
  XOR U2609 ( .A(n1899), .B(Y0[13]), .Z(n788) );
  XNOR U2610 ( .A(n1900), .B(n1901), .Z(n1899) );
  AND U2611 ( .A(n859), .B(n1903), .Z(n1902) );
  XNOR U2612 ( .A(n1897), .B(n1901), .Z(n1903) );
  XNOR U2613 ( .A(n1896), .B(n1901), .Z(n1897) );
  XNOR U2614 ( .A(n1825), .B(n1824), .Z(n1901) );
  XOR U2615 ( .A(n1904), .B(n1809), .Z(n1824) );
  NANDN U2616 ( .B(n1905), .A(n1906), .Z(n1815) );
  XOR U2617 ( .A(n1909), .B(n1822), .Z(n1819) );
  NAND U2618 ( .A(n1910), .B(n924), .Z(n1822) );
  NAND U2619 ( .A(n1911), .B(n1821), .Z(n1909) );
  NANDN U2620 ( .B(n927), .A(n1915), .Z(n1911) );
  XNOR U2621 ( .A(n1808), .B(n1823), .Z(n1904) );
  IV U2622 ( .A(n1810), .Z(n1808) );
  XNOR U2623 ( .A(n1843), .B(n1842), .Z(n1825) );
  XOR U2624 ( .A(n1922), .B(n1853), .Z(n1842) );
  XNOR U2625 ( .A(n1836), .B(n1835), .Z(n1853) );
  XOR U2626 ( .A(n1923), .B(n1831), .Z(n1835) );
  XNOR U2627 ( .A(n1829), .B(n1924), .Z(n1831) );
  ANDN U2628 ( .A(n1404), .B(n1186), .Z(n1924) );
  XOR U2629 ( .A(n1925), .B(n1926), .Z(n1829) );
  AND U2630 ( .A(n1927), .B(n1928), .Z(n1926) );
  XNOR U2631 ( .A(n1929), .B(n1925), .Z(n1928) );
  AND U2632 ( .A(n1184), .B(n1341), .Z(n1833) );
  XNOR U2633 ( .A(n1839), .B(n1840), .Z(n1836) );
  NANDN U2634 ( .B(n1206), .A(n1316), .Z(n1840) );
  XNOR U2635 ( .A(n1838), .B(n1933), .Z(n1839) );
  ANDN U2636 ( .A(n1276), .B(n1318), .Z(n1933) );
  XNOR U2637 ( .A(n1852), .B(n1841), .Z(n1922) );
  XOR U2638 ( .A(n1940), .B(n1863), .Z(n1852) );
  XNOR U2639 ( .A(n1848), .B(n1850), .Z(n1863) );
  NAND U2640 ( .A(n1083), .B(n1575), .Z(n1850) );
  XNOR U2641 ( .A(n1846), .B(n1941), .Z(n1848) );
  ANDN U2642 ( .A(n1582), .B(n1085), .Z(n1941) );
  XOR U2643 ( .A(n1942), .B(n1943), .Z(n1846) );
  AND U2644 ( .A(n1944), .B(n1945), .Z(n1943) );
  XOR U2645 ( .A(n1946), .B(n1942), .Z(n1945) );
  XNOR U2646 ( .A(n1862), .B(n1851), .Z(n1940) );
  XOR U2647 ( .A(n1950), .B(n1858), .Z(n1862) );
  XNOR U2648 ( .A(n1856), .B(n1951), .Z(n1858) );
  ANDN U2649 ( .A(n1766), .B(n1001), .Z(n1951) );
  XOR U2650 ( .A(n1952), .B(n1953), .Z(n1856) );
  AND U2651 ( .A(n1954), .B(n1955), .Z(n1953) );
  XNOR U2652 ( .A(n1956), .B(n1952), .Z(n1955) );
  AND U2653 ( .A(n999), .B(n1759), .Z(n1860) );
  XNOR U2654 ( .A(n1871), .B(n1870), .Z(n1843) );
  XOR U2655 ( .A(n1960), .B(n1879), .Z(n1870) );
  XNOR U2656 ( .A(n1867), .B(n1868), .Z(n1879) );
  NANDN U2657 ( .B(n1019), .A(n1616), .Z(n1868) );
  XNOR U2658 ( .A(n1866), .B(n1961), .Z(n1867) );
  ANDN U2659 ( .A(n1060), .B(n1618), .Z(n1961) );
  XNOR U2660 ( .A(n1878), .B(n1869), .Z(n1960) );
  XOR U2661 ( .A(n1968), .B(n1875), .Z(n1878) );
  XNOR U2662 ( .A(n1874), .B(n1969), .Z(n1875) );
  ANDN U2663 ( .A(n1167), .B(n1459), .Z(n1969) );
  AND U2664 ( .A(n1457), .B(n1113), .Z(n1876) );
  XOR U2665 ( .A(n1887), .B(n1886), .Z(n1871) );
  XOR U2666 ( .A(n1976), .B(n1883), .Z(n1886) );
  XNOR U2667 ( .A(n1882), .B(n1977), .Z(n1883) );
  ANDN U2668 ( .A(n992), .B(n1793), .Z(n1977) );
  AND U2669 ( .A(n1791), .B(n951), .Z(n1884) );
  XOR U2670 ( .A(n1894), .B(n1893), .Z(n1887) );
  NAND U2671 ( .A(n1984), .B(n895), .Z(n1893) );
  XNOR U2672 ( .A(n1892), .B(n1985), .Z(n1894) );
  ANDN U2673 ( .A(n926), .B(n1986), .Z(n1985) );
  NAND U2674 ( .A(n1987), .B(n1988), .Z(n1892) );
  NAND U2675 ( .A(n1989), .B(n1990), .Z(n1987) );
  IV U2676 ( .A(n1895), .Z(n1896) );
  MUX U2677 ( .IN0(Y[11]), .IN1(n785), .SEL(n847), .F(n310) );
  XOR U2678 ( .A(n1995), .B(Y0[12]), .Z(n785) );
  XOR U2679 ( .A(n1996), .B(n1997), .Z(n1995) );
  AND U2680 ( .A(n859), .B(n1999), .Z(n1998) );
  XOR U2681 ( .A(n1993), .B(n1997), .Z(n1999) );
  XOR U2682 ( .A(n1992), .B(n1997), .Z(n1993) );
  XNOR U2683 ( .A(n2000), .B(n1921), .Z(n1917) );
  XOR U2684 ( .A(n1906), .B(n1905), .Z(n1921) );
  NANDN U2685 ( .B(n2001), .A(n2002), .Z(n1905) );
  AND U2686 ( .A(n2004), .B(n2005), .Z(n2003) );
  NANDN U2687 ( .B(n2006), .A(n894), .Z(n2005) );
  NANDN U2688 ( .B(n2007), .A(n2008), .Z(n2004) );
  XNOR U2689 ( .A(n1913), .B(n1914), .Z(n1908) );
  NAND U2690 ( .A(n1910), .B(n955), .Z(n1914) );
  XNOR U2691 ( .A(n1912), .B(n2012), .Z(n1913) );
  ANDN U2692 ( .A(n1915), .B(n957), .Z(n2012) );
  XNOR U2693 ( .A(n1920), .B(n1916), .Z(n2000) );
  IV U2694 ( .A(n1919), .Z(n1920) );
  XNOR U2695 ( .A(n1939), .B(n1938), .Z(n1918) );
  XOR U2696 ( .A(n2022), .B(n1949), .Z(n1938) );
  XNOR U2697 ( .A(n1932), .B(n1931), .Z(n1949) );
  XOR U2698 ( .A(n2023), .B(n1927), .Z(n1931) );
  XNOR U2699 ( .A(n1925), .B(n2024), .Z(n1927) );
  ANDN U2700 ( .A(n1404), .B(n1250), .Z(n2024) );
  AND U2701 ( .A(n1248), .B(n1341), .Z(n1929) );
  XNOR U2702 ( .A(n1935), .B(n1936), .Z(n1932) );
  NANDN U2703 ( .B(n1206), .A(n1383), .Z(n1936) );
  XNOR U2704 ( .A(n1934), .B(n2031), .Z(n1935) );
  ANDN U2705 ( .A(n1276), .B(n1385), .Z(n2031) );
  XNOR U2706 ( .A(n1948), .B(n1937), .Z(n2022) );
  XOR U2707 ( .A(n2038), .B(n1959), .Z(n1948) );
  XNOR U2708 ( .A(n1944), .B(n1946), .Z(n1959) );
  NAND U2709 ( .A(n1125), .B(n1575), .Z(n1946) );
  XNOR U2710 ( .A(n1942), .B(n2039), .Z(n1944) );
  ANDN U2711 ( .A(n1582), .B(n1127), .Z(n2039) );
  XNOR U2712 ( .A(n1958), .B(n1947), .Z(n2038) );
  XOR U2713 ( .A(n2046), .B(n1954), .Z(n1958) );
  XNOR U2714 ( .A(n1952), .B(n2047), .Z(n1954) );
  ANDN U2715 ( .A(n1766), .B(n1041), .Z(n2047) );
  XOR U2716 ( .A(n2048), .B(n2049), .Z(n1952) );
  AND U2717 ( .A(n2050), .B(n2051), .Z(n2049) );
  XNOR U2718 ( .A(n2052), .B(n2048), .Z(n2051) );
  AND U2719 ( .A(n1039), .B(n1759), .Z(n1956) );
  XNOR U2720 ( .A(n1967), .B(n1966), .Z(n1939) );
  XOR U2721 ( .A(n2056), .B(n1975), .Z(n1966) );
  XNOR U2722 ( .A(n1963), .B(n1964), .Z(n1975) );
  NANDN U2723 ( .B(n1019), .A(n1700), .Z(n1964) );
  XNOR U2724 ( .A(n1962), .B(n2057), .Z(n1963) );
  ANDN U2725 ( .A(n1060), .B(n1702), .Z(n2057) );
  XNOR U2726 ( .A(n1974), .B(n1965), .Z(n2056) );
  XOR U2727 ( .A(n2064), .B(n1971), .Z(n1974) );
  XNOR U2728 ( .A(n1970), .B(n2065), .Z(n1971) );
  ANDN U2729 ( .A(n1167), .B(n1537), .Z(n2065) );
  AND U2730 ( .A(n1535), .B(n1113), .Z(n1972) );
  XOR U2731 ( .A(n1983), .B(n1982), .Z(n1967) );
  XOR U2732 ( .A(n2072), .B(n1979), .Z(n1982) );
  XNOR U2733 ( .A(n1978), .B(n2073), .Z(n1979) );
  ANDN U2734 ( .A(n992), .B(n1890), .Z(n2073) );
  AND U2735 ( .A(n1888), .B(n951), .Z(n1980) );
  XOR U2736 ( .A(n1990), .B(n1989), .Z(n1983) );
  NAND U2737 ( .A(n2080), .B(n895), .Z(n1989) );
  XOR U2738 ( .A(n1988), .B(n2081), .Z(n1990) );
  ANDN U2739 ( .A(n926), .B(n2082), .Z(n2081) );
  ANDN U2740 ( .A(n2083), .B(n2084), .Z(n1988) );
  NAND U2741 ( .A(n2085), .B(n2086), .Z(n2083) );
  IV U2742 ( .A(n1991), .Z(n1992) );
  MUX U2743 ( .IN0(Y[10]), .IN1(n782), .SEL(n847), .F(n309) );
  XOR U2744 ( .A(n2091), .B(Y0[11]), .Z(n782) );
  XNOR U2745 ( .A(n2092), .B(n2093), .Z(n2091) );
  AND U2746 ( .A(n859), .B(n2095), .Z(n2094) );
  XNOR U2747 ( .A(n2089), .B(n2093), .Z(n2095) );
  XNOR U2748 ( .A(n2088), .B(n2093), .Z(n2089) );
  XNOR U2749 ( .A(n2018), .B(n2017), .Z(n2093) );
  XOR U2750 ( .A(n2096), .B(n2021), .Z(n2017) );
  XOR U2751 ( .A(n2011), .B(n2010), .Z(n2001) );
  XOR U2752 ( .A(n2104), .B(n2008), .Z(n2100) );
  AND U2753 ( .A(n2105), .B(n924), .Z(n2008) );
  NAND U2754 ( .A(n2106), .B(n2007), .Z(n2104) );
  XOR U2755 ( .A(n2107), .B(n2108), .Z(n2007) );
  AND U2756 ( .A(n2109), .B(n2110), .Z(n2108) );
  XNOR U2757 ( .A(n2111), .B(n2107), .Z(n2110) );
  NANDN U2758 ( .B(n927), .A(n2112), .Z(n2106) );
  XNOR U2759 ( .A(n2014), .B(n2015), .Z(n2011) );
  NAND U2760 ( .A(n1910), .B(n999), .Z(n2015) );
  XNOR U2761 ( .A(n2013), .B(n2113), .Z(n2014) );
  ANDN U2762 ( .A(n1915), .B(n1001), .Z(n2113) );
  XNOR U2763 ( .A(n2020), .B(n2016), .Z(n2096) );
  IV U2764 ( .A(n2019), .Z(n2020) );
  XNOR U2765 ( .A(n2037), .B(n2036), .Z(n2018) );
  XOR U2766 ( .A(n2123), .B(n2045), .Z(n2036) );
  XNOR U2767 ( .A(n2030), .B(n2029), .Z(n2045) );
  XOR U2768 ( .A(n2124), .B(n2026), .Z(n2029) );
  XNOR U2769 ( .A(n2025), .B(n2125), .Z(n2026) );
  ANDN U2770 ( .A(n1404), .B(n1318), .Z(n2125) );
  AND U2771 ( .A(n1316), .B(n1341), .Z(n2027) );
  XNOR U2772 ( .A(n2033), .B(n2034), .Z(n2030) );
  NANDN U2773 ( .B(n1206), .A(n1457), .Z(n2034) );
  XNOR U2774 ( .A(n2032), .B(n2132), .Z(n2033) );
  ANDN U2775 ( .A(n1276), .B(n1459), .Z(n2132) );
  XNOR U2776 ( .A(n2044), .B(n2035), .Z(n2123) );
  XOR U2777 ( .A(n2139), .B(n2055), .Z(n2044) );
  XNOR U2778 ( .A(n2041), .B(n2042), .Z(n2055) );
  NAND U2779 ( .A(n1184), .B(n1575), .Z(n2042) );
  XNOR U2780 ( .A(n2040), .B(n2140), .Z(n2041) );
  ANDN U2781 ( .A(n1582), .B(n1186), .Z(n2140) );
  XNOR U2782 ( .A(n2054), .B(n2043), .Z(n2139) );
  XOR U2783 ( .A(n2147), .B(n2050), .Z(n2054) );
  XNOR U2784 ( .A(n2048), .B(n2148), .Z(n2050) );
  ANDN U2785 ( .A(n1766), .B(n1085), .Z(n2148) );
  XOR U2786 ( .A(n2149), .B(n2150), .Z(n2048) );
  AND U2787 ( .A(n2151), .B(n2152), .Z(n2150) );
  XNOR U2788 ( .A(n2153), .B(n2149), .Z(n2152) );
  AND U2789 ( .A(n1083), .B(n1759), .Z(n2052) );
  XNOR U2790 ( .A(n2063), .B(n2062), .Z(n2037) );
  XOR U2791 ( .A(n2157), .B(n2071), .Z(n2062) );
  XNOR U2792 ( .A(n2059), .B(n2060), .Z(n2071) );
  NANDN U2793 ( .B(n1019), .A(n1791), .Z(n2060) );
  XNOR U2794 ( .A(n2058), .B(n2158), .Z(n2059) );
  ANDN U2795 ( .A(n1060), .B(n1793), .Z(n2158) );
  XNOR U2796 ( .A(n2070), .B(n2061), .Z(n2157) );
  XOR U2797 ( .A(n2165), .B(n2067), .Z(n2070) );
  XNOR U2798 ( .A(n2066), .B(n2166), .Z(n2067) );
  ANDN U2799 ( .A(n1167), .B(n1618), .Z(n2166) );
  AND U2800 ( .A(n1616), .B(n1113), .Z(n2068) );
  XOR U2801 ( .A(n2079), .B(n2078), .Z(n2063) );
  XOR U2802 ( .A(n2173), .B(n2075), .Z(n2078) );
  XNOR U2803 ( .A(n2074), .B(n2174), .Z(n2075) );
  ANDN U2804 ( .A(n992), .B(n1986), .Z(n2174) );
  AND U2805 ( .A(n1984), .B(n951), .Z(n2076) );
  XOR U2806 ( .A(n2086), .B(n2085), .Z(n2079) );
  NAND U2807 ( .A(n2181), .B(n895), .Z(n2085) );
  XNOR U2808 ( .A(n2084), .B(n2182), .Z(n2086) );
  ANDN U2809 ( .A(n926), .B(n2183), .Z(n2182) );
  NAND U2810 ( .A(n2184), .B(n2185), .Z(n2084) );
  NAND U2811 ( .A(n2186), .B(n2187), .Z(n2184) );
  IV U2812 ( .A(n2087), .Z(n2088) );
  MUX U2813 ( .IN0(Y[9]), .IN1(n779), .SEL(n847), .F(n308) );
  XOR U2814 ( .A(n2192), .B(Y0[10]), .Z(n779) );
  XOR U2815 ( .A(n2193), .B(n2194), .Z(n2192) );
  AND U2816 ( .A(n859), .B(n2196), .Z(n2195) );
  XOR U2817 ( .A(n2190), .B(n2194), .Z(n2196) );
  XOR U2818 ( .A(n2189), .B(n2194), .Z(n2190) );
  XNOR U2819 ( .A(n2197), .B(n2122), .Z(n2118) );
  XNOR U2820 ( .A(n2099), .B(n2098), .Z(n2122) );
  XOR U2821 ( .A(n2097), .B(n2198), .Z(n2098) );
  AND U2822 ( .A(n2199), .B(n2200), .Z(n2198) );
  NANDN U2823 ( .B(n2201), .A(n2202), .Z(n2200) );
  AND U2824 ( .A(n2203), .B(n2204), .Z(n2199) );
  NANDN U2825 ( .B(n2205), .A(n894), .Z(n2204) );
  OR U2826 ( .A(n2206), .B(n2207), .Z(n2203) );
  XNOR U2827 ( .A(n2103), .B(n2102), .Z(n2099) );
  XOR U2828 ( .A(n2211), .B(n2109), .Z(n2102) );
  XNOR U2829 ( .A(n2107), .B(n2212), .Z(n2109) );
  ANDN U2830 ( .A(n2112), .B(n957), .Z(n2212) );
  XOR U2831 ( .A(n2213), .B(n2214), .Z(n2107) );
  AND U2832 ( .A(n2215), .B(n2216), .Z(n2214) );
  XNOR U2833 ( .A(n2217), .B(n2213), .Z(n2216) );
  AND U2834 ( .A(n2105), .B(n955), .Z(n2111) );
  XNOR U2835 ( .A(n2115), .B(n2116), .Z(n2103) );
  NAND U2836 ( .A(n1910), .B(n1039), .Z(n2116) );
  XNOR U2837 ( .A(n2114), .B(n2221), .Z(n2115) );
  ANDN U2838 ( .A(n1915), .B(n1041), .Z(n2221) );
  XNOR U2839 ( .A(n2121), .B(n2117), .Z(n2197) );
  IV U2840 ( .A(n2120), .Z(n2121) );
  XNOR U2841 ( .A(n2138), .B(n2137), .Z(n2119) );
  XOR U2842 ( .A(n2231), .B(n2146), .Z(n2137) );
  XNOR U2843 ( .A(n2131), .B(n2130), .Z(n2146) );
  XOR U2844 ( .A(n2232), .B(n2127), .Z(n2130) );
  XNOR U2845 ( .A(n2126), .B(n2233), .Z(n2127) );
  ANDN U2846 ( .A(n1404), .B(n1385), .Z(n2233) );
  AND U2847 ( .A(n1383), .B(n1341), .Z(n2128) );
  XNOR U2848 ( .A(n2134), .B(n2135), .Z(n2131) );
  NANDN U2849 ( .B(n1206), .A(n1535), .Z(n2135) );
  XNOR U2850 ( .A(n2133), .B(n2240), .Z(n2134) );
  ANDN U2851 ( .A(n1276), .B(n1537), .Z(n2240) );
  XNOR U2852 ( .A(n2145), .B(n2136), .Z(n2231) );
  XOR U2853 ( .A(n2247), .B(n2156), .Z(n2145) );
  XNOR U2854 ( .A(n2142), .B(n2143), .Z(n2156) );
  NAND U2855 ( .A(n1248), .B(n1575), .Z(n2143) );
  XNOR U2856 ( .A(n2141), .B(n2248), .Z(n2142) );
  ANDN U2857 ( .A(n1582), .B(n1250), .Z(n2248) );
  XNOR U2858 ( .A(n2155), .B(n2144), .Z(n2247) );
  XOR U2859 ( .A(n2255), .B(n2151), .Z(n2155) );
  XNOR U2860 ( .A(n2149), .B(n2256), .Z(n2151) );
  ANDN U2861 ( .A(n1766), .B(n1127), .Z(n2256) );
  AND U2862 ( .A(n1125), .B(n1759), .Z(n2153) );
  XNOR U2863 ( .A(n2164), .B(n2163), .Z(n2138) );
  XOR U2864 ( .A(n2263), .B(n2172), .Z(n2163) );
  XNOR U2865 ( .A(n2160), .B(n2161), .Z(n2172) );
  NANDN U2866 ( .B(n1019), .A(n1888), .Z(n2161) );
  XNOR U2867 ( .A(n2159), .B(n2264), .Z(n2160) );
  ANDN U2868 ( .A(n1060), .B(n1890), .Z(n2264) );
  XNOR U2869 ( .A(n2171), .B(n2162), .Z(n2263) );
  XOR U2870 ( .A(n2271), .B(n2168), .Z(n2171) );
  XNOR U2871 ( .A(n2167), .B(n2272), .Z(n2168) );
  ANDN U2872 ( .A(n1167), .B(n1702), .Z(n2272) );
  AND U2873 ( .A(n1700), .B(n1113), .Z(n2169) );
  XOR U2874 ( .A(n2180), .B(n2179), .Z(n2164) );
  XOR U2875 ( .A(n2279), .B(n2176), .Z(n2179) );
  XNOR U2876 ( .A(n2175), .B(n2280), .Z(n2176) );
  ANDN U2877 ( .A(n992), .B(n2082), .Z(n2280) );
  AND U2878 ( .A(n2080), .B(n951), .Z(n2177) );
  XOR U2879 ( .A(n2187), .B(n2186), .Z(n2180) );
  NAND U2880 ( .A(n2287), .B(n895), .Z(n2186) );
  XOR U2881 ( .A(n2185), .B(n2288), .Z(n2187) );
  ANDN U2882 ( .A(n926), .B(n2289), .Z(n2288) );
  ANDN U2883 ( .A(n2290), .B(n2291), .Z(n2185) );
  NAND U2884 ( .A(n2292), .B(n2293), .Z(n2290) );
  IV U2885 ( .A(n2188), .Z(n2189) );
  MUX U2886 ( .IN0(Y[8]), .IN1(n776), .SEL(n847), .F(n307) );
  XOR U2887 ( .A(n2298), .B(Y0[9]), .Z(n776) );
  XOR U2888 ( .A(n2299), .B(n2300), .Z(n2298) );
  AND U2889 ( .A(n859), .B(n2302), .Z(n2301) );
  XOR U2890 ( .A(n2296), .B(n2300), .Z(n2302) );
  XOR U2891 ( .A(n2295), .B(n2300), .Z(n2296) );
  XNOR U2892 ( .A(n2303), .B(n2230), .Z(n2226) );
  XNOR U2893 ( .A(n2210), .B(n2209), .Z(n2230) );
  XOR U2894 ( .A(n2304), .B(n2206), .Z(n2209) );
  XNOR U2895 ( .A(n2305), .B(n2202), .Z(n2206) );
  AND U2896 ( .A(n2306), .B(n924), .Z(n2202) );
  NAND U2897 ( .A(n2307), .B(n2201), .Z(n2305) );
  NANDN U2898 ( .B(n927), .A(n2311), .Z(n2307) );
  XNOR U2899 ( .A(n2207), .B(n2208), .Z(n2304) );
  XNOR U2900 ( .A(n2315), .B(n2318), .Z(n2317) );
  XNOR U2901 ( .A(n2220), .B(n2219), .Z(n2210) );
  XOR U2902 ( .A(n2319), .B(n2215), .Z(n2219) );
  XNOR U2903 ( .A(n2213), .B(n2320), .Z(n2215) );
  ANDN U2904 ( .A(n2112), .B(n1001), .Z(n2320) );
  XOR U2905 ( .A(n2321), .B(n2322), .Z(n2213) );
  AND U2906 ( .A(n2323), .B(n2324), .Z(n2322) );
  XNOR U2907 ( .A(n2325), .B(n2321), .Z(n2324) );
  AND U2908 ( .A(n2105), .B(n999), .Z(n2217) );
  XNOR U2909 ( .A(n2223), .B(n2224), .Z(n2220) );
  NAND U2910 ( .A(n1910), .B(n1083), .Z(n2224) );
  XNOR U2911 ( .A(n2222), .B(n2329), .Z(n2223) );
  ANDN U2912 ( .A(n1915), .B(n1085), .Z(n2329) );
  XNOR U2913 ( .A(n2229), .B(n2225), .Z(n2303) );
  IV U2914 ( .A(n2228), .Z(n2229) );
  XNOR U2915 ( .A(n2246), .B(n2245), .Z(n2227) );
  XOR U2916 ( .A(n2338), .B(n2254), .Z(n2245) );
  XNOR U2917 ( .A(n2239), .B(n2238), .Z(n2254) );
  XOR U2918 ( .A(n2339), .B(n2235), .Z(n2238) );
  XNOR U2919 ( .A(n2234), .B(n2340), .Z(n2235) );
  ANDN U2920 ( .A(n1404), .B(n1459), .Z(n2340) );
  AND U2921 ( .A(n1457), .B(n1341), .Z(n2236) );
  XNOR U2922 ( .A(n2242), .B(n2243), .Z(n2239) );
  NANDN U2923 ( .B(n1206), .A(n1616), .Z(n2243) );
  XNOR U2924 ( .A(n2241), .B(n2347), .Z(n2242) );
  ANDN U2925 ( .A(n1276), .B(n1618), .Z(n2347) );
  XNOR U2926 ( .A(n2253), .B(n2244), .Z(n2338) );
  XOR U2927 ( .A(n2354), .B(n2262), .Z(n2253) );
  XNOR U2928 ( .A(n2250), .B(n2251), .Z(n2262) );
  NAND U2929 ( .A(n1316), .B(n1575), .Z(n2251) );
  XNOR U2930 ( .A(n2249), .B(n2355), .Z(n2250) );
  ANDN U2931 ( .A(n1582), .B(n1318), .Z(n2355) );
  XNOR U2932 ( .A(n2261), .B(n2252), .Z(n2354) );
  XOR U2933 ( .A(n2362), .B(n2258), .Z(n2261) );
  XNOR U2934 ( .A(n2257), .B(n2363), .Z(n2258) );
  ANDN U2935 ( .A(n1766), .B(n1186), .Z(n2363) );
  AND U2936 ( .A(n1184), .B(n1759), .Z(n2259) );
  XNOR U2937 ( .A(n2270), .B(n2269), .Z(n2246) );
  XOR U2938 ( .A(n2370), .B(n2278), .Z(n2269) );
  XNOR U2939 ( .A(n2266), .B(n2267), .Z(n2278) );
  NANDN U2940 ( .B(n1019), .A(n1984), .Z(n2267) );
  XNOR U2941 ( .A(n2265), .B(n2371), .Z(n2266) );
  ANDN U2942 ( .A(n1060), .B(n1986), .Z(n2371) );
  XNOR U2943 ( .A(n2277), .B(n2268), .Z(n2370) );
  XOR U2944 ( .A(n2378), .B(n2274), .Z(n2277) );
  XNOR U2945 ( .A(n2273), .B(n2379), .Z(n2274) );
  ANDN U2946 ( .A(n1167), .B(n1793), .Z(n2379) );
  AND U2947 ( .A(n1791), .B(n1113), .Z(n2275) );
  XOR U2948 ( .A(n2286), .B(n2285), .Z(n2270) );
  XOR U2949 ( .A(n2386), .B(n2282), .Z(n2285) );
  XNOR U2950 ( .A(n2281), .B(n2387), .Z(n2282) );
  ANDN U2951 ( .A(n992), .B(n2183), .Z(n2387) );
  AND U2952 ( .A(n2181), .B(n951), .Z(n2283) );
  XOR U2953 ( .A(n2293), .B(n2292), .Z(n2286) );
  NAND U2954 ( .A(n2394), .B(n895), .Z(n2292) );
  XNOR U2955 ( .A(n2291), .B(n2395), .Z(n2293) );
  ANDN U2956 ( .A(n926), .B(n2396), .Z(n2395) );
  NAND U2957 ( .A(n2397), .B(n2398), .Z(n2291) );
  NAND U2958 ( .A(n2399), .B(n2400), .Z(n2397) );
  IV U2959 ( .A(n2294), .Z(n2295) );
  MUX U2960 ( .IN0(Y[7]), .IN1(n773), .SEL(n847), .F(n306) );
  XOR U2961 ( .A(n2405), .B(Y0[8]), .Z(n773) );
  XOR U2962 ( .A(n2406), .B(n2407), .Z(n2405) );
  AND U2963 ( .A(n859), .B(n2409), .Z(n2408) );
  XOR U2964 ( .A(n2403), .B(n2407), .Z(n2409) );
  XOR U2965 ( .A(n2402), .B(n2407), .Z(n2403) );
  XNOR U2966 ( .A(n2410), .B(n2337), .Z(n2334) );
  XNOR U2967 ( .A(n2314), .B(n2313), .Z(n2337) );
  XOR U2968 ( .A(n2411), .B(n2318), .Z(n2313) );
  XNOR U2969 ( .A(n2309), .B(n2310), .Z(n2318) );
  NAND U2970 ( .A(n2306), .B(n955), .Z(n2310) );
  XNOR U2971 ( .A(n2308), .B(n2412), .Z(n2309) );
  ANDN U2972 ( .A(n2311), .B(n957), .Z(n2412) );
  XNOR U2973 ( .A(n2316), .B(n2312), .Z(n2411) );
  XOR U2974 ( .A(n2315), .B(n2419), .Z(n2316) );
  AND U2975 ( .A(n2420), .B(n2421), .Z(n2419) );
  NANDN U2976 ( .B(n2422), .A(n894), .Z(n2421) );
  NANDN U2977 ( .B(n2423), .A(n2424), .Z(n2420) );
  XNOR U2978 ( .A(n2328), .B(n2327), .Z(n2314) );
  XOR U2979 ( .A(n2428), .B(n2323), .Z(n2327) );
  XNOR U2980 ( .A(n2321), .B(n2429), .Z(n2323) );
  ANDN U2981 ( .A(n2112), .B(n1041), .Z(n2429) );
  AND U2982 ( .A(n2105), .B(n1039), .Z(n2325) );
  XNOR U2983 ( .A(n2331), .B(n2332), .Z(n2328) );
  NAND U2984 ( .A(n1910), .B(n1125), .Z(n2332) );
  XNOR U2985 ( .A(n2330), .B(n2436), .Z(n2331) );
  ANDN U2986 ( .A(n1915), .B(n1127), .Z(n2436) );
  XNOR U2987 ( .A(n2353), .B(n2352), .Z(n2335) );
  XOR U2988 ( .A(n2446), .B(n2361), .Z(n2352) );
  XNOR U2989 ( .A(n2346), .B(n2345), .Z(n2361) );
  XOR U2990 ( .A(n2447), .B(n2342), .Z(n2345) );
  XNOR U2991 ( .A(n2341), .B(n2448), .Z(n2342) );
  ANDN U2992 ( .A(n1404), .B(n1537), .Z(n2448) );
  AND U2993 ( .A(n1535), .B(n1341), .Z(n2343) );
  XNOR U2994 ( .A(n2349), .B(n2350), .Z(n2346) );
  NANDN U2995 ( .B(n1206), .A(n1700), .Z(n2350) );
  XNOR U2996 ( .A(n2348), .B(n2455), .Z(n2349) );
  ANDN U2997 ( .A(n1276), .B(n1702), .Z(n2455) );
  XNOR U2998 ( .A(n2360), .B(n2351), .Z(n2446) );
  XOR U2999 ( .A(n2462), .B(n2369), .Z(n2360) );
  XNOR U3000 ( .A(n2357), .B(n2358), .Z(n2369) );
  NAND U3001 ( .A(n1383), .B(n1575), .Z(n2358) );
  XNOR U3002 ( .A(n2356), .B(n2463), .Z(n2357) );
  ANDN U3003 ( .A(n1582), .B(n1385), .Z(n2463) );
  XNOR U3004 ( .A(n2368), .B(n2359), .Z(n2462) );
  XOR U3005 ( .A(n2470), .B(n2365), .Z(n2368) );
  XNOR U3006 ( .A(n2364), .B(n2471), .Z(n2365) );
  ANDN U3007 ( .A(n1766), .B(n1250), .Z(n2471) );
  AND U3008 ( .A(n1248), .B(n1759), .Z(n2366) );
  XNOR U3009 ( .A(n2377), .B(n2376), .Z(n2353) );
  XOR U3010 ( .A(n2478), .B(n2385), .Z(n2376) );
  XNOR U3011 ( .A(n2373), .B(n2374), .Z(n2385) );
  NANDN U3012 ( .B(n1019), .A(n2080), .Z(n2374) );
  XNOR U3013 ( .A(n2372), .B(n2479), .Z(n2373) );
  ANDN U3014 ( .A(n1060), .B(n2082), .Z(n2479) );
  XNOR U3015 ( .A(n2384), .B(n2375), .Z(n2478) );
  XOR U3016 ( .A(n2486), .B(n2381), .Z(n2384) );
  XNOR U3017 ( .A(n2380), .B(n2487), .Z(n2381) );
  ANDN U3018 ( .A(n1167), .B(n1890), .Z(n2487) );
  AND U3019 ( .A(n1888), .B(n1113), .Z(n2382) );
  XOR U3020 ( .A(n2393), .B(n2392), .Z(n2377) );
  XOR U3021 ( .A(n2494), .B(n2389), .Z(n2392) );
  XNOR U3022 ( .A(n2388), .B(n2495), .Z(n2389) );
  ANDN U3023 ( .A(n992), .B(n2289), .Z(n2495) );
  AND U3024 ( .A(n2287), .B(n951), .Z(n2390) );
  XOR U3025 ( .A(n2400), .B(n2399), .Z(n2393) );
  NAND U3026 ( .A(n2502), .B(n895), .Z(n2399) );
  XOR U3027 ( .A(n2398), .B(n2503), .Z(n2400) );
  ANDN U3028 ( .A(n926), .B(n2504), .Z(n2503) );
  ANDN U3029 ( .A(n2505), .B(n2506), .Z(n2398) );
  NAND U3030 ( .A(n2507), .B(n2508), .Z(n2505) );
  IV U3031 ( .A(n2401), .Z(n2402) );
  MUX U3032 ( .IN0(Y[6]), .IN1(n770), .SEL(n847), .F(n305) );
  XOR U3033 ( .A(n2513), .B(Y0[7]), .Z(n770) );
  XOR U3034 ( .A(n2514), .B(n2515), .Z(n2513) );
  AND U3035 ( .A(n859), .B(n2517), .Z(n2516) );
  XOR U3036 ( .A(n2511), .B(n2515), .Z(n2517) );
  XOR U3037 ( .A(n2510), .B(n2515), .Z(n2511) );
  XNOR U3038 ( .A(n2518), .B(n2445), .Z(n2441) );
  XNOR U3039 ( .A(n2418), .B(n2417), .Z(n2445) );
  XOR U3040 ( .A(n2519), .B(n2427), .Z(n2417) );
  XNOR U3041 ( .A(n2414), .B(n2415), .Z(n2427) );
  NAND U3042 ( .A(n2306), .B(n999), .Z(n2415) );
  XNOR U3043 ( .A(n2413), .B(n2520), .Z(n2414) );
  ANDN U3044 ( .A(n2311), .B(n1001), .Z(n2520) );
  XOR U3045 ( .A(n2521), .B(n2522), .Z(n2413) );
  AND U3046 ( .A(n2523), .B(n2524), .Z(n2522) );
  XOR U3047 ( .A(n2525), .B(n2521), .Z(n2524) );
  XNOR U3048 ( .A(n2426), .B(n2416), .Z(n2519) );
  XOR U3049 ( .A(n2533), .B(n2424), .Z(n2529) );
  AND U3050 ( .A(n2534), .B(n924), .Z(n2424) );
  NAND U3051 ( .A(n2535), .B(n2423), .Z(n2533) );
  XOR U3052 ( .A(n2536), .B(n2537), .Z(n2423) );
  AND U3053 ( .A(n2538), .B(n2539), .Z(n2537) );
  XNOR U3054 ( .A(n2540), .B(n2536), .Z(n2539) );
  NANDN U3055 ( .B(n927), .A(n2541), .Z(n2535) );
  XNOR U3056 ( .A(n2435), .B(n2434), .Z(n2418) );
  XOR U3057 ( .A(n2542), .B(n2431), .Z(n2434) );
  XNOR U3058 ( .A(n2430), .B(n2543), .Z(n2431) );
  ANDN U3059 ( .A(n2112), .B(n1085), .Z(n2543) );
  AND U3060 ( .A(n2105), .B(n1083), .Z(n2432) );
  XNOR U3061 ( .A(n2438), .B(n2439), .Z(n2435) );
  NAND U3062 ( .A(n1910), .B(n1184), .Z(n2439) );
  XNOR U3063 ( .A(n2437), .B(n2550), .Z(n2438) );
  ANDN U3064 ( .A(n1915), .B(n1186), .Z(n2550) );
  XNOR U3065 ( .A(n2444), .B(n2440), .Z(n2518) );
  XOR U3066 ( .A(n2561), .B(n2562), .Z(n2557) );
  NANDN U3067 ( .B(n2563), .A(n2564), .Z(n2561) );
  XNOR U3068 ( .A(n2461), .B(n2460), .Z(n2442) );
  XOR U3069 ( .A(n2565), .B(n2469), .Z(n2460) );
  XNOR U3070 ( .A(n2454), .B(n2453), .Z(n2469) );
  XOR U3071 ( .A(n2566), .B(n2450), .Z(n2453) );
  XNOR U3072 ( .A(n2449), .B(n2567), .Z(n2450) );
  ANDN U3073 ( .A(n1404), .B(n1618), .Z(n2567) );
  AND U3074 ( .A(n1616), .B(n1341), .Z(n2451) );
  XNOR U3075 ( .A(n2457), .B(n2458), .Z(n2454) );
  NANDN U3076 ( .B(n1206), .A(n1791), .Z(n2458) );
  XNOR U3077 ( .A(n2456), .B(n2574), .Z(n2457) );
  ANDN U3078 ( .A(n1276), .B(n1793), .Z(n2574) );
  XNOR U3079 ( .A(n2468), .B(n2459), .Z(n2565) );
  XOR U3080 ( .A(n2581), .B(n2477), .Z(n2468) );
  XNOR U3081 ( .A(n2465), .B(n2466), .Z(n2477) );
  NAND U3082 ( .A(n1457), .B(n1575), .Z(n2466) );
  XNOR U3083 ( .A(n2464), .B(n2582), .Z(n2465) );
  ANDN U3084 ( .A(n1582), .B(n1459), .Z(n2582) );
  XNOR U3085 ( .A(n2476), .B(n2467), .Z(n2581) );
  XOR U3086 ( .A(n2589), .B(n2473), .Z(n2476) );
  XNOR U3087 ( .A(n2472), .B(n2590), .Z(n2473) );
  ANDN U3088 ( .A(n1766), .B(n1318), .Z(n2590) );
  AND U3089 ( .A(n1316), .B(n1759), .Z(n2474) );
  XNOR U3090 ( .A(n2485), .B(n2484), .Z(n2461) );
  XOR U3091 ( .A(n2597), .B(n2493), .Z(n2484) );
  XNOR U3092 ( .A(n2481), .B(n2482), .Z(n2493) );
  NANDN U3093 ( .B(n1019), .A(n2181), .Z(n2482) );
  XNOR U3094 ( .A(n2480), .B(n2598), .Z(n2481) );
  ANDN U3095 ( .A(n1060), .B(n2183), .Z(n2598) );
  XNOR U3096 ( .A(n2492), .B(n2483), .Z(n2597) );
  XOR U3097 ( .A(n2605), .B(n2489), .Z(n2492) );
  XNOR U3098 ( .A(n2488), .B(n2606), .Z(n2489) );
  ANDN U3099 ( .A(n1167), .B(n1986), .Z(n2606) );
  AND U3100 ( .A(n1984), .B(n1113), .Z(n2490) );
  XOR U3101 ( .A(n2501), .B(n2500), .Z(n2485) );
  XOR U3102 ( .A(n2613), .B(n2497), .Z(n2500) );
  XNOR U3103 ( .A(n2496), .B(n2614), .Z(n2497) );
  ANDN U3104 ( .A(n992), .B(n2396), .Z(n2614) );
  AND U3105 ( .A(n2394), .B(n951), .Z(n2498) );
  XOR U3106 ( .A(n2508), .B(n2507), .Z(n2501) );
  NAND U3107 ( .A(n2621), .B(n895), .Z(n2507) );
  XNOR U3108 ( .A(n2506), .B(n2622), .Z(n2508) );
  ANDN U3109 ( .A(n926), .B(n2623), .Z(n2622) );
  NAND U3110 ( .A(n2624), .B(n2625), .Z(n2506) );
  NAND U3111 ( .A(n2626), .B(n2627), .Z(n2624) );
  IV U3112 ( .A(n2509), .Z(n2510) );
  MUX U3113 ( .IN0(Y[5]), .IN1(n767), .SEL(n847), .F(n304) );
  XOR U3114 ( .A(n2632), .B(Y0[6]), .Z(n767) );
  XOR U3115 ( .A(n2633), .B(n2634), .Z(n2632) );
  AND U3116 ( .A(n859), .B(n2636), .Z(n2635) );
  XOR U3117 ( .A(n2630), .B(n2634), .Z(n2636) );
  XOR U3118 ( .A(n2629), .B(n2634), .Z(n2630) );
  XNOR U3119 ( .A(n2637), .B(n2560), .Z(n2555) );
  XNOR U3120 ( .A(n2528), .B(n2527), .Z(n2560) );
  XOR U3121 ( .A(n2638), .B(n2532), .Z(n2527) );
  XNOR U3122 ( .A(n2523), .B(n2525), .Z(n2532) );
  NAND U3123 ( .A(n2306), .B(n1039), .Z(n2525) );
  XNOR U3124 ( .A(n2521), .B(n2639), .Z(n2523) );
  ANDN U3125 ( .A(n2311), .B(n1041), .Z(n2639) );
  XNOR U3126 ( .A(n2531), .B(n2526), .Z(n2638) );
  XOR U3127 ( .A(n2646), .B(n2538), .Z(n2531) );
  XNOR U3128 ( .A(n2536), .B(n2647), .Z(n2538) );
  ANDN U3129 ( .A(n2541), .B(n957), .Z(n2647) );
  XOR U3130 ( .A(n2648), .B(n2649), .Z(n2536) );
  AND U3131 ( .A(n2650), .B(n2651), .Z(n2649) );
  XNOR U3132 ( .A(n2652), .B(n2648), .Z(n2651) );
  AND U3133 ( .A(n2534), .B(n955), .Z(n2540) );
  XNOR U3134 ( .A(n2549), .B(n2548), .Z(n2528) );
  XOR U3135 ( .A(n2656), .B(n2545), .Z(n2548) );
  XNOR U3136 ( .A(n2544), .B(n2657), .Z(n2545) );
  ANDN U3137 ( .A(n2112), .B(n1127), .Z(n2657) );
  AND U3138 ( .A(n2105), .B(n1125), .Z(n2546) );
  XNOR U3139 ( .A(n2552), .B(n2553), .Z(n2549) );
  NAND U3140 ( .A(n1910), .B(n1248), .Z(n2553) );
  XNOR U3141 ( .A(n2551), .B(n2664), .Z(n2552) );
  ANDN U3142 ( .A(n1915), .B(n1250), .Z(n2664) );
  XNOR U3143 ( .A(n2559), .B(n2554), .Z(n2637) );
  XOR U3144 ( .A(n2558), .B(n2671), .Z(n2559) );
  AND U3145 ( .A(n2562), .B(n2672), .Z(n2671) );
  AND U3146 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U3147 ( .B(n2675), .A(n894), .Z(n2674) );
  NAND U3148 ( .A(n2676), .B(n2677), .Z(n2673) );
  ANDN U3149 ( .A(n2564), .B(n2563), .Z(n2562) );
  ANDN U3150 ( .A(n2678), .B(n2679), .Z(n2563) );
  OR U3151 ( .A(n2680), .B(n2681), .Z(n2564) );
  XNOR U3152 ( .A(n2580), .B(n2579), .Z(n2556) );
  XOR U3153 ( .A(n2685), .B(n2588), .Z(n2579) );
  XNOR U3154 ( .A(n2573), .B(n2572), .Z(n2588) );
  XOR U3155 ( .A(n2686), .B(n2569), .Z(n2572) );
  XNOR U3156 ( .A(n2568), .B(n2687), .Z(n2569) );
  ANDN U3157 ( .A(n1404), .B(n1702), .Z(n2687) );
  AND U3158 ( .A(n1700), .B(n1341), .Z(n2570) );
  XNOR U3159 ( .A(n2576), .B(n2577), .Z(n2573) );
  NANDN U3160 ( .B(n1206), .A(n1888), .Z(n2577) );
  XNOR U3161 ( .A(n2575), .B(n2694), .Z(n2576) );
  ANDN U3162 ( .A(n1276), .B(n1890), .Z(n2694) );
  XNOR U3163 ( .A(n2587), .B(n2578), .Z(n2685) );
  XOR U3164 ( .A(n2701), .B(n2596), .Z(n2587) );
  XNOR U3165 ( .A(n2584), .B(n2585), .Z(n2596) );
  NAND U3166 ( .A(n1535), .B(n1575), .Z(n2585) );
  XNOR U3167 ( .A(n2583), .B(n2702), .Z(n2584) );
  ANDN U3168 ( .A(n1582), .B(n1537), .Z(n2702) );
  XNOR U3169 ( .A(n2595), .B(n2586), .Z(n2701) );
  XOR U3170 ( .A(n2709), .B(n2592), .Z(n2595) );
  XNOR U3171 ( .A(n2591), .B(n2710), .Z(n2592) );
  ANDN U3172 ( .A(n1766), .B(n1385), .Z(n2710) );
  AND U3173 ( .A(n1383), .B(n1759), .Z(n2593) );
  XNOR U3174 ( .A(n2604), .B(n2603), .Z(n2580) );
  XOR U3175 ( .A(n2717), .B(n2612), .Z(n2603) );
  XNOR U3176 ( .A(n2600), .B(n2601), .Z(n2612) );
  NANDN U3177 ( .B(n1019), .A(n2287), .Z(n2601) );
  XNOR U3178 ( .A(n2599), .B(n2718), .Z(n2600) );
  ANDN U3179 ( .A(n1060), .B(n2289), .Z(n2718) );
  XNOR U3180 ( .A(n2611), .B(n2602), .Z(n2717) );
  XOR U3181 ( .A(n2725), .B(n2608), .Z(n2611) );
  XNOR U3182 ( .A(n2607), .B(n2726), .Z(n2608) );
  ANDN U3183 ( .A(n1167), .B(n2082), .Z(n2726) );
  AND U3184 ( .A(n2080), .B(n1113), .Z(n2609) );
  XOR U3185 ( .A(n2620), .B(n2619), .Z(n2604) );
  XOR U3186 ( .A(n2733), .B(n2616), .Z(n2619) );
  XNOR U3187 ( .A(n2615), .B(n2734), .Z(n2616) );
  ANDN U3188 ( .A(n992), .B(n2504), .Z(n2734) );
  AND U3189 ( .A(n2502), .B(n951), .Z(n2617) );
  XOR U3190 ( .A(n2627), .B(n2626), .Z(n2620) );
  NAND U3191 ( .A(n2741), .B(n895), .Z(n2626) );
  XOR U3192 ( .A(n2625), .B(n2742), .Z(n2627) );
  ANDN U3193 ( .A(n926), .B(n2743), .Z(n2742) );
  ANDN U3194 ( .A(n2744), .B(n2745), .Z(n2625) );
  NAND U3195 ( .A(n2746), .B(n2747), .Z(n2744) );
  IV U3196 ( .A(n2628), .Z(n2629) );
  MUX U3197 ( .IN0(Y[4]), .IN1(n764), .SEL(n847), .F(n303) );
  XOR U3198 ( .A(n2752), .B(Y0[5]), .Z(n764) );
  XOR U3199 ( .A(n2753), .B(n2754), .Z(n2752) );
  AND U3200 ( .A(n859), .B(n2756), .Z(n2755) );
  XOR U3201 ( .A(n2750), .B(n2754), .Z(n2756) );
  XOR U3202 ( .A(n2749), .B(n2754), .Z(n2750) );
  XNOR U3203 ( .A(n2757), .B(n2684), .Z(n2669) );
  XNOR U3204 ( .A(n2645), .B(n2644), .Z(n2684) );
  XOR U3205 ( .A(n2758), .B(n2655), .Z(n2644) );
  XNOR U3206 ( .A(n2641), .B(n2642), .Z(n2655) );
  NAND U3207 ( .A(n2306), .B(n1083), .Z(n2642) );
  XNOR U3208 ( .A(n2640), .B(n2759), .Z(n2641) );
  ANDN U3209 ( .A(n2311), .B(n1085), .Z(n2759) );
  XNOR U3210 ( .A(n2654), .B(n2643), .Z(n2758) );
  XOR U3211 ( .A(n2766), .B(n2650), .Z(n2654) );
  XNOR U3212 ( .A(n2648), .B(n2767), .Z(n2650) );
  ANDN U3213 ( .A(n2541), .B(n1001), .Z(n2767) );
  XOR U3214 ( .A(n2768), .B(n2769), .Z(n2648) );
  AND U3215 ( .A(n2770), .B(n2771), .Z(n2769) );
  XNOR U3216 ( .A(n2772), .B(n2768), .Z(n2771) );
  AND U3217 ( .A(n2534), .B(n999), .Z(n2652) );
  XNOR U3218 ( .A(n2663), .B(n2662), .Z(n2645) );
  XOR U3219 ( .A(n2776), .B(n2659), .Z(n2662) );
  XNOR U3220 ( .A(n2658), .B(n2777), .Z(n2659) );
  ANDN U3221 ( .A(n2112), .B(n1186), .Z(n2777) );
  AND U3222 ( .A(n2105), .B(n1184), .Z(n2660) );
  XNOR U3223 ( .A(n2666), .B(n2667), .Z(n2663) );
  NAND U3224 ( .A(n1910), .B(n1316), .Z(n2667) );
  XNOR U3225 ( .A(n2665), .B(n2784), .Z(n2666) );
  ANDN U3226 ( .A(n1915), .B(n1318), .Z(n2784) );
  XOR U3227 ( .A(n2683), .B(n2668), .Z(n2757) );
  XOR U3228 ( .A(n2791), .B(n2676), .Z(n2683) );
  XOR U3229 ( .A(n2795), .B(n2681), .Z(n2679) );
  NAND U3230 ( .A(n2796), .B(n924), .Z(n2681) );
  NAND U3231 ( .A(n2797), .B(n2680), .Z(n2795) );
  NANDN U3232 ( .B(n927), .A(n2801), .Z(n2797) );
  ANDN U3233 ( .A(n2802), .B(n2803), .Z(n2677) );
  XNOR U3234 ( .A(n2700), .B(n2699), .Z(n2670) );
  XOR U3235 ( .A(n2807), .B(n2708), .Z(n2699) );
  XNOR U3236 ( .A(n2693), .B(n2692), .Z(n2708) );
  XOR U3237 ( .A(n2808), .B(n2689), .Z(n2692) );
  XNOR U3238 ( .A(n2688), .B(n2809), .Z(n2689) );
  ANDN U3239 ( .A(n1404), .B(n1793), .Z(n2809) );
  AND U3240 ( .A(n1791), .B(n1341), .Z(n2690) );
  XNOR U3241 ( .A(n2696), .B(n2697), .Z(n2693) );
  NANDN U3242 ( .B(n1206), .A(n1984), .Z(n2697) );
  XNOR U3243 ( .A(n2695), .B(n2816), .Z(n2696) );
  ANDN U3244 ( .A(n1276), .B(n1986), .Z(n2816) );
  XNOR U3245 ( .A(n2707), .B(n2698), .Z(n2807) );
  XOR U3246 ( .A(n2823), .B(n2716), .Z(n2707) );
  XNOR U3247 ( .A(n2704), .B(n2705), .Z(n2716) );
  NAND U3248 ( .A(n1616), .B(n1575), .Z(n2705) );
  XNOR U3249 ( .A(n2703), .B(n2824), .Z(n2704) );
  ANDN U3250 ( .A(n1582), .B(n1618), .Z(n2824) );
  XNOR U3251 ( .A(n2715), .B(n2706), .Z(n2823) );
  XOR U3252 ( .A(n2831), .B(n2712), .Z(n2715) );
  XNOR U3253 ( .A(n2711), .B(n2832), .Z(n2712) );
  ANDN U3254 ( .A(n1766), .B(n1459), .Z(n2832) );
  AND U3255 ( .A(n1457), .B(n1759), .Z(n2713) );
  XNOR U3256 ( .A(n2724), .B(n2723), .Z(n2700) );
  XOR U3257 ( .A(n2839), .B(n2732), .Z(n2723) );
  XNOR U3258 ( .A(n2720), .B(n2721), .Z(n2732) );
  NANDN U3259 ( .B(n1019), .A(n2394), .Z(n2721) );
  XNOR U3260 ( .A(n2719), .B(n2840), .Z(n2720) );
  ANDN U3261 ( .A(n1060), .B(n2396), .Z(n2840) );
  XNOR U3262 ( .A(n2731), .B(n2722), .Z(n2839) );
  XOR U3263 ( .A(n2847), .B(n2728), .Z(n2731) );
  XNOR U3264 ( .A(n2727), .B(n2848), .Z(n2728) );
  ANDN U3265 ( .A(n1167), .B(n2183), .Z(n2848) );
  AND U3266 ( .A(n2181), .B(n1113), .Z(n2729) );
  XOR U3267 ( .A(n2740), .B(n2739), .Z(n2724) );
  XOR U3268 ( .A(n2855), .B(n2736), .Z(n2739) );
  XNOR U3269 ( .A(n2735), .B(n2856), .Z(n2736) );
  ANDN U3270 ( .A(n992), .B(n2623), .Z(n2856) );
  AND U3271 ( .A(n2621), .B(n951), .Z(n2737) );
  XOR U3272 ( .A(n2747), .B(n2746), .Z(n2740) );
  NAND U3273 ( .A(n2863), .B(n895), .Z(n2746) );
  XNOR U3274 ( .A(n2745), .B(n2864), .Z(n2747) );
  ANDN U3275 ( .A(n926), .B(n2865), .Z(n2864) );
  NAND U3276 ( .A(n2866), .B(n2867), .Z(n2745) );
  NAND U3277 ( .A(n2868), .B(n2869), .Z(n2866) );
  IV U3278 ( .A(n2748), .Z(n2749) );
  MUX U3279 ( .IN0(Y[3]), .IN1(n761), .SEL(n847), .F(n302) );
  XNOR U3280 ( .A(n2873), .B(Y0[4]), .Z(n761) );
  XNOR U3281 ( .A(n2875), .B(n2876), .Z(n2873) );
  XOR U3282 ( .A(n2874), .B(n2877), .Z(n2875) );
  AND U3283 ( .A(n859), .B(n2878), .Z(n2877) );
  XNOR U3284 ( .A(n2871), .B(n2876), .Z(n2878) );
  XOR U3285 ( .A(n2876), .B(n2870), .Z(n2871) );
  NOR U3286 ( .A(n2879), .B(n2880), .Z(n2870) );
  XNOR U3287 ( .A(n2881), .B(n2806), .Z(n2789) );
  XNOR U3288 ( .A(n2765), .B(n2764), .Z(n2806) );
  XOR U3289 ( .A(n2882), .B(n2775), .Z(n2764) );
  XNOR U3290 ( .A(n2761), .B(n2762), .Z(n2775) );
  NAND U3291 ( .A(n2306), .B(n1125), .Z(n2762) );
  XNOR U3292 ( .A(n2760), .B(n2883), .Z(n2761) );
  ANDN U3293 ( .A(n2311), .B(n1127), .Z(n2883) );
  XNOR U3294 ( .A(n2774), .B(n2763), .Z(n2882) );
  XOR U3295 ( .A(n2890), .B(n2770), .Z(n2774) );
  XNOR U3296 ( .A(n2768), .B(n2891), .Z(n2770) );
  ANDN U3297 ( .A(n2541), .B(n1041), .Z(n2891) );
  AND U3298 ( .A(n2534), .B(n1039), .Z(n2772) );
  XNOR U3299 ( .A(n2783), .B(n2782), .Z(n2765) );
  XOR U3300 ( .A(n2898), .B(n2779), .Z(n2782) );
  XNOR U3301 ( .A(n2778), .B(n2899), .Z(n2779) );
  ANDN U3302 ( .A(n2112), .B(n1250), .Z(n2899) );
  AND U3303 ( .A(n2105), .B(n1248), .Z(n2780) );
  XNOR U3304 ( .A(n2786), .B(n2787), .Z(n2783) );
  NAND U3305 ( .A(n1910), .B(n1383), .Z(n2787) );
  XNOR U3306 ( .A(n2785), .B(n2906), .Z(n2786) );
  ANDN U3307 ( .A(n1915), .B(n1385), .Z(n2906) );
  XNOR U3308 ( .A(n2805), .B(n2788), .Z(n2881) );
  XOR U3309 ( .A(n2913), .B(n2803), .Z(n2805) );
  XOR U3310 ( .A(n2794), .B(n2793), .Z(n2803) );
  XNOR U3311 ( .A(n2792), .B(n2914), .Z(n2793) );
  AND U3312 ( .A(n2915), .B(n2916), .Z(n2914) );
  NANDN U3313 ( .B(n2917), .A(n894), .Z(n2916) );
  NANDN U3314 ( .B(n2918), .A(n2919), .Z(n2915) );
  XNOR U3315 ( .A(n2799), .B(n2800), .Z(n2794) );
  NAND U3316 ( .A(n2796), .B(n955), .Z(n2800) );
  XNOR U3317 ( .A(n2798), .B(n2923), .Z(n2799) );
  ANDN U3318 ( .A(n2801), .B(n957), .Z(n2923) );
  NOR U3319 ( .A(n2927), .B(n2928), .Z(n2802) );
  XNOR U3320 ( .A(n2822), .B(n2821), .Z(n2790) );
  XOR U3321 ( .A(n2932), .B(n2830), .Z(n2821) );
  XNOR U3322 ( .A(n2815), .B(n2814), .Z(n2830) );
  XOR U3323 ( .A(n2933), .B(n2811), .Z(n2814) );
  XNOR U3324 ( .A(n2810), .B(n2934), .Z(n2811) );
  ANDN U3325 ( .A(n1404), .B(n1890), .Z(n2934) );
  AND U3326 ( .A(n1888), .B(n1341), .Z(n2812) );
  XNOR U3327 ( .A(n2818), .B(n2819), .Z(n2815) );
  NANDN U3328 ( .B(n1206), .A(n2080), .Z(n2819) );
  XNOR U3329 ( .A(n2817), .B(n2941), .Z(n2818) );
  ANDN U3330 ( .A(n1276), .B(n2082), .Z(n2941) );
  XNOR U3331 ( .A(n2829), .B(n2820), .Z(n2932) );
  XOR U3332 ( .A(n2948), .B(n2838), .Z(n2829) );
  XNOR U3333 ( .A(n2826), .B(n2827), .Z(n2838) );
  NAND U3334 ( .A(n1700), .B(n1575), .Z(n2827) );
  XNOR U3335 ( .A(n2825), .B(n2949), .Z(n2826) );
  ANDN U3336 ( .A(n1582), .B(n1702), .Z(n2949) );
  XNOR U3337 ( .A(n2837), .B(n2828), .Z(n2948) );
  XOR U3338 ( .A(n2956), .B(n2834), .Z(n2837) );
  XNOR U3339 ( .A(n2833), .B(n2957), .Z(n2834) );
  ANDN U3340 ( .A(n1766), .B(n1537), .Z(n2957) );
  AND U3341 ( .A(n1535), .B(n1759), .Z(n2835) );
  XNOR U3342 ( .A(n2846), .B(n2845), .Z(n2822) );
  XOR U3343 ( .A(n2964), .B(n2854), .Z(n2845) );
  XNOR U3344 ( .A(n2842), .B(n2843), .Z(n2854) );
  NANDN U3345 ( .B(n1019), .A(n2502), .Z(n2843) );
  XNOR U3346 ( .A(n2841), .B(n2965), .Z(n2842) );
  ANDN U3347 ( .A(n1060), .B(n2504), .Z(n2965) );
  XNOR U3348 ( .A(n2853), .B(n2844), .Z(n2964) );
  XOR U3349 ( .A(n2972), .B(n2850), .Z(n2853) );
  XNOR U3350 ( .A(n2849), .B(n2973), .Z(n2850) );
  ANDN U3351 ( .A(n1167), .B(n2289), .Z(n2973) );
  AND U3352 ( .A(n2287), .B(n1113), .Z(n2851) );
  XOR U3353 ( .A(n2862), .B(n2861), .Z(n2846) );
  XOR U3354 ( .A(n2980), .B(n2858), .Z(n2861) );
  XNOR U3355 ( .A(n2857), .B(n2981), .Z(n2858) );
  ANDN U3356 ( .A(n992), .B(n2743), .Z(n2981) );
  AND U3357 ( .A(n2741), .B(n951), .Z(n2859) );
  XOR U3358 ( .A(n2869), .B(n2868), .Z(n2862) );
  NAND U3359 ( .A(n2988), .B(n895), .Z(n2868) );
  XOR U3360 ( .A(n2867), .B(n2989), .Z(n2869) );
  ANDN U3361 ( .A(n926), .B(n2990), .Z(n2989) );
  ANDN U3362 ( .A(n2991), .B(n2992), .Z(n2867) );
  NAND U3363 ( .A(n2993), .B(n2994), .Z(n2991) );
  IV U3364 ( .A(n2872), .Z(n2874) );
  MUX U3365 ( .IN0(Y[2]), .IN1(n758), .SEL(n847), .F(n301) );
  IV U3366 ( .A(n2998), .Z(n847) );
  XNOR U3367 ( .A(n2996), .B(Y0[3]), .Z(n758) );
  XNOR U3368 ( .A(n2999), .B(n3000), .Z(n2996) );
  XOR U3369 ( .A(n2997), .B(n3001), .Z(n2999) );
  AND U3370 ( .A(n859), .B(n3002), .Z(n3001) );
  XNOR U3371 ( .A(n2880), .B(n3000), .Z(n3002) );
  NANDN U3372 ( .B(n3003), .A(n3004), .Z(n2879) );
  XNOR U3373 ( .A(n3005), .B(n2931), .Z(n2911) );
  XNOR U3374 ( .A(n2889), .B(n2888), .Z(n2931) );
  XOR U3375 ( .A(n3006), .B(n2897), .Z(n2888) );
  XNOR U3376 ( .A(n2885), .B(n2886), .Z(n2897) );
  NAND U3377 ( .A(n2306), .B(n1184), .Z(n2886) );
  XNOR U3378 ( .A(n2884), .B(n3007), .Z(n2885) );
  ANDN U3379 ( .A(n2311), .B(n1186), .Z(n3007) );
  XNOR U3380 ( .A(n2896), .B(n2887), .Z(n3006) );
  XOR U3381 ( .A(n3014), .B(n2893), .Z(n2896) );
  XNOR U3382 ( .A(n2892), .B(n3015), .Z(n2893) );
  ANDN U3383 ( .A(n2541), .B(n1085), .Z(n3015) );
  AND U3384 ( .A(n2534), .B(n1083), .Z(n2894) );
  XNOR U3385 ( .A(n2905), .B(n2904), .Z(n2889) );
  XOR U3386 ( .A(n3022), .B(n2901), .Z(n2904) );
  XNOR U3387 ( .A(n2900), .B(n3023), .Z(n2901) );
  ANDN U3388 ( .A(n2112), .B(n1318), .Z(n3023) );
  AND U3389 ( .A(n2105), .B(n1316), .Z(n2902) );
  XNOR U3390 ( .A(n2908), .B(n2909), .Z(n2905) );
  NAND U3391 ( .A(n1910), .B(n1457), .Z(n2909) );
  XNOR U3392 ( .A(n2907), .B(n3030), .Z(n2908) );
  ANDN U3393 ( .A(n1915), .B(n1459), .Z(n3030) );
  XNOR U3394 ( .A(n2930), .B(n2910), .Z(n3005) );
  XOR U3395 ( .A(n3037), .B(n2928), .Z(n2930) );
  XOR U3396 ( .A(n2922), .B(n2921), .Z(n2928) );
  XOR U3397 ( .A(n3042), .B(n2919), .Z(n3038) );
  AND U3398 ( .A(n3043), .B(n924), .Z(n2919) );
  NAND U3399 ( .A(n3044), .B(n2918), .Z(n3042) );
  XOR U3400 ( .A(n3045), .B(n3046), .Z(n2918) );
  AND U3401 ( .A(n3047), .B(n3048), .Z(n3046) );
  XNOR U3402 ( .A(n3049), .B(n3045), .Z(n3048) );
  NANDN U3403 ( .B(n927), .A(n3050), .Z(n3044) );
  XNOR U3404 ( .A(n2925), .B(n2926), .Z(n2922) );
  NAND U3405 ( .A(n2796), .B(n999), .Z(n2926) );
  XNOR U3406 ( .A(n2924), .B(n3051), .Z(n2925) );
  ANDN U3407 ( .A(n2801), .B(n1001), .Z(n3051) );
  XOR U3408 ( .A(n3052), .B(n3053), .Z(n2924) );
  AND U3409 ( .A(n3054), .B(n3055), .Z(n3053) );
  XOR U3410 ( .A(n3056), .B(n3052), .Z(n3055) );
  XNOR U3411 ( .A(n2927), .B(n2929), .Z(n3037) );
  XNOR U3412 ( .A(n3060), .B(n3063), .Z(n3062) );
  XNOR U3413 ( .A(n2947), .B(n2946), .Z(n2912) );
  XOR U3414 ( .A(n3064), .B(n2955), .Z(n2946) );
  XNOR U3415 ( .A(n2940), .B(n2939), .Z(n2955) );
  XOR U3416 ( .A(n3065), .B(n2936), .Z(n2939) );
  XNOR U3417 ( .A(n2935), .B(n3066), .Z(n2936) );
  ANDN U3418 ( .A(n1404), .B(n1986), .Z(n3066) );
  AND U3419 ( .A(n1984), .B(n1341), .Z(n2937) );
  XNOR U3420 ( .A(n2943), .B(n2944), .Z(n2940) );
  NANDN U3421 ( .B(n1206), .A(n2181), .Z(n2944) );
  XNOR U3422 ( .A(n2942), .B(n3073), .Z(n2943) );
  ANDN U3423 ( .A(n1276), .B(n2183), .Z(n3073) );
  XNOR U3424 ( .A(n2954), .B(n2945), .Z(n3064) );
  XOR U3425 ( .A(n3080), .B(n2963), .Z(n2954) );
  XNOR U3426 ( .A(n2951), .B(n2952), .Z(n2963) );
  NAND U3427 ( .A(n1791), .B(n1575), .Z(n2952) );
  XNOR U3428 ( .A(n2950), .B(n3081), .Z(n2951) );
  ANDN U3429 ( .A(n1582), .B(n1793), .Z(n3081) );
  XNOR U3430 ( .A(n2962), .B(n2953), .Z(n3080) );
  XOR U3431 ( .A(n3088), .B(n2959), .Z(n2962) );
  XNOR U3432 ( .A(n2958), .B(n3089), .Z(n2959) );
  ANDN U3433 ( .A(n1766), .B(n1618), .Z(n3089) );
  AND U3434 ( .A(n1616), .B(n1759), .Z(n2960) );
  XNOR U3435 ( .A(n2971), .B(n2970), .Z(n2947) );
  XOR U3436 ( .A(n3096), .B(n2979), .Z(n2970) );
  XNOR U3437 ( .A(n2967), .B(n2968), .Z(n2979) );
  NANDN U3438 ( .B(n1019), .A(n2621), .Z(n2968) );
  XNOR U3439 ( .A(n2966), .B(n3097), .Z(n2967) );
  ANDN U3440 ( .A(n1060), .B(n2623), .Z(n3097) );
  XNOR U3441 ( .A(n2978), .B(n2969), .Z(n3096) );
  XOR U3442 ( .A(n3104), .B(n2975), .Z(n2978) );
  XNOR U3443 ( .A(n2974), .B(n3105), .Z(n2975) );
  ANDN U3444 ( .A(n1167), .B(n2396), .Z(n3105) );
  AND U3445 ( .A(n2394), .B(n1113), .Z(n2976) );
  XOR U3446 ( .A(n2987), .B(n2986), .Z(n2971) );
  XOR U3447 ( .A(n3112), .B(n2983), .Z(n2986) );
  XNOR U3448 ( .A(n2982), .B(n3113), .Z(n2983) );
  ANDN U3449 ( .A(n992), .B(n2865), .Z(n3113) );
  AND U3450 ( .A(n2863), .B(n951), .Z(n2984) );
  XOR U3451 ( .A(n2994), .B(n2993), .Z(n2987) );
  NAND U3452 ( .A(n3120), .B(n895), .Z(n2993) );
  XNOR U3453 ( .A(n2992), .B(n3121), .Z(n2994) );
  ANDN U3454 ( .A(n926), .B(n3122), .Z(n3121) );
  NAND U3455 ( .A(n3123), .B(n3124), .Z(n2992) );
  NAND U3456 ( .A(n3125), .B(n3126), .Z(n3123) );
  IV U3457 ( .A(n2995), .Z(n2997) );
  MUX U3458 ( .IN0(n755), .IN1(Y[1]), .SEL(n2998), .F(n300) );
  XNOR U3459 ( .A(n3128), .B(Y0[2]), .Z(n755) );
  XNOR U3460 ( .A(n3129), .B(n3130), .Z(n3128) );
  XNOR U3461 ( .A(n3127), .B(n3131), .Z(n3129) );
  AND U3462 ( .A(n859), .B(n3132), .Z(n3131) );
  XNOR U3463 ( .A(n3003), .B(n3130), .Z(n3132) );
  XOR U3464 ( .A(n3130), .B(n3004), .Z(n3003) );
  ANDN U3465 ( .A(n3133), .B(n3134), .Z(n3004) );
  XNOR U3466 ( .A(n3135), .B(n3059), .Z(n3035) );
  XNOR U3467 ( .A(n3013), .B(n3012), .Z(n3059) );
  XOR U3468 ( .A(n3136), .B(n3021), .Z(n3012) );
  XNOR U3469 ( .A(n3009), .B(n3010), .Z(n3021) );
  NAND U3470 ( .A(n2306), .B(n1248), .Z(n3010) );
  XNOR U3471 ( .A(n3008), .B(n3137), .Z(n3009) );
  ANDN U3472 ( .A(n2311), .B(n1250), .Z(n3137) );
  XNOR U3473 ( .A(n3020), .B(n3011), .Z(n3136) );
  XOR U3474 ( .A(n3144), .B(n3017), .Z(n3020) );
  XNOR U3475 ( .A(n3016), .B(n3145), .Z(n3017) );
  ANDN U3476 ( .A(n2541), .B(n1127), .Z(n3145) );
  AND U3477 ( .A(n2534), .B(n1125), .Z(n3018) );
  XNOR U3478 ( .A(n3029), .B(n3028), .Z(n3013) );
  XOR U3479 ( .A(n3152), .B(n3025), .Z(n3028) );
  XNOR U3480 ( .A(n3024), .B(n3153), .Z(n3025) );
  ANDN U3481 ( .A(n2112), .B(n1385), .Z(n3153) );
  AND U3482 ( .A(n2105), .B(n1383), .Z(n3026) );
  XNOR U3483 ( .A(n3032), .B(n3033), .Z(n3029) );
  NAND U3484 ( .A(n1910), .B(n1535), .Z(n3033) );
  XNOR U3485 ( .A(n3031), .B(n3160), .Z(n3032) );
  ANDN U3486 ( .A(n1915), .B(n1537), .Z(n3160) );
  XOR U3487 ( .A(n3058), .B(n3034), .Z(n3135) );
  XNOR U3488 ( .A(n3167), .B(n3063), .Z(n3058) );
  XNOR U3489 ( .A(n3041), .B(n3040), .Z(n3063) );
  XOR U3490 ( .A(n3168), .B(n3047), .Z(n3040) );
  XNOR U3491 ( .A(n3045), .B(n3169), .Z(n3047) );
  ANDN U3492 ( .A(n3050), .B(n957), .Z(n3169) );
  AND U3493 ( .A(n3043), .B(n955), .Z(n3049) );
  XNOR U3494 ( .A(n3054), .B(n3056), .Z(n3041) );
  NAND U3495 ( .A(n2796), .B(n1039), .Z(n3056) );
  XNOR U3496 ( .A(n3052), .B(n3176), .Z(n3054) );
  ANDN U3497 ( .A(n2801), .B(n1041), .Z(n3176) );
  XNOR U3498 ( .A(n3061), .B(n3057), .Z(n3167) );
  XOR U3499 ( .A(n3060), .B(n3183), .Z(n3061) );
  AND U3500 ( .A(n3184), .B(n3185), .Z(n3183) );
  NANDN U3501 ( .B(n3186), .A(n3187), .Z(n3185) );
  AND U3502 ( .A(n3188), .B(n3189), .Z(n3184) );
  NANDN U3503 ( .B(n3190), .A(n894), .Z(n3189) );
  OR U3504 ( .A(n3191), .B(n3192), .Z(n3188) );
  XNOR U3505 ( .A(n3079), .B(n3078), .Z(n3036) );
  XOR U3506 ( .A(n3196), .B(n3087), .Z(n3078) );
  XNOR U3507 ( .A(n3072), .B(n3071), .Z(n3087) );
  XOR U3508 ( .A(n3197), .B(n3068), .Z(n3071) );
  XNOR U3509 ( .A(n3067), .B(n3198), .Z(n3068) );
  ANDN U3510 ( .A(n1404), .B(n2082), .Z(n3198) );
  AND U3511 ( .A(n2080), .B(n1341), .Z(n3069) );
  XNOR U3512 ( .A(n3075), .B(n3076), .Z(n3072) );
  NANDN U3513 ( .B(n1206), .A(n2287), .Z(n3076) );
  XNOR U3514 ( .A(n3074), .B(n3205), .Z(n3075) );
  ANDN U3515 ( .A(n1276), .B(n2289), .Z(n3205) );
  XNOR U3516 ( .A(n3086), .B(n3077), .Z(n3196) );
  XOR U3517 ( .A(n3212), .B(n3095), .Z(n3086) );
  XNOR U3518 ( .A(n3083), .B(n3084), .Z(n3095) );
  NAND U3519 ( .A(n1888), .B(n1575), .Z(n3084) );
  XNOR U3520 ( .A(n3082), .B(n3213), .Z(n3083) );
  ANDN U3521 ( .A(n1582), .B(n1890), .Z(n3213) );
  XNOR U3522 ( .A(n3094), .B(n3085), .Z(n3212) );
  XOR U3523 ( .A(n3220), .B(n3091), .Z(n3094) );
  XNOR U3524 ( .A(n3090), .B(n3221), .Z(n3091) );
  ANDN U3525 ( .A(n1766), .B(n1702), .Z(n3221) );
  AND U3526 ( .A(n1700), .B(n1759), .Z(n3092) );
  XNOR U3527 ( .A(n3103), .B(n3102), .Z(n3079) );
  XOR U3528 ( .A(n3228), .B(n3111), .Z(n3102) );
  XNOR U3529 ( .A(n3099), .B(n3100), .Z(n3111) );
  NANDN U3530 ( .B(n1019), .A(n2741), .Z(n3100) );
  XNOR U3531 ( .A(n3098), .B(n3229), .Z(n3099) );
  ANDN U3532 ( .A(n1060), .B(n2743), .Z(n3229) );
  XNOR U3533 ( .A(n3110), .B(n3101), .Z(n3228) );
  XOR U3534 ( .A(n3236), .B(n3107), .Z(n3110) );
  XNOR U3535 ( .A(n3106), .B(n3237), .Z(n3107) );
  ANDN U3536 ( .A(n1167), .B(n2504), .Z(n3237) );
  AND U3537 ( .A(n2502), .B(n1113), .Z(n3108) );
  XOR U3538 ( .A(n3119), .B(n3118), .Z(n3103) );
  XOR U3539 ( .A(n3244), .B(n3115), .Z(n3118) );
  XNOR U3540 ( .A(n3114), .B(n3245), .Z(n3115) );
  ANDN U3541 ( .A(n992), .B(n2990), .Z(n3245) );
  AND U3542 ( .A(n2988), .B(n951), .Z(n3116) );
  XOR U3543 ( .A(n3126), .B(n3125), .Z(n3119) );
  NAND U3544 ( .A(n3252), .B(n895), .Z(n3125) );
  XOR U3545 ( .A(n3124), .B(n3253), .Z(n3126) );
  ANDN U3546 ( .A(n926), .B(n3254), .Z(n3253) );
  ANDN U3547 ( .A(n3255), .B(n3256), .Z(n3124) );
  NAND U3548 ( .A(n3257), .B(n3258), .Z(n3255) );
  MUX U3549 ( .IN0(n751), .IN1(Y[0]), .SEL(n2998), .F(n299) );
  NANDN U3550 ( .B(rst), .A(n846), .Z(n2998) );
  AND U3551 ( .A(n3261), .B(n3262), .Z(n846) );
  AND U3552 ( .A(n3263), .B(n3264), .Z(n3262) );
  ANDN U3553 ( .A(n3265), .B(n[7]), .Z(n3264) );
  NOR U3554 ( .A(n[8]), .B(n[9]), .Z(n3265) );
  NOR U3555 ( .A(n[5]), .B(n[6]), .Z(n3263) );
  AND U3556 ( .A(n3266), .B(n3267), .Z(n3261) );
  NOR U3557 ( .A(n[1]), .B(n[2]), .Z(n3267) );
  ANDN U3558 ( .A(n746), .B(n[0]), .Z(n3266) );
  NOR U3559 ( .A(n[3]), .B(n[4]), .Z(n746) );
  XOR U3560 ( .A(n3260), .B(Y0[1]), .Z(n751) );
  XOR U3561 ( .A(n3268), .B(n3269), .Z(n3260) );
  XOR U3562 ( .A(n3270), .B(n3259), .Z(n3268) );
  NAND U3563 ( .A(n3271), .B(n859), .Z(n3270) );
  XOR U3564 ( .A(A[31]), .B(X[31]), .Z(n859) );
  XOR U3565 ( .A(n3133), .B(n3269), .Z(n3271) );
  XOR U3566 ( .A(n3134), .B(n3269), .Z(n3133) );
  XNOR U3567 ( .A(n3272), .B(n3182), .Z(n3165) );
  XNOR U3568 ( .A(n3143), .B(n3142), .Z(n3182) );
  XOR U3569 ( .A(n3273), .B(n3151), .Z(n3142) );
  XNOR U3570 ( .A(n3139), .B(n3140), .Z(n3151) );
  NAND U3571 ( .A(n2306), .B(n1316), .Z(n3140) );
  XNOR U3572 ( .A(n3138), .B(n3274), .Z(n3139) );
  ANDN U3573 ( .A(n2311), .B(n1318), .Z(n3274) );
  XNOR U3574 ( .A(n3150), .B(n3141), .Z(n3273) );
  XOR U3575 ( .A(n3281), .B(n3147), .Z(n3150) );
  XNOR U3576 ( .A(n3146), .B(n3282), .Z(n3147) );
  ANDN U3577 ( .A(n2541), .B(n1186), .Z(n3282) );
  AND U3578 ( .A(n2534), .B(n1184), .Z(n3148) );
  XNOR U3579 ( .A(n3159), .B(n3158), .Z(n3143) );
  XOR U3580 ( .A(n3289), .B(n3155), .Z(n3158) );
  XNOR U3581 ( .A(n3154), .B(n3290), .Z(n3155) );
  ANDN U3582 ( .A(n2112), .B(n1459), .Z(n3290) );
  AND U3583 ( .A(n2105), .B(n1457), .Z(n3156) );
  XNOR U3584 ( .A(n3162), .B(n3163), .Z(n3159) );
  NAND U3585 ( .A(n1910), .B(n1616), .Z(n3163) );
  XNOR U3586 ( .A(n3161), .B(n3297), .Z(n3162) );
  ANDN U3587 ( .A(n1915), .B(n1618), .Z(n3297) );
  XOR U3588 ( .A(n3181), .B(n3164), .Z(n3272) );
  XNOR U3589 ( .A(n3304), .B(n3195), .Z(n3181) );
  XNOR U3590 ( .A(n3175), .B(n3174), .Z(n3195) );
  XOR U3591 ( .A(n3305), .B(n3171), .Z(n3174) );
  XNOR U3592 ( .A(n3170), .B(n3306), .Z(n3171) );
  ANDN U3593 ( .A(n3050), .B(n1001), .Z(n3306) );
  AND U3594 ( .A(n3043), .B(n999), .Z(n3172) );
  XNOR U3595 ( .A(n3178), .B(n3179), .Z(n3175) );
  NAND U3596 ( .A(n2796), .B(n1083), .Z(n3179) );
  XNOR U3597 ( .A(n3177), .B(n3313), .Z(n3178) );
  ANDN U3598 ( .A(n2801), .B(n1085), .Z(n3313) );
  XOR U3599 ( .A(n3194), .B(n3180), .Z(n3304) );
  XNOR U3600 ( .A(n3320), .B(n3191), .Z(n3194) );
  XNOR U3601 ( .A(n3321), .B(n3187), .Z(n3191) );
  AND U3602 ( .A(n3322), .B(n924), .Z(n3187) );
  NAND U3603 ( .A(n3323), .B(n3186), .Z(n3321) );
  NANDN U3604 ( .B(n927), .A(n3327), .Z(n3323) );
  XNOR U3605 ( .A(n3192), .B(n3193), .Z(n3320) );
  XNOR U3606 ( .A(n3331), .B(n3334), .Z(n3333) );
  XNOR U3607 ( .A(n3211), .B(n3210), .Z(n3166) );
  XOR U3608 ( .A(n3335), .B(n3219), .Z(n3210) );
  XNOR U3609 ( .A(n3204), .B(n3203), .Z(n3219) );
  XOR U3610 ( .A(n3336), .B(n3200), .Z(n3203) );
  XNOR U3611 ( .A(n3199), .B(n3337), .Z(n3200) );
  ANDN U3612 ( .A(n1404), .B(n2183), .Z(n3337) );
  AND U3613 ( .A(n2181), .B(n1341), .Z(n3201) );
  XNOR U3614 ( .A(n3207), .B(n3208), .Z(n3204) );
  NANDN U3615 ( .B(n1206), .A(n2394), .Z(n3208) );
  XNOR U3616 ( .A(n3206), .B(n3344), .Z(n3207) );
  ANDN U3617 ( .A(n1276), .B(n2396), .Z(n3344) );
  XNOR U3618 ( .A(n3218), .B(n3209), .Z(n3335) );
  XOR U3619 ( .A(n3351), .B(n3227), .Z(n3218) );
  XNOR U3620 ( .A(n3215), .B(n3216), .Z(n3227) );
  NAND U3621 ( .A(n1984), .B(n1575), .Z(n3216) );
  XNOR U3622 ( .A(n3214), .B(n3352), .Z(n3215) );
  ANDN U3623 ( .A(n1582), .B(n1986), .Z(n3352) );
  XNOR U3624 ( .A(n3226), .B(n3217), .Z(n3351) );
  XOR U3625 ( .A(n3359), .B(n3223), .Z(n3226) );
  XNOR U3626 ( .A(n3222), .B(n3360), .Z(n3223) );
  ANDN U3627 ( .A(n1766), .B(n1793), .Z(n3360) );
  AND U3628 ( .A(n1791), .B(n1759), .Z(n3224) );
  XNOR U3629 ( .A(n3235), .B(n3234), .Z(n3211) );
  XOR U3630 ( .A(n3367), .B(n3243), .Z(n3234) );
  XNOR U3631 ( .A(n3231), .B(n3232), .Z(n3243) );
  NANDN U3632 ( .B(n1019), .A(n2863), .Z(n3232) );
  XNOR U3633 ( .A(n3230), .B(n3368), .Z(n3231) );
  ANDN U3634 ( .A(n1060), .B(n2865), .Z(n3368) );
  XNOR U3635 ( .A(n3242), .B(n3233), .Z(n3367) );
  XOR U3636 ( .A(n3375), .B(n3239), .Z(n3242) );
  XNOR U3637 ( .A(n3238), .B(n3376), .Z(n3239) );
  ANDN U3638 ( .A(n1167), .B(n2623), .Z(n3376) );
  AND U3639 ( .A(n2621), .B(n1113), .Z(n3240) );
  XOR U3640 ( .A(n3251), .B(n3250), .Z(n3235) );
  XOR U3641 ( .A(n3383), .B(n3247), .Z(n3250) );
  XNOR U3642 ( .A(n3246), .B(n3384), .Z(n3247) );
  ANDN U3643 ( .A(n992), .B(n3122), .Z(n3384) );
  AND U3644 ( .A(n3120), .B(n951), .Z(n3248) );
  XOR U3645 ( .A(n3258), .B(n3257), .Z(n3251) );
  NAND U3646 ( .A(n3391), .B(n895), .Z(n3257) );
  XNOR U3647 ( .A(n3256), .B(n3392), .Z(n3258) );
  ANDN U3648 ( .A(n926), .B(n3393), .Z(n3392) );
  NAND U3649 ( .A(n3394), .B(n3395), .Z(n3256) );
  NAND U3650 ( .A(n3396), .B(n3397), .Z(n3394) );
  XNOR U3651 ( .A(n3398), .B(n3319), .Z(n3302) );
  XNOR U3652 ( .A(n3280), .B(n3279), .Z(n3319) );
  XOR U3653 ( .A(n3399), .B(n3288), .Z(n3279) );
  XNOR U3654 ( .A(n3276), .B(n3277), .Z(n3288) );
  NAND U3655 ( .A(n2306), .B(n1383), .Z(n3277) );
  XNOR U3656 ( .A(n3275), .B(n3400), .Z(n3276) );
  ANDN U3657 ( .A(n2311), .B(n1385), .Z(n3400) );
  XOR U3658 ( .A(n3401), .B(n3402), .Z(n3275) );
  AND U3659 ( .A(n3403), .B(n3404), .Z(n3402) );
  XOR U3660 ( .A(n3405), .B(n3401), .Z(n3404) );
  XNOR U3661 ( .A(n3287), .B(n3278), .Z(n3399) );
  XOR U3662 ( .A(n3409), .B(n3284), .Z(n3287) );
  XNOR U3663 ( .A(n3283), .B(n3410), .Z(n3284) );
  ANDN U3664 ( .A(n2541), .B(n1250), .Z(n3410) );
  XOR U3665 ( .A(n3411), .B(n3412), .Z(n3283) );
  AND U3666 ( .A(n3413), .B(n3414), .Z(n3412) );
  XNOR U3667 ( .A(n3415), .B(n3411), .Z(n3414) );
  AND U3668 ( .A(n2534), .B(n1248), .Z(n3285) );
  XNOR U3669 ( .A(n3296), .B(n3295), .Z(n3280) );
  XOR U3670 ( .A(n3419), .B(n3292), .Z(n3295) );
  XNOR U3671 ( .A(n3291), .B(n3420), .Z(n3292) );
  ANDN U3672 ( .A(n2112), .B(n1537), .Z(n3420) );
  AND U3673 ( .A(n2105), .B(n1535), .Z(n3293) );
  XNOR U3674 ( .A(n3299), .B(n3300), .Z(n3296) );
  NAND U3675 ( .A(n1910), .B(n1700), .Z(n3300) );
  XNOR U3676 ( .A(n3298), .B(n3427), .Z(n3299) );
  ANDN U3677 ( .A(n1915), .B(n1702), .Z(n3427) );
  XNOR U3678 ( .A(n3318), .B(n3301), .Z(n3398) );
  XNOR U3679 ( .A(n3431), .B(n3432), .Z(n3301) );
  XNOR U3680 ( .A(n3433), .B(n3330), .Z(n3318) );
  XNOR U3681 ( .A(n3312), .B(n3311), .Z(n3330) );
  XOR U3682 ( .A(n3434), .B(n3308), .Z(n3311) );
  XNOR U3683 ( .A(n3307), .B(n3435), .Z(n3308) );
  ANDN U3684 ( .A(n3050), .B(n1041), .Z(n3435) );
  XOR U3685 ( .A(n3436), .B(n3437), .Z(n3307) );
  AND U3686 ( .A(n3438), .B(n3439), .Z(n3437) );
  XNOR U3687 ( .A(n3440), .B(n3436), .Z(n3439) );
  AND U3688 ( .A(n3043), .B(n1039), .Z(n3309) );
  XNOR U3689 ( .A(n3315), .B(n3316), .Z(n3312) );
  NAND U3690 ( .A(n2796), .B(n1125), .Z(n3316) );
  XNOR U3691 ( .A(n3314), .B(n3444), .Z(n3315) );
  ANDN U3692 ( .A(n2801), .B(n1127), .Z(n3444) );
  XOR U3693 ( .A(n3445), .B(n3446), .Z(n3314) );
  AND U3694 ( .A(n3447), .B(n3448), .Z(n3446) );
  XOR U3695 ( .A(n3449), .B(n3445), .Z(n3448) );
  XNOR U3696 ( .A(n3329), .B(n3317), .Z(n3433) );
  XOR U3697 ( .A(n3450), .B(n3451), .Z(n3317) );
  AND U3698 ( .A(n3452), .B(n3453), .Z(n3451) );
  XOR U3699 ( .A(n3454), .B(n3455), .Z(n3453) );
  XNOR U3700 ( .A(n3456), .B(n3450), .Z(n3454) );
  XNOR U3701 ( .A(n3407), .B(n3457), .Z(n3452) );
  XNOR U3702 ( .A(n3450), .B(n3408), .Z(n3457) );
  XNOR U3703 ( .A(n3426), .B(n3425), .Z(n3408) );
  XOR U3704 ( .A(n3458), .B(n3422), .Z(n3425) );
  XNOR U3705 ( .A(n3421), .B(n3459), .Z(n3422) );
  ANDN U3706 ( .A(n2112), .B(n1618), .Z(n3459) );
  AND U3707 ( .A(n2105), .B(n1616), .Z(n3423) );
  XNOR U3708 ( .A(n3429), .B(n3430), .Z(n3426) );
  NAND U3709 ( .A(n1791), .B(n1910), .Z(n3430) );
  XNOR U3710 ( .A(n3428), .B(n3466), .Z(n3429) );
  ANDN U3711 ( .A(n1915), .B(n1793), .Z(n3466) );
  XOR U3712 ( .A(n3470), .B(n3418), .Z(n3407) );
  XNOR U3713 ( .A(n3403), .B(n3405), .Z(n3418) );
  NAND U3714 ( .A(n2306), .B(n1457), .Z(n3405) );
  XNOR U3715 ( .A(n3401), .B(n3471), .Z(n3403) );
  ANDN U3716 ( .A(n2311), .B(n1459), .Z(n3471) );
  XNOR U3717 ( .A(n3417), .B(n3406), .Z(n3470) );
  XOR U3718 ( .A(n3478), .B(n3413), .Z(n3417) );
  XNOR U3719 ( .A(n3411), .B(n3479), .Z(n3413) );
  ANDN U3720 ( .A(n2541), .B(n1318), .Z(n3479) );
  XOR U3721 ( .A(n3480), .B(n3481), .Z(n3411) );
  AND U3722 ( .A(n3482), .B(n3483), .Z(n3481) );
  XNOR U3723 ( .A(n3484), .B(n3480), .Z(n3483) );
  AND U3724 ( .A(n2534), .B(n1316), .Z(n3415) );
  XOR U3725 ( .A(n3488), .B(n3489), .Z(n3450) );
  AND U3726 ( .A(n3490), .B(n3491), .Z(n3489) );
  XOR U3727 ( .A(n3492), .B(n3493), .Z(n3491) );
  XOR U3728 ( .A(n3488), .B(n3494), .Z(n3493) );
  XNOR U3729 ( .A(n3476), .B(n3495), .Z(n3490) );
  XNOR U3730 ( .A(n3488), .B(n3477), .Z(n3495) );
  XNOR U3731 ( .A(n3465), .B(n3464), .Z(n3477) );
  XOR U3732 ( .A(n3496), .B(n3461), .Z(n3464) );
  XNOR U3733 ( .A(n3460), .B(n3497), .Z(n3461) );
  ANDN U3734 ( .A(n2112), .B(n1702), .Z(n3497) );
  XOR U3735 ( .A(n3498), .B(n3499), .Z(n3460) );
  AND U3736 ( .A(n3500), .B(n3501), .Z(n3499) );
  XNOR U3737 ( .A(n3502), .B(n3498), .Z(n3501) );
  AND U3738 ( .A(n2105), .B(n1700), .Z(n3462) );
  XNOR U3739 ( .A(n3468), .B(n3469), .Z(n3465) );
  NAND U3740 ( .A(n1888), .B(n1910), .Z(n3469) );
  XNOR U3741 ( .A(n3467), .B(n3506), .Z(n3468) );
  ANDN U3742 ( .A(n1915), .B(n1890), .Z(n3506) );
  XOR U3743 ( .A(n3507), .B(n3508), .Z(n3467) );
  AND U3744 ( .A(n3509), .B(n3510), .Z(n3508) );
  XOR U3745 ( .A(n3511), .B(n3507), .Z(n3510) );
  XOR U3746 ( .A(n3512), .B(n3487), .Z(n3476) );
  XNOR U3747 ( .A(n3473), .B(n3474), .Z(n3487) );
  NAND U3748 ( .A(n2306), .B(n1535), .Z(n3474) );
  XNOR U3749 ( .A(n3472), .B(n3513), .Z(n3473) );
  ANDN U3750 ( .A(n2311), .B(n1537), .Z(n3513) );
  XOR U3751 ( .A(n3514), .B(n3515), .Z(n3472) );
  AND U3752 ( .A(n3516), .B(n3517), .Z(n3515) );
  XOR U3753 ( .A(n3518), .B(n3514), .Z(n3517) );
  XNOR U3754 ( .A(n3486), .B(n3475), .Z(n3512) );
  XOR U3755 ( .A(n3522), .B(n3482), .Z(n3486) );
  XNOR U3756 ( .A(n3480), .B(n3523), .Z(n3482) );
  ANDN U3757 ( .A(n2541), .B(n1385), .Z(n3523) );
  XOR U3758 ( .A(n3524), .B(n3525), .Z(n3480) );
  AND U3759 ( .A(n3526), .B(n3527), .Z(n3525) );
  XNOR U3760 ( .A(n3528), .B(n3524), .Z(n3527) );
  XOR U3761 ( .A(n3529), .B(n3484), .Z(n3522) );
  AND U3762 ( .A(n2534), .B(n1383), .Z(n3484) );
  IV U3763 ( .A(n3485), .Z(n3529) );
  XOR U3764 ( .A(n3533), .B(n3534), .Z(n3488) );
  AND U3765 ( .A(n3535), .B(n3536), .Z(n3534) );
  XOR U3766 ( .A(n3537), .B(n3538), .Z(n3536) );
  XOR U3767 ( .A(n3533), .B(n3539), .Z(n3538) );
  XNOR U3768 ( .A(n3520), .B(n3540), .Z(n3535) );
  XNOR U3769 ( .A(n3533), .B(n3521), .Z(n3540) );
  XNOR U3770 ( .A(n3505), .B(n3504), .Z(n3521) );
  XOR U3771 ( .A(n3541), .B(n3500), .Z(n3504) );
  XNOR U3772 ( .A(n3498), .B(n3542), .Z(n3500) );
  ANDN U3773 ( .A(n2112), .B(n1793), .Z(n3542) );
  XOR U3774 ( .A(n3543), .B(n3544), .Z(n3498) );
  AND U3775 ( .A(n3545), .B(n3546), .Z(n3544) );
  XNOR U3776 ( .A(n3547), .B(n3543), .Z(n3546) );
  AND U3777 ( .A(n1791), .B(n2105), .Z(n3502) );
  XNOR U3778 ( .A(n3509), .B(n3511), .Z(n3505) );
  NAND U3779 ( .A(n1984), .B(n1910), .Z(n3511) );
  XNOR U3780 ( .A(n3507), .B(n3551), .Z(n3509) );
  ANDN U3781 ( .A(n1915), .B(n1986), .Z(n3551) );
  XOR U3782 ( .A(n3555), .B(n3532), .Z(n3520) );
  XNOR U3783 ( .A(n3516), .B(n3518), .Z(n3532) );
  NAND U3784 ( .A(n2306), .B(n1616), .Z(n3518) );
  XNOR U3785 ( .A(n3514), .B(n3556), .Z(n3516) );
  ANDN U3786 ( .A(n2311), .B(n1618), .Z(n3556) );
  XOR U3787 ( .A(n3557), .B(n3558), .Z(n3514) );
  AND U3788 ( .A(n3559), .B(n3560), .Z(n3558) );
  XOR U3789 ( .A(n3561), .B(n3557), .Z(n3560) );
  XNOR U3790 ( .A(n3531), .B(n3519), .Z(n3555) );
  XOR U3791 ( .A(n3565), .B(n3526), .Z(n3531) );
  XNOR U3792 ( .A(n3524), .B(n3566), .Z(n3526) );
  ANDN U3793 ( .A(n2541), .B(n1459), .Z(n3566) );
  XOR U3794 ( .A(n3567), .B(n3568), .Z(n3524) );
  AND U3795 ( .A(n3569), .B(n3570), .Z(n3568) );
  XNOR U3796 ( .A(n3571), .B(n3567), .Z(n3570) );
  AND U3797 ( .A(n2534), .B(n1457), .Z(n3528) );
  XOR U3798 ( .A(n3575), .B(n3576), .Z(n3533) );
  AND U3799 ( .A(n3577), .B(n3578), .Z(n3576) );
  XOR U3800 ( .A(n3579), .B(n3580), .Z(n3578) );
  XOR U3801 ( .A(n3575), .B(n3581), .Z(n3580) );
  XNOR U3802 ( .A(n3563), .B(n3582), .Z(n3577) );
  XNOR U3803 ( .A(n3575), .B(n3564), .Z(n3582) );
  XNOR U3804 ( .A(n3550), .B(n3549), .Z(n3564) );
  XOR U3805 ( .A(n3583), .B(n3545), .Z(n3549) );
  XNOR U3806 ( .A(n3543), .B(n3584), .Z(n3545) );
  ANDN U3807 ( .A(n2112), .B(n1890), .Z(n3584) );
  XOR U3808 ( .A(n3585), .B(n3586), .Z(n3543) );
  AND U3809 ( .A(n3587), .B(n3588), .Z(n3586) );
  XNOR U3810 ( .A(n3589), .B(n3585), .Z(n3588) );
  AND U3811 ( .A(n1888), .B(n2105), .Z(n3547) );
  XNOR U3812 ( .A(n3553), .B(n3554), .Z(n3550) );
  NAND U3813 ( .A(n2080), .B(n1910), .Z(n3554) );
  XNOR U3814 ( .A(n3552), .B(n3593), .Z(n3553) );
  ANDN U3815 ( .A(n1915), .B(n2082), .Z(n3593) );
  XOR U3816 ( .A(n3594), .B(n3595), .Z(n3552) );
  AND U3817 ( .A(n3596), .B(n3597), .Z(n3595) );
  XOR U3818 ( .A(n3598), .B(n3594), .Z(n3597) );
  XOR U3819 ( .A(n3599), .B(n3574), .Z(n3563) );
  XNOR U3820 ( .A(n3559), .B(n3561), .Z(n3574) );
  NAND U3821 ( .A(n2306), .B(n1700), .Z(n3561) );
  XNOR U3822 ( .A(n3557), .B(n3600), .Z(n3559) );
  ANDN U3823 ( .A(n2311), .B(n1702), .Z(n3600) );
  XNOR U3824 ( .A(n3573), .B(n3562), .Z(n3599) );
  XOR U3825 ( .A(n3607), .B(n3569), .Z(n3573) );
  XNOR U3826 ( .A(n3567), .B(n3608), .Z(n3569) );
  ANDN U3827 ( .A(n2541), .B(n1537), .Z(n3608) );
  XOR U3828 ( .A(n3609), .B(n3610), .Z(n3567) );
  AND U3829 ( .A(n3611), .B(n3612), .Z(n3610) );
  XNOR U3830 ( .A(n3613), .B(n3609), .Z(n3612) );
  XOR U3831 ( .A(n3614), .B(n3571), .Z(n3607) );
  AND U3832 ( .A(n2534), .B(n1535), .Z(n3571) );
  IV U3833 ( .A(n3572), .Z(n3614) );
  XOR U3834 ( .A(n3618), .B(n3619), .Z(n3575) );
  AND U3835 ( .A(n3620), .B(n3621), .Z(n3619) );
  XOR U3836 ( .A(n3622), .B(n3623), .Z(n3621) );
  XOR U3837 ( .A(n3618), .B(n3624), .Z(n3623) );
  XNOR U3838 ( .A(n3605), .B(n3625), .Z(n3620) );
  XNOR U3839 ( .A(n3618), .B(n3606), .Z(n3625) );
  XNOR U3840 ( .A(n3592), .B(n3591), .Z(n3606) );
  XOR U3841 ( .A(n3626), .B(n3587), .Z(n3591) );
  XNOR U3842 ( .A(n3585), .B(n3627), .Z(n3587) );
  ANDN U3843 ( .A(n2112), .B(n1986), .Z(n3627) );
  XOR U3844 ( .A(n3628), .B(n3629), .Z(n3585) );
  AND U3845 ( .A(n3630), .B(n3631), .Z(n3629) );
  XNOR U3846 ( .A(n3632), .B(n3628), .Z(n3631) );
  AND U3847 ( .A(n1984), .B(n2105), .Z(n3589) );
  XNOR U3848 ( .A(n3596), .B(n3598), .Z(n3592) );
  NAND U3849 ( .A(n2181), .B(n1910), .Z(n3598) );
  XNOR U3850 ( .A(n3594), .B(n3636), .Z(n3596) );
  ANDN U3851 ( .A(n1915), .B(n2183), .Z(n3636) );
  XOR U3852 ( .A(n3640), .B(n3617), .Z(n3605) );
  XNOR U3853 ( .A(n3602), .B(n3603), .Z(n3617) );
  NAND U3854 ( .A(n1791), .B(n2306), .Z(n3603) );
  XNOR U3855 ( .A(n3601), .B(n3641), .Z(n3602) );
  ANDN U3856 ( .A(n2311), .B(n1793), .Z(n3641) );
  XOR U3857 ( .A(n3642), .B(n3643), .Z(n3601) );
  AND U3858 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U3859 ( .A(n3646), .B(n3642), .Z(n3645) );
  XNOR U3860 ( .A(n3616), .B(n3604), .Z(n3640) );
  XOR U3861 ( .A(n3650), .B(n3611), .Z(n3616) );
  XNOR U3862 ( .A(n3609), .B(n3651), .Z(n3611) );
  ANDN U3863 ( .A(n2541), .B(n1618), .Z(n3651) );
  XOR U3864 ( .A(n3652), .B(n3653), .Z(n3609) );
  AND U3865 ( .A(n3654), .B(n3655), .Z(n3653) );
  XNOR U3866 ( .A(n3656), .B(n3652), .Z(n3655) );
  AND U3867 ( .A(n2534), .B(n1616), .Z(n3613) );
  XOR U3868 ( .A(n3660), .B(n3661), .Z(n3618) );
  AND U3869 ( .A(n3662), .B(n3663), .Z(n3661) );
  XOR U3870 ( .A(n3664), .B(n3665), .Z(n3663) );
  XOR U3871 ( .A(n3660), .B(n3666), .Z(n3665) );
  XNOR U3872 ( .A(n3648), .B(n3667), .Z(n3662) );
  XNOR U3873 ( .A(n3660), .B(n3649), .Z(n3667) );
  XNOR U3874 ( .A(n3635), .B(n3634), .Z(n3649) );
  XOR U3875 ( .A(n3668), .B(n3630), .Z(n3634) );
  XNOR U3876 ( .A(n3628), .B(n3669), .Z(n3630) );
  ANDN U3877 ( .A(n2112), .B(n2082), .Z(n3669) );
  XOR U3878 ( .A(n3670), .B(n3671), .Z(n3628) );
  AND U3879 ( .A(n3672), .B(n3673), .Z(n3671) );
  XNOR U3880 ( .A(n3674), .B(n3670), .Z(n3673) );
  XOR U3881 ( .A(n3675), .B(n3632), .Z(n3668) );
  AND U3882 ( .A(n2080), .B(n2105), .Z(n3632) );
  IV U3883 ( .A(n3633), .Z(n3675) );
  XNOR U3884 ( .A(n3638), .B(n3639), .Z(n3635) );
  NAND U3885 ( .A(n2287), .B(n1910), .Z(n3639) );
  XNOR U3886 ( .A(n3637), .B(n3679), .Z(n3638) );
  ANDN U3887 ( .A(n1915), .B(n2289), .Z(n3679) );
  XOR U3888 ( .A(n3680), .B(n3681), .Z(n3637) );
  AND U3889 ( .A(n3682), .B(n3683), .Z(n3681) );
  XOR U3890 ( .A(n3684), .B(n3680), .Z(n3683) );
  XOR U3891 ( .A(n3685), .B(n3659), .Z(n3648) );
  XNOR U3892 ( .A(n3644), .B(n3646), .Z(n3659) );
  NAND U3893 ( .A(n1888), .B(n2306), .Z(n3646) );
  XNOR U3894 ( .A(n3642), .B(n3686), .Z(n3644) );
  ANDN U3895 ( .A(n2311), .B(n1890), .Z(n3686) );
  XOR U3896 ( .A(n3687), .B(n3688), .Z(n3642) );
  AND U3897 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR U3898 ( .A(n3691), .B(n3687), .Z(n3690) );
  XNOR U3899 ( .A(n3658), .B(n3647), .Z(n3685) );
  XOR U3900 ( .A(n3695), .B(n3654), .Z(n3658) );
  XNOR U3901 ( .A(n3652), .B(n3696), .Z(n3654) );
  ANDN U3902 ( .A(n2541), .B(n1702), .Z(n3696) );
  XOR U3903 ( .A(n3697), .B(n3698), .Z(n3652) );
  AND U3904 ( .A(n3699), .B(n3700), .Z(n3698) );
  XNOR U3905 ( .A(n3701), .B(n3697), .Z(n3700) );
  XOR U3906 ( .A(n3702), .B(n3656), .Z(n3695) );
  AND U3907 ( .A(n2534), .B(n1700), .Z(n3656) );
  IV U3908 ( .A(n3657), .Z(n3702) );
  XOR U3909 ( .A(n3706), .B(n3707), .Z(n3660) );
  AND U3910 ( .A(n3708), .B(n3709), .Z(n3707) );
  XOR U3911 ( .A(n3710), .B(n3711), .Z(n3709) );
  XOR U3912 ( .A(n3706), .B(n3712), .Z(n3711) );
  XNOR U3913 ( .A(n3693), .B(n3713), .Z(n3708) );
  XNOR U3914 ( .A(n3706), .B(n3694), .Z(n3713) );
  XNOR U3915 ( .A(n3678), .B(n3677), .Z(n3694) );
  XOR U3916 ( .A(n3714), .B(n3672), .Z(n3677) );
  XNOR U3917 ( .A(n3670), .B(n3715), .Z(n3672) );
  ANDN U3918 ( .A(n2112), .B(n2183), .Z(n3715) );
  XOR U3919 ( .A(n3716), .B(n3717), .Z(n3670) );
  AND U3920 ( .A(n3718), .B(n3719), .Z(n3717) );
  XNOR U3921 ( .A(n3720), .B(n3716), .Z(n3719) );
  XOR U3922 ( .A(n3721), .B(n3674), .Z(n3714) );
  AND U3923 ( .A(n2181), .B(n2105), .Z(n3674) );
  IV U3924 ( .A(n3676), .Z(n3721) );
  XNOR U3925 ( .A(n3682), .B(n3684), .Z(n3678) );
  NAND U3926 ( .A(n2394), .B(n1910), .Z(n3684) );
  XNOR U3927 ( .A(n3680), .B(n3725), .Z(n3682) );
  ANDN U3928 ( .A(n1915), .B(n2396), .Z(n3725) );
  XOR U3929 ( .A(n3726), .B(n3727), .Z(n3680) );
  AND U3930 ( .A(n3728), .B(n3729), .Z(n3727) );
  XOR U3931 ( .A(n3730), .B(n3726), .Z(n3729) );
  XOR U3932 ( .A(n3731), .B(n3705), .Z(n3693) );
  XNOR U3933 ( .A(n3689), .B(n3691), .Z(n3705) );
  NAND U3934 ( .A(n1984), .B(n2306), .Z(n3691) );
  XNOR U3935 ( .A(n3687), .B(n3732), .Z(n3689) );
  ANDN U3936 ( .A(n2311), .B(n1986), .Z(n3732) );
  XNOR U3937 ( .A(n3704), .B(n3692), .Z(n3731) );
  XOR U3938 ( .A(n3739), .B(n3699), .Z(n3704) );
  XNOR U3939 ( .A(n3697), .B(n3740), .Z(n3699) );
  ANDN U3940 ( .A(n2541), .B(n1793), .Z(n3740) );
  XOR U3941 ( .A(n3741), .B(n3742), .Z(n3697) );
  AND U3942 ( .A(n3743), .B(n3744), .Z(n3742) );
  XNOR U3943 ( .A(n3745), .B(n3741), .Z(n3744) );
  XOR U3944 ( .A(n3746), .B(n3701), .Z(n3739) );
  AND U3945 ( .A(n1791), .B(n2534), .Z(n3701) );
  IV U3946 ( .A(n3703), .Z(n3746) );
  XOR U3947 ( .A(n3750), .B(n3751), .Z(n3706) );
  AND U3948 ( .A(n3752), .B(n3753), .Z(n3751) );
  XOR U3949 ( .A(n3754), .B(n3755), .Z(n3753) );
  XOR U3950 ( .A(n3750), .B(n3756), .Z(n3755) );
  XNOR U3951 ( .A(n3737), .B(n3757), .Z(n3752) );
  XNOR U3952 ( .A(n3750), .B(n3738), .Z(n3757) );
  XNOR U3953 ( .A(n3724), .B(n3723), .Z(n3738) );
  XOR U3954 ( .A(n3758), .B(n3718), .Z(n3723) );
  XNOR U3955 ( .A(n3716), .B(n3759), .Z(n3718) );
  ANDN U3956 ( .A(n2112), .B(n2289), .Z(n3759) );
  XOR U3957 ( .A(n3760), .B(n3761), .Z(n3716) );
  AND U3958 ( .A(n3762), .B(n3763), .Z(n3761) );
  XNOR U3959 ( .A(n3764), .B(n3760), .Z(n3763) );
  XOR U3960 ( .A(n3765), .B(n3720), .Z(n3758) );
  AND U3961 ( .A(n2287), .B(n2105), .Z(n3720) );
  IV U3962 ( .A(n3722), .Z(n3765) );
  XNOR U3963 ( .A(n3728), .B(n3730), .Z(n3724) );
  NAND U3964 ( .A(n2502), .B(n1910), .Z(n3730) );
  XNOR U3965 ( .A(n3726), .B(n3769), .Z(n3728) );
  ANDN U3966 ( .A(n1915), .B(n2504), .Z(n3769) );
  XOR U3967 ( .A(n3770), .B(n3771), .Z(n3726) );
  AND U3968 ( .A(n3772), .B(n3773), .Z(n3771) );
  XOR U3969 ( .A(n3774), .B(n3770), .Z(n3773) );
  XOR U3970 ( .A(n3775), .B(n3749), .Z(n3737) );
  XNOR U3971 ( .A(n3734), .B(n3735), .Z(n3749) );
  NAND U3972 ( .A(n2080), .B(n2306), .Z(n3735) );
  XNOR U3973 ( .A(n3733), .B(n3776), .Z(n3734) );
  ANDN U3974 ( .A(n2311), .B(n2082), .Z(n3776) );
  XOR U3975 ( .A(n3777), .B(n3778), .Z(n3733) );
  AND U3976 ( .A(n3779), .B(n3780), .Z(n3778) );
  XOR U3977 ( .A(n3781), .B(n3777), .Z(n3780) );
  XNOR U3978 ( .A(n3748), .B(n3736), .Z(n3775) );
  XOR U3979 ( .A(n3785), .B(n3743), .Z(n3748) );
  XNOR U3980 ( .A(n3741), .B(n3786), .Z(n3743) );
  ANDN U3981 ( .A(n2541), .B(n1890), .Z(n3786) );
  XOR U3982 ( .A(n3787), .B(n3788), .Z(n3741) );
  AND U3983 ( .A(n3789), .B(n3790), .Z(n3788) );
  XNOR U3984 ( .A(n3791), .B(n3787), .Z(n3790) );
  XOR U3985 ( .A(n3792), .B(n3745), .Z(n3785) );
  AND U3986 ( .A(n1888), .B(n2534), .Z(n3745) );
  IV U3987 ( .A(n3747), .Z(n3792) );
  XOR U3988 ( .A(n3796), .B(n3797), .Z(n3750) );
  AND U3989 ( .A(n3798), .B(n3799), .Z(n3797) );
  XOR U3990 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U3991 ( .A(n3796), .B(n3802), .Z(n3801) );
  XNOR U3992 ( .A(n3783), .B(n3803), .Z(n3798) );
  XNOR U3993 ( .A(n3796), .B(n3784), .Z(n3803) );
  XNOR U3994 ( .A(n3768), .B(n3767), .Z(n3784) );
  XOR U3995 ( .A(n3804), .B(n3762), .Z(n3767) );
  XNOR U3996 ( .A(n3760), .B(n3805), .Z(n3762) );
  ANDN U3997 ( .A(n2112), .B(n2396), .Z(n3805) );
  XOR U3998 ( .A(n3806), .B(n3807), .Z(n3760) );
  AND U3999 ( .A(n3808), .B(n3809), .Z(n3807) );
  XNOR U4000 ( .A(n3810), .B(n3806), .Z(n3809) );
  XOR U4001 ( .A(n3811), .B(n3764), .Z(n3804) );
  AND U4002 ( .A(n2394), .B(n2105), .Z(n3764) );
  IV U4003 ( .A(n3766), .Z(n3811) );
  XNOR U4004 ( .A(n3772), .B(n3774), .Z(n3768) );
  NAND U4005 ( .A(n2621), .B(n1910), .Z(n3774) );
  XNOR U4006 ( .A(n3770), .B(n3815), .Z(n3772) );
  ANDN U4007 ( .A(n1915), .B(n2623), .Z(n3815) );
  XOR U4008 ( .A(n3816), .B(n3817), .Z(n3770) );
  AND U4009 ( .A(n3818), .B(n3819), .Z(n3817) );
  XOR U4010 ( .A(n3820), .B(n3816), .Z(n3819) );
  XOR U4011 ( .A(n3821), .B(n3795), .Z(n3783) );
  XNOR U4012 ( .A(n3779), .B(n3781), .Z(n3795) );
  NAND U4013 ( .A(n2181), .B(n2306), .Z(n3781) );
  XNOR U4014 ( .A(n3777), .B(n3822), .Z(n3779) );
  ANDN U4015 ( .A(n2311), .B(n2183), .Z(n3822) );
  XOR U4016 ( .A(n3823), .B(n3824), .Z(n3777) );
  AND U4017 ( .A(n3825), .B(n3826), .Z(n3824) );
  XOR U4018 ( .A(n3827), .B(n3823), .Z(n3826) );
  XNOR U4019 ( .A(n3794), .B(n3782), .Z(n3821) );
  XOR U4020 ( .A(n3831), .B(n3789), .Z(n3794) );
  XNOR U4021 ( .A(n3787), .B(n3832), .Z(n3789) );
  ANDN U4022 ( .A(n2541), .B(n1986), .Z(n3832) );
  XOR U4023 ( .A(n3833), .B(n3834), .Z(n3787) );
  AND U4024 ( .A(n3835), .B(n3836), .Z(n3834) );
  XNOR U4025 ( .A(n3837), .B(n3833), .Z(n3836) );
  XOR U4026 ( .A(n3838), .B(n3791), .Z(n3831) );
  AND U4027 ( .A(n1984), .B(n2534), .Z(n3791) );
  IV U4028 ( .A(n3793), .Z(n3838) );
  XOR U4029 ( .A(n3842), .B(n3843), .Z(n3796) );
  AND U4030 ( .A(n3844), .B(n3845), .Z(n3843) );
  XOR U4031 ( .A(n3846), .B(n3847), .Z(n3845) );
  XOR U4032 ( .A(n3842), .B(n3848), .Z(n3847) );
  XNOR U4033 ( .A(n3829), .B(n3849), .Z(n3844) );
  XNOR U4034 ( .A(n3842), .B(n3830), .Z(n3849) );
  XNOR U4035 ( .A(n3814), .B(n3813), .Z(n3830) );
  XOR U4036 ( .A(n3850), .B(n3808), .Z(n3813) );
  XNOR U4037 ( .A(n3806), .B(n3851), .Z(n3808) );
  ANDN U4038 ( .A(n2112), .B(n2504), .Z(n3851) );
  XOR U4039 ( .A(n3852), .B(n3853), .Z(n3806) );
  AND U4040 ( .A(n3854), .B(n3855), .Z(n3853) );
  XNOR U4041 ( .A(n3856), .B(n3852), .Z(n3855) );
  XOR U4042 ( .A(n3857), .B(n3810), .Z(n3850) );
  AND U4043 ( .A(n2502), .B(n2105), .Z(n3810) );
  IV U4044 ( .A(n3812), .Z(n3857) );
  XNOR U4045 ( .A(n3818), .B(n3820), .Z(n3814) );
  NAND U4046 ( .A(n2741), .B(n1910), .Z(n3820) );
  XNOR U4047 ( .A(n3816), .B(n3861), .Z(n3818) );
  ANDN U4048 ( .A(n1915), .B(n2743), .Z(n3861) );
  XOR U4049 ( .A(n3862), .B(n3863), .Z(n3816) );
  AND U4050 ( .A(n3864), .B(n3865), .Z(n3863) );
  XOR U4051 ( .A(n3866), .B(n3862), .Z(n3865) );
  XOR U4052 ( .A(n3867), .B(n3841), .Z(n3829) );
  XNOR U4053 ( .A(n3825), .B(n3827), .Z(n3841) );
  NAND U4054 ( .A(n2287), .B(n2306), .Z(n3827) );
  XNOR U4055 ( .A(n3823), .B(n3868), .Z(n3825) );
  ANDN U4056 ( .A(n2311), .B(n2289), .Z(n3868) );
  XOR U4057 ( .A(n3869), .B(n3870), .Z(n3823) );
  AND U4058 ( .A(n3871), .B(n3872), .Z(n3870) );
  XOR U4059 ( .A(n3873), .B(n3869), .Z(n3872) );
  XNOR U4060 ( .A(n3840), .B(n3828), .Z(n3867) );
  XOR U4061 ( .A(n3877), .B(n3835), .Z(n3840) );
  XNOR U4062 ( .A(n3833), .B(n3878), .Z(n3835) );
  ANDN U4063 ( .A(n2541), .B(n2082), .Z(n3878) );
  XOR U4064 ( .A(n3879), .B(n3880), .Z(n3833) );
  AND U4065 ( .A(n3881), .B(n3882), .Z(n3880) );
  XNOR U4066 ( .A(n3883), .B(n3879), .Z(n3882) );
  XOR U4067 ( .A(n3884), .B(n3837), .Z(n3877) );
  AND U4068 ( .A(n2080), .B(n2534), .Z(n3837) );
  IV U4069 ( .A(n3839), .Z(n3884) );
  XOR U4070 ( .A(n3888), .B(n3889), .Z(n3842) );
  AND U4071 ( .A(n3890), .B(n3891), .Z(n3889) );
  XOR U4072 ( .A(n3892), .B(n3893), .Z(n3891) );
  XOR U4073 ( .A(n3888), .B(n3894), .Z(n3893) );
  XNOR U4074 ( .A(n3875), .B(n3895), .Z(n3890) );
  XNOR U4075 ( .A(n3888), .B(n3876), .Z(n3895) );
  XNOR U4076 ( .A(n3860), .B(n3859), .Z(n3876) );
  XOR U4077 ( .A(n3896), .B(n3854), .Z(n3859) );
  XNOR U4078 ( .A(n3852), .B(n3897), .Z(n3854) );
  ANDN U4079 ( .A(n2112), .B(n2623), .Z(n3897) );
  XOR U4080 ( .A(n3898), .B(n3899), .Z(n3852) );
  AND U4081 ( .A(n3900), .B(n3901), .Z(n3899) );
  XNOR U4082 ( .A(n3902), .B(n3898), .Z(n3901) );
  XOR U4083 ( .A(n3903), .B(n3856), .Z(n3896) );
  AND U4084 ( .A(n2621), .B(n2105), .Z(n3856) );
  IV U4085 ( .A(n3858), .Z(n3903) );
  XNOR U4086 ( .A(n3864), .B(n3866), .Z(n3860) );
  NAND U4087 ( .A(n2863), .B(n1910), .Z(n3866) );
  XNOR U4088 ( .A(n3862), .B(n3907), .Z(n3864) );
  ANDN U4089 ( .A(n1915), .B(n2865), .Z(n3907) );
  XOR U4090 ( .A(n3911), .B(n3887), .Z(n3875) );
  XNOR U4091 ( .A(n3871), .B(n3873), .Z(n3887) );
  NAND U4092 ( .A(n2394), .B(n2306), .Z(n3873) );
  XNOR U4093 ( .A(n3869), .B(n3912), .Z(n3871) );
  ANDN U4094 ( .A(n2311), .B(n2396), .Z(n3912) );
  XOR U4095 ( .A(n3913), .B(n3914), .Z(n3869) );
  AND U4096 ( .A(n3915), .B(n3916), .Z(n3914) );
  XOR U4097 ( .A(n3917), .B(n3913), .Z(n3916) );
  XNOR U4098 ( .A(n3886), .B(n3874), .Z(n3911) );
  XOR U4099 ( .A(n3921), .B(n3881), .Z(n3886) );
  XNOR U4100 ( .A(n3879), .B(n3922), .Z(n3881) );
  ANDN U4101 ( .A(n2541), .B(n2183), .Z(n3922) );
  XOR U4102 ( .A(n3923), .B(n3924), .Z(n3879) );
  AND U4103 ( .A(n3925), .B(n3926), .Z(n3924) );
  XNOR U4104 ( .A(n3927), .B(n3923), .Z(n3926) );
  XOR U4105 ( .A(n3928), .B(n3883), .Z(n3921) );
  AND U4106 ( .A(n2181), .B(n2534), .Z(n3883) );
  IV U4107 ( .A(n3885), .Z(n3928) );
  XOR U4108 ( .A(n3932), .B(n3933), .Z(n3888) );
  AND U4109 ( .A(n3934), .B(n3935), .Z(n3933) );
  XOR U4110 ( .A(n3936), .B(n3937), .Z(n3935) );
  XOR U4111 ( .A(n3932), .B(n3938), .Z(n3937) );
  XNOR U4112 ( .A(n3919), .B(n3939), .Z(n3934) );
  XNOR U4113 ( .A(n3932), .B(n3920), .Z(n3939) );
  XNOR U4114 ( .A(n3906), .B(n3905), .Z(n3920) );
  XOR U4115 ( .A(n3940), .B(n3900), .Z(n3905) );
  XNOR U4116 ( .A(n3898), .B(n3941), .Z(n3900) );
  ANDN U4117 ( .A(n2112), .B(n2743), .Z(n3941) );
  XOR U4118 ( .A(n3942), .B(n3943), .Z(n3898) );
  AND U4119 ( .A(n3944), .B(n3945), .Z(n3943) );
  XNOR U4120 ( .A(n3946), .B(n3942), .Z(n3945) );
  XOR U4121 ( .A(n3947), .B(n3902), .Z(n3940) );
  AND U4122 ( .A(n2741), .B(n2105), .Z(n3902) );
  IV U4123 ( .A(n3904), .Z(n3947) );
  XNOR U4124 ( .A(n3909), .B(n3910), .Z(n3906) );
  NAND U4125 ( .A(n2988), .B(n1910), .Z(n3910) );
  XNOR U4126 ( .A(n3908), .B(n3951), .Z(n3909) );
  ANDN U4127 ( .A(n1915), .B(n2990), .Z(n3951) );
  XOR U4128 ( .A(n3952), .B(n3953), .Z(n3908) );
  AND U4129 ( .A(n3954), .B(n3955), .Z(n3953) );
  XOR U4130 ( .A(n3956), .B(n3952), .Z(n3955) );
  XOR U4131 ( .A(n3957), .B(n3931), .Z(n3919) );
  XNOR U4132 ( .A(n3915), .B(n3917), .Z(n3931) );
  NAND U4133 ( .A(n2502), .B(n2306), .Z(n3917) );
  XNOR U4134 ( .A(n3913), .B(n3958), .Z(n3915) );
  ANDN U4135 ( .A(n2311), .B(n2504), .Z(n3958) );
  XOR U4136 ( .A(n3959), .B(n3960), .Z(n3913) );
  AND U4137 ( .A(n3961), .B(n3962), .Z(n3960) );
  XOR U4138 ( .A(n3963), .B(n3959), .Z(n3962) );
  XNOR U4139 ( .A(n3930), .B(n3918), .Z(n3957) );
  XOR U4140 ( .A(n3967), .B(n3925), .Z(n3930) );
  XNOR U4141 ( .A(n3923), .B(n3968), .Z(n3925) );
  ANDN U4142 ( .A(n2541), .B(n2289), .Z(n3968) );
  XOR U4143 ( .A(n3969), .B(n3970), .Z(n3923) );
  AND U4144 ( .A(n3971), .B(n3972), .Z(n3970) );
  XNOR U4145 ( .A(n3973), .B(n3969), .Z(n3972) );
  XOR U4146 ( .A(n3974), .B(n3927), .Z(n3967) );
  AND U4147 ( .A(n2287), .B(n2534), .Z(n3927) );
  IV U4148 ( .A(n3929), .Z(n3974) );
  XOR U4149 ( .A(n3978), .B(n3979), .Z(n3932) );
  AND U4150 ( .A(n3980), .B(n3981), .Z(n3979) );
  XOR U4151 ( .A(n3982), .B(n3983), .Z(n3981) );
  XOR U4152 ( .A(n3978), .B(n3984), .Z(n3983) );
  XNOR U4153 ( .A(n3965), .B(n3985), .Z(n3980) );
  XNOR U4154 ( .A(n3978), .B(n3966), .Z(n3985) );
  XNOR U4155 ( .A(n3950), .B(n3949), .Z(n3966) );
  XOR U4156 ( .A(n3986), .B(n3944), .Z(n3949) );
  XNOR U4157 ( .A(n3942), .B(n3987), .Z(n3944) );
  ANDN U4158 ( .A(n2112), .B(n2865), .Z(n3987) );
  XOR U4159 ( .A(n3988), .B(n3989), .Z(n3942) );
  AND U4160 ( .A(n3990), .B(n3991), .Z(n3989) );
  XNOR U4161 ( .A(n3992), .B(n3988), .Z(n3991) );
  XOR U4162 ( .A(n3993), .B(n3946), .Z(n3986) );
  AND U4163 ( .A(n2863), .B(n2105), .Z(n3946) );
  IV U4164 ( .A(n3948), .Z(n3993) );
  XNOR U4165 ( .A(n3954), .B(n3956), .Z(n3950) );
  NAND U4166 ( .A(n3120), .B(n1910), .Z(n3956) );
  XNOR U4167 ( .A(n3952), .B(n3997), .Z(n3954) );
  ANDN U4168 ( .A(n1915), .B(n3122), .Z(n3997) );
  XOR U4169 ( .A(n3998), .B(n3999), .Z(n3952) );
  AND U4170 ( .A(n4000), .B(n4001), .Z(n3999) );
  XOR U4171 ( .A(n4002), .B(n3998), .Z(n4001) );
  XOR U4172 ( .A(n4003), .B(n3977), .Z(n3965) );
  XNOR U4173 ( .A(n3961), .B(n3963), .Z(n3977) );
  NAND U4174 ( .A(n2621), .B(n2306), .Z(n3963) );
  XNOR U4175 ( .A(n3959), .B(n4004), .Z(n3961) );
  ANDN U4176 ( .A(n2311), .B(n2623), .Z(n4004) );
  XOR U4177 ( .A(n4005), .B(n4006), .Z(n3959) );
  AND U4178 ( .A(n4007), .B(n4008), .Z(n4006) );
  XOR U4179 ( .A(n4009), .B(n4005), .Z(n4008) );
  XNOR U4180 ( .A(n3976), .B(n3964), .Z(n4003) );
  XOR U4181 ( .A(n4013), .B(n3971), .Z(n3976) );
  XNOR U4182 ( .A(n3969), .B(n4014), .Z(n3971) );
  ANDN U4183 ( .A(n2541), .B(n2396), .Z(n4014) );
  XOR U4184 ( .A(n4015), .B(n4016), .Z(n3969) );
  AND U4185 ( .A(n4017), .B(n4018), .Z(n4016) );
  XNOR U4186 ( .A(n4019), .B(n4015), .Z(n4018) );
  XOR U4187 ( .A(n4020), .B(n3973), .Z(n4013) );
  AND U4188 ( .A(n2394), .B(n2534), .Z(n3973) );
  IV U4189 ( .A(n3975), .Z(n4020) );
  XOR U4190 ( .A(n4024), .B(n4025), .Z(n3978) );
  AND U4191 ( .A(n4026), .B(n4027), .Z(n4025) );
  XOR U4192 ( .A(n4028), .B(n4029), .Z(n4027) );
  XOR U4193 ( .A(n4024), .B(n4030), .Z(n4029) );
  XNOR U4194 ( .A(n4011), .B(n4031), .Z(n4026) );
  XNOR U4195 ( .A(n4024), .B(n4012), .Z(n4031) );
  XNOR U4196 ( .A(n3996), .B(n3995), .Z(n4012) );
  XOR U4197 ( .A(n4032), .B(n3990), .Z(n3995) );
  XNOR U4198 ( .A(n3988), .B(n4033), .Z(n3990) );
  ANDN U4199 ( .A(n2112), .B(n2990), .Z(n4033) );
  XOR U4200 ( .A(n4034), .B(n4035), .Z(n3988) );
  AND U4201 ( .A(n4036), .B(n4037), .Z(n4035) );
  XNOR U4202 ( .A(n4038), .B(n4034), .Z(n4037) );
  XOR U4203 ( .A(n4039), .B(n3992), .Z(n4032) );
  AND U4204 ( .A(n2988), .B(n2105), .Z(n3992) );
  IV U4205 ( .A(n3994), .Z(n4039) );
  XNOR U4206 ( .A(n4000), .B(n4002), .Z(n3996) );
  NAND U4207 ( .A(n3252), .B(n1910), .Z(n4002) );
  XNOR U4208 ( .A(n3998), .B(n4043), .Z(n4000) );
  ANDN U4209 ( .A(n1915), .B(n3254), .Z(n4043) );
  XOR U4210 ( .A(n4044), .B(n4045), .Z(n3998) );
  AND U4211 ( .A(n4046), .B(n4047), .Z(n4045) );
  XOR U4212 ( .A(n4048), .B(n4044), .Z(n4047) );
  XOR U4213 ( .A(n4049), .B(n4023), .Z(n4011) );
  XNOR U4214 ( .A(n4007), .B(n4009), .Z(n4023) );
  NAND U4215 ( .A(n2741), .B(n2306), .Z(n4009) );
  XNOR U4216 ( .A(n4005), .B(n4050), .Z(n4007) );
  ANDN U4217 ( .A(n2311), .B(n2743), .Z(n4050) );
  XOR U4218 ( .A(n4051), .B(n4052), .Z(n4005) );
  AND U4219 ( .A(n4053), .B(n4054), .Z(n4052) );
  XOR U4220 ( .A(n4055), .B(n4051), .Z(n4054) );
  XNOR U4221 ( .A(n4022), .B(n4010), .Z(n4049) );
  XOR U4222 ( .A(n4059), .B(n4017), .Z(n4022) );
  XNOR U4223 ( .A(n4015), .B(n4060), .Z(n4017) );
  ANDN U4224 ( .A(n2541), .B(n2504), .Z(n4060) );
  XOR U4225 ( .A(n4061), .B(n4062), .Z(n4015) );
  AND U4226 ( .A(n4063), .B(n4064), .Z(n4062) );
  XNOR U4227 ( .A(n4065), .B(n4061), .Z(n4064) );
  XOR U4228 ( .A(n4066), .B(n4019), .Z(n4059) );
  AND U4229 ( .A(n2502), .B(n2534), .Z(n4019) );
  IV U4230 ( .A(n4021), .Z(n4066) );
  XOR U4231 ( .A(n4070), .B(n4071), .Z(n4024) );
  AND U4232 ( .A(n4072), .B(n4073), .Z(n4071) );
  XOR U4233 ( .A(n4074), .B(n4075), .Z(n4073) );
  XOR U4234 ( .A(n4070), .B(n4076), .Z(n4075) );
  XNOR U4235 ( .A(n4057), .B(n4077), .Z(n4072) );
  XNOR U4236 ( .A(n4070), .B(n4058), .Z(n4077) );
  XNOR U4237 ( .A(n4042), .B(n4041), .Z(n4058) );
  XOR U4238 ( .A(n4078), .B(n4036), .Z(n4041) );
  XNOR U4239 ( .A(n4034), .B(n4079), .Z(n4036) );
  ANDN U4240 ( .A(n2112), .B(n3122), .Z(n4079) );
  XOR U4241 ( .A(n4083), .B(n4038), .Z(n4078) );
  AND U4242 ( .A(n3120), .B(n2105), .Z(n4038) );
  IV U4243 ( .A(n4040), .Z(n4083) );
  XNOR U4244 ( .A(n4046), .B(n4048), .Z(n4042) );
  NAND U4245 ( .A(n3391), .B(n1910), .Z(n4048) );
  XNOR U4246 ( .A(n4044), .B(n4087), .Z(n4046) );
  ANDN U4247 ( .A(n1915), .B(n3393), .Z(n4087) );
  XOR U4248 ( .A(n4091), .B(n4069), .Z(n4057) );
  XNOR U4249 ( .A(n4053), .B(n4055), .Z(n4069) );
  NAND U4250 ( .A(n2863), .B(n2306), .Z(n4055) );
  XNOR U4251 ( .A(n4051), .B(n4092), .Z(n4053) );
  ANDN U4252 ( .A(n2311), .B(n2865), .Z(n4092) );
  XOR U4253 ( .A(n4093), .B(n4094), .Z(n4051) );
  AND U4254 ( .A(n4095), .B(n4096), .Z(n4094) );
  XOR U4255 ( .A(n4097), .B(n4093), .Z(n4096) );
  XNOR U4256 ( .A(n4068), .B(n4056), .Z(n4091) );
  XOR U4257 ( .A(n4101), .B(n4063), .Z(n4068) );
  XNOR U4258 ( .A(n4061), .B(n4102), .Z(n4063) );
  ANDN U4259 ( .A(n2541), .B(n2623), .Z(n4102) );
  XOR U4260 ( .A(n4103), .B(n4104), .Z(n4061) );
  AND U4261 ( .A(n4105), .B(n4106), .Z(n4104) );
  XNOR U4262 ( .A(n4107), .B(n4103), .Z(n4106) );
  XOR U4263 ( .A(n4108), .B(n4065), .Z(n4101) );
  AND U4264 ( .A(n2621), .B(n2534), .Z(n4065) );
  IV U4265 ( .A(n4067), .Z(n4108) );
  XOR U4266 ( .A(n4113), .B(n4114), .Z(n3432) );
  XOR U4267 ( .A(n4115), .B(n4112), .Z(n4113) );
  XNOR U4268 ( .A(n4100), .B(n4099), .Z(n3431) );
  XOR U4269 ( .A(n4116), .B(n4111), .Z(n4099) );
  XNOR U4270 ( .A(n4095), .B(n4097), .Z(n4111) );
  NAND U4271 ( .A(n2988), .B(n2306), .Z(n4097) );
  XNOR U4272 ( .A(n4093), .B(n4117), .Z(n4095) );
  ANDN U4273 ( .A(n2311), .B(n2990), .Z(n4117) );
  XOR U4274 ( .A(n4110), .B(n4098), .Z(n4116) );
  XOR U4275 ( .A(n4121), .B(n4122), .Z(n4098) );
  XOR U4276 ( .A(n4123), .B(n4105), .Z(n4110) );
  XNOR U4277 ( .A(n4103), .B(n4124), .Z(n4105) );
  ANDN U4278 ( .A(n2541), .B(n2743), .Z(n4124) );
  AND U4279 ( .A(n2741), .B(n2534), .Z(n4107) );
  XNOR U4280 ( .A(n4128), .B(n4129), .Z(n4109) );
  AND U4281 ( .A(n4130), .B(n4131), .Z(n4129) );
  XNOR U4282 ( .A(n4126), .B(n4132), .Z(n4131) );
  XNOR U4283 ( .A(n4127), .B(n4128), .Z(n4132) );
  AND U4284 ( .A(n2863), .B(n2534), .Z(n4127) );
  XOR U4285 ( .A(n4125), .B(n4133), .Z(n4126) );
  ANDN U4286 ( .A(n2541), .B(n2865), .Z(n4133) );
  XNOR U4287 ( .A(n4119), .B(n4137), .Z(n4130) );
  XNOR U4288 ( .A(n4120), .B(n4128), .Z(n4137) );
  AND U4289 ( .A(n3120), .B(n2306), .Z(n4120) );
  XOR U4290 ( .A(n4118), .B(n4138), .Z(n4119) );
  ANDN U4291 ( .A(n2311), .B(n3122), .Z(n4138) );
  XOR U4292 ( .A(n4142), .B(n4143), .Z(n4128) );
  AND U4293 ( .A(n4144), .B(n4145), .Z(n4143) );
  XNOR U4294 ( .A(n4135), .B(n4146), .Z(n4145) );
  XNOR U4295 ( .A(n4136), .B(n4142), .Z(n4146) );
  AND U4296 ( .A(n2988), .B(n2534), .Z(n4136) );
  XOR U4297 ( .A(n4134), .B(n4147), .Z(n4135) );
  ANDN U4298 ( .A(n2541), .B(n2990), .Z(n4147) );
  XNOR U4299 ( .A(n4140), .B(n4151), .Z(n4144) );
  XNOR U4300 ( .A(n4141), .B(n4142), .Z(n4151) );
  AND U4301 ( .A(n3252), .B(n2306), .Z(n4141) );
  XOR U4302 ( .A(n4139), .B(n4152), .Z(n4140) );
  ANDN U4303 ( .A(n2311), .B(n3254), .Z(n4152) );
  XOR U4304 ( .A(n4156), .B(n4157), .Z(n4142) );
  AND U4305 ( .A(n4158), .B(n4159), .Z(n4157) );
  XNOR U4306 ( .A(n4149), .B(n4160), .Z(n4159) );
  XNOR U4307 ( .A(n4150), .B(n4156), .Z(n4160) );
  AND U4308 ( .A(n3120), .B(n2534), .Z(n4150) );
  XOR U4309 ( .A(n4148), .B(n4161), .Z(n4149) );
  ANDN U4310 ( .A(n2541), .B(n3122), .Z(n4161) );
  XNOR U4311 ( .A(n4154), .B(n4165), .Z(n4158) );
  XNOR U4312 ( .A(n4155), .B(n4156), .Z(n4165) );
  AND U4313 ( .A(n3391), .B(n2306), .Z(n4155) );
  XOR U4314 ( .A(n4153), .B(n4166), .Z(n4154) );
  ANDN U4315 ( .A(n2311), .B(n3393), .Z(n4166) );
  XNOR U4316 ( .A(n4171), .B(n4163), .Z(n4122) );
  XNOR U4317 ( .A(n4162), .B(n4172), .Z(n4163) );
  ANDN U4318 ( .A(n2541), .B(n3254), .Z(n4172) );
  XNOR U4319 ( .A(n4175), .B(n4173), .Z(n4174) );
  ANDN U4320 ( .A(n2541), .B(n3393), .Z(n4175) );
  XNOR U4321 ( .A(n4170), .B(n4164), .Z(n4171) );
  AND U4322 ( .A(n3252), .B(n2534), .Z(n4164) );
  XNOR U4323 ( .A(n4168), .B(n4169), .Z(n4121) );
  NAND U4324 ( .A(n4179), .B(n2306), .Z(n4169) );
  XNOR U4325 ( .A(n4167), .B(n4180), .Z(n4168) );
  ANDN U4326 ( .A(n2311), .B(n4181), .Z(n4180) );
  NAND U4327 ( .A(A[0]), .B(n4182), .Z(n4167) );
  NANDN U4328 ( .B(n2306), .A(n4183), .Z(n4182) );
  NANDN U4329 ( .B(n4184), .A(n2311), .Z(n4183) );
  IV U4330 ( .A(n2205), .Z(n2306) );
  XNOR U4331 ( .A(n4177), .B(n4178), .Z(n4170) );
  NAND U4332 ( .A(n4179), .B(n2534), .Z(n4178) );
  XNOR U4333 ( .A(n4176), .B(n4187), .Z(n4177) );
  ANDN U4334 ( .A(n2541), .B(n4181), .Z(n4187) );
  NAND U4335 ( .A(A[0]), .B(n4188), .Z(n4176) );
  NANDN U4336 ( .B(n2534), .A(n4189), .Z(n4188) );
  NANDN U4337 ( .B(n4184), .A(n2541), .Z(n4189) );
  IV U4338 ( .A(n2422), .Z(n2534) );
  XNOR U4339 ( .A(n4086), .B(n4085), .Z(n4100) );
  XOR U4340 ( .A(n4192), .B(n4081), .Z(n4085) );
  XNOR U4341 ( .A(n4080), .B(n4193), .Z(n4081) );
  ANDN U4342 ( .A(n2112), .B(n3254), .Z(n4193) );
  XNOR U4343 ( .A(n4196), .B(n4194), .Z(n4195) );
  ANDN U4344 ( .A(n2112), .B(n3393), .Z(n4196) );
  XNOR U4345 ( .A(n4084), .B(n4082), .Z(n4192) );
  AND U4346 ( .A(n3252), .B(n2105), .Z(n4082) );
  XNOR U4347 ( .A(n4198), .B(n4199), .Z(n4084) );
  NAND U4348 ( .A(n4179), .B(n2105), .Z(n4199) );
  XNOR U4349 ( .A(n4197), .B(n4200), .Z(n4198) );
  ANDN U4350 ( .A(n2112), .B(n4181), .Z(n4200) );
  NAND U4351 ( .A(A[0]), .B(n4201), .Z(n4197) );
  NANDN U4352 ( .B(n2105), .A(n4202), .Z(n4201) );
  NANDN U4353 ( .B(n4184), .A(n2112), .Z(n4202) );
  IV U4354 ( .A(n2006), .Z(n2105) );
  XNOR U4355 ( .A(n4089), .B(n4090), .Z(n4086) );
  NAND U4356 ( .A(n4179), .B(n1910), .Z(n4090) );
  XNOR U4357 ( .A(n4088), .B(n4205), .Z(n4089) );
  ANDN U4358 ( .A(n1915), .B(n4181), .Z(n4205) );
  NAND U4359 ( .A(A[0]), .B(n4206), .Z(n4088) );
  NANDN U4360 ( .B(n1910), .A(n4207), .Z(n4206) );
  NANDN U4361 ( .B(n4184), .A(n1915), .Z(n4207) );
  IV U4362 ( .A(n1814), .Z(n1910) );
  XNOR U4363 ( .A(n4210), .B(n4211), .Z(n4112) );
  XOR U4364 ( .A(n4212), .B(n3334), .Z(n3329) );
  XNOR U4365 ( .A(n3325), .B(n3326), .Z(n3334) );
  NAND U4366 ( .A(n3322), .B(n955), .Z(n3326) );
  XNOR U4367 ( .A(n3324), .B(n4213), .Z(n3325) );
  ANDN U4368 ( .A(n3327), .B(n957), .Z(n4213) );
  XOR U4369 ( .A(n4214), .B(n4215), .Z(n3324) );
  AND U4370 ( .A(n4216), .B(n4217), .Z(n4215) );
  XOR U4371 ( .A(n4218), .B(n4214), .Z(n4217) );
  XNOR U4372 ( .A(n3332), .B(n3328), .Z(n4212) );
  XNOR U4373 ( .A(n3443), .B(n3442), .Z(n3455) );
  XOR U4374 ( .A(n4220), .B(n3438), .Z(n3442) );
  XNOR U4375 ( .A(n3436), .B(n4221), .Z(n3438) );
  ANDN U4376 ( .A(n3050), .B(n1085), .Z(n4221) );
  XOR U4377 ( .A(n4222), .B(n4223), .Z(n3436) );
  AND U4378 ( .A(n4224), .B(n4225), .Z(n4223) );
  XNOR U4379 ( .A(n4226), .B(n4222), .Z(n4225) );
  AND U4380 ( .A(n3043), .B(n1083), .Z(n3440) );
  XNOR U4381 ( .A(n3447), .B(n3449), .Z(n3443) );
  NAND U4382 ( .A(n2796), .B(n1184), .Z(n3449) );
  XNOR U4383 ( .A(n3445), .B(n4230), .Z(n3447) );
  ANDN U4384 ( .A(n2801), .B(n1186), .Z(n4230) );
  XOR U4385 ( .A(n4231), .B(n4232), .Z(n3445) );
  AND U4386 ( .A(n4233), .B(n4234), .Z(n4232) );
  XOR U4387 ( .A(n4235), .B(n4231), .Z(n4234) );
  XOR U4388 ( .A(n4236), .B(n4237), .Z(n3456) );
  XNOR U4389 ( .A(n4238), .B(n4219), .Z(n4236) );
  XOR U4390 ( .A(n4240), .B(n4241), .Z(n3494) );
  XOR U4391 ( .A(n4242), .B(n4239), .Z(n4240) );
  XNOR U4392 ( .A(n4229), .B(n4228), .Z(n3492) );
  XOR U4393 ( .A(n4243), .B(n4224), .Z(n4228) );
  XNOR U4394 ( .A(n4222), .B(n4244), .Z(n4224) );
  ANDN U4395 ( .A(n3050), .B(n1127), .Z(n4244) );
  XOR U4396 ( .A(n4245), .B(n4246), .Z(n4222) );
  AND U4397 ( .A(n4247), .B(n4248), .Z(n4246) );
  XNOR U4398 ( .A(n4249), .B(n4245), .Z(n4248) );
  XOR U4399 ( .A(n4250), .B(n4226), .Z(n4243) );
  AND U4400 ( .A(n3043), .B(n1125), .Z(n4226) );
  IV U4401 ( .A(n4227), .Z(n4250) );
  XNOR U4402 ( .A(n4233), .B(n4235), .Z(n4229) );
  NAND U4403 ( .A(n2796), .B(n1248), .Z(n4235) );
  XNOR U4404 ( .A(n4231), .B(n4254), .Z(n4233) );
  ANDN U4405 ( .A(n2801), .B(n1250), .Z(n4254) );
  XOR U4406 ( .A(n4255), .B(n4256), .Z(n4231) );
  AND U4407 ( .A(n4257), .B(n4258), .Z(n4256) );
  XOR U4408 ( .A(n4259), .B(n4255), .Z(n4258) );
  XOR U4409 ( .A(n4261), .B(n4262), .Z(n3539) );
  XOR U4410 ( .A(n4263), .B(n4260), .Z(n4261) );
  XNOR U4411 ( .A(n4253), .B(n4252), .Z(n3537) );
  XOR U4412 ( .A(n4264), .B(n4247), .Z(n4252) );
  XNOR U4413 ( .A(n4245), .B(n4265), .Z(n4247) );
  ANDN U4414 ( .A(n3050), .B(n1186), .Z(n4265) );
  XOR U4415 ( .A(n4266), .B(n4267), .Z(n4245) );
  AND U4416 ( .A(n4268), .B(n4269), .Z(n4267) );
  XNOR U4417 ( .A(n4270), .B(n4266), .Z(n4269) );
  XOR U4418 ( .A(n4271), .B(n4249), .Z(n4264) );
  AND U4419 ( .A(n3043), .B(n1184), .Z(n4249) );
  IV U4420 ( .A(n4251), .Z(n4271) );
  XNOR U4421 ( .A(n4257), .B(n4259), .Z(n4253) );
  NAND U4422 ( .A(n2796), .B(n1316), .Z(n4259) );
  XNOR U4423 ( .A(n4255), .B(n4275), .Z(n4257) );
  ANDN U4424 ( .A(n2801), .B(n1318), .Z(n4275) );
  XOR U4425 ( .A(n4276), .B(n4277), .Z(n4255) );
  AND U4426 ( .A(n4278), .B(n4279), .Z(n4277) );
  XOR U4427 ( .A(n4280), .B(n4276), .Z(n4279) );
  XOR U4428 ( .A(n4282), .B(n4283), .Z(n3581) );
  XOR U4429 ( .A(n4284), .B(n4281), .Z(n4282) );
  XNOR U4430 ( .A(n4274), .B(n4273), .Z(n3579) );
  XOR U4431 ( .A(n4285), .B(n4268), .Z(n4273) );
  XNOR U4432 ( .A(n4266), .B(n4286), .Z(n4268) );
  ANDN U4433 ( .A(n3050), .B(n1250), .Z(n4286) );
  XOR U4434 ( .A(n4287), .B(n4288), .Z(n4266) );
  AND U4435 ( .A(n4289), .B(n4290), .Z(n4288) );
  XNOR U4436 ( .A(n4291), .B(n4287), .Z(n4290) );
  AND U4437 ( .A(n3043), .B(n1248), .Z(n4270) );
  XNOR U4438 ( .A(n4278), .B(n4280), .Z(n4274) );
  NAND U4439 ( .A(n2796), .B(n1383), .Z(n4280) );
  XNOR U4440 ( .A(n4276), .B(n4295), .Z(n4278) );
  ANDN U4441 ( .A(n2801), .B(n1385), .Z(n4295) );
  XOR U4442 ( .A(n4296), .B(n4297), .Z(n4276) );
  AND U4443 ( .A(n4298), .B(n4299), .Z(n4297) );
  XOR U4444 ( .A(n4300), .B(n4296), .Z(n4299) );
  XOR U4445 ( .A(n4302), .B(n4303), .Z(n3624) );
  XOR U4446 ( .A(n4304), .B(n4301), .Z(n4302) );
  XNOR U4447 ( .A(n4294), .B(n4293), .Z(n3622) );
  XOR U4448 ( .A(n4305), .B(n4289), .Z(n4293) );
  XNOR U4449 ( .A(n4287), .B(n4306), .Z(n4289) );
  ANDN U4450 ( .A(n3050), .B(n1318), .Z(n4306) );
  XOR U4451 ( .A(n4307), .B(n4308), .Z(n4287) );
  AND U4452 ( .A(n4309), .B(n4310), .Z(n4308) );
  XNOR U4453 ( .A(n4311), .B(n4307), .Z(n4310) );
  XOR U4454 ( .A(n4312), .B(n4291), .Z(n4305) );
  AND U4455 ( .A(n3043), .B(n1316), .Z(n4291) );
  IV U4456 ( .A(n4292), .Z(n4312) );
  XNOR U4457 ( .A(n4298), .B(n4300), .Z(n4294) );
  NAND U4458 ( .A(n2796), .B(n1457), .Z(n4300) );
  XNOR U4459 ( .A(n4296), .B(n4316), .Z(n4298) );
  ANDN U4460 ( .A(n2801), .B(n1459), .Z(n4316) );
  XOR U4461 ( .A(n4317), .B(n4318), .Z(n4296) );
  AND U4462 ( .A(n4319), .B(n4320), .Z(n4318) );
  XOR U4463 ( .A(n4321), .B(n4317), .Z(n4320) );
  XOR U4464 ( .A(n4323), .B(n4324), .Z(n3666) );
  XOR U4465 ( .A(n4325), .B(n4322), .Z(n4323) );
  XNOR U4466 ( .A(n4315), .B(n4314), .Z(n3664) );
  XOR U4467 ( .A(n4326), .B(n4309), .Z(n4314) );
  XNOR U4468 ( .A(n4307), .B(n4327), .Z(n4309) );
  ANDN U4469 ( .A(n3050), .B(n1385), .Z(n4327) );
  XOR U4470 ( .A(n4328), .B(n4329), .Z(n4307) );
  AND U4471 ( .A(n4330), .B(n4331), .Z(n4329) );
  XNOR U4472 ( .A(n4332), .B(n4328), .Z(n4331) );
  XOR U4473 ( .A(n4333), .B(n4311), .Z(n4326) );
  AND U4474 ( .A(n3043), .B(n1383), .Z(n4311) );
  IV U4475 ( .A(n4313), .Z(n4333) );
  XNOR U4476 ( .A(n4319), .B(n4321), .Z(n4315) );
  NAND U4477 ( .A(n2796), .B(n1535), .Z(n4321) );
  XNOR U4478 ( .A(n4317), .B(n4337), .Z(n4319) );
  ANDN U4479 ( .A(n2801), .B(n1537), .Z(n4337) );
  XOR U4480 ( .A(n4338), .B(n4339), .Z(n4317) );
  AND U4481 ( .A(n4340), .B(n4341), .Z(n4339) );
  XOR U4482 ( .A(n4342), .B(n4338), .Z(n4341) );
  XOR U4483 ( .A(n4344), .B(n4345), .Z(n3712) );
  XOR U4484 ( .A(n4346), .B(n4343), .Z(n4344) );
  XNOR U4485 ( .A(n4336), .B(n4335), .Z(n3710) );
  XOR U4486 ( .A(n4347), .B(n4330), .Z(n4335) );
  XNOR U4487 ( .A(n4328), .B(n4348), .Z(n4330) );
  ANDN U4488 ( .A(n3050), .B(n1459), .Z(n4348) );
  XOR U4489 ( .A(n4349), .B(n4350), .Z(n4328) );
  AND U4490 ( .A(n4351), .B(n4352), .Z(n4350) );
  XNOR U4491 ( .A(n4353), .B(n4349), .Z(n4352) );
  XOR U4492 ( .A(n4354), .B(n4332), .Z(n4347) );
  AND U4493 ( .A(n3043), .B(n1457), .Z(n4332) );
  IV U4494 ( .A(n4334), .Z(n4354) );
  XNOR U4495 ( .A(n4340), .B(n4342), .Z(n4336) );
  NAND U4496 ( .A(n2796), .B(n1616), .Z(n4342) );
  XNOR U4497 ( .A(n4338), .B(n4358), .Z(n4340) );
  ANDN U4498 ( .A(n2801), .B(n1618), .Z(n4358) );
  XOR U4499 ( .A(n4359), .B(n4360), .Z(n4338) );
  AND U4500 ( .A(n4361), .B(n4362), .Z(n4360) );
  XOR U4501 ( .A(n4363), .B(n4359), .Z(n4362) );
  XOR U4502 ( .A(n4365), .B(n4366), .Z(n3756) );
  XOR U4503 ( .A(n4367), .B(n4364), .Z(n4365) );
  XNOR U4504 ( .A(n4357), .B(n4356), .Z(n3754) );
  XOR U4505 ( .A(n4368), .B(n4351), .Z(n4356) );
  XNOR U4506 ( .A(n4349), .B(n4369), .Z(n4351) );
  ANDN U4507 ( .A(n3050), .B(n1537), .Z(n4369) );
  XOR U4508 ( .A(n4370), .B(n4371), .Z(n4349) );
  AND U4509 ( .A(n4372), .B(n4373), .Z(n4371) );
  XNOR U4510 ( .A(n4374), .B(n4370), .Z(n4373) );
  XOR U4511 ( .A(n4375), .B(n4353), .Z(n4368) );
  AND U4512 ( .A(n3043), .B(n1535), .Z(n4353) );
  IV U4513 ( .A(n4355), .Z(n4375) );
  XNOR U4514 ( .A(n4361), .B(n4363), .Z(n4357) );
  NAND U4515 ( .A(n2796), .B(n1700), .Z(n4363) );
  XNOR U4516 ( .A(n4359), .B(n4379), .Z(n4361) );
  ANDN U4517 ( .A(n2801), .B(n1702), .Z(n4379) );
  XOR U4518 ( .A(n4380), .B(n4381), .Z(n4359) );
  AND U4519 ( .A(n4382), .B(n4383), .Z(n4381) );
  XOR U4520 ( .A(n4384), .B(n4380), .Z(n4383) );
  XOR U4521 ( .A(n4386), .B(n4387), .Z(n3802) );
  XOR U4522 ( .A(n4388), .B(n4385), .Z(n4386) );
  XNOR U4523 ( .A(n4378), .B(n4377), .Z(n3800) );
  XOR U4524 ( .A(n4389), .B(n4372), .Z(n4377) );
  XNOR U4525 ( .A(n4370), .B(n4390), .Z(n4372) );
  ANDN U4526 ( .A(n3050), .B(n1618), .Z(n4390) );
  XOR U4527 ( .A(n4391), .B(n4392), .Z(n4370) );
  AND U4528 ( .A(n4393), .B(n4394), .Z(n4392) );
  XNOR U4529 ( .A(n4395), .B(n4391), .Z(n4394) );
  XOR U4530 ( .A(n4396), .B(n4374), .Z(n4389) );
  AND U4531 ( .A(n3043), .B(n1616), .Z(n4374) );
  IV U4532 ( .A(n4376), .Z(n4396) );
  XNOR U4533 ( .A(n4382), .B(n4384), .Z(n4378) );
  NAND U4534 ( .A(n2796), .B(n1791), .Z(n4384) );
  XNOR U4535 ( .A(n4380), .B(n4400), .Z(n4382) );
  ANDN U4536 ( .A(n2801), .B(n1793), .Z(n4400) );
  XOR U4537 ( .A(n4401), .B(n4402), .Z(n4380) );
  AND U4538 ( .A(n4403), .B(n4404), .Z(n4402) );
  XOR U4539 ( .A(n4405), .B(n4401), .Z(n4404) );
  XOR U4540 ( .A(n4407), .B(n4408), .Z(n3848) );
  XOR U4541 ( .A(n4409), .B(n4406), .Z(n4407) );
  XNOR U4542 ( .A(n4399), .B(n4398), .Z(n3846) );
  XOR U4543 ( .A(n4410), .B(n4393), .Z(n4398) );
  XNOR U4544 ( .A(n4391), .B(n4411), .Z(n4393) );
  ANDN U4545 ( .A(n3050), .B(n1702), .Z(n4411) );
  XOR U4546 ( .A(n4412), .B(n4413), .Z(n4391) );
  AND U4547 ( .A(n4414), .B(n4415), .Z(n4413) );
  XNOR U4548 ( .A(n4416), .B(n4412), .Z(n4415) );
  XOR U4549 ( .A(n4417), .B(n4395), .Z(n4410) );
  AND U4550 ( .A(n3043), .B(n1700), .Z(n4395) );
  IV U4551 ( .A(n4397), .Z(n4417) );
  XNOR U4552 ( .A(n4403), .B(n4405), .Z(n4399) );
  NAND U4553 ( .A(n2796), .B(n1888), .Z(n4405) );
  XNOR U4554 ( .A(n4401), .B(n4421), .Z(n4403) );
  ANDN U4555 ( .A(n2801), .B(n1890), .Z(n4421) );
  XOR U4556 ( .A(n4422), .B(n4423), .Z(n4401) );
  AND U4557 ( .A(n4424), .B(n4425), .Z(n4423) );
  XOR U4558 ( .A(n4426), .B(n4422), .Z(n4425) );
  XOR U4559 ( .A(n4428), .B(n4429), .Z(n3894) );
  XOR U4560 ( .A(n4430), .B(n4427), .Z(n4428) );
  XNOR U4561 ( .A(n4420), .B(n4419), .Z(n3892) );
  XOR U4562 ( .A(n4431), .B(n4414), .Z(n4419) );
  XNOR U4563 ( .A(n4412), .B(n4432), .Z(n4414) );
  ANDN U4564 ( .A(n3050), .B(n1793), .Z(n4432) );
  XOR U4565 ( .A(n4433), .B(n4434), .Z(n4412) );
  AND U4566 ( .A(n4435), .B(n4436), .Z(n4434) );
  XNOR U4567 ( .A(n4437), .B(n4433), .Z(n4436) );
  XOR U4568 ( .A(n4438), .B(n4416), .Z(n4431) );
  AND U4569 ( .A(n3043), .B(n1791), .Z(n4416) );
  IV U4570 ( .A(n4418), .Z(n4438) );
  XNOR U4571 ( .A(n4424), .B(n4426), .Z(n4420) );
  NAND U4572 ( .A(n2796), .B(n1984), .Z(n4426) );
  XNOR U4573 ( .A(n4422), .B(n4442), .Z(n4424) );
  ANDN U4574 ( .A(n2801), .B(n1986), .Z(n4442) );
  XOR U4575 ( .A(n4443), .B(n4444), .Z(n4422) );
  AND U4576 ( .A(n4445), .B(n4446), .Z(n4444) );
  XOR U4577 ( .A(n4447), .B(n4443), .Z(n4446) );
  XOR U4578 ( .A(n4449), .B(n4450), .Z(n3938) );
  XOR U4579 ( .A(n4451), .B(n4448), .Z(n4449) );
  XNOR U4580 ( .A(n4441), .B(n4440), .Z(n3936) );
  XOR U4581 ( .A(n4452), .B(n4435), .Z(n4440) );
  XNOR U4582 ( .A(n4433), .B(n4453), .Z(n4435) );
  ANDN U4583 ( .A(n3050), .B(n1890), .Z(n4453) );
  XOR U4584 ( .A(n4454), .B(n4455), .Z(n4433) );
  AND U4585 ( .A(n4456), .B(n4457), .Z(n4455) );
  XNOR U4586 ( .A(n4458), .B(n4454), .Z(n4457) );
  XOR U4587 ( .A(n4459), .B(n4437), .Z(n4452) );
  AND U4588 ( .A(n3043), .B(n1888), .Z(n4437) );
  IV U4589 ( .A(n4439), .Z(n4459) );
  XNOR U4590 ( .A(n4445), .B(n4447), .Z(n4441) );
  NAND U4591 ( .A(n2796), .B(n2080), .Z(n4447) );
  XNOR U4592 ( .A(n4443), .B(n4463), .Z(n4445) );
  ANDN U4593 ( .A(n2801), .B(n2082), .Z(n4463) );
  XOR U4594 ( .A(n4464), .B(n4465), .Z(n4443) );
  AND U4595 ( .A(n4466), .B(n4467), .Z(n4465) );
  XOR U4596 ( .A(n4468), .B(n4464), .Z(n4467) );
  XOR U4597 ( .A(n4470), .B(n4471), .Z(n3984) );
  XOR U4598 ( .A(n4472), .B(n4469), .Z(n4470) );
  XNOR U4599 ( .A(n4462), .B(n4461), .Z(n3982) );
  XOR U4600 ( .A(n4473), .B(n4456), .Z(n4461) );
  XNOR U4601 ( .A(n4454), .B(n4474), .Z(n4456) );
  ANDN U4602 ( .A(n3050), .B(n1986), .Z(n4474) );
  XOR U4603 ( .A(n4475), .B(n4476), .Z(n4454) );
  AND U4604 ( .A(n4477), .B(n4478), .Z(n4476) );
  XNOR U4605 ( .A(n4479), .B(n4475), .Z(n4478) );
  XOR U4606 ( .A(n4480), .B(n4458), .Z(n4473) );
  AND U4607 ( .A(n3043), .B(n1984), .Z(n4458) );
  IV U4608 ( .A(n4460), .Z(n4480) );
  XNOR U4609 ( .A(n4466), .B(n4468), .Z(n4462) );
  NAND U4610 ( .A(n2796), .B(n2181), .Z(n4468) );
  XNOR U4611 ( .A(n4464), .B(n4484), .Z(n4466) );
  ANDN U4612 ( .A(n2801), .B(n2183), .Z(n4484) );
  XOR U4613 ( .A(n4485), .B(n4486), .Z(n4464) );
  AND U4614 ( .A(n4487), .B(n4488), .Z(n4486) );
  XOR U4615 ( .A(n4489), .B(n4485), .Z(n4488) );
  XOR U4616 ( .A(n4491), .B(n4492), .Z(n4030) );
  XOR U4617 ( .A(n4493), .B(n4490), .Z(n4491) );
  XNOR U4618 ( .A(n4483), .B(n4482), .Z(n4028) );
  XOR U4619 ( .A(n4494), .B(n4477), .Z(n4482) );
  XNOR U4620 ( .A(n4475), .B(n4495), .Z(n4477) );
  ANDN U4621 ( .A(n3050), .B(n2082), .Z(n4495) );
  XOR U4622 ( .A(n4496), .B(n4497), .Z(n4475) );
  AND U4623 ( .A(n4498), .B(n4499), .Z(n4497) );
  XNOR U4624 ( .A(n4500), .B(n4496), .Z(n4499) );
  XOR U4625 ( .A(n4501), .B(n4479), .Z(n4494) );
  AND U4626 ( .A(n3043), .B(n2080), .Z(n4479) );
  IV U4627 ( .A(n4481), .Z(n4501) );
  XNOR U4628 ( .A(n4487), .B(n4489), .Z(n4483) );
  NAND U4629 ( .A(n2796), .B(n2287), .Z(n4489) );
  XNOR U4630 ( .A(n4485), .B(n4505), .Z(n4487) );
  ANDN U4631 ( .A(n2801), .B(n2289), .Z(n4505) );
  XOR U4632 ( .A(n4506), .B(n4507), .Z(n4485) );
  AND U4633 ( .A(n4508), .B(n4509), .Z(n4507) );
  XOR U4634 ( .A(n4510), .B(n4506), .Z(n4509) );
  XOR U4635 ( .A(n4512), .B(n4513), .Z(n4076) );
  XOR U4636 ( .A(n4514), .B(n4511), .Z(n4512) );
  XNOR U4637 ( .A(n4504), .B(n4503), .Z(n4074) );
  XOR U4638 ( .A(n4515), .B(n4498), .Z(n4503) );
  XNOR U4639 ( .A(n4496), .B(n4516), .Z(n4498) );
  ANDN U4640 ( .A(n3050), .B(n2183), .Z(n4516) );
  XOR U4641 ( .A(n4517), .B(n4518), .Z(n4496) );
  AND U4642 ( .A(n4519), .B(n4520), .Z(n4518) );
  XNOR U4643 ( .A(n4521), .B(n4517), .Z(n4520) );
  XOR U4644 ( .A(n4522), .B(n4500), .Z(n4515) );
  AND U4645 ( .A(n3043), .B(n2181), .Z(n4500) );
  IV U4646 ( .A(n4502), .Z(n4522) );
  XNOR U4647 ( .A(n4508), .B(n4510), .Z(n4504) );
  NAND U4648 ( .A(n2796), .B(n2394), .Z(n4510) );
  XNOR U4649 ( .A(n4506), .B(n4526), .Z(n4508) );
  ANDN U4650 ( .A(n2801), .B(n2396), .Z(n4526) );
  XOR U4651 ( .A(n4527), .B(n4528), .Z(n4506) );
  AND U4652 ( .A(n4529), .B(n4530), .Z(n4528) );
  XOR U4653 ( .A(n4531), .B(n4527), .Z(n4530) );
  XOR U4654 ( .A(n4533), .B(n4534), .Z(n4115) );
  XOR U4655 ( .A(n4535), .B(n4532), .Z(n4533) );
  XNOR U4656 ( .A(n4525), .B(n4524), .Z(n4114) );
  XOR U4657 ( .A(n4536), .B(n4519), .Z(n4524) );
  XNOR U4658 ( .A(n4517), .B(n4537), .Z(n4519) );
  ANDN U4659 ( .A(n3050), .B(n2289), .Z(n4537) );
  AND U4660 ( .A(n3043), .B(n2287), .Z(n4521) );
  XNOR U4661 ( .A(n4529), .B(n4531), .Z(n4525) );
  NAND U4662 ( .A(n2796), .B(n2502), .Z(n4531) );
  XNOR U4663 ( .A(n4527), .B(n4544), .Z(n4529) );
  ANDN U4664 ( .A(n2801), .B(n2504), .Z(n4544) );
  XOR U4665 ( .A(n4548), .B(n4549), .Z(n4532) );
  AND U4666 ( .A(n4550), .B(n4551), .Z(n4549) );
  XOR U4667 ( .A(n4552), .B(n4553), .Z(n4551) );
  XNOR U4668 ( .A(n4548), .B(n4554), .Z(n4553) );
  XNOR U4669 ( .A(n4542), .B(n4555), .Z(n4550) );
  XNOR U4670 ( .A(n4548), .B(n4543), .Z(n4555) );
  XNOR U4671 ( .A(n4546), .B(n4547), .Z(n4543) );
  NAND U4672 ( .A(n2621), .B(n2796), .Z(n4547) );
  XNOR U4673 ( .A(n4545), .B(n4556), .Z(n4546) );
  ANDN U4674 ( .A(n2801), .B(n2623), .Z(n4556) );
  XOR U4675 ( .A(n4560), .B(n4539), .Z(n4542) );
  XNOR U4676 ( .A(n4538), .B(n4561), .Z(n4539) );
  ANDN U4677 ( .A(n3050), .B(n2396), .Z(n4561) );
  AND U4678 ( .A(n3043), .B(n2394), .Z(n4540) );
  XOR U4679 ( .A(n4568), .B(n4569), .Z(n4548) );
  AND U4680 ( .A(n4570), .B(n4571), .Z(n4569) );
  XOR U4681 ( .A(n4572), .B(n4573), .Z(n4571) );
  XNOR U4682 ( .A(n4568), .B(n4574), .Z(n4573) );
  XNOR U4683 ( .A(n4566), .B(n4575), .Z(n4570) );
  XNOR U4684 ( .A(n4568), .B(n4567), .Z(n4575) );
  XNOR U4685 ( .A(n4558), .B(n4559), .Z(n4567) );
  NAND U4686 ( .A(n2741), .B(n2796), .Z(n4559) );
  XNOR U4687 ( .A(n4557), .B(n4576), .Z(n4558) );
  ANDN U4688 ( .A(n2801), .B(n2743), .Z(n4576) );
  XOR U4689 ( .A(n4580), .B(n4563), .Z(n4566) );
  XNOR U4690 ( .A(n4562), .B(n4581), .Z(n4563) );
  ANDN U4691 ( .A(n3050), .B(n2504), .Z(n4581) );
  AND U4692 ( .A(n3043), .B(n2502), .Z(n4564) );
  XOR U4693 ( .A(n4588), .B(n4589), .Z(n4568) );
  AND U4694 ( .A(n4590), .B(n4591), .Z(n4589) );
  XOR U4695 ( .A(n4592), .B(n4593), .Z(n4591) );
  XNOR U4696 ( .A(n4588), .B(n4594), .Z(n4593) );
  XNOR U4697 ( .A(n4586), .B(n4595), .Z(n4590) );
  XNOR U4698 ( .A(n4588), .B(n4587), .Z(n4595) );
  XNOR U4699 ( .A(n4578), .B(n4579), .Z(n4587) );
  NAND U4700 ( .A(n2863), .B(n2796), .Z(n4579) );
  XNOR U4701 ( .A(n4577), .B(n4596), .Z(n4578) );
  ANDN U4702 ( .A(n2801), .B(n2865), .Z(n4596) );
  XOR U4703 ( .A(n4600), .B(n4583), .Z(n4586) );
  XNOR U4704 ( .A(n4582), .B(n4601), .Z(n4583) );
  ANDN U4705 ( .A(n3050), .B(n2623), .Z(n4601) );
  AND U4706 ( .A(n2621), .B(n3043), .Z(n4584) );
  XOR U4707 ( .A(n4608), .B(n4609), .Z(n4588) );
  AND U4708 ( .A(n4610), .B(n4611), .Z(n4609) );
  XOR U4709 ( .A(n4612), .B(n4613), .Z(n4611) );
  XNOR U4710 ( .A(n4608), .B(n4614), .Z(n4613) );
  XNOR U4711 ( .A(n4606), .B(n4615), .Z(n4610) );
  XNOR U4712 ( .A(n4608), .B(n4607), .Z(n4615) );
  XNOR U4713 ( .A(n4598), .B(n4599), .Z(n4607) );
  NAND U4714 ( .A(n2988), .B(n2796), .Z(n4599) );
  XNOR U4715 ( .A(n4597), .B(n4616), .Z(n4598) );
  ANDN U4716 ( .A(n2801), .B(n2990), .Z(n4616) );
  XOR U4717 ( .A(n4620), .B(n4603), .Z(n4606) );
  XNOR U4718 ( .A(n4602), .B(n4621), .Z(n4603) );
  ANDN U4719 ( .A(n3050), .B(n2743), .Z(n4621) );
  AND U4720 ( .A(n2741), .B(n3043), .Z(n4604) );
  XOR U4721 ( .A(n4628), .B(n4629), .Z(n4608) );
  AND U4722 ( .A(n4630), .B(n4631), .Z(n4629) );
  XOR U4723 ( .A(n4632), .B(n4633), .Z(n4631) );
  XNOR U4724 ( .A(n4628), .B(n4634), .Z(n4633) );
  XNOR U4725 ( .A(n4626), .B(n4635), .Z(n4630) );
  XNOR U4726 ( .A(n4628), .B(n4627), .Z(n4635) );
  XNOR U4727 ( .A(n4618), .B(n4619), .Z(n4627) );
  NAND U4728 ( .A(n3120), .B(n2796), .Z(n4619) );
  XNOR U4729 ( .A(n4617), .B(n4636), .Z(n4618) );
  ANDN U4730 ( .A(n2801), .B(n3122), .Z(n4636) );
  XOR U4731 ( .A(n4640), .B(n4623), .Z(n4626) );
  XNOR U4732 ( .A(n4622), .B(n4641), .Z(n4623) );
  ANDN U4733 ( .A(n3050), .B(n2865), .Z(n4641) );
  AND U4734 ( .A(n2863), .B(n3043), .Z(n4624) );
  XOR U4735 ( .A(n4648), .B(n4649), .Z(n4628) );
  AND U4736 ( .A(n4650), .B(n4651), .Z(n4649) );
  XOR U4737 ( .A(n4652), .B(n4653), .Z(n4651) );
  XNOR U4738 ( .A(n4648), .B(n4654), .Z(n4653) );
  XNOR U4739 ( .A(n4646), .B(n4655), .Z(n4650) );
  XNOR U4740 ( .A(n4648), .B(n4647), .Z(n4655) );
  XNOR U4741 ( .A(n4638), .B(n4639), .Z(n4647) );
  NAND U4742 ( .A(n3252), .B(n2796), .Z(n4639) );
  XNOR U4743 ( .A(n4637), .B(n4656), .Z(n4638) );
  ANDN U4744 ( .A(n2801), .B(n3254), .Z(n4656) );
  XOR U4745 ( .A(n4657), .B(n4658), .Z(n4637) );
  AND U4746 ( .A(n4659), .B(n4660), .Z(n4658) );
  XOR U4747 ( .A(n4661), .B(n4657), .Z(n4660) );
  XOR U4748 ( .A(n4662), .B(n4643), .Z(n4646) );
  XNOR U4749 ( .A(n4642), .B(n4663), .Z(n4643) );
  ANDN U4750 ( .A(n3050), .B(n2990), .Z(n4663) );
  XOR U4751 ( .A(n4664), .B(n4665), .Z(n4642) );
  AND U4752 ( .A(n4666), .B(n4667), .Z(n4665) );
  XNOR U4753 ( .A(n4668), .B(n4664), .Z(n4667) );
  AND U4754 ( .A(n2988), .B(n3043), .Z(n4644) );
  XOR U4755 ( .A(n4672), .B(n4673), .Z(n4648) );
  AND U4756 ( .A(n4674), .B(n4675), .Z(n4673) );
  XOR U4757 ( .A(n4676), .B(n4677), .Z(n4675) );
  XNOR U4758 ( .A(n4672), .B(n4678), .Z(n4677) );
  XNOR U4759 ( .A(n4670), .B(n4679), .Z(n4674) );
  XNOR U4760 ( .A(n4672), .B(n4671), .Z(n4679) );
  XNOR U4761 ( .A(n4659), .B(n4661), .Z(n4671) );
  NAND U4762 ( .A(n3391), .B(n2796), .Z(n4661) );
  XNOR U4763 ( .A(n4657), .B(n4680), .Z(n4659) );
  ANDN U4764 ( .A(n2801), .B(n3393), .Z(n4680) );
  XOR U4765 ( .A(n4684), .B(n4666), .Z(n4670) );
  XNOR U4766 ( .A(n4664), .B(n4685), .Z(n4666) );
  ANDN U4767 ( .A(n3050), .B(n3122), .Z(n4685) );
  XOR U4768 ( .A(n4686), .B(n4687), .Z(n4664) );
  AND U4769 ( .A(n4688), .B(n4689), .Z(n4687) );
  XNOR U4770 ( .A(n4690), .B(n4686), .Z(n4689) );
  AND U4771 ( .A(n3120), .B(n3043), .Z(n4668) );
  XOR U4772 ( .A(n4695), .B(n4696), .Z(n4211) );
  XNOR U4773 ( .A(n4693), .B(n4692), .Z(n4210) );
  XOR U4774 ( .A(n4698), .B(n4688), .Z(n4692) );
  XNOR U4775 ( .A(n4686), .B(n4699), .Z(n4688) );
  ANDN U4776 ( .A(n3050), .B(n3254), .Z(n4699) );
  XNOR U4777 ( .A(n4702), .B(n4700), .Z(n4701) );
  ANDN U4778 ( .A(n3050), .B(n3393), .Z(n4702) );
  XNOR U4779 ( .A(n4691), .B(n4690), .Z(n4698) );
  AND U4780 ( .A(n3252), .B(n3043), .Z(n4690) );
  XNOR U4781 ( .A(n4704), .B(n4705), .Z(n4691) );
  NAND U4782 ( .A(n4179), .B(n3043), .Z(n4705) );
  XNOR U4783 ( .A(n4703), .B(n4706), .Z(n4704) );
  ANDN U4784 ( .A(n3050), .B(n4181), .Z(n4706) );
  NAND U4785 ( .A(A[0]), .B(n4707), .Z(n4703) );
  NANDN U4786 ( .B(n3043), .A(n4708), .Z(n4707) );
  NANDN U4787 ( .B(n4184), .A(n3050), .Z(n4708) );
  IV U4788 ( .A(n2917), .Z(n3043) );
  XNOR U4789 ( .A(n4682), .B(n4683), .Z(n4693) );
  NAND U4790 ( .A(n4179), .B(n2796), .Z(n4683) );
  XNOR U4791 ( .A(n4681), .B(n4711), .Z(n4682) );
  ANDN U4792 ( .A(n2801), .B(n4181), .Z(n4711) );
  NAND U4793 ( .A(A[0]), .B(n4712), .Z(n4681) );
  NANDN U4794 ( .B(n2796), .A(n4713), .Z(n4712) );
  NANDN U4795 ( .B(n4184), .A(n2801), .Z(n4713) );
  IV U4796 ( .A(n2675), .Z(n2796) );
  XOR U4797 ( .A(n4716), .B(n4717), .Z(n4694) );
  XOR U4798 ( .A(n3331), .B(n4718), .Z(n3332) );
  AND U4799 ( .A(n4719), .B(n4720), .Z(n4718) );
  NANDN U4800 ( .B(n4721), .A(n894), .Z(n4720) );
  NANDN U4801 ( .B(n4722), .A(n4723), .Z(n4719) );
  XNOR U4802 ( .A(n4216), .B(n4218), .Z(n4237) );
  NAND U4803 ( .A(n3322), .B(n999), .Z(n4218) );
  XNOR U4804 ( .A(n4214), .B(n4725), .Z(n4216) );
  ANDN U4805 ( .A(n3327), .B(n1001), .Z(n4725) );
  XOR U4806 ( .A(n4726), .B(n4727), .Z(n4214) );
  AND U4807 ( .A(n4728), .B(n4729), .Z(n4727) );
  XOR U4808 ( .A(n4730), .B(n4726), .Z(n4729) );
  XNOR U4809 ( .A(n4731), .B(n4732), .Z(n4238) );
  IV U4810 ( .A(n4724), .Z(n4732) );
  XOR U4811 ( .A(n4733), .B(n4723), .Z(n4731) );
  AND U4812 ( .A(n4734), .B(n924), .Z(n4723) );
  IV U4813 ( .A(n957), .Z(n924) );
  NAND U4814 ( .A(n4735), .B(n4722), .Z(n4733) );
  XOR U4815 ( .A(n4736), .B(n4737), .Z(n4722) );
  AND U4816 ( .A(n4738), .B(n4739), .Z(n4737) );
  XNOR U4817 ( .A(n4740), .B(n4736), .Z(n4739) );
  NANDN U4818 ( .B(n927), .A(X[0]), .Z(n4735) );
  IV U4819 ( .A(n894), .Z(n927) );
  AND U4820 ( .A(n4741), .B(n4742), .Z(n894) );
  AND U4821 ( .A(A[31]), .B(n4743), .Z(n4741) );
  XNOR U4822 ( .A(n4728), .B(n4730), .Z(n4241) );
  NAND U4823 ( .A(n3322), .B(n1039), .Z(n4730) );
  XNOR U4824 ( .A(n4726), .B(n4745), .Z(n4728) );
  ANDN U4825 ( .A(n3327), .B(n1041), .Z(n4745) );
  XOR U4826 ( .A(n4746), .B(n4747), .Z(n4726) );
  AND U4827 ( .A(n4748), .B(n4749), .Z(n4747) );
  XOR U4828 ( .A(n4750), .B(n4746), .Z(n4749) );
  XNOR U4829 ( .A(n4751), .B(n4738), .Z(n4242) );
  XNOR U4830 ( .A(n4736), .B(n4752), .Z(n4738) );
  ANDN U4831 ( .A(X[0]), .B(n957), .Z(n4752) );
  XOR U4832 ( .A(n4743), .B(A[30]), .Z(n4742) );
  ANDN U4833 ( .A(n4753), .B(n4754), .Z(n4743) );
  XOR U4834 ( .A(n4755), .B(n4756), .Z(n4736) );
  AND U4835 ( .A(n4757), .B(n4758), .Z(n4756) );
  XNOR U4836 ( .A(n4759), .B(n4755), .Z(n4758) );
  XOR U4837 ( .A(n4760), .B(n4740), .Z(n4751) );
  AND U4838 ( .A(n4734), .B(n955), .Z(n4740) );
  IV U4839 ( .A(n1001), .Z(n955) );
  IV U4840 ( .A(n4744), .Z(n4760) );
  XNOR U4841 ( .A(n4748), .B(n4750), .Z(n4262) );
  NAND U4842 ( .A(n3322), .B(n1083), .Z(n4750) );
  XNOR U4843 ( .A(n4746), .B(n4762), .Z(n4748) );
  ANDN U4844 ( .A(n3327), .B(n1085), .Z(n4762) );
  XOR U4845 ( .A(n4763), .B(n4764), .Z(n4746) );
  AND U4846 ( .A(n4765), .B(n4766), .Z(n4764) );
  XOR U4847 ( .A(n4767), .B(n4763), .Z(n4766) );
  XNOR U4848 ( .A(n4768), .B(n4757), .Z(n4263) );
  XNOR U4849 ( .A(n4755), .B(n4769), .Z(n4757) );
  ANDN U4850 ( .A(X[0]), .B(n1001), .Z(n4769) );
  ANDN U4851 ( .A(n4770), .B(n4771), .Z(n4753) );
  XOR U4852 ( .A(n4772), .B(n4773), .Z(n4755) );
  AND U4853 ( .A(n4774), .B(n4775), .Z(n4773) );
  XNOR U4854 ( .A(n4776), .B(n4772), .Z(n4775) );
  XOR U4855 ( .A(n4777), .B(n4759), .Z(n4768) );
  AND U4856 ( .A(n4734), .B(n999), .Z(n4759) );
  IV U4857 ( .A(n1041), .Z(n999) );
  IV U4858 ( .A(n4761), .Z(n4777) );
  XNOR U4859 ( .A(n4765), .B(n4767), .Z(n4283) );
  NAND U4860 ( .A(n3322), .B(n1125), .Z(n4767) );
  XNOR U4861 ( .A(n4763), .B(n4779), .Z(n4765) );
  ANDN U4862 ( .A(n3327), .B(n1127), .Z(n4779) );
  XOR U4863 ( .A(n4780), .B(n4781), .Z(n4763) );
  AND U4864 ( .A(n4782), .B(n4783), .Z(n4781) );
  XOR U4865 ( .A(n4784), .B(n4780), .Z(n4783) );
  XNOR U4866 ( .A(n4785), .B(n4774), .Z(n4284) );
  XNOR U4867 ( .A(n4772), .B(n4786), .Z(n4774) );
  ANDN U4868 ( .A(X[0]), .B(n1041), .Z(n4786) );
  XNOR U4869 ( .A(n4770), .B(A[28]), .Z(n4771) );
  ANDN U4870 ( .A(n4787), .B(n4788), .Z(n4770) );
  XOR U4871 ( .A(n4789), .B(n4790), .Z(n4772) );
  AND U4872 ( .A(n4791), .B(n4792), .Z(n4790) );
  XNOR U4873 ( .A(n4793), .B(n4789), .Z(n4792) );
  AND U4874 ( .A(n4734), .B(n1039), .Z(n4776) );
  IV U4875 ( .A(n1085), .Z(n1039) );
  XNOR U4876 ( .A(n4782), .B(n4784), .Z(n4303) );
  NAND U4877 ( .A(n3322), .B(n1184), .Z(n4784) );
  XNOR U4878 ( .A(n4780), .B(n4795), .Z(n4782) );
  ANDN U4879 ( .A(n3327), .B(n1186), .Z(n4795) );
  XOR U4880 ( .A(n4796), .B(n4797), .Z(n4780) );
  AND U4881 ( .A(n4798), .B(n4799), .Z(n4797) );
  XOR U4882 ( .A(n4800), .B(n4796), .Z(n4799) );
  XNOR U4883 ( .A(n4801), .B(n4791), .Z(n4304) );
  XNOR U4884 ( .A(n4789), .B(n4802), .Z(n4791) );
  ANDN U4885 ( .A(X[0]), .B(n1085), .Z(n4802) );
  ANDN U4886 ( .A(n4803), .B(n4804), .Z(n4787) );
  XOR U4887 ( .A(n4805), .B(n4806), .Z(n4789) );
  AND U4888 ( .A(n4807), .B(n4808), .Z(n4806) );
  XNOR U4889 ( .A(n4809), .B(n4805), .Z(n4808) );
  AND U4890 ( .A(n4734), .B(n1083), .Z(n4793) );
  IV U4891 ( .A(n1127), .Z(n1083) );
  XNOR U4892 ( .A(n4798), .B(n4800), .Z(n4324) );
  NAND U4893 ( .A(n3322), .B(n1248), .Z(n4800) );
  XNOR U4894 ( .A(n4796), .B(n4811), .Z(n4798) );
  ANDN U4895 ( .A(n3327), .B(n1250), .Z(n4811) );
  XOR U4896 ( .A(n4812), .B(n4813), .Z(n4796) );
  AND U4897 ( .A(n4814), .B(n4815), .Z(n4813) );
  XOR U4898 ( .A(n4816), .B(n4812), .Z(n4815) );
  XNOR U4899 ( .A(n4817), .B(n4807), .Z(n4325) );
  XNOR U4900 ( .A(n4805), .B(n4818), .Z(n4807) );
  ANDN U4901 ( .A(X[0]), .B(n1127), .Z(n4818) );
  XNOR U4902 ( .A(n4803), .B(A[26]), .Z(n4804) );
  ANDN U4903 ( .A(n4819), .B(n4820), .Z(n4803) );
  XOR U4904 ( .A(n4821), .B(n4822), .Z(n4805) );
  AND U4905 ( .A(n4823), .B(n4824), .Z(n4822) );
  XNOR U4906 ( .A(n4825), .B(n4821), .Z(n4824) );
  XOR U4907 ( .A(n4826), .B(n4809), .Z(n4817) );
  AND U4908 ( .A(n4734), .B(n1125), .Z(n4809) );
  IV U4909 ( .A(n1186), .Z(n1125) );
  IV U4910 ( .A(n4810), .Z(n4826) );
  XNOR U4911 ( .A(n4814), .B(n4816), .Z(n4345) );
  NAND U4912 ( .A(n3322), .B(n1316), .Z(n4816) );
  XNOR U4913 ( .A(n4812), .B(n4828), .Z(n4814) );
  ANDN U4914 ( .A(n3327), .B(n1318), .Z(n4828) );
  XOR U4915 ( .A(n4829), .B(n4830), .Z(n4812) );
  AND U4916 ( .A(n4831), .B(n4832), .Z(n4830) );
  XOR U4917 ( .A(n4833), .B(n4829), .Z(n4832) );
  XNOR U4918 ( .A(n4834), .B(n4823), .Z(n4346) );
  XNOR U4919 ( .A(n4821), .B(n4835), .Z(n4823) );
  ANDN U4920 ( .A(X[0]), .B(n1186), .Z(n4835) );
  ANDN U4921 ( .A(n4836), .B(n4837), .Z(n4819) );
  XOR U4922 ( .A(n4838), .B(n4839), .Z(n4821) );
  AND U4923 ( .A(n4840), .B(n4841), .Z(n4839) );
  XNOR U4924 ( .A(n4842), .B(n4838), .Z(n4841) );
  XOR U4925 ( .A(n4843), .B(n4825), .Z(n4834) );
  AND U4926 ( .A(n4734), .B(n1184), .Z(n4825) );
  IV U4927 ( .A(n1250), .Z(n1184) );
  IV U4928 ( .A(n4827), .Z(n4843) );
  XNOR U4929 ( .A(n4831), .B(n4833), .Z(n4366) );
  NAND U4930 ( .A(n3322), .B(n1383), .Z(n4833) );
  XNOR U4931 ( .A(n4829), .B(n4845), .Z(n4831) );
  ANDN U4932 ( .A(n3327), .B(n1385), .Z(n4845) );
  XOR U4933 ( .A(n4846), .B(n4847), .Z(n4829) );
  AND U4934 ( .A(n4848), .B(n4849), .Z(n4847) );
  XOR U4935 ( .A(n4850), .B(n4846), .Z(n4849) );
  XNOR U4936 ( .A(n4851), .B(n4840), .Z(n4367) );
  XNOR U4937 ( .A(n4838), .B(n4852), .Z(n4840) );
  ANDN U4938 ( .A(X[0]), .B(n1250), .Z(n4852) );
  XNOR U4939 ( .A(n4836), .B(A[24]), .Z(n4837) );
  ANDN U4940 ( .A(n4853), .B(n4854), .Z(n4836) );
  XOR U4941 ( .A(n4855), .B(n4856), .Z(n4838) );
  AND U4942 ( .A(n4857), .B(n4858), .Z(n4856) );
  XNOR U4943 ( .A(n4859), .B(n4855), .Z(n4858) );
  XOR U4944 ( .A(n4860), .B(n4842), .Z(n4851) );
  AND U4945 ( .A(n4734), .B(n1248), .Z(n4842) );
  IV U4946 ( .A(n1318), .Z(n1248) );
  IV U4947 ( .A(n4844), .Z(n4860) );
  XNOR U4948 ( .A(n4848), .B(n4850), .Z(n4387) );
  NAND U4949 ( .A(n3322), .B(n1457), .Z(n4850) );
  XNOR U4950 ( .A(n4846), .B(n4862), .Z(n4848) );
  ANDN U4951 ( .A(n3327), .B(n1459), .Z(n4862) );
  XOR U4952 ( .A(n4863), .B(n4864), .Z(n4846) );
  AND U4953 ( .A(n4865), .B(n4866), .Z(n4864) );
  XOR U4954 ( .A(n4867), .B(n4863), .Z(n4866) );
  XNOR U4955 ( .A(n4868), .B(n4857), .Z(n4388) );
  XNOR U4956 ( .A(n4855), .B(n4869), .Z(n4857) );
  ANDN U4957 ( .A(X[0]), .B(n1318), .Z(n4869) );
  ANDN U4958 ( .A(n4870), .B(n4871), .Z(n4853) );
  XOR U4959 ( .A(n4872), .B(n4873), .Z(n4855) );
  AND U4960 ( .A(n4874), .B(n4875), .Z(n4873) );
  XNOR U4961 ( .A(n4876), .B(n4872), .Z(n4875) );
  XOR U4962 ( .A(n4877), .B(n4859), .Z(n4868) );
  AND U4963 ( .A(n4734), .B(n1316), .Z(n4859) );
  IV U4964 ( .A(n1385), .Z(n1316) );
  IV U4965 ( .A(n4861), .Z(n4877) );
  XNOR U4966 ( .A(n4865), .B(n4867), .Z(n4408) );
  NAND U4967 ( .A(n3322), .B(n1535), .Z(n4867) );
  XNOR U4968 ( .A(n4863), .B(n4879), .Z(n4865) );
  ANDN U4969 ( .A(n3327), .B(n1537), .Z(n4879) );
  XOR U4970 ( .A(n4880), .B(n4881), .Z(n4863) );
  AND U4971 ( .A(n4882), .B(n4883), .Z(n4881) );
  XOR U4972 ( .A(n4884), .B(n4880), .Z(n4883) );
  XNOR U4973 ( .A(n4885), .B(n4874), .Z(n4409) );
  XNOR U4974 ( .A(n4872), .B(n4886), .Z(n4874) );
  ANDN U4975 ( .A(X[0]), .B(n1385), .Z(n4886) );
  XNOR U4976 ( .A(n4870), .B(A[22]), .Z(n4871) );
  ANDN U4977 ( .A(n4887), .B(n4888), .Z(n4870) );
  XOR U4978 ( .A(n4889), .B(n4890), .Z(n4872) );
  AND U4979 ( .A(n4891), .B(n4892), .Z(n4890) );
  XNOR U4980 ( .A(n4893), .B(n4889), .Z(n4892) );
  XOR U4981 ( .A(n4894), .B(n4876), .Z(n4885) );
  AND U4982 ( .A(n4734), .B(n1383), .Z(n4876) );
  IV U4983 ( .A(n1459), .Z(n1383) );
  IV U4984 ( .A(n4878), .Z(n4894) );
  XNOR U4985 ( .A(n4882), .B(n4884), .Z(n4429) );
  NAND U4986 ( .A(n3322), .B(n1616), .Z(n4884) );
  XNOR U4987 ( .A(n4880), .B(n4896), .Z(n4882) );
  ANDN U4988 ( .A(n3327), .B(n1618), .Z(n4896) );
  XOR U4989 ( .A(n4897), .B(n4898), .Z(n4880) );
  AND U4990 ( .A(n4899), .B(n4900), .Z(n4898) );
  XOR U4991 ( .A(n4901), .B(n4897), .Z(n4900) );
  XNOR U4992 ( .A(n4902), .B(n4891), .Z(n4430) );
  XNOR U4993 ( .A(n4889), .B(n4903), .Z(n4891) );
  ANDN U4994 ( .A(X[0]), .B(n1459), .Z(n4903) );
  ANDN U4995 ( .A(n4904), .B(n4905), .Z(n4887) );
  XOR U4996 ( .A(n4906), .B(n4907), .Z(n4889) );
  AND U4997 ( .A(n4908), .B(n4909), .Z(n4907) );
  XNOR U4998 ( .A(n4910), .B(n4906), .Z(n4909) );
  XOR U4999 ( .A(n4911), .B(n4893), .Z(n4902) );
  AND U5000 ( .A(n4734), .B(n1457), .Z(n4893) );
  IV U5001 ( .A(n1537), .Z(n1457) );
  IV U5002 ( .A(n4895), .Z(n4911) );
  XNOR U5003 ( .A(n4899), .B(n4901), .Z(n4450) );
  NAND U5004 ( .A(n3322), .B(n1700), .Z(n4901) );
  XNOR U5005 ( .A(n4897), .B(n4913), .Z(n4899) );
  ANDN U5006 ( .A(n3327), .B(n1702), .Z(n4913) );
  XOR U5007 ( .A(n4914), .B(n4915), .Z(n4897) );
  AND U5008 ( .A(n4916), .B(n4917), .Z(n4915) );
  XOR U5009 ( .A(n4918), .B(n4914), .Z(n4917) );
  XNOR U5010 ( .A(n4919), .B(n4908), .Z(n4451) );
  XNOR U5011 ( .A(n4906), .B(n4920), .Z(n4908) );
  ANDN U5012 ( .A(X[0]), .B(n1537), .Z(n4920) );
  XNOR U5013 ( .A(n4904), .B(A[20]), .Z(n4905) );
  ANDN U5014 ( .A(n4921), .B(n4922), .Z(n4904) );
  XOR U5015 ( .A(n4923), .B(n4924), .Z(n4906) );
  AND U5016 ( .A(n4925), .B(n4926), .Z(n4924) );
  XNOR U5017 ( .A(n4927), .B(n4923), .Z(n4926) );
  XOR U5018 ( .A(n4928), .B(n4910), .Z(n4919) );
  AND U5019 ( .A(n4734), .B(n1535), .Z(n4910) );
  IV U5020 ( .A(n1618), .Z(n1535) );
  IV U5021 ( .A(n4912), .Z(n4928) );
  XNOR U5022 ( .A(n4916), .B(n4918), .Z(n4471) );
  NAND U5023 ( .A(n3322), .B(n1791), .Z(n4918) );
  XNOR U5024 ( .A(n4914), .B(n4930), .Z(n4916) );
  ANDN U5025 ( .A(n3327), .B(n1793), .Z(n4930) );
  XOR U5026 ( .A(n4931), .B(n4932), .Z(n4914) );
  AND U5027 ( .A(n4933), .B(n4934), .Z(n4932) );
  XOR U5028 ( .A(n4935), .B(n4931), .Z(n4934) );
  XNOR U5029 ( .A(n4936), .B(n4925), .Z(n4472) );
  XNOR U5030 ( .A(n4923), .B(n4937), .Z(n4925) );
  ANDN U5031 ( .A(X[0]), .B(n1618), .Z(n4937) );
  ANDN U5032 ( .A(n4938), .B(n4939), .Z(n4921) );
  XOR U5033 ( .A(n4940), .B(n4941), .Z(n4923) );
  AND U5034 ( .A(n4942), .B(n4943), .Z(n4941) );
  XNOR U5035 ( .A(n4944), .B(n4940), .Z(n4943) );
  XOR U5036 ( .A(n4945), .B(n4927), .Z(n4936) );
  AND U5037 ( .A(n4734), .B(n1616), .Z(n4927) );
  IV U5038 ( .A(n1702), .Z(n1616) );
  IV U5039 ( .A(n4929), .Z(n4945) );
  XNOR U5040 ( .A(n4933), .B(n4935), .Z(n4492) );
  NAND U5041 ( .A(n3322), .B(n1888), .Z(n4935) );
  XNOR U5042 ( .A(n4931), .B(n4947), .Z(n4933) );
  ANDN U5043 ( .A(n3327), .B(n1890), .Z(n4947) );
  XOR U5044 ( .A(n4948), .B(n4949), .Z(n4931) );
  AND U5045 ( .A(n4950), .B(n4951), .Z(n4949) );
  XOR U5046 ( .A(n4952), .B(n4948), .Z(n4951) );
  XNOR U5047 ( .A(n4953), .B(n4942), .Z(n4493) );
  XNOR U5048 ( .A(n4940), .B(n4954), .Z(n4942) );
  ANDN U5049 ( .A(X[0]), .B(n1702), .Z(n4954) );
  XNOR U5050 ( .A(n4938), .B(A[18]), .Z(n4939) );
  ANDN U5051 ( .A(n4955), .B(n4956), .Z(n4938) );
  XOR U5052 ( .A(n4957), .B(n4958), .Z(n4940) );
  AND U5053 ( .A(n4959), .B(n4960), .Z(n4958) );
  XNOR U5054 ( .A(n4961), .B(n4957), .Z(n4960) );
  XOR U5055 ( .A(n4962), .B(n4944), .Z(n4953) );
  AND U5056 ( .A(n4734), .B(n1700), .Z(n4944) );
  IV U5057 ( .A(n1793), .Z(n1700) );
  IV U5058 ( .A(n4946), .Z(n4962) );
  XNOR U5059 ( .A(n4950), .B(n4952), .Z(n4513) );
  NAND U5060 ( .A(n3322), .B(n1984), .Z(n4952) );
  XNOR U5061 ( .A(n4948), .B(n4964), .Z(n4950) );
  ANDN U5062 ( .A(n3327), .B(n1986), .Z(n4964) );
  XOR U5063 ( .A(n4965), .B(n4966), .Z(n4948) );
  AND U5064 ( .A(n4967), .B(n4968), .Z(n4966) );
  XOR U5065 ( .A(n4969), .B(n4965), .Z(n4968) );
  XNOR U5066 ( .A(n4970), .B(n4959), .Z(n4514) );
  XNOR U5067 ( .A(n4957), .B(n4971), .Z(n4959) );
  ANDN U5068 ( .A(X[0]), .B(n1793), .Z(n4971) );
  ANDN U5069 ( .A(n4972), .B(n4973), .Z(n4955) );
  XOR U5070 ( .A(n4974), .B(n4975), .Z(n4957) );
  AND U5071 ( .A(n4976), .B(n4977), .Z(n4975) );
  XNOR U5072 ( .A(n4978), .B(n4974), .Z(n4977) );
  XOR U5073 ( .A(n4979), .B(n4961), .Z(n4970) );
  AND U5074 ( .A(n4734), .B(n1791), .Z(n4961) );
  IV U5075 ( .A(n1890), .Z(n1791) );
  IV U5076 ( .A(n4963), .Z(n4979) );
  XNOR U5077 ( .A(n4967), .B(n4969), .Z(n4534) );
  NAND U5078 ( .A(n3322), .B(n2080), .Z(n4969) );
  XNOR U5079 ( .A(n4965), .B(n4981), .Z(n4967) );
  ANDN U5080 ( .A(n3327), .B(n2082), .Z(n4981) );
  XNOR U5081 ( .A(n4985), .B(n4976), .Z(n4535) );
  XNOR U5082 ( .A(n4974), .B(n4986), .Z(n4976) );
  ANDN U5083 ( .A(X[0]), .B(n1890), .Z(n4986) );
  AND U5084 ( .A(n4734), .B(n1888), .Z(n4978) );
  XNOR U5085 ( .A(n4983), .B(n4984), .Z(n4552) );
  NAND U5086 ( .A(n3322), .B(n2181), .Z(n4984) );
  XNOR U5087 ( .A(n4982), .B(n4991), .Z(n4983) );
  ANDN U5088 ( .A(n3327), .B(n2183), .Z(n4991) );
  XNOR U5089 ( .A(n4995), .B(n4988), .Z(n4554) );
  XNOR U5090 ( .A(n4987), .B(n4996), .Z(n4988) );
  ANDN U5091 ( .A(X[0]), .B(n1986), .Z(n4996) );
  AND U5092 ( .A(n4734), .B(n1984), .Z(n4989) );
  XNOR U5093 ( .A(n4993), .B(n4994), .Z(n4572) );
  NAND U5094 ( .A(n3322), .B(n2287), .Z(n4994) );
  XNOR U5095 ( .A(n4992), .B(n5001), .Z(n4993) );
  ANDN U5096 ( .A(n3327), .B(n2289), .Z(n5001) );
  XNOR U5097 ( .A(n5005), .B(n4998), .Z(n4574) );
  XNOR U5098 ( .A(n4997), .B(n5006), .Z(n4998) );
  ANDN U5099 ( .A(X[0]), .B(n2082), .Z(n5006) );
  AND U5100 ( .A(n4734), .B(n2080), .Z(n4999) );
  XNOR U5101 ( .A(n5003), .B(n5004), .Z(n4592) );
  NAND U5102 ( .A(n3322), .B(n2394), .Z(n5004) );
  XNOR U5103 ( .A(n5002), .B(n5011), .Z(n5003) );
  ANDN U5104 ( .A(n3327), .B(n2396), .Z(n5011) );
  XNOR U5105 ( .A(n5015), .B(n5008), .Z(n4594) );
  XNOR U5106 ( .A(n5007), .B(n5016), .Z(n5008) );
  ANDN U5107 ( .A(X[0]), .B(n2183), .Z(n5016) );
  XOR U5108 ( .A(n5017), .B(n5018), .Z(n5007) );
  AND U5109 ( .A(n5019), .B(n5020), .Z(n5018) );
  XNOR U5110 ( .A(n5021), .B(n5017), .Z(n5020) );
  AND U5111 ( .A(n4734), .B(n2181), .Z(n5009) );
  XNOR U5112 ( .A(n5013), .B(n5014), .Z(n4612) );
  NAND U5113 ( .A(n3322), .B(n2502), .Z(n5014) );
  XNOR U5114 ( .A(n5012), .B(n5023), .Z(n5013) );
  ANDN U5115 ( .A(n3327), .B(n2504), .Z(n5023) );
  XOR U5116 ( .A(n5024), .B(n5025), .Z(n5012) );
  AND U5117 ( .A(n5026), .B(n5027), .Z(n5025) );
  XOR U5118 ( .A(n5028), .B(n5024), .Z(n5027) );
  XNOR U5119 ( .A(n5029), .B(n5019), .Z(n4614) );
  XNOR U5120 ( .A(n5017), .B(n5030), .Z(n5019) );
  ANDN U5121 ( .A(X[0]), .B(n2289), .Z(n5030) );
  XOR U5122 ( .A(n5031), .B(n5032), .Z(n5017) );
  AND U5123 ( .A(n5033), .B(n5034), .Z(n5032) );
  XNOR U5124 ( .A(n5035), .B(n5031), .Z(n5034) );
  XOR U5125 ( .A(n5036), .B(n5021), .Z(n5029) );
  AND U5126 ( .A(n4734), .B(n2287), .Z(n5021) );
  IV U5127 ( .A(n5022), .Z(n5036) );
  XNOR U5128 ( .A(n5026), .B(n5028), .Z(n4632) );
  NAND U5129 ( .A(n3322), .B(n2621), .Z(n5028) );
  XNOR U5130 ( .A(n5024), .B(n5038), .Z(n5026) );
  ANDN U5131 ( .A(n3327), .B(n2623), .Z(n5038) );
  XOR U5132 ( .A(n5039), .B(n5040), .Z(n5024) );
  AND U5133 ( .A(n5041), .B(n5042), .Z(n5040) );
  XOR U5134 ( .A(n5043), .B(n5039), .Z(n5042) );
  XNOR U5135 ( .A(n5044), .B(n5033), .Z(n4634) );
  XNOR U5136 ( .A(n5031), .B(n5045), .Z(n5033) );
  ANDN U5137 ( .A(X[0]), .B(n2396), .Z(n5045) );
  XOR U5138 ( .A(n5046), .B(n5047), .Z(n5031) );
  AND U5139 ( .A(n5048), .B(n5049), .Z(n5047) );
  XNOR U5140 ( .A(n5050), .B(n5046), .Z(n5049) );
  XOR U5141 ( .A(n5051), .B(n5035), .Z(n5044) );
  AND U5142 ( .A(n4734), .B(n2394), .Z(n5035) );
  IV U5143 ( .A(n5037), .Z(n5051) );
  XNOR U5144 ( .A(n5041), .B(n5043), .Z(n4652) );
  NAND U5145 ( .A(n3322), .B(n2741), .Z(n5043) );
  XNOR U5146 ( .A(n5039), .B(n5053), .Z(n5041) );
  ANDN U5147 ( .A(n3327), .B(n2743), .Z(n5053) );
  XNOR U5148 ( .A(n5057), .B(n5048), .Z(n4654) );
  XNOR U5149 ( .A(n5046), .B(n5058), .Z(n5048) );
  ANDN U5150 ( .A(X[0]), .B(n2504), .Z(n5058) );
  XOR U5151 ( .A(n5059), .B(n5060), .Z(n5046) );
  AND U5152 ( .A(n5061), .B(n5062), .Z(n5060) );
  XNOR U5153 ( .A(n5063), .B(n5059), .Z(n5062) );
  AND U5154 ( .A(n4734), .B(n2502), .Z(n5050) );
  XNOR U5155 ( .A(n5055), .B(n5056), .Z(n4676) );
  NAND U5156 ( .A(n3322), .B(n2863), .Z(n5056) );
  XNOR U5157 ( .A(n5054), .B(n5065), .Z(n5055) );
  ANDN U5158 ( .A(n3327), .B(n2865), .Z(n5065) );
  XNOR U5159 ( .A(n5069), .B(n5061), .Z(n4678) );
  XNOR U5160 ( .A(n5059), .B(n5070), .Z(n5061) );
  ANDN U5161 ( .A(X[0]), .B(n2623), .Z(n5070) );
  XOR U5162 ( .A(n5071), .B(n5072), .Z(n5059) );
  AND U5163 ( .A(n5073), .B(n5074), .Z(n5072) );
  XNOR U5164 ( .A(n5075), .B(n5071), .Z(n5074) );
  AND U5165 ( .A(n4734), .B(n2621), .Z(n5063) );
  XNOR U5166 ( .A(n5067), .B(n5068), .Z(n4696) );
  NAND U5167 ( .A(n3322), .B(n2988), .Z(n5068) );
  XNOR U5168 ( .A(n5066), .B(n5077), .Z(n5067) );
  ANDN U5169 ( .A(n3327), .B(n2990), .Z(n5077) );
  XNOR U5170 ( .A(n5081), .B(n5073), .Z(n4697) );
  XNOR U5171 ( .A(n5071), .B(n5082), .Z(n5073) );
  ANDN U5172 ( .A(X[0]), .B(n2743), .Z(n5082) );
  AND U5173 ( .A(n4734), .B(n2741), .Z(n5075) );
  XNOR U5174 ( .A(n5086), .B(n5087), .Z(n5076) );
  AND U5175 ( .A(n5088), .B(n5089), .Z(n5087) );
  XNOR U5176 ( .A(n5084), .B(n5090), .Z(n5089) );
  XNOR U5177 ( .A(n5085), .B(n5086), .Z(n5090) );
  AND U5178 ( .A(n4734), .B(n2863), .Z(n5085) );
  XOR U5179 ( .A(n5083), .B(n5091), .Z(n5084) );
  ANDN U5180 ( .A(X[0]), .B(n2865), .Z(n5091) );
  XNOR U5181 ( .A(n5079), .B(n5095), .Z(n5088) );
  XNOR U5182 ( .A(n5080), .B(n5086), .Z(n5095) );
  AND U5183 ( .A(n3120), .B(n3322), .Z(n5080) );
  XOR U5184 ( .A(n5078), .B(n5096), .Z(n5079) );
  ANDN U5185 ( .A(n3327), .B(n3122), .Z(n5096) );
  XOR U5186 ( .A(n5100), .B(n5101), .Z(n5086) );
  AND U5187 ( .A(n5102), .B(n5103), .Z(n5101) );
  XNOR U5188 ( .A(n5093), .B(n5104), .Z(n5103) );
  XNOR U5189 ( .A(n5094), .B(n5100), .Z(n5104) );
  AND U5190 ( .A(n4734), .B(n2988), .Z(n5094) );
  XOR U5191 ( .A(n5092), .B(n5105), .Z(n5093) );
  ANDN U5192 ( .A(X[0]), .B(n2990), .Z(n5105) );
  XNOR U5193 ( .A(n5098), .B(n5109), .Z(n5102) );
  XNOR U5194 ( .A(n5099), .B(n5100), .Z(n5109) );
  AND U5195 ( .A(n3252), .B(n3322), .Z(n5099) );
  XOR U5196 ( .A(n5097), .B(n5110), .Z(n5098) );
  ANDN U5197 ( .A(n3327), .B(n3254), .Z(n5110) );
  XOR U5198 ( .A(n5111), .B(n5112), .Z(n5097) );
  ANDN U5199 ( .A(n5113), .B(n5114), .Z(n5112) );
  XNOR U5200 ( .A(n5115), .B(n5111), .Z(n5113) );
  XOR U5201 ( .A(n5116), .B(n5117), .Z(n5100) );
  AND U5202 ( .A(n5118), .B(n5119), .Z(n5117) );
  XNOR U5203 ( .A(n5107), .B(n5120), .Z(n5119) );
  XNOR U5204 ( .A(n5108), .B(n5116), .Z(n5120) );
  AND U5205 ( .A(n4734), .B(n3120), .Z(n5108) );
  XOR U5206 ( .A(n5106), .B(n5121), .Z(n5107) );
  ANDN U5207 ( .A(X[0]), .B(n3122), .Z(n5121) );
  XNOR U5208 ( .A(n5114), .B(n5125), .Z(n5118) );
  XNOR U5209 ( .A(n5115), .B(n5116), .Z(n5125) );
  AND U5210 ( .A(n3391), .B(n3322), .Z(n5115) );
  XOR U5211 ( .A(n5111), .B(n5126), .Z(n5114) );
  ANDN U5212 ( .A(n3327), .B(n3393), .Z(n5126) );
  XNOR U5213 ( .A(n5131), .B(n5123), .Z(n4717) );
  XNOR U5214 ( .A(n5122), .B(n5132), .Z(n5123) );
  ANDN U5215 ( .A(X[0]), .B(n3254), .Z(n5132) );
  XNOR U5216 ( .A(n5135), .B(n5133), .Z(n5134) );
  ANDN U5217 ( .A(X[0]), .B(n3393), .Z(n5135) );
  ANDN U5218 ( .A(n4734), .B(n4181), .Z(n5136) );
  XNOR U5219 ( .A(n5130), .B(n5124), .Z(n5131) );
  AND U5220 ( .A(n4734), .B(n3252), .Z(n5124) );
  XNOR U5221 ( .A(n5128), .B(n5129), .Z(n4716) );
  NAND U5222 ( .A(n4179), .B(n3322), .Z(n5129) );
  XNOR U5223 ( .A(n5127), .B(n5140), .Z(n5128) );
  ANDN U5224 ( .A(n3327), .B(n4181), .Z(n5140) );
  NAND U5225 ( .A(A[0]), .B(n5141), .Z(n5127) );
  NANDN U5226 ( .B(n3322), .A(n5142), .Z(n5141) );
  NANDN U5227 ( .B(n4184), .A(n3327), .Z(n5142) );
  IV U5228 ( .A(n3190), .Z(n3322) );
  XNOR U5229 ( .A(n5138), .B(n5139), .Z(n5130) );
  NAND U5230 ( .A(n4179), .B(n4734), .Z(n5139) );
  XNOR U5231 ( .A(n5137), .B(n5145), .Z(n5138) );
  ANDN U5232 ( .A(X[0]), .B(n4181), .Z(n5145) );
  NAND U5233 ( .A(A[0]), .B(n5146), .Z(n5137) );
  NANDN U5234 ( .B(n4734), .A(n5147), .Z(n5146) );
  NANDN U5235 ( .B(n4184), .A(X[0]), .Z(n5147) );
  IV U5236 ( .A(n4721), .Z(n4734) );
  XNOR U5237 ( .A(n3350), .B(n3349), .Z(n3303) );
  XOR U5238 ( .A(n5149), .B(n3358), .Z(n3349) );
  XNOR U5239 ( .A(n3343), .B(n3342), .Z(n3358) );
  XOR U5240 ( .A(n5150), .B(n3339), .Z(n3342) );
  XNOR U5241 ( .A(n3338), .B(n5151), .Z(n3339) );
  ANDN U5242 ( .A(n1404), .B(n2289), .Z(n5151) );
  AND U5243 ( .A(n2287), .B(n1341), .Z(n3340) );
  XNOR U5244 ( .A(n3346), .B(n3347), .Z(n3343) );
  NANDN U5245 ( .B(n1206), .A(n2502), .Z(n3347) );
  XNOR U5246 ( .A(n3345), .B(n5158), .Z(n3346) );
  ANDN U5247 ( .A(n1276), .B(n2504), .Z(n5158) );
  XOR U5248 ( .A(n3357), .B(n3348), .Z(n5149) );
  XNOR U5249 ( .A(n5162), .B(n5163), .Z(n3348) );
  XOR U5250 ( .A(n5164), .B(n3366), .Z(n3357) );
  XNOR U5251 ( .A(n3354), .B(n3355), .Z(n3366) );
  NAND U5252 ( .A(n2080), .B(n1575), .Z(n3355) );
  XNOR U5253 ( .A(n3353), .B(n5165), .Z(n3354) );
  ANDN U5254 ( .A(n1582), .B(n2082), .Z(n5165) );
  XNOR U5255 ( .A(n3365), .B(n3356), .Z(n5164) );
  XOR U5256 ( .A(n5169), .B(n5170), .Z(n3356) );
  AND U5257 ( .A(n5171), .B(n5172), .Z(n5170) );
  XOR U5258 ( .A(n5173), .B(n5174), .Z(n5172) );
  XNOR U5259 ( .A(n5169), .B(n5175), .Z(n5174) );
  XNOR U5260 ( .A(n5156), .B(n5176), .Z(n5171) );
  XNOR U5261 ( .A(n5169), .B(n5157), .Z(n5176) );
  XNOR U5262 ( .A(n5160), .B(n5161), .Z(n5157) );
  NANDN U5263 ( .B(n1206), .A(n2621), .Z(n5161) );
  XNOR U5264 ( .A(n5159), .B(n5177), .Z(n5160) );
  ANDN U5265 ( .A(n1276), .B(n2623), .Z(n5177) );
  XOR U5266 ( .A(n5181), .B(n5153), .Z(n5156) );
  XNOR U5267 ( .A(n5152), .B(n5182), .Z(n5153) );
  ANDN U5268 ( .A(n1404), .B(n2396), .Z(n5182) );
  AND U5269 ( .A(n2394), .B(n1341), .Z(n5154) );
  XOR U5270 ( .A(n5189), .B(n5190), .Z(n5169) );
  AND U5271 ( .A(n5191), .B(n5192), .Z(n5190) );
  XOR U5272 ( .A(n5193), .B(n5194), .Z(n5192) );
  XNOR U5273 ( .A(n5189), .B(n5195), .Z(n5194) );
  XNOR U5274 ( .A(n5187), .B(n5196), .Z(n5191) );
  XNOR U5275 ( .A(n5189), .B(n5188), .Z(n5196) );
  XNOR U5276 ( .A(n5179), .B(n5180), .Z(n5188) );
  NANDN U5277 ( .B(n1206), .A(n2741), .Z(n5180) );
  XNOR U5278 ( .A(n5178), .B(n5197), .Z(n5179) );
  ANDN U5279 ( .A(n1276), .B(n2743), .Z(n5197) );
  XOR U5280 ( .A(n5201), .B(n5184), .Z(n5187) );
  XNOR U5281 ( .A(n5183), .B(n5202), .Z(n5184) );
  ANDN U5282 ( .A(n1404), .B(n2504), .Z(n5202) );
  AND U5283 ( .A(n2502), .B(n1341), .Z(n5185) );
  XOR U5284 ( .A(n5209), .B(n5210), .Z(n5189) );
  AND U5285 ( .A(n5211), .B(n5212), .Z(n5210) );
  XOR U5286 ( .A(n5213), .B(n5214), .Z(n5212) );
  XNOR U5287 ( .A(n5209), .B(n5215), .Z(n5214) );
  XNOR U5288 ( .A(n5207), .B(n5216), .Z(n5211) );
  XNOR U5289 ( .A(n5209), .B(n5208), .Z(n5216) );
  XNOR U5290 ( .A(n5199), .B(n5200), .Z(n5208) );
  NANDN U5291 ( .B(n1206), .A(n2863), .Z(n5200) );
  XNOR U5292 ( .A(n5198), .B(n5217), .Z(n5199) );
  ANDN U5293 ( .A(n1276), .B(n2865), .Z(n5217) );
  XOR U5294 ( .A(n5221), .B(n5204), .Z(n5207) );
  XNOR U5295 ( .A(n5203), .B(n5222), .Z(n5204) );
  ANDN U5296 ( .A(n1404), .B(n2623), .Z(n5222) );
  AND U5297 ( .A(n2621), .B(n1341), .Z(n5205) );
  XOR U5298 ( .A(n5229), .B(n5230), .Z(n5209) );
  AND U5299 ( .A(n5231), .B(n5232), .Z(n5230) );
  XOR U5300 ( .A(n5233), .B(n5234), .Z(n5232) );
  XNOR U5301 ( .A(n5229), .B(n5235), .Z(n5234) );
  XNOR U5302 ( .A(n5227), .B(n5236), .Z(n5231) );
  XNOR U5303 ( .A(n5229), .B(n5228), .Z(n5236) );
  XNOR U5304 ( .A(n5219), .B(n5220), .Z(n5228) );
  NANDN U5305 ( .B(n1206), .A(n2988), .Z(n5220) );
  XNOR U5306 ( .A(n5218), .B(n5237), .Z(n5219) );
  ANDN U5307 ( .A(n1276), .B(n2990), .Z(n5237) );
  XOR U5308 ( .A(n5241), .B(n5224), .Z(n5227) );
  XNOR U5309 ( .A(n5223), .B(n5242), .Z(n5224) );
  ANDN U5310 ( .A(n1404), .B(n2743), .Z(n5242) );
  AND U5311 ( .A(n2741), .B(n1341), .Z(n5225) );
  XOR U5312 ( .A(n5249), .B(n5250), .Z(n5229) );
  AND U5313 ( .A(n5251), .B(n5252), .Z(n5250) );
  XOR U5314 ( .A(n5253), .B(n5254), .Z(n5252) );
  XNOR U5315 ( .A(n5249), .B(n5255), .Z(n5254) );
  XNOR U5316 ( .A(n5247), .B(n5256), .Z(n5251) );
  XNOR U5317 ( .A(n5249), .B(n5248), .Z(n5256) );
  XNOR U5318 ( .A(n5239), .B(n5240), .Z(n5248) );
  NANDN U5319 ( .B(n1206), .A(n3120), .Z(n5240) );
  XNOR U5320 ( .A(n5238), .B(n5257), .Z(n5239) );
  ANDN U5321 ( .A(n1276), .B(n3122), .Z(n5257) );
  XOR U5322 ( .A(n5261), .B(n5244), .Z(n5247) );
  XNOR U5323 ( .A(n5243), .B(n5262), .Z(n5244) );
  ANDN U5324 ( .A(n1404), .B(n2865), .Z(n5262) );
  XOR U5325 ( .A(n5263), .B(n5264), .Z(n5243) );
  AND U5326 ( .A(n5265), .B(n5266), .Z(n5264) );
  XNOR U5327 ( .A(n5267), .B(n5263), .Z(n5266) );
  AND U5328 ( .A(n2863), .B(n1341), .Z(n5245) );
  XOR U5329 ( .A(n5271), .B(n5272), .Z(n5249) );
  AND U5330 ( .A(n5273), .B(n5274), .Z(n5272) );
  XOR U5331 ( .A(n5275), .B(n5276), .Z(n5274) );
  XNOR U5332 ( .A(n5271), .B(n5277), .Z(n5276) );
  XNOR U5333 ( .A(n5269), .B(n5278), .Z(n5273) );
  XNOR U5334 ( .A(n5271), .B(n5270), .Z(n5278) );
  XNOR U5335 ( .A(n5259), .B(n5260), .Z(n5270) );
  NANDN U5336 ( .B(n1206), .A(n3252), .Z(n5260) );
  XNOR U5337 ( .A(n5258), .B(n5279), .Z(n5259) );
  ANDN U5338 ( .A(n1276), .B(n3254), .Z(n5279) );
  XOR U5339 ( .A(n5280), .B(n5281), .Z(n5258) );
  AND U5340 ( .A(n5282), .B(n5283), .Z(n5281) );
  XOR U5341 ( .A(n5284), .B(n5280), .Z(n5283) );
  XOR U5342 ( .A(n5285), .B(n5265), .Z(n5269) );
  XNOR U5343 ( .A(n5263), .B(n5286), .Z(n5265) );
  ANDN U5344 ( .A(n1404), .B(n2990), .Z(n5286) );
  XOR U5345 ( .A(n5287), .B(n5288), .Z(n5263) );
  AND U5346 ( .A(n5289), .B(n5290), .Z(n5288) );
  XNOR U5347 ( .A(n5291), .B(n5287), .Z(n5290) );
  AND U5348 ( .A(n2988), .B(n1341), .Z(n5267) );
  XOR U5349 ( .A(n5295), .B(n5296), .Z(n5271) );
  AND U5350 ( .A(n5297), .B(n5298), .Z(n5296) );
  XOR U5351 ( .A(n5299), .B(n5300), .Z(n5298) );
  XNOR U5352 ( .A(n5295), .B(n5301), .Z(n5300) );
  XNOR U5353 ( .A(n5293), .B(n5302), .Z(n5297) );
  XNOR U5354 ( .A(n5295), .B(n5294), .Z(n5302) );
  XNOR U5355 ( .A(n5282), .B(n5284), .Z(n5294) );
  NANDN U5356 ( .B(n1206), .A(n3391), .Z(n5284) );
  XNOR U5357 ( .A(n5280), .B(n5303), .Z(n5282) );
  ANDN U5358 ( .A(n1276), .B(n3393), .Z(n5303) );
  XOR U5359 ( .A(n5307), .B(n5289), .Z(n5293) );
  XNOR U5360 ( .A(n5287), .B(n5308), .Z(n5289) );
  ANDN U5361 ( .A(n1404), .B(n3122), .Z(n5308) );
  AND U5362 ( .A(n3120), .B(n1341), .Z(n5291) );
  XOR U5363 ( .A(n5316), .B(n5317), .Z(n5163) );
  XNOR U5364 ( .A(n5314), .B(n5313), .Z(n5162) );
  XOR U5365 ( .A(n5319), .B(n5310), .Z(n5313) );
  XNOR U5366 ( .A(n5309), .B(n5320), .Z(n5310) );
  ANDN U5367 ( .A(n1404), .B(n3254), .Z(n5320) );
  XNOR U5368 ( .A(n5323), .B(n5321), .Z(n5322) );
  ANDN U5369 ( .A(n1404), .B(n3393), .Z(n5323) );
  XNOR U5370 ( .A(n5312), .B(n5311), .Z(n5319) );
  AND U5371 ( .A(n3252), .B(n1341), .Z(n5311) );
  XNOR U5372 ( .A(n5326), .B(n5327), .Z(n5312) );
  NAND U5373 ( .A(n4179), .B(n1341), .Z(n5327) );
  XNOR U5374 ( .A(n5325), .B(n5328), .Z(n5326) );
  ANDN U5375 ( .A(n1404), .B(n4181), .Z(n5328) );
  NAND U5376 ( .A(A[0]), .B(n5329), .Z(n5325) );
  NANDN U5377 ( .B(n1341), .A(n5330), .Z(n5329) );
  NANDN U5378 ( .B(n4184), .A(n1404), .Z(n5330) );
  IV U5379 ( .A(n5324), .Z(n1341) );
  XNOR U5380 ( .A(n5305), .B(n5306), .Z(n5314) );
  NANDN U5381 ( .B(n1206), .A(n4179), .Z(n5306) );
  XNOR U5382 ( .A(n5304), .B(n5333), .Z(n5305) );
  ANDN U5383 ( .A(n1276), .B(n4181), .Z(n5333) );
  NAND U5384 ( .A(A[0]), .B(n5334), .Z(n5304) );
  NAND U5385 ( .A(n5335), .B(n1206), .Z(n5334) );
  NANDN U5386 ( .B(n4184), .A(n1276), .Z(n5335) );
  XOR U5387 ( .A(n5338), .B(n5339), .Z(n5315) );
  XOR U5388 ( .A(n5340), .B(n3362), .Z(n3365) );
  XNOR U5389 ( .A(n3361), .B(n5341), .Z(n3362) );
  ANDN U5390 ( .A(n1766), .B(n1890), .Z(n5341) );
  XNOR U5391 ( .A(n4972), .B(A[16]), .Z(n4973) );
  ANDN U5392 ( .A(n5342), .B(n5343), .Z(n4972) );
  AND U5393 ( .A(n1888), .B(n1759), .Z(n3363) );
  IV U5394 ( .A(n1986), .Z(n1888) );
  XNOR U5395 ( .A(n5167), .B(n5168), .Z(n5173) );
  NAND U5396 ( .A(n2181), .B(n1575), .Z(n5168) );
  XNOR U5397 ( .A(n5166), .B(n5348), .Z(n5167) );
  ANDN U5398 ( .A(n1582), .B(n2183), .Z(n5348) );
  XNOR U5399 ( .A(n5352), .B(n5345), .Z(n5175) );
  XNOR U5400 ( .A(n5344), .B(n5353), .Z(n5345) );
  ANDN U5401 ( .A(n1766), .B(n1986), .Z(n5353) );
  ANDN U5402 ( .A(n5354), .B(n5355), .Z(n5342) );
  AND U5403 ( .A(n1984), .B(n1759), .Z(n5346) );
  IV U5404 ( .A(n2082), .Z(n1984) );
  XNOR U5405 ( .A(n5350), .B(n5351), .Z(n5193) );
  NAND U5406 ( .A(n2287), .B(n1575), .Z(n5351) );
  XNOR U5407 ( .A(n5349), .B(n5360), .Z(n5350) );
  ANDN U5408 ( .A(n1582), .B(n2289), .Z(n5360) );
  XNOR U5409 ( .A(n5364), .B(n5357), .Z(n5195) );
  XNOR U5410 ( .A(n5356), .B(n5365), .Z(n5357) );
  ANDN U5411 ( .A(n1766), .B(n2082), .Z(n5365) );
  XNOR U5412 ( .A(n5354), .B(A[14]), .Z(n5355) );
  ANDN U5413 ( .A(n5366), .B(n5367), .Z(n5354) );
  AND U5414 ( .A(n2080), .B(n1759), .Z(n5358) );
  IV U5415 ( .A(n2183), .Z(n2080) );
  XNOR U5416 ( .A(n5362), .B(n5363), .Z(n5213) );
  NAND U5417 ( .A(n2394), .B(n1575), .Z(n5363) );
  XNOR U5418 ( .A(n5361), .B(n5372), .Z(n5362) );
  ANDN U5419 ( .A(n1582), .B(n2396), .Z(n5372) );
  XNOR U5420 ( .A(n5376), .B(n5369), .Z(n5215) );
  XNOR U5421 ( .A(n5368), .B(n5377), .Z(n5369) );
  ANDN U5422 ( .A(n1766), .B(n2183), .Z(n5377) );
  ANDN U5423 ( .A(n5378), .B(n5379), .Z(n5366) );
  AND U5424 ( .A(n2181), .B(n1759), .Z(n5370) );
  IV U5425 ( .A(n2289), .Z(n2181) );
  XNOR U5426 ( .A(n5374), .B(n5375), .Z(n5233) );
  NAND U5427 ( .A(n2502), .B(n1575), .Z(n5375) );
  XNOR U5428 ( .A(n5373), .B(n5384), .Z(n5374) );
  ANDN U5429 ( .A(n1582), .B(n2504), .Z(n5384) );
  XNOR U5430 ( .A(n5388), .B(n5381), .Z(n5235) );
  XNOR U5431 ( .A(n5380), .B(n5389), .Z(n5381) );
  ANDN U5432 ( .A(n1766), .B(n2289), .Z(n5389) );
  XNOR U5433 ( .A(n5378), .B(A[12]), .Z(n5379) );
  ANDN U5434 ( .A(n5390), .B(n5391), .Z(n5378) );
  AND U5435 ( .A(n2287), .B(n1759), .Z(n5382) );
  IV U5436 ( .A(n2396), .Z(n2287) );
  XNOR U5437 ( .A(n5386), .B(n5387), .Z(n5253) );
  NAND U5438 ( .A(n2621), .B(n1575), .Z(n5387) );
  XNOR U5439 ( .A(n5385), .B(n5396), .Z(n5386) );
  ANDN U5440 ( .A(n1582), .B(n2623), .Z(n5396) );
  XOR U5441 ( .A(n5397), .B(n5398), .Z(n5385) );
  AND U5442 ( .A(n5399), .B(n5400), .Z(n5398) );
  XOR U5443 ( .A(n5401), .B(n5397), .Z(n5400) );
  XNOR U5444 ( .A(n5402), .B(n5393), .Z(n5255) );
  XNOR U5445 ( .A(n5392), .B(n5403), .Z(n5393) );
  ANDN U5446 ( .A(n1766), .B(n2396), .Z(n5403) );
  ANDN U5447 ( .A(n5404), .B(n5405), .Z(n5390) );
  AND U5448 ( .A(n2394), .B(n1759), .Z(n5394) );
  IV U5449 ( .A(n2504), .Z(n2394) );
  XNOR U5450 ( .A(n5399), .B(n5401), .Z(n5275) );
  NAND U5451 ( .A(n2741), .B(n1575), .Z(n5401) );
  XNOR U5452 ( .A(n5397), .B(n5410), .Z(n5399) );
  ANDN U5453 ( .A(n1582), .B(n2743), .Z(n5410) );
  XOR U5454 ( .A(n5411), .B(n5412), .Z(n5397) );
  AND U5455 ( .A(n5413), .B(n5414), .Z(n5412) );
  XOR U5456 ( .A(n5415), .B(n5411), .Z(n5414) );
  XNOR U5457 ( .A(n5416), .B(n5407), .Z(n5277) );
  XNOR U5458 ( .A(n5406), .B(n5417), .Z(n5407) );
  ANDN U5459 ( .A(n1766), .B(n2504), .Z(n5417) );
  XNOR U5460 ( .A(n5404), .B(A[10]), .Z(n5405) );
  ANDN U5461 ( .A(n5418), .B(n5419), .Z(n5404) );
  XOR U5462 ( .A(n5420), .B(n5421), .Z(n5406) );
  AND U5463 ( .A(n5422), .B(n5423), .Z(n5421) );
  XNOR U5464 ( .A(n5424), .B(n5420), .Z(n5423) );
  XOR U5465 ( .A(n5425), .B(n5408), .Z(n5416) );
  AND U5466 ( .A(n2502), .B(n1759), .Z(n5408) );
  IV U5467 ( .A(n2623), .Z(n2502) );
  IV U5468 ( .A(n5409), .Z(n5425) );
  XNOR U5469 ( .A(n5413), .B(n5415), .Z(n5299) );
  NAND U5470 ( .A(n2863), .B(n1575), .Z(n5415) );
  XNOR U5471 ( .A(n5411), .B(n5427), .Z(n5413) );
  ANDN U5472 ( .A(n1582), .B(n2865), .Z(n5427) );
  XNOR U5473 ( .A(n5431), .B(n5422), .Z(n5301) );
  XNOR U5474 ( .A(n5420), .B(n5432), .Z(n5422) );
  ANDN U5475 ( .A(n1766), .B(n2623), .Z(n5432) );
  ANDN U5476 ( .A(n5433), .B(n5434), .Z(n5418) );
  XOR U5477 ( .A(n5435), .B(n5436), .Z(n5420) );
  AND U5478 ( .A(n5437), .B(n5438), .Z(n5436) );
  XNOR U5479 ( .A(n5439), .B(n5435), .Z(n5438) );
  AND U5480 ( .A(n2621), .B(n1759), .Z(n5424) );
  IV U5481 ( .A(n2743), .Z(n2621) );
  XNOR U5482 ( .A(n5429), .B(n5430), .Z(n5317) );
  NAND U5483 ( .A(n2988), .B(n1575), .Z(n5430) );
  XNOR U5484 ( .A(n5428), .B(n5441), .Z(n5429) );
  ANDN U5485 ( .A(n1582), .B(n2990), .Z(n5441) );
  XNOR U5486 ( .A(n5445), .B(n5437), .Z(n5318) );
  XNOR U5487 ( .A(n5435), .B(n5446), .Z(n5437) );
  ANDN U5488 ( .A(n1766), .B(n2743), .Z(n5446) );
  AND U5489 ( .A(n2741), .B(n1759), .Z(n5439) );
  XNOR U5490 ( .A(n5450), .B(n5451), .Z(n5440) );
  AND U5491 ( .A(n5452), .B(n5453), .Z(n5451) );
  XNOR U5492 ( .A(n5448), .B(n5454), .Z(n5453) );
  XNOR U5493 ( .A(n5449), .B(n5450), .Z(n5454) );
  AND U5494 ( .A(n2863), .B(n1759), .Z(n5449) );
  XOR U5495 ( .A(n5447), .B(n5455), .Z(n5448) );
  ANDN U5496 ( .A(n1766), .B(n2865), .Z(n5455) );
  XNOR U5497 ( .A(n5443), .B(n5459), .Z(n5452) );
  XNOR U5498 ( .A(n5444), .B(n5450), .Z(n5459) );
  AND U5499 ( .A(n3120), .B(n1575), .Z(n5444) );
  XOR U5500 ( .A(n5442), .B(n5460), .Z(n5443) );
  ANDN U5501 ( .A(n1582), .B(n3122), .Z(n5460) );
  XOR U5502 ( .A(n5464), .B(n5465), .Z(n5450) );
  AND U5503 ( .A(n5466), .B(n5467), .Z(n5465) );
  XNOR U5504 ( .A(n5457), .B(n5468), .Z(n5467) );
  XNOR U5505 ( .A(n5458), .B(n5464), .Z(n5468) );
  AND U5506 ( .A(n2988), .B(n1759), .Z(n5458) );
  XOR U5507 ( .A(n5456), .B(n5469), .Z(n5457) );
  ANDN U5508 ( .A(n1766), .B(n2990), .Z(n5469) );
  XNOR U5509 ( .A(n5462), .B(n5473), .Z(n5466) );
  XNOR U5510 ( .A(n5463), .B(n5464), .Z(n5473) );
  AND U5511 ( .A(n3252), .B(n1575), .Z(n5463) );
  XOR U5512 ( .A(n5461), .B(n5474), .Z(n5462) );
  ANDN U5513 ( .A(n1582), .B(n3254), .Z(n5474) );
  XOR U5514 ( .A(n5475), .B(n5476), .Z(n5461) );
  ANDN U5515 ( .A(n5477), .B(n5478), .Z(n5476) );
  XNOR U5516 ( .A(n5479), .B(n5475), .Z(n5477) );
  XOR U5517 ( .A(n5480), .B(n5481), .Z(n5464) );
  AND U5518 ( .A(n5482), .B(n5483), .Z(n5481) );
  XNOR U5519 ( .A(n5471), .B(n5484), .Z(n5483) );
  XNOR U5520 ( .A(n5472), .B(n5480), .Z(n5484) );
  AND U5521 ( .A(n3120), .B(n1759), .Z(n5472) );
  XOR U5522 ( .A(n5470), .B(n5485), .Z(n5471) );
  ANDN U5523 ( .A(n1766), .B(n3122), .Z(n5485) );
  XNOR U5524 ( .A(n5478), .B(n5489), .Z(n5482) );
  XNOR U5525 ( .A(n5479), .B(n5480), .Z(n5489) );
  AND U5526 ( .A(n3391), .B(n1575), .Z(n5479) );
  XOR U5527 ( .A(n5475), .B(n5490), .Z(n5478) );
  ANDN U5528 ( .A(n1582), .B(n3393), .Z(n5490) );
  XNOR U5529 ( .A(n5495), .B(n5487), .Z(n5339) );
  XNOR U5530 ( .A(n5486), .B(n5496), .Z(n5487) );
  ANDN U5531 ( .A(n1766), .B(n3254), .Z(n5496) );
  XNOR U5532 ( .A(n5499), .B(n5497), .Z(n5498) );
  ANDN U5533 ( .A(n1766), .B(n3393), .Z(n5499) );
  XNOR U5534 ( .A(n5494), .B(n5488), .Z(n5495) );
  AND U5535 ( .A(n3252), .B(n1759), .Z(n5488) );
  XNOR U5536 ( .A(n5492), .B(n5493), .Z(n5338) );
  NAND U5537 ( .A(n4179), .B(n1575), .Z(n5493) );
  XNOR U5538 ( .A(n5491), .B(n5503), .Z(n5492) );
  ANDN U5539 ( .A(n1582), .B(n4181), .Z(n5503) );
  NAND U5540 ( .A(A[0]), .B(n5504), .Z(n5491) );
  NANDN U5541 ( .B(n1575), .A(n5505), .Z(n5504) );
  NANDN U5542 ( .B(n4184), .A(n1582), .Z(n5505) );
  IV U5543 ( .A(n1501), .Z(n1575) );
  XNOR U5544 ( .A(n5501), .B(n5502), .Z(n5494) );
  NAND U5545 ( .A(n4179), .B(n1759), .Z(n5502) );
  XNOR U5546 ( .A(n5500), .B(n5508), .Z(n5501) );
  ANDN U5547 ( .A(n1766), .B(n4181), .Z(n5508) );
  NAND U5548 ( .A(A[0]), .B(n5509), .Z(n5500) );
  NANDN U5549 ( .B(n1759), .A(n5510), .Z(n5509) );
  NANDN U5550 ( .B(n4184), .A(n1766), .Z(n5510) );
  IV U5551 ( .A(n1666), .Z(n1759) );
  XNOR U5552 ( .A(n3374), .B(n3373), .Z(n3350) );
  XOR U5553 ( .A(n5513), .B(n3382), .Z(n3373) );
  XNOR U5554 ( .A(n3370), .B(n3371), .Z(n3382) );
  NANDN U5555 ( .B(n1019), .A(n2988), .Z(n3371) );
  XNOR U5556 ( .A(n3369), .B(n5514), .Z(n3370) );
  ANDN U5557 ( .A(n1060), .B(n2990), .Z(n5514) );
  XOR U5558 ( .A(n3381), .B(n3372), .Z(n5513) );
  XOR U5559 ( .A(n5518), .B(n5519), .Z(n3372) );
  XOR U5560 ( .A(n5520), .B(n3378), .Z(n3381) );
  XNOR U5561 ( .A(n3377), .B(n5521), .Z(n3378) );
  ANDN U5562 ( .A(n1167), .B(n2743), .Z(n5521) );
  XNOR U5563 ( .A(n5433), .B(A[8]), .Z(n5434) );
  ANDN U5564 ( .A(n5522), .B(n5523), .Z(n5433) );
  AND U5565 ( .A(n2741), .B(n1113), .Z(n3379) );
  IV U5566 ( .A(n2865), .Z(n2741) );
  XNOR U5567 ( .A(n5527), .B(n5528), .Z(n3380) );
  AND U5568 ( .A(n5529), .B(n5530), .Z(n5528) );
  XNOR U5569 ( .A(n5525), .B(n5531), .Z(n5530) );
  XNOR U5570 ( .A(n5526), .B(n5527), .Z(n5531) );
  AND U5571 ( .A(n2863), .B(n1113), .Z(n5526) );
  IV U5572 ( .A(n2990), .Z(n2863) );
  XOR U5573 ( .A(n5524), .B(n5532), .Z(n5525) );
  ANDN U5574 ( .A(n1167), .B(n2865), .Z(n5532) );
  ANDN U5575 ( .A(n5533), .B(n5534), .Z(n5522) );
  XNOR U5576 ( .A(n5516), .B(n5538), .Z(n5529) );
  XNOR U5577 ( .A(n5517), .B(n5527), .Z(n5538) );
  ANDN U5578 ( .A(n3120), .B(n1019), .Z(n5517) );
  XOR U5579 ( .A(n5515), .B(n5539), .Z(n5516) );
  ANDN U5580 ( .A(n1060), .B(n3122), .Z(n5539) );
  XOR U5581 ( .A(n5543), .B(n5544), .Z(n5527) );
  AND U5582 ( .A(n5545), .B(n5546), .Z(n5544) );
  XNOR U5583 ( .A(n5536), .B(n5547), .Z(n5546) );
  XNOR U5584 ( .A(n5537), .B(n5543), .Z(n5547) );
  AND U5585 ( .A(n2988), .B(n1113), .Z(n5537) );
  IV U5586 ( .A(n3122), .Z(n2988) );
  XOR U5587 ( .A(n5535), .B(n5548), .Z(n5536) );
  ANDN U5588 ( .A(n1167), .B(n2990), .Z(n5548) );
  XNOR U5589 ( .A(n5533), .B(A[6]), .Z(n5534) );
  ANDN U5590 ( .A(n5549), .B(n5550), .Z(n5533) );
  XNOR U5591 ( .A(n5541), .B(n5554), .Z(n5545) );
  XNOR U5592 ( .A(n5542), .B(n5543), .Z(n5554) );
  ANDN U5593 ( .A(n3252), .B(n1019), .Z(n5542) );
  XOR U5594 ( .A(n5540), .B(n5555), .Z(n5541) );
  ANDN U5595 ( .A(n1060), .B(n3254), .Z(n5555) );
  XOR U5596 ( .A(n5556), .B(n5557), .Z(n5540) );
  ANDN U5597 ( .A(n5558), .B(n5559), .Z(n5557) );
  XNOR U5598 ( .A(n5560), .B(n5556), .Z(n5558) );
  XOR U5599 ( .A(n5561), .B(n5562), .Z(n5543) );
  AND U5600 ( .A(n5563), .B(n5564), .Z(n5562) );
  XNOR U5601 ( .A(n5552), .B(n5565), .Z(n5564) );
  XNOR U5602 ( .A(n5553), .B(n5561), .Z(n5565) );
  AND U5603 ( .A(n3120), .B(n1113), .Z(n5553) );
  XOR U5604 ( .A(n5551), .B(n5566), .Z(n5552) );
  ANDN U5605 ( .A(n1167), .B(n3122), .Z(n5566) );
  ANDN U5606 ( .A(n5567), .B(n5568), .Z(n5549) );
  XNOR U5607 ( .A(n5559), .B(n5572), .Z(n5563) );
  XNOR U5608 ( .A(n5560), .B(n5561), .Z(n5572) );
  ANDN U5609 ( .A(n3391), .B(n1019), .Z(n5560) );
  XOR U5610 ( .A(n5556), .B(n5573), .Z(n5559) );
  ANDN U5611 ( .A(n1060), .B(n3393), .Z(n5573) );
  XNOR U5612 ( .A(n5578), .B(n5570), .Z(n5519) );
  XNOR U5613 ( .A(n5569), .B(n5579), .Z(n5570) );
  ANDN U5614 ( .A(n1167), .B(n3254), .Z(n5579) );
  XNOR U5615 ( .A(n5582), .B(n5580), .Z(n5581) );
  ANDN U5616 ( .A(n1167), .B(n3393), .Z(n5582) );
  XNOR U5617 ( .A(n5577), .B(n5571), .Z(n5578) );
  AND U5618 ( .A(n3252), .B(n1113), .Z(n5571) );
  XNOR U5619 ( .A(n5575), .B(n5576), .Z(n5518) );
  NANDN U5620 ( .B(n1019), .A(n4179), .Z(n5576) );
  XNOR U5621 ( .A(n5574), .B(n5587), .Z(n5575) );
  ANDN U5622 ( .A(n1060), .B(n4181), .Z(n5587) );
  NAND U5623 ( .A(A[0]), .B(n5588), .Z(n5574) );
  NAND U5624 ( .A(n5589), .B(n1019), .Z(n5588) );
  NANDN U5625 ( .B(n4184), .A(n1060), .Z(n5589) );
  XNOR U5626 ( .A(n5585), .B(n5586), .Z(n5577) );
  NAND U5627 ( .A(n4179), .B(n1113), .Z(n5586) );
  XNOR U5628 ( .A(n5584), .B(n5592), .Z(n5585) );
  ANDN U5629 ( .A(n1167), .B(n4181), .Z(n5592) );
  NAND U5630 ( .A(A[0]), .B(n5593), .Z(n5584) );
  NANDN U5631 ( .B(n1113), .A(n5594), .Z(n5593) );
  NANDN U5632 ( .B(n4184), .A(n1167), .Z(n5594) );
  IV U5633 ( .A(n5583), .Z(n1113) );
  XOR U5634 ( .A(n3390), .B(n3389), .Z(n3374) );
  XOR U5635 ( .A(n5597), .B(n3386), .Z(n3389) );
  XNOR U5636 ( .A(n3385), .B(n5598), .Z(n3386) );
  ANDN U5637 ( .A(n992), .B(n3254), .Z(n5598) );
  IV U5638 ( .A(n3120), .Z(n3254) );
  XNOR U5639 ( .A(n5567), .B(A[4]), .Z(n5568) );
  ANDN U5640 ( .A(n5599), .B(n5600), .Z(n5567) );
  XNOR U5641 ( .A(n5603), .B(n5601), .Z(n5602) );
  ANDN U5642 ( .A(n992), .B(n3393), .Z(n5603) );
  IV U5643 ( .A(n3252), .Z(n3393) );
  IV U5644 ( .A(n4181), .Z(n3391) );
  XNOR U5645 ( .A(n3388), .B(n3387), .Z(n5597) );
  AND U5646 ( .A(n3252), .B(n951), .Z(n3387) );
  ANDN U5647 ( .A(n5608), .B(n5609), .Z(n5599) );
  XNOR U5648 ( .A(n5606), .B(n5607), .Z(n3388) );
  NAND U5649 ( .A(n4179), .B(n951), .Z(n5607) );
  XNOR U5650 ( .A(n5605), .B(n5610), .Z(n5606) );
  ANDN U5651 ( .A(n992), .B(n4181), .Z(n5610) );
  NAND U5652 ( .A(A[0]), .B(n5611), .Z(n5605) );
  NANDN U5653 ( .B(n951), .A(n5612), .Z(n5611) );
  NANDN U5654 ( .B(n4184), .A(n992), .Z(n5612) );
  IV U5655 ( .A(n5604), .Z(n951) );
  XOR U5656 ( .A(n3397), .B(n3396), .Z(n3390) );
  NAND U5657 ( .A(n4179), .B(n895), .Z(n3396) );
  IV U5658 ( .A(n4184), .Z(n4179) );
  XOR U5659 ( .A(n3395), .B(n5615), .Z(n3397) );
  ANDN U5660 ( .A(n926), .B(n4181), .Z(n5615) );
  XNOR U5661 ( .A(n5608), .B(A[2]), .Z(n5609) );
  NOR U5662 ( .A(A[0]), .B(n5616), .Z(n5608) );
  NANDN U5663 ( .B(n895), .A(n5618), .Z(n5617) );
  NANDN U5664 ( .B(n4184), .A(n926), .Z(n5618) );
  XOR U5665 ( .A(A[0]), .B(A[1]), .Z(n5616) );
  AND U5666 ( .A(n5620), .B(n5619), .Z(n895) );
  ANDN U5667 ( .A(X[31]), .B(n5621), .Z(n5620) );
  NANDN U5668 ( .B(n5622), .A(n5614), .Z(n5621) );
  XNOR U5669 ( .A(n5622), .B(X[29]), .Z(n5614) );
  NAND U5670 ( .A(n5613), .B(n5623), .Z(n5622) );
  XOR U5671 ( .A(n5623), .B(X[28]), .Z(n5613) );
  ANDN U5672 ( .A(n5590), .B(n5624), .Z(n5623) );
  XNOR U5673 ( .A(n5624), .B(X[27]), .Z(n5590) );
  NAND U5674 ( .A(n5591), .B(n5625), .Z(n5624) );
  XOR U5675 ( .A(n5625), .B(X[26]), .Z(n5591) );
  ANDN U5676 ( .A(n5596), .B(n5626), .Z(n5625) );
  XNOR U5677 ( .A(n5626), .B(X[25]), .Z(n5596) );
  NAND U5678 ( .A(n5595), .B(n5627), .Z(n5626) );
  XOR U5679 ( .A(n5627), .B(X[24]), .Z(n5595) );
  ANDN U5680 ( .A(n5336), .B(n5628), .Z(n5627) );
  XNOR U5681 ( .A(n5628), .B(X[23]), .Z(n5336) );
  NAND U5682 ( .A(n5337), .B(n5629), .Z(n5628) );
  XOR U5683 ( .A(n5629), .B(X[22]), .Z(n5337) );
  ANDN U5684 ( .A(n5332), .B(n5630), .Z(n5629) );
  XNOR U5685 ( .A(n5630), .B(X[21]), .Z(n5332) );
  NAND U5686 ( .A(n5331), .B(n5631), .Z(n5630) );
  XOR U5687 ( .A(n5631), .B(X[20]), .Z(n5331) );
  ANDN U5688 ( .A(n5507), .B(n5632), .Z(n5631) );
  XNOR U5689 ( .A(n5632), .B(X[19]), .Z(n5507) );
  NAND U5690 ( .A(n5506), .B(n5633), .Z(n5632) );
  XOR U5691 ( .A(n5633), .B(X[18]), .Z(n5506) );
  ANDN U5692 ( .A(n5512), .B(n5634), .Z(n5633) );
  XNOR U5693 ( .A(n5634), .B(X[17]), .Z(n5512) );
  NAND U5694 ( .A(n5511), .B(n5635), .Z(n5634) );
  XOR U5695 ( .A(n5635), .B(X[16]), .Z(n5511) );
  ANDN U5696 ( .A(n4209), .B(n5636), .Z(n5635) );
  XNOR U5697 ( .A(n5636), .B(X[15]), .Z(n4209) );
  NAND U5698 ( .A(n4208), .B(n5637), .Z(n5636) );
  XOR U5699 ( .A(n5637), .B(X[14]), .Z(n4208) );
  ANDN U5700 ( .A(n4204), .B(n5638), .Z(n5637) );
  XNOR U5701 ( .A(n5638), .B(X[13]), .Z(n4204) );
  NAND U5702 ( .A(n4203), .B(n5639), .Z(n5638) );
  XOR U5703 ( .A(n5639), .B(X[12]), .Z(n4203) );
  ANDN U5704 ( .A(n4186), .B(n5640), .Z(n5639) );
  XNOR U5705 ( .A(n5640), .B(X[11]), .Z(n4186) );
  NAND U5706 ( .A(n4185), .B(n5641), .Z(n5640) );
  XOR U5707 ( .A(n5641), .B(X[10]), .Z(n4185) );
  ANDN U5708 ( .A(n4191), .B(n5642), .Z(n5641) );
  XNOR U5709 ( .A(n5642), .B(X[9]), .Z(n4191) );
  NAND U5710 ( .A(n4190), .B(n5643), .Z(n5642) );
  XOR U5711 ( .A(n5643), .B(X[8]), .Z(n4190) );
  ANDN U5712 ( .A(n4715), .B(n5644), .Z(n5643) );
  XNOR U5713 ( .A(n5644), .B(X[7]), .Z(n4715) );
  NAND U5714 ( .A(n4714), .B(n5645), .Z(n5644) );
  XOR U5715 ( .A(n5645), .B(X[6]), .Z(n4714) );
  ANDN U5716 ( .A(n4710), .B(n5646), .Z(n5645) );
  XNOR U5717 ( .A(n5646), .B(X[5]), .Z(n4710) );
  NAND U5718 ( .A(n4709), .B(n5647), .Z(n5646) );
  XOR U5719 ( .A(n5647), .B(X[4]), .Z(n4709) );
  ANDN U5720 ( .A(n5144), .B(n5648), .Z(n5647) );
  XNOR U5721 ( .A(n5648), .B(X[3]), .Z(n5144) );
  NAND U5722 ( .A(n5143), .B(n5649), .Z(n5648) );
  XOR U5723 ( .A(n5649), .B(X[2]), .Z(n5143) );
  NOR U5724 ( .A(n5148), .B(X[0]), .Z(n5649) );
  XOR U5725 ( .A(X[0]), .B(X[1]), .Z(n5148) );
endmodule

